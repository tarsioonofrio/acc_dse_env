-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        -- replace ADDR_WIDHT, INPUT_SIZE and ADDRESS_SIZE generics with constants using python
        ADDR_WIDHT      : integer := 10;
        INPUT_SIZE      : integer := 8;
        ADDRESS_SIZE    : integer := 12;

        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(ADDRESS_SIZE-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(4-1 downto 0);
    signal bram_addr     : std_logic_vector(10-1 downto 0);

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(10-1 downto 0);
          

    MEM_IFMAP_LAYER0_ENTITY0 : if BRAM_NAME = "ifmap_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000a20000009c000000a0000000a6000000a50000009f0000009e",
            INIT_01 => X"000000aa000000a9000000a6000000a1000000a0000000a10000009f0000009e",
            INIT_02 => X"0000009400000096000000950000009c000000a0000000a0000000a2000000a7",
            INIT_03 => X"000000740000007e000000890000008f0000008d0000008c0000008f00000095",
            INIT_04 => X"000000a2000000a4000000a0000000a2000000a60000009f0000009700000098",
            INIT_05 => X"000000ab000000ab000000aa000000a30000009f0000009b0000009c000000a3",
            INIT_06 => X"0000008d0000008c0000008b00000091000000970000009a000000a0000000a9",
            INIT_07 => X"000000770000007d000000880000008f0000008e000000910000009300000095",
            INIT_08 => X"000000a5000000a5000000a3000000a0000000a70000009e0000009700000097",
            INIT_09 => X"000000a9000000a7000000a6000000a10000009d0000009e000000a2000000a3",
            INIT_0A => X"0000007200000065000000620000006e00000079000000910000009f000000aa",
            INIT_0B => X"00000078000000820000008b0000008e0000008c0000008f0000008600000078",
            INIT_0C => X"000000a9000000a9000000a7000000a7000000ae000000a00000009b0000009b",
            INIT_0D => X"000000a4000000a20000009d000000b1000000bf000000a7000000a5000000a5",
            INIT_0E => X"0000004a000000500000005c000000620000006700000068000000950000009e",
            INIT_0F => X"0000007f000000880000008c0000008c00000084000000710000005300000056",
            INIT_10 => X"000000a6000000a9000000a3000000a9000000aa000000a10000009c0000009b",
            INIT_11 => X"0000008e0000009200000097000000c3000000f6000000ad000000a4000000a4",
            INIT_12 => X"0000005d000000610000006a0000007000000071000000550000004e0000006f",
            INIT_13 => X"00000081000000850000008a000000800000006900000055000000540000004a",
            INIT_14 => X"000000a7000000a7000000a5000000a100000093000000820000008500000094",
            INIT_15 => X"0000004200000061000000800000009d000000b4000000a3000000a5000000a3",
            INIT_16 => X"0000005e00000072000000770000007a00000076000000590000004200000045",
            INIT_17 => X"000000860000008a0000008c0000006c000000430000003a0000005b00000063",
            INIT_18 => X"000000aa000000a8000000aa00000099000000580000002f0000006d0000007f",
            INIT_19 => X"00000044000000640000007f0000008100000093000000a4000000a6000000a9",
            INIT_1A => X"0000006b000000690000007c000000920000008400000053000000480000004e",
            INIT_1B => X"000000860000008d000000840000004f0000002e0000003f0000005500000073",
            INIT_1C => X"000000a8000000a5000000a70000008f000000460000002a0000006300000083",
            INIT_1D => X"00000058000000740000009000000082000000780000008c000000a1000000ab",
            INIT_1E => X"0000006a0000006600000088000000a30000007c0000004d000000550000005b",
            INIT_1F => X"000000880000008a0000006b0000003900000031000000360000005500000064",
            INIT_20 => X"000000a6000000a3000000a1000000990000007c0000003600000067000000aa",
            INIT_21 => X"00000056000000790000009c0000009d0000007d00000071000000ae000000a5",
            INIT_22 => X"0000005700000071000000920000008a00000051000000500000005400000052",
            INIT_23 => X"00000089000000850000004a0000002800000038000000470000005600000053",
            INIT_24 => X"000000990000009c0000009e000000ae0000009a0000005e00000086000000b4",
            INIT_25 => X"0000005d0000007d00000094000000ae0000009c000000cf000000ed000000cf",
            INIT_26 => X"0000006a000000850000008f000000890000004c0000003b0000004a00000056",
            INIT_27 => X"000000840000005f00000028000000320000004b000000540000005700000056",
            INIT_28 => X"0000007a0000009f0000009b000000b1000000a50000008e0000006c000000b7",
            INIT_29 => X"000000780000007d0000009c000000b7000000a4000000dc000000ed000000d5",
            INIT_2A => X"0000006b0000009b0000009d000000af0000005b0000002d000000500000004e",
            INIT_2B => X"000000680000003b000000290000003b0000004e000000580000006700000057",
            INIT_2C => X"00000086000000ad000000a6000000bb000000aa0000008700000064000000bc",
            INIT_2D => X"0000007500000086000000bd000000b9000000aa000000c7000000c200000075",
            INIT_2E => X"0000005d00000092000000a0000000d20000007d000000260000005400000066",
            INIT_2F => X"0000004c0000003e000000370000004900000055000000680000005e00000053",
            INIT_30 => X"0000009f000000b2000000a6000000ae000000af0000007f0000005a000000bd",
            INIT_31 => X"0000007b000000a0000000d8000000ba00000089000000a8000000a800000061",
            INIT_32 => X"0000005b0000007b0000009b000000c200000096000000320000007300000078",
            INIT_33 => X"000000490000004f0000004900000054000000560000005f0000005400000054",
            INIT_34 => X"000000a7000000ad0000008800000077000000b9000000980000005d000000bd",
            INIT_35 => X"0000008d000000b4000000e2000000bd000000a7000000910000009300000067",
            INIT_36 => X"000000570000007200000095000000ba0000009a00000047000000750000007e",
            INIT_37 => X"0000005e000000610000005a0000006400000063000000500000004800000050",
            INIT_38 => X"000000a70000009c0000006300000069000000ba000000a80000006c000000c2",
            INIT_39 => X"0000009a00000091000000ac000000be000000c60000008a0000007300000064",
            INIT_3A => X"0000006e0000008200000089000000b300000098000000470000006700000092",
            INIT_3B => X"000000750000006100000064000000730000006d0000005f0000005b00000055",
            INIT_3C => X"0000009b0000008c0000004e00000082000000b8000000ac00000084000000c5",
            INIT_3D => X"000000830000008700000091000000f2000000e60000008f0000008200000073",
            INIT_3E => X"000000570000007000000098000000a8000000900000005f0000006c00000079",
            INIT_3F => X"0000008800000079000000670000007800000070000000690000005700000047",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008a0000007e0000004e000000a8000000bf000000a800000092000000cb",
            INIT_41 => X"00000071000000710000008c000000a2000000ad0000009a000000600000008a",
            INIT_42 => X"0000006d00000087000000940000009c000000ab000000700000006900000065",
            INIT_43 => X"00000090000000970000007d0000006b000000650000005e0000004f0000004e",
            INIT_44 => X"0000009c000000600000005e000000b0000000b7000000a4000000a3000000d6",
            INIT_45 => X"0000007300000066000000740000007200000076000000810000006a00000094",
            INIT_46 => X"0000004b00000085000000800000004400000076000000900000006500000056",
            INIT_47 => X"0000008c000000960000008f0000007400000066000000470000003a0000003c",
            INIT_48 => X"0000008d000000560000007c000000b0000000ad000000a7000000b2000000d4",
            INIT_49 => X"00000093000000810000007c000000860000004d000000680000008700000099",
            INIT_4A => X"000000400000004b0000006b0000007500000084000000960000005c00000055",
            INIT_4B => X"000000970000009a000000a00000009b0000008500000056000000410000002c",
            INIT_4C => X"000000770000005600000090000000b1000000ae000000ab000000bb000000c7",
            INIT_4D => X"000000b8000000910000006c000000810000004600000090000000890000007a",
            INIT_4E => X"0000003400000033000000590000008600000089000000830000004900000074",
            INIT_4F => X"000000950000009e000000a4000000ab000000a3000000790000005a0000002f",
            INIT_50 => X"000000830000006300000098000000b5000000b1000000b3000000c3000000a5",
            INIT_51 => X"000000bf000000b20000007a0000005d000000500000005d00000067000000ab",
            INIT_52 => X"00000018000000260000002e0000003c00000057000000590000006400000096",
            INIT_53 => X"000000780000007f0000008000000090000000900000006c0000003c0000002e",
            INIT_54 => X"00000096000000530000008a000000b5000000b2000000b1000000c300000075",
            INIT_55 => X"000000c2000000be000000b0000000950000008600000085000000db000000f5",
            INIT_56 => X"0000003a0000003100000022000000230000003d0000006e0000007d000000a8",
            INIT_57 => X"000000370000003b000000450000004e00000048000000450000003a0000003d",
            INIT_58 => X"000000d30000006d0000008c000000b1000000b0000000ae000000af0000004f",
            INIT_59 => X"0000007a000000740000007c000000720000007c000000d0000000fc000000fd",
            INIT_5A => X"000000380000003300000032000000340000003c000000440000004400000068",
            INIT_5B => X"0000002a0000002b000000300000003b000000330000002b0000003300000038",
            INIT_5C => X"000000f6000000a5000000a5000000b2000000a8000000900000006000000029",
            INIT_5D => X"000000300000003100000031000000350000003c0000006e000000e3000000fd",
            INIT_5E => X"0000002b0000002e0000002e000000260000002a0000002e0000002a0000002d",
            INIT_5F => X"0000002d000000330000003500000037000000320000002e0000002e0000002a",
            INIT_60 => X"000000fe000000c200000084000000a6000000830000003b0000001d0000001d",
            INIT_61 => X"00000032000000310000003300000032000000320000003d0000008d000000f1",
            INIT_62 => X"0000002a00000026000000270000002300000022000000270000002a0000002f",
            INIT_63 => X"000000330000002e00000032000000380000003b0000003e000000380000002d",
            INIT_64 => X"00000100000000d7000000800000008000000049000000220000001e00000030",
            INIT_65 => X"0000002d0000002e0000003400000034000000320000003600000042000000bb",
            INIT_66 => X"0000002e0000002b00000028000000280000002700000024000000290000002b",
            INIT_67 => X"000000530000004600000032000000360000003b000000400000003e0000003b",
            INIT_68 => X"000000f0000000e00000008000000042000000290000001f0000002300000034",
            INIT_69 => X"0000002f0000002c0000002c0000003600000038000000310000003a0000007c",
            INIT_6A => X"0000003a000000360000002d0000002c0000002c0000002b0000002b0000002e",
            INIT_6B => X"0000004c000000550000004900000033000000240000002b0000002e00000036",
            INIT_6C => X"000000d3000000ca0000004e0000002c000000230000001d0000002300000032",
            INIT_6D => X"0000002d00000028000000300000003a00000030000000360000004100000061",
            INIT_6E => X"000000300000002700000027000000330000002e0000002f000000300000002f",
            INIT_6F => X"000000330000002e0000004300000043000000280000001c000000270000002f",
            INIT_70 => X"000000aa000000680000002e0000002900000021000000200000002300000032",
            INIT_71 => X"0000002d000000360000003a0000003d00000035000000340000003600000040",
            INIT_72 => X"00000027000000280000002a0000002e000000310000002e000000290000002a",
            INIT_73 => X"000000330000000f0000001f0000002f0000003f0000002c0000002800000025",
            INIT_74 => X"000000470000002a0000002b00000025000000260000001f0000002a00000044",
            INIT_75 => X"000000350000003a0000003800000031000000260000001b0000001f00000031",
            INIT_76 => X"00000021000000270000002d0000003200000035000000390000003c00000038",
            INIT_77 => X"000000280000000d0000002600000038000000490000004f0000003e0000002a",
            INIT_78 => X"000000280000002c0000002a000000270000002b00000023000000310000003d",
            INIT_79 => X"0000002f000000240000001d0000001b0000001e000000170000001b0000002a",
            INIT_7A => X"0000002b0000002b00000031000000450000004b000000420000003e00000038",
            INIT_7B => X"000000140000001d0000001a0000003c0000005d0000006d000000550000003c",
            INIT_7C => X"000000260000002800000028000000280000002b0000002d0000003800000036",
            INIT_7D => X"00000012000000130000001d000000190000001d000000160000001a00000024",
            INIT_7E => X"0000002d0000003400000035000000420000004a0000003d0000002f00000020",
            INIT_7F => X"0000001500000022000000180000003000000059000000690000005900000043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY1 : if BRAM_NAME = "ifmap_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000071000000730000006d0000007000000076000000740000006f00000070",
            INIT_01 => X"0000007700000075000000750000006f0000006f00000074000000710000006f",
            INIT_02 => X"0000006a0000006b0000006b0000006d000000700000006f0000007100000075",
            INIT_03 => X"000000550000005b0000005f000000610000006100000062000000650000006b",
            INIT_04 => X"0000007200000075000000710000007000000074000000720000006e00000070",
            INIT_05 => X"000000730000007500000077000000710000006e0000006f0000006e00000074",
            INIT_06 => X"0000006400000066000000680000006e00000073000000700000006f00000073",
            INIT_07 => X"000000580000005b0000005f0000006200000061000000660000006600000069",
            INIT_08 => X"0000007500000075000000730000006a0000006f0000006f0000006d0000006e",
            INIT_09 => X"0000007100000072000000730000006f0000006d000000720000007300000073",
            INIT_0A => X"000000550000004d0000004e0000005a000000600000006f0000007200000074",
            INIT_0B => X"000000590000005f000000620000006300000063000000670000006000000056",
            INIT_0C => X"0000007700000078000000750000006e000000700000006d0000006e0000006b",
            INIT_0D => X"00000072000000730000006f00000082000000920000007b0000007500000073",
            INIT_0E => X"0000003f0000004b0000005a0000005a00000057000000500000006f00000070",
            INIT_0F => X"0000005e00000063000000650000006600000062000000550000003e00000046",
            INIT_10 => X"000000740000007800000071000000720000007200000073000000720000006b",
            INIT_11 => X"0000006c0000006f000000720000009c000000d6000000800000007400000071",
            INIT_12 => X"0000005e00000066000000720000006e00000067000000450000003500000050",
            INIT_13 => X"0000005d0000005e000000650000006000000053000000490000004e00000048",
            INIT_14 => X"000000730000007400000071000000730000007000000064000000680000006d",
            INIT_15 => X"000000320000004b000000660000007a0000008a00000076000000740000006f",
            INIT_16 => X"00000060000000740000007a000000790000007100000053000000380000003a",
            INIT_17 => X"0000005f0000006200000069000000540000003a0000003a0000005b00000064",
            INIT_18 => X"000000760000007300000076000000750000004a000000250000005f00000064",
            INIT_19 => X"00000043000000570000006c000000620000006b000000780000007400000075",
            INIT_1A => X"0000006600000063000000760000008e00000082000000540000004b00000053",
            INIT_1B => X"0000005d00000063000000620000003d0000002f00000047000000530000006f",
            INIT_1C => X"0000007400000072000000750000006f000000400000002b0000006000000073",
            INIT_1D => X"000000570000006a000000830000006e0000005e0000006d0000007100000077",
            INIT_1E => X"000000620000005d0000007c00000099000000760000004d000000580000005f",
            INIT_1F => X"0000006100000067000000530000002f000000350000003c000000510000005d",
            INIT_20 => X"0000007a00000075000000710000007c000000790000003a00000069000000a1",
            INIT_21 => X"000000500000006f0000008f0000008d00000069000000590000008700000079",
            INIT_22 => X"0000004f00000067000000870000007d000000470000004e0000005500000051",
            INIT_23 => X"000000670000006a0000003b000000230000003900000049000000520000004d",
            INIT_24 => X"000000760000007400000074000000950000009a000000640000008b000000b0",
            INIT_25 => X"000000550000006e000000830000009900000083000000b4000000d6000000b4",
            INIT_26 => X"000000620000007c000000850000007d00000044000000390000004a00000054",
            INIT_27 => X"000000670000004b0000001e000000310000004c000000550000005500000051",
            INIT_28 => X"0000005900000076000000700000009c000000a90000009700000074000000b7",
            INIT_29 => X"0000006f0000006c000000890000009f00000087000000bf000000e0000000c5",
            INIT_2A => X"000000640000009300000093000000a5000000550000002c000000500000004c",
            INIT_2B => X"000000510000002e000000240000003b0000004f000000580000006600000053",
            INIT_2C => X"0000005d0000007b00000078000000a7000000af000000900000006c000000bf",
            INIT_2D => X"0000006b00000077000000ab000000a10000008e000000ab000000b60000005f",
            INIT_2E => X"000000590000008b00000098000000c900000079000000260000005400000062",
            INIT_2F => X"0000003800000037000000350000004b00000057000000680000005d00000050",
            INIT_30 => X"0000006d0000007b0000007b0000009c000000b40000008600000060000000c2",
            INIT_31 => X"0000007100000095000000ca000000a600000072000000900000009a00000044",
            INIT_32 => X"000000580000007600000095000000bb00000093000000320000007200000072",
            INIT_33 => X"000000370000004a0000004900000057000000570000005f0000005400000053",
            INIT_34 => X"000000740000007c0000006a0000006e000000bc0000009a0000005f000000c0",
            INIT_35 => X"00000083000000ac000000d8000000ae000000950000007d0000008400000048",
            INIT_36 => X"000000550000006e00000090000000b500000098000000470000007200000075",
            INIT_37 => X"0000004900000059000000580000006500000064000000500000004900000050",
            INIT_38 => X"0000007a00000077000000590000006d000000ba000000a70000006b000000c4",
            INIT_39 => X"0000008f0000008c000000a5000000b4000000b90000007b0000006a0000004a",
            INIT_3A => X"0000006d0000008000000085000000af00000098000000470000006400000088",
            INIT_3B => X"0000005f0000005500000060000000740000006e000000600000005d00000056",
            INIT_3C => X"0000007d000000780000005300000089000000b2000000a700000081000000c5",
            INIT_3D => X"00000079000000820000008a000000ec000000dd00000083000000780000005e",
            INIT_3E => X"000000550000006c000000930000009f00000086000000580000006800000070",
            INIT_3F => X"0000006800000060000000560000006e0000006d000000680000005800000048",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007e0000007d00000056000000aa000000b6000000a400000092000000cb",
            INIT_41 => X"0000006a0000006a0000008400000098000000a30000008f0000005000000079",
            INIT_42 => X"00000069000000820000008d0000008a0000008f0000005a0000006500000065",
            INIT_43 => X"000000680000006c00000058000000530000005b0000005d0000004f0000004c",
            INIT_44 => X"000000950000006000000066000000b6000000b8000000a7000000a6000000d7",
            INIT_45 => X"0000006e0000005b000000690000006600000069000000740000005d00000089",
            INIT_46 => X"000000450000007e00000078000000380000006000000080000000670000005b",
            INIT_47 => X"0000006e00000074000000700000005e0000005d000000460000003800000038",
            INIT_48 => X"0000008b0000005800000083000000b8000000b5000000af000000b8000000d3",
            INIT_49 => X"0000008f000000750000006f00000079000000400000005a0000008000000094",
            INIT_4A => X"0000003b00000044000000630000006d000000750000008b000000600000005c",
            INIT_4B => X"0000006f00000073000000780000007700000069000000450000003e00000029",
            INIT_4C => X"000000790000005a00000095000000b6000000b3000000b0000000bd000000c0",
            INIT_4D => X"000000b00000008600000061000000760000003b00000086000000880000007c",
            INIT_4E => X"000000330000003100000056000000810000007c000000770000004b00000076",
            INIT_4F => X"0000006b0000006f0000007100000079000000760000005b0000005a00000031",
            INIT_50 => X"00000087000000670000009d000000b5000000ad000000b2000000c10000009c",
            INIT_51 => X"000000b6000000ad000000760000005a0000004d0000005a00000069000000af",
            INIT_52 => X"000000210000002e000000340000003d0000004d0000004e0000006400000094",
            INIT_53 => X"00000069000000710000006d0000007b0000007d000000640000004700000039",
            INIT_54 => X"000000990000005700000090000000b3000000a9000000b2000000c800000078",
            INIT_55 => X"000000c0000000c4000000b60000009c0000008d0000008c000000de000000f7",
            INIT_56 => X"000000510000004600000036000000310000003e0000006d00000085000000ac",
            INIT_57 => X"0000005a0000005c000000600000006800000065000000630000005400000055",
            INIT_58 => X"000000d30000007000000092000000b1000000ac000000b7000000c500000069",
            INIT_59 => X"00000085000000850000008d000000840000008f000000e0000000fd000000fc",
            INIT_5A => X"0000005d00000055000000540000005400000052000000570000005d0000007c",
            INIT_5B => X"0000005f00000061000000610000006c00000068000000600000005b0000005e",
            INIT_5C => X"000000f5000000a6000000aa000000b6000000ae000000a80000008900000059",
            INIT_5D => X"000000480000004b0000004c000000500000005800000088000000e7000000fb",
            INIT_5E => X"00000057000000590000005a000000560000005200000051000000510000004f",
            INIT_5F => X"0000005a0000005f0000005e00000060000000600000005e0000005d00000059",
            INIT_60 => X"000000fa000000bd00000088000000b30000009900000066000000570000005b",
            INIT_61 => X"00000054000000530000005500000054000000540000005e0000009f000000f5",
            INIT_62 => X"000000590000005500000056000000530000004f000000520000005400000056",
            INIT_63 => X"000000670000005e00000063000000660000006500000067000000670000005c",
            INIT_64 => X"000000fd000000d500000088000000940000006a000000550000005e0000006f",
            INIT_65 => X"00000052000000530000005a0000005a000000580000005b0000005d000000c6",
            INIT_66 => X"0000005f0000005c000000590000005600000053000000500000005100000052",
            INIT_67 => X"000000890000007b000000690000006c0000006c0000006d0000006e0000006c",
            INIT_68 => X"000000f5000000e5000000910000005f00000053000000560000006300000072",
            INIT_69 => X"0000005300000052000000520000005c0000005e000000570000005c0000008f",
            INIT_6A => X"0000006e0000006a000000610000005a00000058000000560000005300000054",
            INIT_6B => X"0000007d0000008a000000820000006c0000005b0000005f0000006100000069",
            INIT_6C => X"000000e4000000db0000006a000000530000005600000059000000620000006e",
            INIT_6D => X"00000052000000500000005700000061000000570000005e000000680000007e",
            INIT_6E => X"000000660000005d0000005c0000006100000059000000590000005700000054",
            INIT_6F => X"00000060000000620000007e0000008100000065000000550000005d00000065",
            INIT_70 => X"000000c5000000850000005400000058000000580000005c000000610000006c",
            INIT_71 => X"000000530000006000000064000000670000005f0000005e0000006100000064",
            INIT_72 => X"0000005c0000005d0000005f0000005c0000005c00000058000000500000004f",
            INIT_73 => X"0000005d0000003c0000005a0000006e0000007d000000660000005d0000005a",
            INIT_74 => X"0000006b0000004f00000059000000570000005b00000058000000640000007c",
            INIT_75 => X"0000005c00000066000000640000005d00000052000000470000004d00000059",
            INIT_76 => X"00000053000000580000005e0000005f0000006100000063000000630000005e",
            INIT_77 => X"000000550000004000000061000000740000008300000084000000700000005b",
            INIT_78 => X"00000051000000580000005c0000005a0000005b000000550000006600000074",
            INIT_79 => X"000000560000005000000049000000470000004a000000430000004800000055",
            INIT_7A => X"00000058000000580000005f00000071000000770000006d000000650000005f",
            INIT_7B => X"00000040000000520000005200000073000000910000009c0000008200000069",
            INIT_7C => X"00000051000000570000005c000000590000005600000059000000690000006b",
            INIT_7D => X"0000003a0000003f00000049000000450000004900000042000000450000004f",
            INIT_7E => X"000000570000005f000000600000006f00000077000000680000005700000046",
            INIT_7F => X"00000043000000540000004d000000630000008700000092000000830000006d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY1;


    MEM_IFMAP_LAYER0_ENTITY2 : if BRAM_NAME = "ifmap_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d0000002f000000290000002e00000035000000330000002f00000031",
            INIT_01 => X"0000002c0000002d00000029000000310000003400000029000000290000002c",
            INIT_02 => X"0000002b0000002d0000002d0000002c0000002b000000270000002600000028",
            INIT_03 => X"00000021000000240000002400000026000000290000002b000000270000002c",
            INIT_04 => X"0000002d0000002f0000002b00000031000000380000002d0000002800000033",
            INIT_05 => X"000000210000002800000029000000340000003600000029000000260000002e",
            INIT_06 => X"000000300000003400000037000000350000003200000029000000210000001e",
            INIT_07 => X"00000022000000200000001f00000022000000260000002d0000002e00000032",
            INIT_08 => X"0000002d0000002d0000002c0000002a0000003000000024000000210000002f",
            INIT_09 => X"0000002300000025000000260000003300000039000000300000002b0000002b",
            INIT_0A => X"000000320000002f000000320000003400000031000000360000002f00000027",
            INIT_0B => X"0000002100000022000000220000002300000027000000330000003700000030",
            INIT_0C => X"00000030000000300000002e0000002b0000002c0000001f0000002000000028",
            INIT_0D => X"000000360000002f000000290000004b0000005f000000390000002d0000002c",
            INIT_0E => X"0000003200000042000000540000004c000000410000002f000000430000003a",
            INIT_0F => X"0000002400000027000000270000002b0000002e0000002d0000002700000034",
            INIT_10 => X"0000002c0000002f000000280000002b0000002f000000310000003000000029",
            INIT_11 => X"000000470000003c000000380000006b000000a40000003b0000002a00000029",
            INIT_12 => X"0000005d00000069000000760000006f00000062000000380000001f00000032",
            INIT_13 => X"00000024000000240000002e000000300000002d0000002f0000004600000043",
            INIT_14 => X"0000002900000029000000270000002c00000035000000390000004000000036",
            INIT_15 => X"0000001f0000002b0000003a0000004e000000550000002a0000002700000025",
            INIT_16 => X"00000060000000740000007a000000780000006e0000004c0000002d0000002b",
            INIT_17 => X"000000280000002c0000003a00000031000000250000002f0000005600000061",
            INIT_18 => X"0000002b000000280000002b000000300000001c000000110000005000000039",
            INIT_19 => X"00000039000000460000004b0000003b0000003400000027000000250000002a",
            INIT_1A => X"0000005e0000005a0000006c00000084000000790000004a0000004000000048",
            INIT_1B => X"00000027000000300000003a0000002400000027000000450000004d00000067",
            INIT_1C => X"00000027000000240000002a0000003800000029000000260000005c0000005a",
            INIT_1D => X"0000004f0000005d0000006b0000004d00000031000000330000003300000031",
            INIT_1E => X"0000005800000051000000700000008c0000006b000000450000005200000058",
            INIT_1F => X"00000027000000330000003200000020000000310000003a0000004a00000054",
            INIT_20 => X"00000032000000290000002b00000052000000710000003b0000006900000090",
            INIT_21 => X"0000004a0000006500000080000000790000004e0000003b0000005f00000042",
            INIT_22 => X"000000460000005d0000007b000000700000003d00000049000000520000004d",
            INIT_23 => X"0000002d0000003b000000230000001b00000035000000430000004c00000045",
            INIT_24 => X"0000003c0000002f000000330000007000000095000000690000008f000000a3",
            INIT_25 => X"0000004f0000006b0000007d0000009100000077000000a6000000c600000092",
            INIT_26 => X"00000059000000720000007a000000700000003a00000035000000470000004f",
            INIT_27 => X"000000390000002c0000000f0000002b000000470000004e0000004e0000004a",
            INIT_28 => X"0000002f00000033000000320000007a000000a80000009e0000007a000000af",
            INIT_29 => X"0000006800000068000000840000009b00000083000000bc000000e2000000b3",
            INIT_2A => X"0000005c0000008a000000890000009a0000004d000000280000004d00000045",
            INIT_2B => X"0000002e0000001f000000210000003b000000490000004f000000600000004d",
            INIT_2C => X"0000002c000000370000003b00000088000000b20000009900000074000000bd",
            INIT_2D => X"0000005f0000006a0000009f0000009700000085000000a4000000bc00000050",
            INIT_2E => X"00000052000000820000008e000000c000000071000000220000004f00000059",
            INIT_2F => X"0000001a00000030000000370000004e000000510000005e000000580000004b",
            INIT_30 => X"0000002f000000350000004400000085000000b90000009000000069000000c2",
            INIT_31 => X"0000006200000081000000b7000000940000005e0000007e000000980000002c",
            INIT_32 => X"000000530000006f0000008c000000b20000008c0000002f0000006d00000069",
            INIT_33 => X"000000180000004000000049000000590000005100000055000000500000004f",
            INIT_34 => X"000000320000003a0000004200000062000000c0000000a300000067000000c1",
            INIT_35 => X"000000750000009d000000c80000009b0000007f000000670000007800000027",
            INIT_36 => X"000000500000006800000088000000ae00000093000000440000006d0000006b",
            INIT_37 => X"000000220000004500000051000000630000005e00000048000000460000004c",
            INIT_38 => X"000000370000003e000000430000006d000000bc000000ac00000070000000c4",
            INIT_39 => X"000000860000008c0000009f000000a9000000a9000000670000005800000022",
            INIT_3A => X"000000690000007a0000007f000000aa00000095000000460000005f0000007d",
            INIT_3B => X"0000002f00000035000000500000006f000000680000005a0000005b00000053",
            INIT_3C => X"0000004d000000580000004d0000008e000000b5000000ae00000088000000c5",
            INIT_3D => X"000000700000008200000089000000e6000000d3000000740000005d00000034",
            INIT_3E => X"00000050000000650000008a00000092000000760000004b0000005f00000065",
            INIT_3F => X"0000003000000030000000360000005d00000063000000630000005700000044",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000710000007e0000005a000000ac000000bc000000b2000000a0000000cc",
            INIT_41 => X"0000005a00000058000000750000008d0000009b000000850000002500000052",
            INIT_42 => X"00000061000000760000007e0000006d000000680000003a000000570000005c",
            INIT_43 => X"0000002e000000370000002d00000037000000520000005e0000004d00000048",
            INIT_44 => X"000000910000006600000069000000ba000000c2000000b8000000b4000000d7",
            INIT_45 => X"000000620000004900000059000000590000005f000000690000003d0000006f",
            INIT_46 => X"0000003d00000073000000690000002000000040000000660000005f00000058",
            INIT_47 => X"000000360000004000000044000000400000004e000000410000003500000033",
            INIT_48 => X"0000008f0000006000000085000000bc000000c1000000bd000000c0000000cd",
            INIT_49 => X"0000008500000064000000600000006c00000037000000500000006f0000008d",
            INIT_4A => X"000000340000003a000000560000005c0000005d000000780000005d0000005d",
            INIT_4B => X"0000002e0000002d000000360000003e0000003b000000280000003c00000027",
            INIT_4C => X"000000840000006300000098000000b8000000b9000000b5000000bb000000b4",
            INIT_4D => X"000000a80000007b000000560000006c000000330000007e0000008700000082",
            INIT_4E => X"000000320000002c0000004e0000007600000069000000670000004900000076",
            INIT_4F => X"0000002e000000320000003400000040000000440000003c0000005d00000034",
            INIT_50 => X"000000920000006f000000a0000000b4000000ac000000af000000bb00000092",
            INIT_51 => X"000000b1000000ad000000740000005600000049000000570000006f000000b9",
            INIT_52 => X"000000290000003300000036000000390000003f000000420000006500000094",
            INIT_53 => X"0000003f000000450000003d0000004c000000520000004b0000005300000045",
            INIT_54 => X"0000009f0000005b00000093000000b3000000a8000000b0000000c80000007c",
            INIT_55 => X"000000c5000000d0000000c0000000a40000009300000090000000e1000000fa",
            INIT_56 => X"0000006600000057000000440000003a0000003e0000006d0000008f000000b5",
            INIT_57 => X"00000073000000700000007000000078000000770000007a0000006f0000006e",
            INIT_58 => X"000000d10000007100000096000000b6000000b1000000c0000000d500000085",
            INIT_59 => X"000000980000009c000000a2000000950000009d000000e8000000fc000000f7",
            INIT_5A => X"0000007d000000730000006e0000006f00000065000000680000007700000094",
            INIT_5B => X"0000008400000089000000840000008e0000008d000000870000008200000083",
            INIT_5C => X"000000ed000000a4000000ae000000c0000000bc000000bc000000a800000087",
            INIT_5D => X"000000650000006b00000069000000690000006f00000099000000e4000000f1",
            INIT_5E => X"000000800000007e0000007d0000007d00000074000000710000007800000073",
            INIT_5F => X"000000850000008b000000860000008700000089000000890000008b00000084",
            INIT_60 => X"000000f2000000b500000089000000bf000000b000000086000000820000008d",
            INIT_61 => X"00000074000000780000007900000077000000760000007f000000af000000f5",
            INIT_62 => X"000000820000007d0000007d0000007800000071000000730000007500000075",
            INIT_63 => X"000000950000008c00000090000000920000008e0000008e0000009100000086",
            INIT_64 => X"000000f9000000d10000008f000000a7000000880000007c0000008c000000a2",
            INIT_65 => X"00000073000000790000007f0000007f0000007d0000008000000076000000cd",
            INIT_66 => X"0000008a00000086000000830000007b00000075000000710000007000000071",
            INIT_67 => X"000000b6000000a7000000980000009a00000095000000930000009800000096",
            INIT_68 => X"000000f7000000ea000000a40000007e0000007a0000008200000093000000a5",
            INIT_69 => X"00000077000000770000007700000081000000830000007b0000007200000099",
            INIT_6A => X"0000009a000000960000008d000000830000007f0000007b0000007700000077",
            INIT_6B => X"000000a9000000b6000000b20000009e0000008a0000008c0000008d00000096",
            INIT_6C => X"000000ea000000e90000008a0000007e000000850000008a00000095000000a2",
            INIT_6D => X"00000077000000740000007b000000850000007c000000810000007e0000008c",
            INIT_6E => X"000000940000008b0000008a0000008c00000084000000820000007e0000007a",
            INIT_6F => X"0000008b0000008e000000b0000000b600000099000000850000008b00000093",
            INIT_70 => X"000000d30000009f0000007d0000008a0000008d0000008f00000093000000a1",
            INIT_71 => X"0000007800000083000000870000008b00000082000000800000007900000077",
            INIT_72 => X"000000880000008a0000008b0000008800000087000000820000007800000076",
            INIT_73 => X"00000088000000670000008c000000a4000000b2000000970000008a00000087",
            INIT_74 => X"0000008500000071000000840000008b000000920000008900000094000000b1",
            INIT_75 => X"0000008000000089000000870000008000000075000000690000006900000072",
            INIT_76 => X"0000007d0000008300000088000000890000008a0000008b0000008900000083",
            INIT_77 => X"0000007f0000006c00000092000000a8000000b5000000b30000009a00000085",
            INIT_78 => X"000000700000007d000000860000008b0000008f0000008400000094000000a8",
            INIT_79 => X"00000078000000730000006c0000006a0000006d000000660000006800000073",
            INIT_7A => X"0000007f0000007f00000086000000980000009c000000900000008700000080",
            INIT_7B => X"0000006b0000007e00000082000000a4000000be000000c5000000aa00000090",
            INIT_7C => X"000000730000007b0000008400000086000000860000008400000095000000a0",
            INIT_7D => X"00000059000000620000006c000000680000006c000000650000006900000072",
            INIT_7E => X"0000007b00000082000000830000009100000098000000890000007600000064",
            INIT_7F => X"0000006e000000810000007c00000091000000af000000b6000000a700000091",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY2;


    MEM_IFMAP_LAYER0_ENTITY3 : if BRAM_NAME = "ifmap_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e8000000e8000000e8000000e8000000e8000000e8000000e7000000eb",
            INIT_01 => X"000000e9000000e9000000e9000000e9000000e9000000e9000000e8000000e8",
            INIT_02 => X"000000e9000000e8000000e8000000e8000000e6000000e7000000e8000000e9",
            INIT_03 => X"000000e8000000e9000000e9000000e8000000e8000000e8000000e9000000e8",
            INIT_04 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_05 => X"000000ec000000ec000000ec000000ec000000ec000000ec000000eb000000eb",
            INIT_06 => X"000000ec000000eb000000ea000000ea000000ea000000ec000000ec000000ed",
            INIT_07 => X"000000eb000000ec000000ec000000eb000000eb000000eb000000ec000000ec",
            INIT_08 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000ea000000ed",
            INIT_09 => X"000000eb000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0A => X"000000ea000000e7000000e7000000e3000000ea000000eb000000ec000000ec",
            INIT_0B => X"000000ea000000eb000000eb000000ea000000ea000000ea000000ea000000ea",
            INIT_0C => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_0D => X"000000eb000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0E => X"000000e4000000cf000000d1000000ba000000df000000e4000000e8000000e9",
            INIT_0F => X"000000eb000000eb000000eb000000ea000000ea000000ea000000ea000000ec",
            INIT_10 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000ea000000ed",
            INIT_11 => X"000000eb000000eb000000ea000000ea000000eb000000eb000000ea000000ea",
            INIT_12 => X"000000e6000000d6000000c3000000a3000000cb000000db000000e9000000ec",
            INIT_13 => X"000000ec000000ec000000ec000000eb000000eb000000eb000000eb000000ed",
            INIT_14 => X"000000eb000000eb000000ec000000ec000000ec000000ec000000ec000000ef",
            INIT_15 => X"000000e5000000eb000000e8000000ea000000ed000000ed000000eb000000ea",
            INIT_16 => X"000000e2000000cf000000b8000000a5000000ae000000b9000000c2000000d0",
            INIT_17 => X"000000ed000000ed000000ed000000ec000000ec000000ec000000ec000000ec",
            INIT_18 => X"000000ec000000ed000000ed000000ea000000e7000000e8000000e4000000e4",
            INIT_19 => X"000000dd000000e9000000e0000000e1000000ef000000ef000000ed000000ed",
            INIT_1A => X"000000c60000009c0000008f000000900000009a0000009f000000a1000000b7",
            INIT_1B => X"000000ef000000ed000000ec000000eb000000eb000000eb000000ec000000e9",
            INIT_1C => X"000000ee000000ed000000ea000000e5000000e3000000e6000000e0000000d4",
            INIT_1D => X"000000d6000000e9000000db000000c9000000f0000000ef000000ef000000ef",
            INIT_1E => X"000000ba000000a20000009f000000a5000000ad000000b8000000b9000000c1",
            INIT_1F => X"000000ee000000ed000000ec000000ea000000e9000000e9000000ea000000e5",
            INIT_20 => X"000000ee000000ec000000e7000000e3000000e1000000e1000000dd000000d8",
            INIT_21 => X"000000e6000000e9000000dc000000c5000000ef000000ed000000ee000000ee",
            INIT_22 => X"000000da000000d9000000d2000000d1000000d0000000db000000d1000000d1",
            INIT_23 => X"000000ee000000ed000000eb000000e6000000e6000000e4000000e4000000e1",
            INIT_24 => X"000000ed000000eb000000e1000000ac000000880000007c0000007700000076",
            INIT_25 => X"000000ec000000e8000000e2000000d6000000e9000000eb000000eb000000ec",
            INIT_26 => X"000000b9000000c9000000d9000000e1000000e1000000e7000000e3000000e4",
            INIT_27 => X"000000ee000000ec000000eb000000df000000ba000000a7000000a7000000ac",
            INIT_28 => X"000000e5000000e3000000de000000920000006f0000006c000000670000006d",
            INIT_29 => X"000000e6000000e8000000e7000000e5000000e6000000e7000000ea000000ec",
            INIT_2A => X"0000008900000092000000a4000000bf000000df000000e5000000e7000000e7",
            INIT_2B => X"000000ed000000eb000000ea000000d800000095000000790000008000000086",
            INIT_2C => X"000000d3000000d5000000df000000d1000000c8000000c7000000bc000000c3",
            INIT_2D => X"000000dc000000d8000000d3000000d1000000d2000000db000000dc000000d8",
            INIT_2E => X"000000b2000000b5000000af000000b7000000da000000e1000000e2000000e1",
            INIT_2F => X"000000ec000000ea000000e7000000db000000b90000008e000000aa000000ba",
            INIT_30 => X"000000ab000000cb000000d6000000df000000d6000000ca000000bf000000c1",
            INIT_31 => X"0000007a0000006f000000650000005d00000062000000ae000000cf000000b1",
            INIT_32 => X"000000d9000000df000000dc000000da000000df000000ca0000009900000089",
            INIT_33 => X"000000eb000000e8000000dd000000db000000de000000c4000000d4000000dd",
            INIT_34 => X"000000be000000bf000000aa0000008a0000007d000000710000006f00000071",
            INIT_35 => X"0000004200000035000000310000002d000000360000009e000000d8000000d0",
            INIT_36 => X"000000cf000000df000000e3000000e9000000ea000000dd0000009f00000066",
            INIT_37 => X"000000dd000000d3000000bc000000b3000000c7000000d4000000d3000000ca",
            INIT_38 => X"000000c3000000970000008b0000007b000000440000003f000000450000003d",
            INIT_39 => X"000000b50000008a000000650000005f00000067000000a3000000ce000000d6",
            INIT_3A => X"00000083000000930000009e000000b7000000cd000000db000000dd000000cf",
            INIT_3B => X"000000c5000000b60000008a000000800000008500000088000000820000007d",
            INIT_3C => X"000000a30000007700000060000000840000007f000000550000003a00000028",
            INIT_3D => X"000000c8000000da000000c6000000b7000000b5000000b6000000b8000000ad",
            INIT_3E => X"000000630000005e000000620000007400000084000000910000009f000000ae",
            INIT_3F => X"000000b9000000bc0000009d000000960000008a0000007a0000006b00000069",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac0000008d000000760000008a000000ce000000860000001a0000000d",
            INIT_41 => X"000000b0000000e2000000e6000000e0000000e4000000dc000000cf000000b5",
            INIT_42 => X"0000009a00000095000000950000009a000000910000008e0000008a00000090",
            INIT_43 => X"0000009d000000a5000000b2000000be000000bb000000ad000000a00000009d",
            INIT_44 => X"000000e2000000d4000000c7000000c5000000e1000000c80000003a00000005",
            INIT_45 => X"000000d2000000dd000000df000000d1000000e6000000e8000000e9000000e5",
            INIT_46 => X"000000b8000000c0000000c2000000bd000000bc000000c1000000b4000000c6",
            INIT_47 => X"0000008a00000080000000830000008800000090000000a1000000ab000000ac",
            INIT_48 => X"000000c2000000c2000000c0000000b8000000ba000000be0000009100000027",
            INIT_49 => X"000000930000009a000000b4000000b1000000be000000c0000000bf000000c2",
            INIT_4A => X"0000006f0000007e000000840000007200000071000000920000009c00000091",
            INIT_4B => X"000000810000008100000079000000690000005e0000005d0000005b0000005c",
            INIT_4C => X"000000820000007f0000008000000083000000890000008f000000a20000007a",
            INIT_4D => X"00000064000000680000007c00000081000000810000007f0000008000000083",
            INIT_4E => X"00000053000000570000005e0000005e0000005e000000700000007600000066",
            INIT_4F => X"0000008200000079000000730000006c000000650000005d0000005300000050",
            INIT_50 => X"0000005a000000570000005700000054000000500000004d0000004c00000049",
            INIT_51 => X"00000078000000760000007600000073000000710000006b000000660000005e",
            INIT_52 => X"000000500000004f000000550000005f000000640000006a0000006e00000073",
            INIT_53 => X"000000880000007d000000710000005c00000052000000500000004d00000050",
            INIT_54 => X"000000160000001400000015000000120000001200000009000000030000000d",
            INIT_55 => X"00000046000000420000003c00000034000000300000002a000000220000001a",
            INIT_56 => X"000000390000003500000035000000370000003c000000430000004800000047",
            INIT_57 => X"0000008900000082000000780000006800000057000000480000003900000039",
            INIT_58 => X"0000000300000008000000160000002400000020000000080000000b00000024",
            INIT_59 => X"0000000300000001000000050000000600000000000000000000000000000001",
            INIT_5A => X"000000270000001e00000016000000150000001500000015000000180000000d",
            INIT_5B => X"00000099000000860000007a000000740000007b000000710000005500000039",
            INIT_5C => X"0000001b0000003100000046000000470000001b0000000d0000001a00000023",
            INIT_5D => X"0000000a0000001f00000039000000110000000000000002000000050000000f",
            INIT_5E => X"000000560000003e00000029000000190000000e000000070000000400000004",
            INIT_5F => X"000000ac0000009200000084000000750000007200000084000000900000007a",
            INIT_60 => X"0000002400000036000000410000002d00000003000000040000000d00000010",
            INIT_61 => X"00000083000000a1000000760000000700000000000000020000000400000012",
            INIT_62 => X"000000970000009a0000008a000000760000006d000000690000006900000070",
            INIT_63 => X"000000b8000000a40000008e00000081000000780000006a000000690000007f",
            INIT_64 => X"00000015000000200000001e0000000c00000000000000000000000c00000028",
            INIT_65 => X"000000cd000000b6000000440000000000000003000000020000000200000007",
            INIT_66 => X"000000670000007b00000096000000ac000000bb000000c3000000c2000000c4",
            INIT_67 => X"000000b9000000ab0000009800000084000000810000007a000000680000005f",
            INIT_68 => X"0000000c000000120000000c0000000400000001000000010000001a00000045",
            INIT_69 => X"000000cb00000099000000200000000100000004000000020000000200000004",
            INIT_6A => X"0000005e000000510000005b000000770000009b000000b3000000bf000000c3",
            INIT_6B => X"000000b8000000ad000000a200000090000000810000007d0000007d00000075",
            INIT_6C => X"0000000400000007000000050000000200000002000000010000002f00000053",
            INIT_6D => X"000000cd0000008e0000001b0000000100000003000000010000000100000001",
            INIT_6E => X"0000007900000066000000550000004a0000005500000079000000a9000000c6",
            INIT_6F => X"000000ba000000b0000000a50000009300000084000000790000007a00000080",
            INIT_70 => X"000000010000000100000001000000020000000300000006000000360000005c",
            INIT_71 => X"0000009d000000660000000f0000000000000001000000010000000100000001",
            INIT_72 => X"0000007c0000007a00000073000000630000004a000000380000004a00000075",
            INIT_73 => X"000000bc000000b1000000a20000009400000088000000800000007d0000007b",
            INIT_74 => X"000000020000000200000005000000080000000b000000130000002b00000057",
            INIT_75 => X"000000470000002a000000040000000000000002000000030000000300000003",
            INIT_76 => X"000000740000007b000000860000008400000071000000500000003900000035",
            INIT_77 => X"000000bc000000b6000000a90000009c0000008f0000008b0000008300000078",
            INIT_78 => X"0000001000000011000000160000001b0000001f000000240000002e00000052",
            INIT_79 => X"0000004000000025000000170000001300000013000000140000001300000012",
            INIT_7A => X"0000007300000075000000830000008b00000080000000740000006800000057",
            INIT_7B => X"000000bb000000b9000000ae0000009f000000940000008b000000830000007b",
            INIT_7C => X"000000300000002e0000002f00000033000000370000003a0000003e00000055",
            INIT_7D => X"0000006800000051000000440000003b00000037000000350000003300000031",
            INIT_7E => X"0000007a00000072000000760000007f0000007f000000850000007f00000074",
            INIT_7F => X"000000ba000000b4000000a80000009e000000950000008d0000008800000081",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY3;


    MEM_IFMAP_LAYER0_ENTITY4 : if BRAM_NAME = "ifmap_layer0_entity4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e8000000e8000000e8000000e8000000e8000000e8000000e7000000eb",
            INIT_01 => X"000000e8000000e9000000e9000000e9000000e9000000e9000000e8000000e8",
            INIT_02 => X"000000e9000000e8000000e7000000e8000000e9000000e9000000e7000000e7",
            INIT_03 => X"000000e8000000e9000000e9000000e8000000e8000000e8000000e9000000e9",
            INIT_04 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_05 => X"000000ec000000ec000000ec000000ec000000ec000000ec000000eb000000eb",
            INIT_06 => X"000000ec000000ec000000ea000000eb000000ec000000ec000000ea000000ea",
            INIT_07 => X"000000eb000000ec000000ec000000eb000000eb000000eb000000ec000000ec",
            INIT_08 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000ea000000ed",
            INIT_09 => X"000000ea000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0A => X"000000ea000000e9000000eb000000e6000000eb000000eb000000ea000000e9",
            INIT_0B => X"000000ea000000eb000000eb000000ea000000ea000000ea000000ea000000ea",
            INIT_0C => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_0D => X"000000eb000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0E => X"000000e4000000d2000000d8000000c0000000e2000000e6000000e8000000e9",
            INIT_0F => X"000000eb000000eb000000eb000000ea000000ea000000ea000000ea000000eb",
            INIT_10 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000ea000000ed",
            INIT_11 => X"000000eb000000eb000000ea000000ea000000eb000000eb000000ea000000ea",
            INIT_12 => X"000000e5000000da000000cd000000ac000000d2000000e1000000ed000000ee",
            INIT_13 => X"000000ec000000ec000000ec000000ec000000eb000000eb000000eb000000eb",
            INIT_14 => X"000000eb000000ec000000eb000000eb000000eb000000eb000000eb000000ef",
            INIT_15 => X"000000e7000000ed000000e9000000eb000000ec000000ec000000eb000000ea",
            INIT_16 => X"000000e4000000d7000000c4000000b3000000bc000000c6000000cd000000d8",
            INIT_17 => X"000000ed000000ed000000ed000000ec000000ec000000ec000000ec000000eb",
            INIT_18 => X"000000ed000000ed000000ec000000e8000000e4000000e6000000e3000000e5",
            INIT_19 => X"000000e2000000ed000000e4000000e5000000ed000000ec000000eb000000eb",
            INIT_1A => X"000000ce000000a90000009f000000a3000000b0000000b4000000b4000000c5",
            INIT_1B => X"000000ed000000ed000000ee000000ec000000eb000000ec000000ed000000ee",
            INIT_1C => X"000000ed000000ee000000ed000000ea000000e8000000ea000000e6000000dc",
            INIT_1D => X"000000da000000ec000000de000000cc000000ee000000ec000000ed000000ed",
            INIT_1E => X"000000c7000000b0000000ae000000b6000000bf000000c9000000c9000000cc",
            INIT_1F => X"000000ee000000ef000000ef000000ef000000ee000000ee000000ef000000ef",
            INIT_20 => X"000000ec000000ed000000ee000000f0000000ef000000ee000000ec000000ea",
            INIT_21 => X"000000e7000000ea000000dd000000c6000000ef000000ed000000ec000000ec",
            INIT_22 => X"000000eb000000e9000000e0000000dd000000da000000e4000000d8000000d5",
            INIT_23 => X"000000ee000000f0000000f0000000f0000000f0000000ef000000ee000000f0",
            INIT_24 => X"000000ea000000ec000000ea000000bc0000009b0000008e0000008a0000008c",
            INIT_25 => X"000000ed000000ea000000e4000000d8000000ed000000ed000000eb000000e9",
            INIT_26 => X"000000cc000000db000000e9000000ed000000e8000000ec000000e6000000e6",
            INIT_27 => X"000000f0000000f0000000f1000000eb000000c7000000b4000000b3000000bd",
            INIT_28 => X"000000e2000000e4000000e50000009f0000007f0000007d0000007900000082",
            INIT_29 => X"000000eb000000ed000000eb000000ea000000ed000000ec000000ea000000e8",
            INIT_2A => X"0000009c000000a5000000b8000000ce000000e8000000ed000000ed000000ec",
            INIT_2B => X"000000f0000000f0000000f1000000e4000000a2000000850000008c00000095",
            INIT_2C => X"000000d1000000d5000000e3000000d9000000d3000000d3000000ca000000d4",
            INIT_2D => X"000000e5000000e1000000dd000000db000000dd000000e2000000de000000d5",
            INIT_2E => X"000000c2000000c8000000c6000000cc000000e7000000ed000000ec000000ea",
            INIT_2F => X"000000f0000000f1000000f0000000e6000000c300000097000000b2000000c5",
            INIT_30 => X"000000ae000000d0000000db000000e1000000d9000000d3000000ca000000cf",
            INIT_31 => X"0000008a00000081000000790000007200000070000000b8000000d5000000b4",
            INIT_32 => X"000000e2000000ea000000e9000000e8000000ec000000d8000000a700000098",
            INIT_33 => X"000000f1000000ef000000e6000000e3000000e6000000cb000000db000000e4",
            INIT_34 => X"000000c7000000c9000000b600000091000000830000007d0000007d00000082",
            INIT_35 => X"0000005400000049000000490000004600000047000000ac000000e6000000db",
            INIT_36 => X"000000d3000000e4000000e7000000ed000000ef000000e3000000a800000072",
            INIT_37 => X"000000e7000000dd000000c5000000ba000000ce000000db000000da000000d0",
            INIT_38 => X"000000c80000009d0000009b0000008d000000550000004f0000005600000051",
            INIT_39 => X"000000c000000097000000750000007000000079000000b4000000df000000e4",
            INIT_3A => X"0000008a0000009a000000a6000000ba000000cb000000db000000de000000d4",
            INIT_3B => X"000000d4000000c500000099000000890000008e000000920000008b00000085",
            INIT_3C => X"0000009e000000730000006b0000009700000090000000620000004600000035",
            INIT_3D => X"000000d2000000e4000000d1000000c2000000c1000000c2000000c2000000b4",
            INIT_3E => X"0000006f0000006a0000006f0000007d0000008800000096000000a5000000b5",
            INIT_3F => X"000000cb000000ce000000ae000000a400000097000000870000007900000076",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a2000000850000007b00000096000000d80000008c0000001d0000000f",
            INIT_41 => X"000000bd000000ee000000f1000000ea000000ea000000e0000000d1000000b5",
            INIT_42 => X"000000ab000000a5000000a5000000ab000000a30000009e0000009a0000009f",
            INIT_43 => X"000000af000000b7000000c4000000cf000000cc000000be000000b1000000ae",
            INIT_44 => X"000000e0000000d4000000cf000000cd000000e8000000cf0000003e00000005",
            INIT_45 => X"000000e4000000ee000000ee000000dd000000ee000000ee000000ec000000e6",
            INIT_46 => X"000000cc000000d4000000d6000000d4000000d5000000d8000000c8000000d9",
            INIT_47 => X"0000009a0000008f000000920000009c000000a5000000b5000000bf000000c1",
            INIT_48 => X"000000d0000000d3000000d3000000c5000000c4000000cc0000009b0000002d",
            INIT_49 => X"000000a9000000b0000000c6000000c1000000cf000000cf000000cb000000ce",
            INIT_4A => X"00000087000000960000009d0000008900000085000000a3000000ab000000a1",
            INIT_4B => X"0000008e0000008d000000850000007d00000074000000720000007000000073",
            INIT_4C => X"000000960000009600000098000000980000009a000000a0000000b300000087",
            INIT_4D => X"0000007a0000007e000000910000009500000095000000930000009300000096",
            INIT_4E => X"000000670000007000000075000000700000006d000000800000008600000078",
            INIT_4F => X"00000090000000850000007d00000079000000750000006f0000006700000061",
            INIT_50 => X"000000690000006600000066000000620000005d0000005a0000005a00000057",
            INIT_51 => X"00000085000000840000008800000089000000830000007c000000770000006f",
            INIT_52 => X"0000005c00000061000000650000006d000000770000007f0000008500000088",
            INIT_53 => X"000000950000008700000077000000680000006200000064000000640000005e",
            INIT_54 => X"0000001e00000019000000190000001a0000001a000000100000000b00000019",
            INIT_55 => X"0000004f0000004d0000004b000000450000003b000000330000002b00000024",
            INIT_56 => X"0000004500000045000000440000004300000048000000510000005800000057",
            INIT_57 => X"00000092000000880000007c0000007100000064000000590000004e00000047",
            INIT_58 => X"000000080000000b000000190000002d0000002c0000000d000000100000002e",
            INIT_59 => X"0000001700000013000000120000000d00000004000000020000000200000004",
            INIT_5A => X"0000003a000000320000002c000000260000001f00000021000000260000001d",
            INIT_5B => X"000000a00000008b0000007b000000730000007b000000730000005a00000046",
            INIT_5C => X"0000001f00000032000000460000005100000029000000130000001b00000029",
            INIT_5D => X"000000240000003200000040000000110000000000000002000000050000000f",
            INIT_5E => X"0000006100000047000000370000002b000000230000001e0000001e0000001e",
            INIT_5F => X"000000b300000098000000860000006f0000006900000078000000830000007c",
            INIT_60 => X"000000210000002b000000340000002c0000000c0000000a0000000a0000000f",
            INIT_61 => X"000000800000009e000000750000000800000001000000020000000400000012",
            INIT_62 => X"0000007e0000007e000000730000006b00000069000000670000006900000070",
            INIT_63 => X"000000c2000000ac0000009300000082000000740000005e000000560000006a",
            INIT_64 => X"0000000a0000000c0000000c0000000600000004000000030000000a00000028",
            INIT_65 => X"00000082000000800000003a0000000000000002000000010000000100000006",
            INIT_66 => X"000000420000004b000000600000006e00000071000000770000007b0000007f",
            INIT_67 => X"000000c5000000b6000000a20000008d00000084000000760000005d00000047",
            INIT_68 => X"0000000200000003000000020000000100000001000000010000001d0000004d",
            INIT_69 => X"0000002f0000002d0000000c0000000100000000000000000000000000000001",
            INIT_6A => X"0000004d00000030000000260000002a0000003100000032000000300000002e",
            INIT_6B => X"000000c6000000bb000000b00000009900000087000000800000007e0000006e",
            INIT_6C => X"000000000000000100000001000000000000000100000001000000340000005e",
            INIT_6D => X"0000002000000019000000030000000200000000000000000000000000000000",
            INIT_6E => X"000000710000005c00000042000000290000001d000000190000001900000019",
            INIT_6F => X"000000c9000000bf000000b30000009d0000008b0000007f0000007e0000007c",
            INIT_70 => X"0000000200000003000000030000000200000002000000070000003c00000066",
            INIT_71 => X"0000001f00000013000000010000000300000001000000000000000000000001",
            INIT_72 => X"0000007c0000007e000000730000005a0000003a0000001b0000000d00000011",
            INIT_73 => X"000000ca000000c0000000b00000009f0000009100000087000000820000007b",
            INIT_74 => X"000000070000000a0000000b0000000a0000000c000000170000003300000063",
            INIT_75 => X"000000150000000d000000050000000600000003000000040000000400000004",
            INIT_76 => X"0000007d0000007e0000007e00000071000000620000004d000000320000001b",
            INIT_77 => X"000000ca000000c5000000b8000000a80000009a000000940000008a00000080",
            INIT_78 => X"000000170000001a0000001c0000001e000000230000002c0000003900000060",
            INIT_79 => X"00000037000000280000001f0000001b00000017000000160000001500000015",
            INIT_7A => X"0000007f0000007a0000007a0000007900000070000000660000005800000046",
            INIT_7B => X"000000ca000000c8000000bd000000ac000000a0000000950000008b00000085",
            INIT_7C => X"000000370000003500000035000000380000003d000000430000004b00000065",
            INIT_7D => X"000000600000005400000047000000430000003e0000003a0000003800000037",
            INIT_7E => X"000000830000007d0000007c0000007f00000079000000740000006d00000067",
            INIT_7F => X"000000c8000000c3000000b7000000ab000000a2000000980000009100000088",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY4;


    MEM_IFMAP_LAYER0_ENTITY5 : if BRAM_NAME = "ifmap_layer0_entity5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e8000000e8000000e8000000e8000000e8000000e8000000e7000000eb",
            INIT_01 => X"000000e9000000e9000000e9000000e9000000e9000000e9000000e8000000e8",
            INIT_02 => X"000000e6000000e8000000ea000000ea000000e8000000e9000000e9000000e9",
            INIT_03 => X"000000e8000000e9000000e9000000e8000000e8000000e8000000e9000000e7",
            INIT_04 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_05 => X"000000ec000000ec000000ec000000ec000000ec000000ec000000eb000000eb",
            INIT_06 => X"000000eb000000ed000000ee000000ed000000ea000000ea000000e9000000e9",
            INIT_07 => X"000000eb000000ec000000ec000000eb000000eb000000eb000000ec000000ea",
            INIT_08 => X"000000ea000000ea000000ea000000ea000000ea000000ea000000ea000000ed",
            INIT_09 => X"000000ea000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0A => X"000000ea000000eb000000ee000000e9000000ec000000ea000000e7000000e7",
            INIT_0B => X"000000ea000000eb000000eb000000ea000000ea000000ea000000ea000000ea",
            INIT_0C => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_0D => X"000000ea000000eb000000ea000000ea000000ea000000ea000000ea000000ea",
            INIT_0E => X"000000e6000000d5000000db000000c5000000e7000000e8000000e7000000e6",
            INIT_0F => X"000000eb000000eb000000eb000000ea000000ea000000ea000000ea000000eb",
            INIT_10 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000ea000000ed",
            INIT_11 => X"000000eb000000eb000000ea000000ea000000eb000000eb000000ea000000ea",
            INIT_12 => X"000000e8000000dd000000d0000000b3000000db000000e6000000ed000000ec",
            INIT_13 => X"000000ec000000ec000000ec000000ec000000eb000000eb000000eb000000ed",
            INIT_14 => X"000000eb000000eb000000eb000000eb000000eb000000eb000000eb000000ee",
            INIT_15 => X"000000e8000000ed000000ea000000ec000000ec000000ec000000eb000000ea",
            INIT_16 => X"000000e8000000dc000000ca000000bd000000c8000000cf000000d2000000da",
            INIT_17 => X"000000ed000000ed000000ed000000ec000000eb000000eb000000eb000000ed",
            INIT_18 => X"000000eb000000eb000000ec000000e9000000e6000000e7000000e4000000e5",
            INIT_19 => X"000000e4000000ee000000e5000000e6000000ee000000ed000000ec000000ec",
            INIT_1A => X"000000d3000000b1000000ab000000b1000000be000000bf000000be000000cc",
            INIT_1B => X"000000ee000000ed000000ed000000ec000000eb000000e9000000ea000000ef",
            INIT_1C => X"000000ec000000eb000000ec000000ea000000ea000000ee000000e9000000de",
            INIT_1D => X"000000da000000eb000000dd000000cb000000ef000000ed000000ee000000ee",
            INIT_1E => X"000000cc000000b9000000bb000000c4000000cb000000d3000000d2000000d2",
            INIT_1F => X"000000ee000000ee000000ee000000ee000000ee000000ed000000ee000000f0",
            INIT_20 => X"000000eb000000eb000000ed000000f0000000f3000000f6000000f3000000f1",
            INIT_21 => X"000000e5000000e7000000da000000c4000000ef000000ed000000ed000000ed",
            INIT_22 => X"000000f1000000f0000000eb000000ea000000e3000000eb000000de000000d9",
            INIT_23 => X"000000ee000000ef000000ef000000ef000000f0000000f0000000f0000000f3",
            INIT_24 => X"000000e8000000e9000000e9000000bf000000a1000000990000009400000095",
            INIT_25 => X"000000ec000000e8000000e2000000d6000000eb000000ec000000eb000000ea",
            INIT_26 => X"000000d3000000e2000000f3000000f7000000ef000000f1000000eb000000e8",
            INIT_27 => X"000000ef000000ef000000ef000000eb000000c9000000b9000000ba000000c3",
            INIT_28 => X"000000e0000000e1000000e7000000a50000008900000089000000850000008d",
            INIT_29 => X"000000ec000000ee000000ec000000eb000000eb000000ea000000ea000000e9",
            INIT_2A => X"000000a3000000ac000000bf000000d5000000ee000000f1000000f0000000ee",
            INIT_2B => X"000000ef000000ee000000ef000000e5000000a60000008f000000990000009f",
            INIT_2C => X"000000ce000000d3000000e7000000e3000000df000000e0000000d7000000e0",
            INIT_2D => X"000000e9000000e6000000e1000000df000000db000000e1000000de000000d6",
            INIT_2E => X"000000ca000000cf000000cb000000d0000000ed000000f1000000ef000000ed",
            INIT_2F => X"000000ef000000ef000000ee000000e9000000ca000000a4000000c4000000d3",
            INIT_30 => X"000000ae000000d0000000e3000000f1000000ea000000e0000000d9000000de",
            INIT_31 => X"000000930000008b000000840000007e00000079000000bc000000d6000000b7",
            INIT_32 => X"000000e9000000f0000000ee000000eb000000ed000000dc000000ae000000a1",
            INIT_33 => X"000000f2000000f2000000e9000000ea000000ed000000d4000000e5000000ed",
            INIT_34 => X"000000cc000000cd000000c1000000a5000000970000008d0000009300000098",
            INIT_35 => X"000000620000005a0000005b0000005b0000005c000000b7000000ea000000e2",
            INIT_36 => X"000000d9000000e9000000ed000000f1000000f1000000e9000000b300000081",
            INIT_37 => X"000000ea000000e3000000cd000000c4000000d6000000df000000dc000000d4",
            INIT_38 => X"000000cf000000a4000000a40000009b0000006600000064000000720000006c",
            INIT_39 => X"000000cf000000a800000087000000830000008a000000be000000e4000000ea",
            INIT_3A => X"00000093000000a3000000ae000000c3000000d4000000e3000000e8000000df",
            INIT_3B => X"000000d8000000cb000000a0000000930000009700000098000000900000008c",
            INIT_3C => X"000000a1000000760000006e0000009c00000099000000740000005e0000004d",
            INIT_3D => X"000000d9000000ec000000d9000000ca000000c8000000c6000000c5000000b6",
            INIT_3E => X"0000007b000000760000007b0000008a000000950000009f000000ac000000ba",
            INIT_3F => X"000000d0000000d5000000b8000000ae000000a1000000910000008200000080",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a2000000860000007b00000096000000dc000000970000002f00000023",
            INIT_41 => X"000000be000000ee000000f0000000e8000000e9000000e1000000d3000000b4",
            INIT_42 => X"000000bb000000b6000000b6000000bb000000b1000000aa000000a2000000a3",
            INIT_43 => X"000000b7000000c1000000d0000000da000000d9000000cc000000bf000000bd",
            INIT_44 => X"000000e5000000da000000d3000000d4000000ef000000d90000004f00000018",
            INIT_45 => X"000000ea000000f1000000ef000000dc000000ef000000f5000000f6000000ed",
            INIT_46 => X"000000e0000000e8000000ea000000e7000000e5000000e6000000d6000000e4",
            INIT_47 => X"000000a50000009e000000a1000000a9000000b3000000c5000000d1000000d4",
            INIT_48 => X"000000e3000000e6000000e5000000d9000000d8000000de000000b300000047",
            INIT_49 => X"000000bc000000c1000000d7000000cf000000dd000000e4000000e4000000e3",
            INIT_4A => X"0000009e000000ad000000b4000000a10000009c000000ba000000c3000000b8",
            INIT_4B => X"0000009c0000009e000000970000008c0000008300000085000000870000008a",
            INIT_4C => X"000000c1000000c0000000be000000bb000000bd000000c2000000cf000000a1",
            INIT_4D => X"0000009a000000a3000000ba000000bc000000bd000000bd000000be000000c0",
            INIT_4E => X"0000008800000090000000990000009400000091000000a3000000aa0000009a",
            INIT_4F => X"0000009c0000009400000092000000900000008d0000008b0000008600000082",
            INIT_50 => X"00000096000000930000008e000000860000007f0000007a000000710000006d",
            INIT_51 => X"000000af000000b4000000ba000000b5000000ac000000a5000000a000000098",
            INIT_52 => X"0000007f000000840000008b000000940000009b000000a3000000a8000000ac",
            INIT_53 => X"0000009c000000920000008a0000007e0000007a000000810000008500000081",
            INIT_54 => X"0000003d0000003a000000380000003400000030000000230000001900000029",
            INIT_55 => X"0000007e0000007e000000790000006a000000570000004d000000460000003e",
            INIT_56 => X"0000006600000067000000680000006a00000070000000780000007e0000007f",
            INIT_57 => X"000000950000008d000000880000008000000077000000730000006e00000069",
            INIT_58 => X"000000180000001e000000290000003a00000035000000130000001400000037",
            INIT_59 => X"0000003e0000003c000000380000002a000000140000000f0000000f00000011",
            INIT_5A => X"0000005a000000530000004f0000004e0000004c0000004d0000005100000047",
            INIT_5B => X"0000009e00000089000000800000007d0000008a0000008a0000007600000065",
            INIT_5C => X"00000025000000390000004c0000005400000029000000120000001a0000002d",
            INIT_5D => X"0000003e0000004e0000005b0000002300000007000000070000000b00000015",
            INIT_5E => X"0000007b00000063000000530000004a000000450000003f0000003e0000003c",
            INIT_5F => X"000000af00000092000000850000007400000072000000870000009500000092",
            INIT_60 => X"000000230000002f000000390000002e0000000b000000080000000900000011",
            INIT_61 => X"00000094000000b3000000860000000f00000003000000040000000700000014",
            INIT_62 => X"0000008d00000090000000850000007e0000007f0000007c0000007d00000083",
            INIT_63 => X"000000be000000a5000000900000008100000074000000610000005b00000074",
            INIT_64 => X"0000000c00000011000000110000000700000004000000030000000700000023",
            INIT_65 => X"0000009400000092000000400000000200000003000000020000000300000007",
            INIT_66 => X"00000045000000530000006a0000007a00000081000000890000008d00000090",
            INIT_67 => X"000000c2000000b00000009e000000870000007e000000710000005800000046",
            INIT_68 => X"0000000500000009000000050000000000000002000000010000001500000040",
            INIT_69 => X"000000440000003b0000000b0000000100000001000000000000000000000002",
            INIT_6A => X"000000470000002e0000002a000000310000003b000000430000004500000043",
            INIT_6B => X"000000c4000000b7000000ab0000009300000080000000780000007400000066",
            INIT_6C => X"0000000200000005000000020000000000000002000000010000002b00000052",
            INIT_6D => X"0000003600000026000000020000000000000000000000000000000000000000",
            INIT_6E => X"0000006900000052000000380000002700000022000000240000002b0000002e",
            INIT_6F => X"000000c7000000bb000000ae0000009600000083000000760000007300000073",
            INIT_70 => X"000000020000000300000001000000000000000100000003000000320000005d",
            INIT_71 => X"0000002f0000001c000000000000000200000001000000000000000000000001",
            INIT_72 => X"000000700000006f000000630000005100000037000000160000000c00000017",
            INIT_73 => X"000000c9000000bc000000ab00000097000000890000007e0000007700000071",
            INIT_74 => X"00000002000000040000000400000002000000040000000b0000002500000059",
            INIT_75 => X"000000180000000d000000020000000600000002000000010000000100000001",
            INIT_76 => X"0000006f000000700000007100000065000000520000003e0000002900000019",
            INIT_77 => X"000000c9000000c1000000b3000000a100000091000000890000007e00000073",
            INIT_78 => X"0000000c0000000d0000000f0000000f00000011000000160000002400000052",
            INIT_79 => X"0000002d0000001b00000015000000140000000f0000000e0000000d0000000c",
            INIT_7A => X"000000700000006b0000006e0000006900000058000000550000005100000043",
            INIT_7B => X"000000c8000000c4000000b7000000a4000000970000008a0000007f00000077",
            INIT_7C => X"0000002600000022000000210000002300000025000000260000003000000053",
            INIT_7D => X"0000004a0000003b000000300000002d0000002e0000002c0000002900000028",
            INIT_7E => X"000000750000006c0000006a0000006b00000061000000610000005c00000053",
            INIT_7F => X"000000c7000000bf000000b2000000a3000000990000008d000000850000007b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY5;


    MEM_IFMAP_LAYER0_ENTITY6 : if BRAM_NAME = "ifmap_layer0_entity6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c1000000bb000000b6000000a6000000840000008b0000009e0000009e",
            INIT_01 => X"000000e6000000e3000000df000000da000000ce000000d1000000cd000000c7",
            INIT_02 => X"000000ea000000ea000000e8000000ec000000eb000000e7000000e2000000d5",
            INIT_03 => X"000000ee000000ed000000e4000000e8000000ee000000e6000000e2000000ec",
            INIT_04 => X"000000c7000000c5000000c1000000ae0000008900000097000000ac000000aa",
            INIT_05 => X"000000ed000000e9000000e7000000e1000000d2000000d9000000d7000000ce",
            INIT_06 => X"000000f2000000ec000000ea000000f5000000f2000000e8000000e4000000db",
            INIT_07 => X"000000f6000000f6000000e8000000e9000000f3000000eb000000e4000000f1",
            INIT_08 => X"000000c7000000ce000000c9000000b50000008e0000009d000000b0000000ae",
            INIT_09 => X"000000ef000000e6000000e6000000e0000000d4000000da000000df000000d1",
            INIT_0A => X"000000f3000000ec000000d5000000e8000000ef000000e9000000e4000000dd",
            INIT_0B => X"000000f5000000fa000000e6000000ed000000f8000000ee000000e7000000f5",
            INIT_0C => X"000000cf000000d4000000cb000000ba00000093000000a0000000b2000000b4",
            INIT_0D => X"000000f0000000df000000e7000000dc000000d6000000dd000000e4000000d6",
            INIT_0E => X"000000f3000000e6000000ac000000b1000000e4000000e9000000e4000000e0",
            INIT_0F => X"000000f4000000f9000000e4000000ee000000fa000000ee000000e8000000f8",
            INIT_10 => X"000000cf000000d9000000cc000000bd00000093000000a5000000b9000000ba",
            INIT_11 => X"000000eb000000d3000000e7000000da000000d6000000de000000e7000000d3",
            INIT_12 => X"000000ed000000e0000000a80000009f000000d4000000e8000000e0000000e2",
            INIT_13 => X"000000f2000000f8000000ea000000e8000000f6000000eb000000e7000000f7",
            INIT_14 => X"000000d3000000db000000cb000000bf0000008e000000aa000000be000000c1",
            INIT_15 => X"000000cd000000c7000000e4000000d6000000d6000000dd000000ea000000d7",
            INIT_16 => X"000000e6000000de0000009e00000070000000c1000000eb000000ce000000cf",
            INIT_17 => X"000000eb000000f3000000e7000000e4000000f1000000e2000000e5000000f5",
            INIT_18 => X"000000d9000000de000000ca000000bf00000085000000ac000000bf000000c4",
            INIT_19 => X"000000b0000000bc000000e3000000d7000000d6000000da000000eb000000df",
            INIT_1A => X"000000b7000000ac0000008900000078000000bb000000cd000000ba000000bb",
            INIT_1B => X"000000eb000000f0000000e1000000e2000000eb000000d8000000df000000db",
            INIT_1C => X"000000e0000000e0000000da000000cb0000008c000000ae000000c5000000cc",
            INIT_1D => X"000000cd000000c9000000dd000000dc000000dc000000dc000000ed000000e8",
            INIT_1E => X"0000003c000000410000003e0000004700000053000000640000008a000000ac",
            INIT_1F => X"000000ec000000ef000000d4000000da000000e4000000d1000000b600000068",
            INIT_20 => X"000000c5000000af000000ba000000b0000000890000009d000000aa000000af",
            INIT_21 => X"000000c1000000c1000000c9000000d4000000d2000000ce000000d4000000d1",
            INIT_22 => X"000000450000005e00000053000000540000005b00000059000000690000008e",
            INIT_23 => X"000000c3000000cf000000a3000000ae000000b7000000a2000000790000004e",
            INIT_24 => X"000000800000006f0000006b0000006900000068000000710000007300000072",
            INIT_25 => X"0000009600000097000000930000009d0000009b00000097000000920000008b",
            INIT_26 => X"0000005300000056000000560000005500000063000000630000006400000076",
            INIT_27 => X"0000007b000000840000006d00000076000000990000009a000000800000008b",
            INIT_28 => X"0000005a000000540000005a00000053000000440000004b0000004c00000042",
            INIT_29 => X"0000006c000000720000006b0000006a00000067000000660000006a0000005d",
            INIT_2A => X"000000720000005f0000004200000048000000550000005b0000005a0000005a",
            INIT_2B => X"0000005e0000005c000000670000007d000000c7000000930000006e00000080",
            INIT_2C => X"00000046000000550000006a0000006f0000004d0000004b0000004100000035",
            INIT_2D => X"000000610000006b000000730000006c0000005d0000005f000000710000005d",
            INIT_2E => X"000000bb00000095000000550000005a00000061000000620000005f00000062",
            INIT_2F => X"00000055000000570000005f0000009a000000cc0000007000000092000000b3",
            INIT_30 => X"000000550000004d00000064000000640000004a0000005e000000560000003a",
            INIT_31 => X"00000057000000620000006e000000690000006c0000007f0000008500000078",
            INIT_32 => X"000000c3000000aa000000700000005f0000005f000000570000005100000051",
            INIT_33 => X"0000004f0000005500000050000000b2000000ad0000007f000000c1000000d0",
            INIT_34 => X"000000500000004700000044000000520000004b00000057000000590000004a",
            INIT_35 => X"00000062000000690000006a000000650000006f000000760000006700000059",
            INIT_36 => X"000000b8000000b40000008e000000720000006d000000620000006200000060",
            INIT_37 => X"000000430000003c00000050000000aa00000084000000a0000000c0000000bf",
            INIT_38 => X"0000005600000046000000480000004f0000004e000000520000004f0000004d",
            INIT_39 => X"000000830000008700000088000000890000008500000081000000790000006d",
            INIT_3A => X"000000b5000000b3000000a30000009400000096000000920000009400000092",
            INIT_3B => X"0000003b00000037000000490000005a00000065000000aa000000b0000000b9",
            INIT_3C => X"0000008a00000084000000830000006d000000680000006a0000005e00000060",
            INIT_3D => X"000000940000009e0000009b0000009b0000009a0000009b0000009800000090",
            INIT_3E => X"000000a9000000920000008200000077000000920000009c0000009d00000096",
            INIT_3F => X"0000004800000056000000620000004500000069000000a7000000a8000000b1",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008f0000009000000087000000810000008300000073000000650000006a",
            INIT_41 => X"0000009000000097000000990000009a0000009a0000009a0000009600000092",
            INIT_42 => X"0000009f00000092000000750000005e0000007f0000008b0000008600000082",
            INIT_43 => X"000000690000009a000000c00000009000000084000000a2000000a3000000a7",
            INIT_44 => X"00000091000000810000005d0000005f0000006d000000760000006c0000005f",
            INIT_45 => X"0000007b0000007a0000007e0000008600000090000000960000009700000095",
            INIT_46 => X"0000009c000000a20000009300000083000000940000009b000000850000007a",
            INIT_47 => X"000000940000009d000000a40000009f0000009500000099000000970000009d",
            INIT_48 => X"0000008c0000007b0000006f0000005600000046000000490000005900000066",
            INIT_49 => X"0000008d000000850000007e000000780000007500000078000000810000008f",
            INIT_4A => X"000000a1000000a50000009d000000970000009f000000990000008e00000096",
            INIT_4B => X"000000950000007d0000007900000083000000900000009a0000009800000099",
            INIT_4C => X"0000007b000000820000008a000000800000006e000000470000003d00000056",
            INIT_4D => X"000000990000009c000000980000008f00000084000000760000006c00000076",
            INIT_4E => X"000000a4000000a00000009a000000990000009a000000910000008900000095",
            INIT_4F => X"00000084000000560000004b0000005c000000690000007d0000009000000098",
            INIT_50 => X"000000760000007b0000007400000073000000720000006b0000006700000068",
            INIT_51 => X"00000075000000850000008d0000008f000000900000008d0000008600000074",
            INIT_52 => X"00000091000000980000009a0000009700000096000000820000005900000062",
            INIT_53 => X"00000041000000490000004700000041000000500000005a0000006000000075",
            INIT_54 => X"0000007e0000007d00000077000000720000006f0000006f0000006b00000063",
            INIT_55 => X"0000003d0000005b0000008200000083000000810000007d0000007d00000075",
            INIT_56 => X"0000005f00000072000000820000008b00000094000000730000003800000039",
            INIT_57 => X"0000001b000000330000004b0000003c0000003a000000490000005300000056",
            INIT_58 => X"0000005b0000006600000075000000740000007200000074000000680000003e",
            INIT_59 => X"0000004c000000600000008200000085000000700000004e0000005100000054",
            INIT_5A => X"000000510000005300000058000000600000006c0000006b0000005600000053",
            INIT_5B => X"000000180000001e0000002e000000340000002d000000330000003d00000046",
            INIT_5C => X"0000003500000041000000680000006b000000690000006a0000006000000039",
            INIT_5D => X"000000620000007300000085000000870000006e00000044000000400000003b",
            INIT_5E => X"00000037000000460000005000000051000000500000004e0000004f00000058",
            INIT_5F => X"000000180000001b0000001e00000022000000290000002d000000310000002c",
            INIT_60 => X"000000490000004f0000006d0000006d00000069000000680000005a00000041",
            INIT_61 => X"000000410000004400000053000000620000006a000000620000005800000055",
            INIT_62 => X"0000002c00000029000000330000004800000052000000510000004a00000046",
            INIT_63 => X"000000190000001b0000001e000000200000002300000027000000370000003d",
            INIT_64 => X"0000005100000058000000630000006600000067000000690000005700000043",
            INIT_65 => X"00000046000000420000003f0000003a000000390000003b000000450000004c",
            INIT_66 => X"0000002c000000310000002f0000002e000000360000003e0000004400000048",
            INIT_67 => X"0000001e00000018000000190000001d0000001c0000001e0000002e00000038",
            INIT_68 => X"0000002c0000002d00000032000000370000003a000000410000003a00000036",
            INIT_69 => X"0000003a0000003e000000400000003e0000003a00000037000000330000002e",
            INIT_6A => X"000000260000002a000000300000003100000030000000250000002600000033",
            INIT_6B => X"0000001f0000001c000000190000001b0000001c0000001b0000002000000029",
            INIT_6C => X"0000002700000021000000200000001f0000001b0000001a0000001d0000001e",
            INIT_6D => X"0000002800000026000000280000002e00000033000000350000003400000031",
            INIT_6E => X"0000002500000024000000250000002900000037000000420000002c00000026",
            INIT_6F => X"00000017000000210000001e0000001c0000001b0000001a0000001b0000001f",
            INIT_70 => X"000000200000001f0000001e0000001c0000001c0000001b0000001f00000021",
            INIT_71 => X"0000002d0000002900000027000000220000001e0000001e0000002100000023",
            INIT_72 => X"0000002000000026000000230000001e0000003100000049000000340000002a",
            INIT_73 => X"0000000d0000001a000000260000001e0000001d0000001b0000001a0000001b",
            INIT_74 => X"0000001b0000001a00000019000000190000001a0000001a0000001e0000001f",
            INIT_75 => X"0000002a00000028000000290000002a0000002800000025000000200000001d",
            INIT_76 => X"0000001d0000001e000000240000001c00000026000000400000002e00000027",
            INIT_77 => X"000000040000000900000025000000210000001c0000001b000000190000001a",
            INIT_78 => X"0000002500000022000000200000001e0000001c000000190000001b00000017",
            INIT_79 => X"000000210000001e000000230000002600000027000000280000002700000027",
            INIT_7A => X"0000001d0000001d0000001d0000001e0000002400000039000000240000001c",
            INIT_7B => X"000000050000000400000013000000240000001b000000170000001800000018",
            INIT_7C => X"0000002500000023000000220000002100000022000000200000001e0000001c",
            INIT_7D => X"0000000c0000000f000000180000001e00000022000000240000002600000026",
            INIT_7E => X"0000001c0000001b0000001b00000019000000200000002d0000001300000008",
            INIT_7F => X"0000000700000004000000050000001900000022000000140000001500000018",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY6;


    MEM_IFMAP_LAYER0_ENTITY7 : if BRAM_NAME = "ifmap_layer0_entity7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d8000000d3000000d0000000c10000009e000000a6000000bb000000be",
            INIT_01 => X"000000ed000000eb000000e8000000e5000000da000000de000000dd000000db",
            INIT_02 => X"000000f1000000f1000000ef000000f1000000ef000000ee000000e9000000dc",
            INIT_03 => X"000000f1000000ef000000e7000000ed000000f3000000eb000000e7000000f2",
            INIT_04 => X"000000da000000da000000d9000000c7000000a0000000b0000000c7000000c8",
            INIT_05 => X"000000f3000000ef000000ee000000e9000000db000000e5000000e5000000df",
            INIT_06 => X"000000f5000000ef000000ed000000f7000000f5000000ee000000ea000000e1",
            INIT_07 => X"000000f7000000f6000000e8000000ec000000f8000000ef000000e9000000f5",
            INIT_08 => X"000000d6000000df000000dc000000c9000000a2000000b3000000c8000000c9",
            INIT_09 => X"000000f4000000ea000000ea000000e5000000db000000e2000000e9000000dd",
            INIT_0A => X"000000f1000000ea000000d6000000eb000000f3000000ee000000e9000000e2",
            INIT_0B => X"000000f4000000f9000000e5000000ee000000fa000000f0000000e9000000f7",
            INIT_0C => X"000000d9000000e1000000d9000000c9000000a4000000b3000000c7000000cb",
            INIT_0D => X"000000f4000000e2000000e8000000dd000000d9000000e3000000eb000000df",
            INIT_0E => X"000000f1000000e4000000af000000b8000000eb000000ed000000e7000000e4",
            INIT_0F => X"000000f2000000f7000000e3000000ed000000fa000000ee000000e8000000f8",
            INIT_10 => X"000000d5000000e1000000d6000000c9000000a1000000b5000000cc000000cf",
            INIT_11 => X"000000ec000000d4000000e5000000d9000000d7000000e2000000ed000000d7",
            INIT_12 => X"000000ec000000e0000000ae000000aa000000e1000000ec000000e1000000e3",
            INIT_13 => X"000000ef000000f5000000e7000000e7000000f6000000eb000000e7000000f7",
            INIT_14 => X"000000d7000000e2000000d4000000c90000009a000000b7000000cd000000d0",
            INIT_15 => X"000000cd000000c7000000e5000000d7000000d7000000df000000ee000000da",
            INIT_16 => X"000000e9000000e3000000a70000007c000000cc000000ef000000d0000000d1",
            INIT_17 => X"000000e8000000f1000000e6000000e2000000ef000000e1000000e5000000f6",
            INIT_18 => X"000000d5000000dd000000cb000000c20000008b000000b3000000c7000000cc",
            INIT_19 => X"000000b0000000bc000000e6000000d8000000d4000000d8000000e9000000db",
            INIT_1A => X"000000be000000b70000009700000081000000c0000000d4000000c0000000be",
            INIT_1B => X"000000e0000000eb000000de000000db000000e5000000d6000000e0000000e0",
            INIT_1C => X"000000cc000000ce000000cb000000c00000008a000000af000000c6000000cd",
            INIT_1D => X"000000ce000000c7000000d8000000d5000000d2000000d0000000df000000d4",
            INIT_1E => X"000000450000005000000050000000550000005d0000007100000095000000b2",
            INIT_1F => X"000000d4000000dd000000c5000000d0000000de000000ce000000b70000006c",
            INIT_20 => X"000000b3000000a0000000ac000000a5000000850000009a000000a8000000ad",
            INIT_21 => X"000000c6000000c1000000bf000000c7000000c3000000bd000000c2000000be",
            INIT_22 => X"0000004f0000006e00000068000000680000006c0000006b0000007900000098",
            INIT_23 => X"000000af000000be00000095000000a3000000af0000009f0000007a00000052",
            INIT_24 => X"0000007f000000700000006e0000006d00000069000000720000007400000073",
            INIT_25 => X"000000a10000009e0000008f00000097000000930000008c0000008800000087",
            INIT_26 => X"0000005c000000660000006c0000006c00000078000000780000007700000086",
            INIT_27 => X"00000078000000820000006a0000006e0000009100000097000000800000008f",
            INIT_28 => X"000000640000006100000069000000630000005200000056000000570000004e",
            INIT_29 => X"0000007f0000008400000076000000720000006f0000006a0000006d00000065",
            INIT_2A => X"000000770000006c00000057000000600000006b0000006e0000006d0000006d",
            INIT_2B => X"00000068000000660000006f00000078000000bf000000900000006f00000084",
            INIT_2C => X"00000051000000620000007a00000080000000620000005f000000550000004a",
            INIT_2D => X"0000007b000000860000008b0000008400000073000000710000008100000068",
            INIT_2E => X"000000bd0000009e000000680000007100000077000000740000007300000078",
            INIT_2F => X"00000063000000630000006700000095000000c50000006d00000094000000b7",
            INIT_30 => X"000000660000005d00000073000000750000005d000000710000006b00000051",
            INIT_31 => X"000000710000007d000000880000008200000083000000950000009800000089",
            INIT_32 => X"000000c2000000af0000007f000000760000007b000000720000006c0000006c",
            INIT_33 => X"000000650000006200000050000000a7000000a200000076000000bd000000ce",
            INIT_34 => X"000000640000005900000054000000620000005d0000006a0000006e00000061",
            INIT_35 => X"0000007c00000082000000830000007e000000860000008a0000007b0000006e",
            INIT_36 => X"000000b4000000b50000009900000086000000870000007e0000007f0000007b",
            INIT_37 => X"00000059000000480000004d000000a00000007a00000097000000b7000000b8",
            INIT_38 => X"0000006b00000058000000580000005f00000061000000660000006500000066",
            INIT_39 => X"0000009d000000a1000000a4000000a30000009e000000970000008e00000082",
            INIT_3A => X"000000ae000000b1000000a9000000a2000000a9000000aa000000ad000000ab",
            INIT_3B => X"0000004b0000003f000000460000005700000062000000a4000000a8000000b0",
            INIT_3C => X"000000a000000098000000940000007e0000007c0000007f000000760000007b",
            INIT_3D => X"000000ae000000b9000000b8000000b7000000b4000000b3000000af000000a7",
            INIT_3E => X"000000a10000008e0000008500000080000000a0000000af000000b2000000ad",
            INIT_3F => X"00000052000000590000005f000000460000006c000000a6000000a2000000a9",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a7000000a60000009a00000094000000980000008a0000007d00000085",
            INIT_41 => X"000000ab000000b5000000b9000000b9000000b6000000b3000000ae000000aa",
            INIT_42 => X"0000009b0000009000000078000000660000008b0000009a0000009800000098",
            INIT_43 => X"0000006c00000099000000bb0000009100000088000000a3000000a2000000a5",
            INIT_44 => X"000000aa000000980000007200000074000000830000008d000000850000007c",
            INIT_45 => X"000000970000009a000000a0000000a7000000ad000000b0000000af000000af",
            INIT_46 => X"0000009e000000a5000000980000008c000000a0000000a80000009600000090",
            INIT_47 => X"00000093000000980000009e0000009e000000970000009c0000009b000000a3",
            INIT_48 => X"000000a400000094000000870000006e0000005d000000600000007100000081",
            INIT_49 => X"000000a50000009f000000990000009400000092000000960000009f000000a9",
            INIT_4A => X"000000a4000000a8000000a4000000a1000000ac000000a8000000a0000000aa",
            INIT_4B => X"000000960000007d0000007900000084000000920000009e0000009e000000a0",
            INIT_4C => X"000000930000009c000000a50000009b00000087000000600000005500000070",
            INIT_4D => X"000000ab000000ae000000ad000000a7000000a0000000970000008d0000008e",
            INIT_4E => X"000000a6000000a3000000a1000000a3000000a8000000a20000009b000000a7",
            INIT_4F => X"0000008a0000005c00000052000000620000006f00000082000000970000009e",
            INIT_50 => X"0000008e000000960000008f0000008f0000008f000000870000008400000085",
            INIT_51 => X"0000008600000097000000a5000000a9000000ab000000a9000000a10000008a",
            INIT_52 => X"000000980000009f000000a3000000a3000000a4000000940000006b00000074",
            INIT_53 => X"00000048000000500000004e0000004b0000005b000000660000006c00000080",
            INIT_54 => X"000000960000009700000093000000900000008f000000900000008c00000084",
            INIT_55 => X"0000004e0000006e0000009c0000009f0000009a00000094000000920000008b",
            INIT_56 => X"0000006d0000007e0000008f00000099000000a3000000840000004a0000004b",
            INIT_57 => X"0000002100000039000000520000004b0000004c0000005a0000006400000067",
            INIT_58 => X"000000730000008100000091000000920000009200000094000000890000005e",
            INIT_59 => X"0000005d000000720000009a0000009d0000008700000063000000660000006a",
            INIT_5A => X"00000065000000660000006a000000710000007c0000007d0000006800000065",
            INIT_5B => X"0000001f0000002500000035000000430000003f000000450000004f00000058",
            INIT_5C => X"0000004d0000005c000000850000008900000086000000860000007d00000056",
            INIT_5D => X"00000073000000840000009600000099000000830000005c0000005900000052",
            INIT_5E => X"0000004f0000005f00000065000000630000006100000060000000610000006a",
            INIT_5F => X"0000001f00000022000000260000002f000000390000003c000000400000003c",
            INIT_60 => X"000000610000006a0000008a000000890000008300000081000000740000005a",
            INIT_61 => X"00000053000000540000005f000000710000007e0000007c000000740000006c",
            INIT_62 => X"00000045000000430000004a0000005c00000064000000620000005c00000059",
            INIT_63 => X"0000002000000023000000260000002b0000002e00000033000000420000004a",
            INIT_64 => X"000000660000006e000000780000007c0000007f00000082000000700000005c",
            INIT_65 => X"0000005b00000054000000500000004b0000004c000000500000005a00000061",
            INIT_66 => X"0000003d0000004300000041000000410000004900000051000000590000005f",
            INIT_67 => X"0000002500000023000000280000002a000000280000002a0000003a00000045",
            INIT_68 => X"0000003f00000040000000450000004a0000004e000000560000004f0000004c",
            INIT_69 => X"000000500000005100000052000000510000004d0000004a0000004600000041",
            INIT_6A => X"00000032000000360000003f0000004300000044000000370000003b00000049",
            INIT_6B => X"0000002500000027000000280000002900000028000000280000002d00000036",
            INIT_6C => X"0000003a0000003500000034000000310000002a000000280000002b0000002d",
            INIT_6D => X"0000003b0000003a0000003b0000004100000046000000480000004700000044",
            INIT_6E => X"0000002f0000002f000000330000003900000049000000550000003f00000038",
            INIT_6F => X"0000001d0000002a0000002a000000290000002800000027000000280000002c",
            INIT_70 => X"0000003200000031000000300000002c0000002600000024000000280000002b",
            INIT_71 => X"0000003d0000003e0000003b0000003500000031000000310000003400000035",
            INIT_72 => X"000000280000002f0000002e0000002c000000420000005e0000004500000037",
            INIT_73 => X"00000012000000200000002e000000290000002a000000280000002700000027",
            INIT_74 => X"0000002b00000029000000290000002700000024000000230000002700000028",
            INIT_75 => X"000000370000003c0000003d0000003d0000003a00000038000000330000002e",
            INIT_76 => X"00000024000000250000002e0000002800000036000000550000003c0000002e",
            INIT_77 => X"000000070000000d000000280000002b0000002a000000280000002600000026",
            INIT_78 => X"00000033000000310000002f0000002c00000028000000240000002600000022",
            INIT_79 => X"0000002b000000330000003700000039000000390000003b0000003900000036",
            INIT_7A => X"00000023000000230000002500000029000000320000004e000000300000001f",
            INIT_7B => X"0000000700000006000000140000002d00000029000000240000002500000025",
            INIT_7C => X"000000310000003000000030000000300000002f0000002d0000002b00000029",
            INIT_7D => X"000000110000001a00000022000000280000002d000000310000003300000032",
            INIT_7E => X"000000230000002200000022000000210000002c0000003f0000001b00000008",
            INIT_7F => X"0000000800000005000000060000001f0000002c000000220000002200000023",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY7;


    MEM_IFMAP_LAYER0_ENTITY8 : if BRAM_NAME = "ifmap_layer0_entity8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000f1000000ee000000ec000000de000000ba000000c2000000da000000de",
            INIT_01 => X"000000f5000000f2000000f1000000f0000000eb000000f4000000f5000000f3",
            INIT_02 => X"000000f3000000f3000000f3000000f9000000f8000000f5000000f0000000e3",
            INIT_03 => X"000000f6000000f3000000ea000000f1000000f7000000ef000000eb000000f5",
            INIT_04 => X"000000ee000000f0000000f0000000df000000b8000000c9000000e2000000e5",
            INIT_05 => X"000000f8000000f5000000f5000000f3000000e8000000f5000000f7000000f3",
            INIT_06 => X"000000f4000000ee000000ee000000fb000000fb000000f3000000ef000000e6",
            INIT_07 => X"000000fb000000fa000000ec000000f0000000fc000000f3000000ec000000f8",
            INIT_08 => X"000000e4000000ef000000ee000000db000000b5000000c7000000de000000e1",
            INIT_09 => X"000000f7000000ee000000ef000000eb000000e4000000ec000000f4000000eb",
            INIT_0A => X"000000ef000000e8000000d7000000ec000000f6000000f1000000ec000000e5",
            INIT_0B => X"000000f7000000fb000000e8000000f1000000fc000000f2000000eb000000f8",
            INIT_0C => X"000000e1000000eb000000e4000000d6000000b3000000c2000000d8000000de",
            INIT_0D => X"000000f7000000e6000000ec000000e1000000dd000000e6000000ef000000e5",
            INIT_0E => X"000000f1000000e5000000b0000000ba000000ee000000f0000000ea000000e6",
            INIT_0F => X"000000f3000000f8000000e4000000ee000000fb000000ef000000e9000000f8",
            INIT_10 => X"000000d9000000e7000000dd000000d2000000ac000000c1000000d9000000df",
            INIT_11 => X"000000ee000000d6000000e8000000db000000d7000000e1000000eb000000da",
            INIT_12 => X"000000ef000000e5000000b2000000b0000000e4000000ee000000e3000000e5",
            INIT_13 => X"000000f0000000f6000000e8000000e7000000f5000000ea000000e7000000f7",
            INIT_14 => X"000000d5000000e1000000d5000000ce000000a4000000bf000000d5000000dc",
            INIT_15 => X"000000ce000000c8000000e3000000d6000000d6000000da000000e6000000d6",
            INIT_16 => X"000000e9000000e6000000ad00000082000000cf000000ed000000ce000000d0",
            INIT_17 => X"000000e6000000f2000000e7000000dd000000e8000000db000000e1000000f4",
            INIT_18 => X"000000d0000000d9000000c9000000c400000096000000b9000000ca000000d4",
            INIT_19 => X"000000af000000b9000000dd000000d4000000d3000000d0000000db000000d3",
            INIT_1A => X"000000bb000000b80000009d00000089000000c5000000d2000000bd000000bb",
            INIT_1B => X"000000d8000000e7000000db000000d1000000da000000ce000000dc000000dd",
            INIT_1C => X"000000cb000000ce000000cc000000c500000093000000b3000000c9000000d3",
            INIT_1D => X"000000cb000000c0000000ce000000ce000000cd000000c6000000d2000000d0",
            INIT_1E => X"00000049000000580000005e000000640000006a0000007a0000009b000000b3",
            INIT_1F => X"000000c1000000ce000000b9000000c6000000d7000000ca000000b70000006f",
            INIT_20 => X"000000b3000000a1000000af000000aa0000008c000000a0000000ad000000b3",
            INIT_21 => X"000000c4000000ba000000b9000000c3000000bd000000b4000000b8000000bb",
            INIT_22 => X"0000005a000000800000007e0000007e0000008000000080000000890000009f",
            INIT_23 => X"0000009f000000b0000000890000009c000000ac0000009e0000007c00000058",
            INIT_24 => X"00000080000000720000007200000072000000700000007b0000007e0000007b",
            INIT_25 => X"000000a7000000a0000000920000009800000090000000890000008600000086",
            INIT_26 => X"000000680000007800000083000000820000008c000000900000008b00000093",
            INIT_27 => X"0000007500000080000000690000006a0000008d000000960000008300000095",
            INIT_28 => X"0000006a00000068000000730000006b00000058000000620000006600000059",
            INIT_29 => X"0000009200000097000000860000007b0000007300000071000000760000006b",
            INIT_2A => X"000000800000007a000000680000006f000000780000007f0000007f00000080",
            INIT_2B => X"000000700000006d0000007500000072000000b60000008b0000006e00000086",
            INIT_2C => X"0000005e00000071000000890000008e0000006a0000006e0000006800000058",
            INIT_2D => X"00000097000000a5000000a5000000940000007d0000007f0000009200000074",
            INIT_2E => X"000000bf000000a5000000720000007b0000007f0000007f000000820000008e",
            INIT_2F => X"0000006c0000006c0000006d0000008c000000b8000000640000008e000000b4",
            INIT_30 => X"000000760000006d000000820000008100000068000000840000008200000064",
            INIT_31 => X"0000008b0000009a000000a50000009b00000097000000a8000000ab0000009a",
            INIT_32 => X"000000c1000000b300000089000000860000008c000000810000007d00000082",
            INIT_33 => X"0000006d0000006900000054000000a00000009800000070000000b9000000cb",
            INIT_34 => X"000000790000006c00000065000000710000006a0000007e0000008600000078",
            INIT_35 => X"000000950000009e000000a1000000990000009f000000a10000009100000083",
            INIT_36 => X"000000b1000000b6000000a1000000960000009b000000910000009300000092",
            INIT_37 => X"000000600000004e000000500000009d0000007600000094000000b5000000b5",
            INIT_38 => X"00000086000000730000007100000074000000720000007d000000800000007f",
            INIT_39 => X"000000b9000000be000000bf000000be000000b8000000b0000000a80000009f",
            INIT_3A => X"000000a8000000af000000ad000000ac000000b8000000be000000c4000000c5",
            INIT_3B => X"0000005100000043000000470000005700000063000000a3000000a5000000ab",
            INIT_3C => X"000000c1000000b8000000b300000099000000910000009a0000009500000097",
            INIT_3D => X"000000c8000000d4000000d2000000d1000000d0000000cf000000cd000000c9",
            INIT_3E => X"0000009b0000008b0000008700000086000000ab000000c3000000c9000000c6",
            INIT_3F => X"000000560000005a0000005c0000004900000071000000a8000000a1000000a5",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000c9000000c6000000b9000000af000000b0000000a70000009f000000a5",
            INIT_41 => X"000000be000000c9000000d0000000d2000000d2000000d2000000d0000000cd",
            INIT_42 => X"000000990000008e0000007a0000006c00000094000000a9000000aa000000aa",
            INIT_43 => X"0000006f00000098000000b5000000930000008e000000a7000000a5000000a7",
            INIT_44 => X"000000ca000000b60000008f0000008d0000009d000000ae000000aa0000009d",
            INIT_45 => X"000000a2000000a7000000b5000000bf000000ca000000d1000000d3000000d0",
            INIT_46 => X"000000a0000000a70000009d00000093000000a9000000b2000000a00000009b",
            INIT_47 => X"0000009400000096000000960000009e0000009c000000a1000000a2000000a9",
            INIT_48 => X"000000c2000000b1000000a40000008a000000790000008000000094000000a2",
            INIT_49 => X"000000b0000000ac000000ac000000aa000000ab000000b2000000bc000000c7",
            INIT_4A => X"000000ac000000af000000ad000000aa000000b5000000b0000000a8000000b4",
            INIT_4B => X"000000990000007d000000760000008500000096000000a3000000a5000000a8",
            INIT_4C => X"000000b0000000ba000000c5000000bc000000a60000007f000000750000008f",
            INIT_4D => X"000000ba000000bf000000be000000b9000000b2000000ab000000a3000000a9",
            INIT_4E => X"000000b2000000af000000ac000000ad000000b1000000ac000000a5000000b4",
            INIT_4F => X"0000009000000062000000570000006700000074000000880000009c000000a4",
            INIT_50 => X"000000aa000000b3000000ae000000b0000000b0000000a8000000a5000000a6",
            INIT_51 => X"00000096000000a8000000b5000000b9000000bd000000be000000b8000000a4",
            INIT_52 => X"000000a2000000ab000000ad000000ad000000ad0000009d0000007600000081",
            INIT_53 => X"0000004e0000005600000054000000500000005f0000006a0000007000000085",
            INIT_54 => X"000000b0000000b3000000b0000000ae000000af000000b1000000ac000000a5",
            INIT_55 => X"0000005e0000007e000000ab000000af000000ad000000ab000000ab000000a4",
            INIT_56 => X"000000750000008800000098000000a2000000ac0000008e0000005500000058",
            INIT_57 => X"000000270000003f000000580000004f000000500000005e000000680000006c",
            INIT_58 => X"0000008b0000009a000000ad000000af000000af000000b2000000a60000007c",
            INIT_59 => X"0000006c00000083000000a9000000ae0000009a0000007a0000007e00000082",
            INIT_5A => X"0000006c0000006d000000710000007900000085000000860000007200000072",
            INIT_5B => X"000000260000002b0000003b00000049000000450000004b000000560000005f",
            INIT_5C => X"00000064000000740000009e000000a30000009f000000a0000000960000006f",
            INIT_5D => X"0000008300000095000000a8000000ac00000097000000730000007000000068",
            INIT_5E => X"00000054000000640000006c0000006a0000006a0000006a0000006b00000077",
            INIT_5F => X"00000025000000280000002c0000003700000041000000440000004900000045",
            INIT_60 => X"0000007700000080000000a2000000a10000009a000000970000008a00000071",
            INIT_61 => X"0000006200000065000000720000008400000092000000900000008800000081",
            INIT_62 => X"0000004b0000004800000050000000630000006c0000006d0000006700000065",
            INIT_63 => X"00000027000000290000002d000000340000003a0000003d0000004d00000055",
            INIT_64 => X"0000007c000000840000008f00000094000000970000009a0000008800000074",
            INIT_65 => X"00000065000000630000005b00000056000000570000005b0000006700000076",
            INIT_66 => X"000000450000004a0000004800000048000000520000005e0000006300000065",
            INIT_67 => X"000000300000002f00000030000000330000003200000034000000440000004e",
            INIT_68 => X"0000005100000052000000560000005c000000630000006a0000006400000060",
            INIT_69 => X"000000580000005e0000005b0000005700000054000000510000004f00000052",
            INIT_6A => X"0000003b00000040000000480000004a0000004c00000044000000440000004d",
            INIT_6B => X"000000300000003400000030000000310000003200000031000000360000003f",
            INIT_6C => X"000000440000003e0000003d0000003c0000003700000036000000390000003b",
            INIT_6D => X"000000420000004500000044000000480000004d0000004f0000004f0000004e",
            INIT_6E => X"00000039000000380000003c000000410000005200000061000000470000003d",
            INIT_6F => X"0000002300000032000000320000003200000031000000300000003100000035",
            INIT_70 => X"000000370000003500000035000000310000002d0000002c0000003000000032",
            INIT_71 => X"0000004400000047000000420000003c00000038000000380000003b0000003a",
            INIT_72 => X"000000330000003a00000038000000350000004b000000680000004b0000003b",
            INIT_73 => X"0000001400000025000000350000003200000033000000310000003000000031",
            INIT_74 => X"000000300000002e0000002e0000002c00000029000000280000002c0000002d",
            INIT_75 => X"0000003d000000440000004400000044000000410000003f0000003900000033",
            INIT_76 => X"0000002f0000003000000038000000310000003f0000005d0000004200000032",
            INIT_77 => X"000000050000000e0000002e0000003400000033000000310000002f0000002f",
            INIT_78 => X"0000003b0000003800000036000000320000002d000000290000002b00000027",
            INIT_79 => X"000000310000003a0000003d000000400000004000000042000000400000003e",
            INIT_7A => X"0000002f0000002f00000030000000320000003b000000550000003500000024",
            INIT_7B => X"00000003000000030000001800000036000000320000002d0000002e0000002e",
            INIT_7C => X"0000003a0000003800000038000000380000003600000034000000320000002f",
            INIT_7D => X"000000140000001e000000270000002d0000003200000035000000370000003a",
            INIT_7E => X"0000002e0000002d0000002d0000002c0000003600000048000000210000000b",
            INIT_7F => X"00000007000000030000000800000025000000340000002b0000002c0000002c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY8;


    MEM_IFMAP_LAYER0_ENTITY9 : if BRAM_NAME = "ifmap_layer0_entity9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a6000000a8000000a6000000b1000000be000000b0000000a70000009b",
            INIT_01 => X"000000b8000000b8000000bb000000bb000000bb000000bb000000b3000000aa",
            INIT_02 => X"000000bd000000bc000000bb000000bb000000ba000000b8000000b4000000b6",
            INIT_03 => X"000000c0000000ca000000c9000000c9000000c3000000bc000000bb000000bb",
            INIT_04 => X"0000009f0000009a0000009b000000b3000000bb000000ab000000a300000099",
            INIT_05 => X"000000a5000000a2000000ab000000a9000000af000000ab000000a50000009f",
            INIT_06 => X"000000a8000000a9000000ad000000a7000000a5000000a6000000a4000000aa",
            INIT_07 => X"000000bd000000cb000000ca000000cc000000ca000000be000000ad000000a9",
            INIT_08 => X"000000bc000000b0000000ae000000bb000000b8000000a8000000a00000009b",
            INIT_09 => X"000000b9000000bc000000c2000000c0000000be000000b1000000b3000000b6",
            INIT_0A => X"000000bf000000c1000000c5000000c3000000c2000000c1000000c2000000c1",
            INIT_0B => X"000000bd000000cc000000ce000000d0000000cf000000ce000000c5000000bf",
            INIT_0C => X"000000c5000000c7000000b9000000b4000000b1000000a60000009d00000097",
            INIT_0D => X"000000cb000000c4000000c5000000d2000000c6000000cd000000cc000000b6",
            INIT_0E => X"000000cc000000c5000000d2000000cf000000cb000000d2000000cf000000cd",
            INIT_0F => X"000000c0000000ce000000cf000000d1000000c9000000cc000000c6000000d0",
            INIT_10 => X"000000c4000000bf000000b5000000b1000000ae000000a80000009e00000097",
            INIT_11 => X"000000ca000000b9000000b9000000c4000000b9000000bd000000c2000000b7",
            INIT_12 => X"000000bc000000be000000c7000000c3000000c0000000c8000000c7000000c7",
            INIT_13 => X"000000c4000000cf000000cc000000ce000000c4000000c9000000c7000000c9",
            INIT_14 => X"000000c3000000c4000000ae000000ab000000ae000000a70000009c00000094",
            INIT_15 => X"000000bf000000bd000000bd000000bb000000b8000000bd000000be000000c0",
            INIT_16 => X"000000c1000000c0000000bc000000c0000000c6000000bb000000c3000000be",
            INIT_17 => X"000000c4000000d1000000d0000000d4000000d1000000cb000000ce000000cd",
            INIT_18 => X"000000c3000000cb000000b0000000a8000000ae000000a50000009900000094",
            INIT_19 => X"000000c3000000c5000000c2000000b6000000be000000bb000000bc000000bc",
            INIT_1A => X"000000c9000000c5000000c5000000c6000000cd000000c8000000c1000000c4",
            INIT_1B => X"000000c3000000cf000000cb000000c5000000c3000000c6000000c8000000c5",
            INIT_1C => X"000000d1000000c7000000bc000000ac000000ac000000a30000009b00000099",
            INIT_1D => X"000000c4000000bb000000bc000000c1000000bf000000bd000000be000000c4",
            INIT_1E => X"000000c8000000c4000000c9000000c2000000ce000000c4000000c2000000ca",
            INIT_1F => X"000000bd000000c7000000c4000000c8000000c9000000c8000000bb000000b5",
            INIT_20 => X"000000be000000b0000000b0000000ae000000ac000000a30000009f000000a0",
            INIT_21 => X"000000b6000000ac000000aa000000b5000000b0000000b0000000af000000b4",
            INIT_22 => X"000000bb000000b4000000bc000000b1000000bb000000b5000000b2000000bb",
            INIT_23 => X"000000b8000000c2000000c0000000c5000000bc000000bc000000c4000000c7",
            INIT_24 => X"000000b0000000b4000000ab000000aa000000ac000000a2000000a7000000ab",
            INIT_25 => X"0000009e0000009900000092000000960000009c000000960000009c0000009b",
            INIT_26 => X"000000a60000009c000000a20000009d0000009d000000a4000000a6000000a6",
            INIT_27 => X"000000b6000000c2000000c1000000c5000000bd000000bc000000c7000000c8",
            INIT_28 => X"000000ae000000b6000000b1000000ad000000b0000000a8000000b4000000af",
            INIT_29 => X"000000ad000000a8000000a30000009f0000009a0000009f000000a00000009c",
            INIT_2A => X"000000ac000000a7000000a8000000a0000000a2000000a0000000a4000000aa",
            INIT_2B => X"000000b7000000c1000000bf000000c5000000c4000000c4000000c3000000c2",
            INIT_2C => X"000000b6000000ae000000aa000000b7000000bb000000b2000000bb000000b5",
            INIT_2D => X"000000c1000000c1000000bb000000b8000000b5000000b4000000b3000000b3",
            INIT_2E => X"000000c0000000c0000000ba000000b8000000b9000000bc000000c0000000c1",
            INIT_2F => X"000000ba000000c4000000bf000000be000000bd000000c0000000bc000000bb",
            INIT_30 => X"000000c1000000950000008400000099000000ab000000ba000000be000000b9",
            INIT_31 => X"000000c4000000c3000000c1000000bf000000bc000000ba000000bf000000c6",
            INIT_32 => X"000000bf000000c0000000be000000bc000000bc000000be000000c0000000c3",
            INIT_33 => X"000000c1000000cc000000ca000000ca000000c5000000c3000000c1000000bf",
            INIT_34 => X"0000006d0000005e00000074000000840000009e000000bc000000c2000000ba",
            INIT_35 => X"000000c7000000c4000000c1000000bf000000c2000000c2000000b100000091",
            INIT_36 => X"000000c6000000c7000000c4000000c4000000c6000000c8000000c7000000c7",
            INIT_37 => X"000000b9000000c6000000c5000000c6000000c4000000c4000000c4000000c5",
            INIT_38 => X"0000005c0000008d000000b8000000c2000000c6000000c4000000c5000000ba",
            INIT_39 => X"000000cc000000cc000000c9000000c3000000b30000008e0000006800000054",
            INIT_3A => X"000000bf000000c2000000c2000000c2000000c7000000cc000000cc000000cc",
            INIT_3B => X"000000b5000000c0000000be000000bf000000be000000be000000be000000bd",
            INIT_3C => X"000000b1000000c9000000c8000000c5000000c8000000c6000000c7000000b8",
            INIT_3D => X"000000cd000000d0000000ca000000ad000000800000005d0000005400000075",
            INIT_3E => X"000000c3000000c5000000c4000000c3000000c7000000c7000000c8000000ca",
            INIT_3F => X"000000b2000000be000000bd000000bf000000bf000000c2000000c3000000c1",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d6000000d0000000ce000000cd000000d0000000cb000000c9000000b9",
            INIT_41 => X"000000cb000000b50000008c000000690000005b0000004c0000005c000000af",
            INIT_42 => X"000000c2000000c2000000c2000000c1000000c2000000c5000000ca000000ce",
            INIT_43 => X"000000b4000000be000000be000000c1000000bf000000c1000000c3000000c2",
            INIT_44 => X"000000d0000000d3000000d4000000d4000000d6000000cf000000cc000000bb",
            INIT_45 => X"0000008400000063000000540000005400000057000000470000007c000000cb",
            INIT_46 => X"000000c4000000c5000000c0000000c3000000cb000000cb000000be000000a7",
            INIT_47 => X"000000b7000000c0000000bf000000c1000000bf000000c0000000c2000000c2",
            INIT_48 => X"000000d0000000d3000000d3000000d4000000d6000000cf000000cf000000be",
            INIT_49 => X"00000053000000560000005400000053000000570000004800000089000000d3",
            INIT_4A => X"000000cc000000cb000000b6000000a30000009b000000830000006b00000059",
            INIT_4B => X"000000b6000000bf000000c0000000c1000000bf000000c2000000c6000000ca",
            INIT_4C => X"000000d5000000d4000000d4000000d5000000d7000000d1000000d2000000bf",
            INIT_4D => X"0000005d000000570000004c0000003f0000003a0000002f00000071000000cc",
            INIT_4E => X"0000009f0000007a0000004d0000003a0000003e00000046000000500000005a",
            INIT_4F => X"000000b9000000c4000000c4000000c8000000c8000000c9000000c2000000b4",
            INIT_50 => X"000000d4000000d1000000d2000000d1000000d3000000cf000000d0000000bf",
            INIT_51 => X"000000580000004a00000044000000330000002500000041000000650000009d",
            INIT_52 => X"000000480000003e0000002e000000370000004900000055000000560000005b",
            INIT_53 => X"000000ba000000c4000000c3000000b80000009e000000850000006b0000004e",
            INIT_54 => X"000000c8000000d1000000ce000000cf000000d1000000cb000000ca000000ba",
            INIT_55 => X"0000006000000032000000350000002d00000064000000970000008c00000095",
            INIT_56 => X"000000420000005900000070000000620000004800000080000000a00000009c",
            INIT_57 => X"000000b2000000bc000000b7000000ad000000a3000000a60000008300000043",
            INIT_58 => X"000000d1000000d1000000d0000000d2000000d2000000ca000000c9000000b9",
            INIT_59 => X"000000a8000000940000009200000090000000bd000000d7000000d3000000d2",
            INIT_5A => X"0000009f000000b1000000b2000000a30000009a000000c0000000ce000000ca",
            INIT_5B => X"000000b0000000bc000000c1000000c4000000c2000000bf000000b20000009c",
            INIT_5C => X"000000b7000000b9000000bc000000c0000000c4000000c0000000bc000000b0",
            INIT_5D => X"000000ad000000ab000000aa000000aa000000ad000000b3000000b2000000b6",
            INIT_5E => X"000000aa000000a5000000a1000000a5000000a7000000a1000000a0000000a9",
            INIT_5F => X"0000009c000000a4000000a30000009d0000009600000098000000a0000000aa",
            INIT_60 => X"0000005d0000005e00000061000000660000006b0000006e0000006300000072",
            INIT_61 => X"00000065000000530000004e0000004d00000050000000580000005500000058",
            INIT_62 => X"000000710000006f0000006e0000006c0000006b0000006a0000006c00000071",
            INIT_63 => X"0000007c0000007a000000790000007800000077000000780000007700000075",
            INIT_64 => X"0000007100000072000000700000007300000075000000710000006d0000007a",
            INIT_65 => X"0000006c0000006e0000006d0000006e0000006d0000006f000000700000006f",
            INIT_66 => X"00000068000000650000006a0000006c0000006b000000690000007000000073",
            INIT_67 => X"000000650000005e00000066000000670000006d0000006d0000006b0000006a",
            INIT_68 => X"0000005e00000062000000680000006d000000700000006b0000006100000078",
            INIT_69 => X"0000004e000000500000004f0000005200000056000000580000005d0000005e",
            INIT_6A => X"0000004100000041000000420000004300000045000000480000004f00000050",
            INIT_6B => X"0000004d000000350000003f0000004300000040000000420000004100000040",
            INIT_6C => X"0000003d0000003f00000042000000420000004500000041000000370000005b",
            INIT_6D => X"0000003f0000003d0000003c00000039000000390000003c0000004000000042",
            INIT_6E => X"0000003c0000003b00000039000000380000003a00000040000000420000003f",
            INIT_6F => X"0000005c0000004b00000031000000340000003900000038000000390000003a",
            INIT_70 => X"0000004100000040000000430000004300000044000000420000003c0000005d",
            INIT_71 => X"0000003d0000003c0000003b0000003b0000003b0000003e0000004100000045",
            INIT_72 => X"00000038000000380000003700000037000000380000003a0000003f00000040",
            INIT_73 => X"00000051000000610000005d0000004100000035000000380000003a00000039",
            INIT_74 => X"0000003b000000390000003b00000039000000390000003d0000003900000059",
            INIT_75 => X"0000003d0000003b0000003d0000003c00000036000000380000003a0000003c",
            INIT_76 => X"0000003d0000003d0000003c0000003c000000390000003a0000003d00000041",
            INIT_77 => X"000000430000003b000000590000006100000046000000390000003e00000042",
            INIT_78 => X"0000003f0000003e0000003e0000003e0000003e0000003f0000003c00000059",
            INIT_79 => X"000000510000004e000000510000005400000052000000410000003d0000003e",
            INIT_7A => X"0000004000000042000000430000005000000053000000550000005400000058",
            INIT_7B => X"0000004b0000003d000000390000004c00000067000000560000003800000034",
            INIT_7C => X"0000004100000043000000420000003f0000003c0000003d0000003c0000005c",
            INIT_7D => X"0000004600000048000000490000004900000048000000410000004300000042",
            INIT_7E => X"0000003e00000040000000400000004b0000004b0000004b0000004a00000049",
            INIT_7F => X"00000049000000400000003c0000003900000040000000580000005600000041",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY9;


    MEM_IFMAP_LAYER0_ENTITY10 : if BRAM_NAME = "ifmap_layer0_entity10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ad000000ad000000ab000000b9000000c0000000b3000000b00000009c",
            INIT_01 => X"000000b5000000b6000000b8000000b9000000b8000000b6000000b3000000af",
            INIT_02 => X"000000bd000000bb000000ba000000ba000000b9000000b7000000b3000000b3",
            INIT_03 => X"000000b7000000ca000000c4000000c5000000c3000000bc000000bb000000bb",
            INIT_04 => X"000000a40000009f000000a2000000be000000c3000000b8000000b30000009b",
            INIT_05 => X"000000a7000000a4000000ae000000ab000000b0000000a9000000a5000000a3",
            INIT_06 => X"000000a9000000ab000000af000000a9000000a6000000a8000000a6000000ac",
            INIT_07 => X"000000be000000d7000000d0000000ce000000cc000000bf000000ae000000aa",
            INIT_08 => X"000000a8000000b2000000c1000000cb000000c4000000b9000000b20000009a",
            INIT_09 => X"000000bc000000be000000c5000000c3000000c4000000be000000af000000a0",
            INIT_0A => X"000000bf000000c1000000c6000000c4000000c3000000c2000000c3000000c4",
            INIT_0B => X"000000bf000000d7000000d0000000ce000000cd000000cd000000c4000000c0",
            INIT_0C => X"00000080000000bc000000c5000000ca000000c3000000bc000000b20000009a",
            INIT_0D => X"0000009400000095000000950000009e0000009b0000009a000000980000006c",
            INIT_0E => X"0000009f000000ae000000a3000000a8000000ad000000a3000000a1000000a7",
            INIT_0F => X"000000bc000000d4000000cd000000cc000000ce000000cc000000d0000000bc",
            INIT_10 => X"0000007e000000bd000000c4000000c6000000bf000000bb000000b10000009a",
            INIT_11 => X"000000710000007600000078000000730000006b0000006a0000008b00000080",
            INIT_12 => X"000000700000008800000070000000760000007e000000720000007200000077",
            INIT_13 => X"000000be000000d6000000cd000000ce000000ce000000c9000000cb000000a0",
            INIT_14 => X"00000093000000b7000000c8000000c5000000bd000000bb000000ae00000097",
            INIT_15 => X"0000009d0000009500000092000000aa000000a500000091000000a8000000a9",
            INIT_16 => X"000000b1000000bc000000b3000000b0000000bd000000b0000000b2000000b4",
            INIT_17 => X"000000be000000d8000000d1000000d0000000d0000000cf000000d0000000c4",
            INIT_18 => X"0000006000000093000000c6000000c2000000bd000000b9000000ac00000098",
            INIT_19 => X"0000008b00000080000000790000009800000098000000900000009700000095",
            INIT_1A => X"000000a400000096000000ad00000096000000a2000000aa000000970000009c",
            INIT_1B => X"000000bc000000d4000000cf000000d3000000d2000000cc000000a60000009c",
            INIT_1C => X"0000006500000077000000b5000000c2000000bb000000b6000000ac0000009b",
            INIT_1D => X"0000007f0000008700000087000000920000007800000083000000830000007b",
            INIT_1E => X"0000009f0000007b000000840000006d0000007b000000830000007b0000007b",
            INIT_1F => X"000000ba000000d0000000c9000000c9000000c7000000bf000000840000007b",
            INIT_20 => X"000000af000000ab000000ba000000c0000000b9000000b4000000af000000a1",
            INIT_21 => X"000000aa000000ad000000ac000000af000000a6000000ac000000a5000000a2",
            INIT_22 => X"000000be000000b2000000ac000000a3000000af000000b2000000b2000000ac",
            INIT_23 => X"000000b9000000d1000000c9000000c8000000cd000000c8000000b0000000ac",
            INIT_24 => X"000000b7000000c2000000c0000000be000000ba000000b4000000b7000000ac",
            INIT_25 => X"000000a2000000a40000009e0000009f000000a3000000a2000000a5000000a0",
            INIT_26 => X"000000b6000000a5000000a3000000a0000000a2000000ac000000ae000000a7",
            INIT_27 => X"000000b8000000d0000000ca000000ca000000cd000000ca000000c6000000c8",
            INIT_28 => X"000000b7000000c1000000c1000000c0000000be000000ba000000c4000000b1",
            INIT_29 => X"000000ac000000aa000000a6000000a40000009f000000a5000000a7000000a3",
            INIT_2A => X"000000b2000000ab000000ad000000a8000000ab000000a6000000a6000000a8",
            INIT_2B => X"000000b8000000d0000000c8000000c8000000c7000000c7000000c6000000c7",
            INIT_2C => X"000000c6000000be000000bb000000c9000000c8000000c3000000cc000000b7",
            INIT_2D => X"000000c6000000c6000000c2000000c1000000c1000000c1000000c1000000c2",
            INIT_2E => X"000000c5000000c4000000c4000000c5000000c6000000c3000000c3000000c6",
            INIT_2F => X"000000bb000000d1000000c8000000ca000000c9000000c9000000cb000000c9",
            INIT_30 => X"000000c40000009a0000008d000000a6000000b2000000c6000000cd000000b9",
            INIT_31 => X"000000ca000000c9000000c7000000c5000000c5000000c7000000ca000000ca",
            INIT_32 => X"000000c6000000c7000000c6000000c4000000c4000000c6000000c7000000c9",
            INIT_33 => X"000000bd000000d4000000ce000000cf000000ce000000cb000000ca000000c7",
            INIT_34 => X"0000006b0000005f0000007c00000090000000a5000000c8000000d0000000ba",
            INIT_35 => X"000000cc000000c9000000c6000000c5000000c7000000c7000000b30000008f",
            INIT_36 => X"000000cd000000cd000000c9000000c9000000cc000000ce000000cd000000cc",
            INIT_37 => X"000000b7000000cf000000ca000000ca000000cb000000cb000000cb000000cc",
            INIT_38 => X"0000005b0000008f000000c1000000ce000000cc000000d0000000d4000000ba",
            INIT_39 => X"000000cf000000cf000000cc000000c6000000b50000008e0000006500000051",
            INIT_3A => X"000000c5000000c6000000c5000000c5000000ca000000cf000000cf000000cf",
            INIT_3B => X"000000b5000000cc000000c5000000c4000000c5000000c5000000c5000000c5",
            INIT_3C => X"000000b3000000cf000000d4000000d1000000ce000000d2000000d6000000b8",
            INIT_3D => X"000000ce000000d2000000cb000000ae000000800000005d0000005300000074",
            INIT_3E => X"000000c9000000c9000000c7000000c6000000c9000000ca000000ca000000cc",
            INIT_3F => X"000000b4000000cb000000c6000000c6000000c7000000c9000000ca000000c8",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d9000000d4000000d6000000d6000000d5000000d6000000d7000000ba",
            INIT_41 => X"000000cc000000b50000008a0000006500000056000000490000005b000000af",
            INIT_42 => X"000000c8000000c9000000c9000000c7000000c6000000c7000000cb000000d0",
            INIT_43 => X"000000b6000000cc000000c8000000ca000000c9000000c9000000ca000000c8",
            INIT_44 => X"000000d3000000d6000000d9000000db000000d9000000d8000000d8000000bb",
            INIT_45 => X"0000008200000061000000510000004f00000052000000440000007b000000cc",
            INIT_46 => X"000000c6000000c7000000c1000000c4000000ca000000c9000000bc000000a5",
            INIT_47 => X"000000b6000000cc000000c7000000c9000000c8000000c8000000c7000000c6",
            INIT_48 => X"000000d2000000d6000000d8000000d8000000d6000000d5000000d9000000bc",
            INIT_49 => X"0000004d00000050000000500000004e000000530000004600000088000000d4",
            INIT_4A => X"000000cc000000c9000000b20000009f000000970000007e0000006600000053",
            INIT_4B => X"000000b4000000c9000000c5000000c7000000c6000000c8000000c9000000cb",
            INIT_4C => X"000000d8000000d7000000d8000000d7000000d5000000d6000000da000000bb",
            INIT_4D => X"000000510000004d000000450000003a000000370000002d00000070000000cc",
            INIT_4E => X"000000a00000007c0000004f0000003b0000003e000000460000004d00000050",
            INIT_4F => X"000000b4000000ca000000c8000000cb000000cd000000cd000000c4000000b5",
            INIT_50 => X"000000d4000000d4000000d6000000d3000000d1000000d2000000d8000000bc",
            INIT_51 => X"0000004d000000410000003e00000030000000210000003a0000005f0000009a",
            INIT_52 => X"000000480000003f0000002f0000003800000048000000540000005400000052",
            INIT_53 => X"000000b6000000ca000000c1000000b50000009e000000840000006b0000004e",
            INIT_54 => X"000000c8000000d4000000d3000000d1000000cf000000ce000000d2000000b8",
            INIT_55 => X"0000005a0000002e000000320000002d000000610000008f0000008500000091",
            INIT_56 => X"00000041000000580000007000000061000000470000007f0000009e00000096",
            INIT_57 => X"000000b0000000c5000000b5000000a8000000a2000000a50000008200000043",
            INIT_58 => X"000000d2000000d5000000d4000000d3000000d0000000cd000000d2000000b7",
            INIT_59 => X"000000a6000000930000009300000094000000bf000000d4000000d1000000d1",
            INIT_5A => X"000000a2000000b4000000b5000000a60000009d000000c3000000d0000000c8",
            INIT_5B => X"000000b1000000c7000000c1000000c3000000c5000000c1000000b40000009f",
            INIT_5C => X"000000b9000000bb000000be000000c2000000c2000000c3000000c4000000ae",
            INIT_5D => X"000000ad000000ae000000b0000000b2000000b5000000b7000000b5000000b8",
            INIT_5E => X"000000b0000000aa000000a6000000aa000000ac000000a6000000a4000000aa",
            INIT_5F => X"0000009e000000af000000a30000009d0000009b0000009d000000a5000000af",
            INIT_60 => X"0000006000000061000000640000006700000069000000700000006c00000070",
            INIT_61 => X"00000067000000570000005300000054000000570000005e0000005a0000005c",
            INIT_62 => X"00000076000000740000007300000071000000700000006f0000007000000073",
            INIT_63 => X"0000007c000000840000007a000000790000007b0000007c0000007b0000007a",
            INIT_64 => X"00000071000000710000006f0000007100000070000000710000007300000075",
            INIT_65 => X"0000006b0000006e0000006d0000006e0000006e0000006f000000700000006f",
            INIT_66 => X"0000006b000000680000006d0000006f0000006e0000006c0000007300000073",
            INIT_67 => X"00000065000000620000005f0000006400000070000000700000006e0000006d",
            INIT_68 => X"0000005d00000061000000660000006a0000006a000000690000006600000071",
            INIT_69 => X"0000004e0000004f0000004e0000005200000055000000590000005e0000005f",
            INIT_6A => X"0000004100000041000000410000004300000044000000470000004f00000050",
            INIT_6B => X"0000006400000047000000370000003c00000041000000420000004200000041",
            INIT_6C => X"0000003c0000003e000000400000004000000040000000410000003c00000054",
            INIT_6D => X"0000003f0000003d0000003c00000039000000380000003d0000004000000042",
            INIT_6E => X"0000003c0000003b0000003a000000380000003b000000410000004300000040",
            INIT_6F => X"000000800000007500000048000000380000003800000038000000390000003a",
            INIT_70 => X"0000003f0000003d000000410000003f0000003e0000003f0000003b00000053",
            INIT_71 => X"0000003d0000003c0000003a0000003a000000390000003c0000003e00000043",
            INIT_72 => X"0000003d0000003e0000003c0000003d0000003e000000400000004400000041",
            INIT_73 => X"0000006300000089000000880000005b000000410000003d0000003a0000003a",
            INIT_74 => X"0000003c0000003a0000003b00000037000000390000003d000000350000004f",
            INIT_75 => X"0000003f0000003d0000003e0000003c00000037000000390000003c0000003d",
            INIT_76 => X"0000003f000000400000003e0000003e0000003b0000003c0000003f00000043",
            INIT_77 => X"0000004a0000004f000000770000008e0000006e000000470000003c0000003e",
            INIT_78 => X"0000003e0000003e0000003e0000003f00000041000000420000003a00000052",
            INIT_79 => X"0000004d0000004a0000004c0000004f0000004f000000410000003e0000003f",
            INIT_7A => X"000000410000003e0000003f0000004c0000004e000000500000005000000054",
            INIT_7B => X"000000450000004000000042000000660000008d0000007c0000005600000042",
            INIT_7C => X"000000390000003b0000003a0000003a0000003a0000003a000000340000004e",
            INIT_7D => X"00000045000000460000004700000047000000450000003a0000003b0000003a",
            INIT_7E => X"000000440000003f0000003f000000490000004a000000490000004800000048",
            INIT_7F => X"00000044000000410000003f000000420000005800000080000000800000005a",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY10;


    MEM_IFMAP_LAYER0_ENTITY11 : if BRAM_NAME = "ifmap_layer0_entity11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b4000000b5000000b7000000ca000000cd000000c1000000bb00000095",
            INIT_01 => X"000000bd000000bd000000c0000000c0000000c0000000c1000000bd000000b6",
            INIT_02 => X"000000be000000c0000000c1000000c1000000c0000000bd000000b9000000ba",
            INIT_03 => X"000000ab000000d4000000d1000000ca000000c3000000bc000000bb000000bb",
            INIT_04 => X"000000b3000000b3000000be000000e0000000e3000000d7000000cc0000009d",
            INIT_05 => X"000000b7000000b4000000be000000bb000000c3000000c3000000bb000000b3",
            INIT_06 => X"000000bc000000bc000000bf000000b9000000b7000000b8000000b7000000bc",
            INIT_07 => X"000000b7000000e3000000de000000df000000e0000000d3000000c2000000be",
            INIT_08 => X"000000b8000000c4000000d5000000df000000db000000d5000000c900000099",
            INIT_09 => X"000000ca000000cc000000d2000000d0000000d4000000d3000000c3000000b1",
            INIT_0A => X"000000d0000000d0000000d4000000d2000000d1000000d0000000d1000000d1",
            INIT_0B => X"000000b8000000e0000000d7000000da000000df000000de000000d5000000d0",
            INIT_0C => X"00000083000000c9000000dc000000e2000000de000000d3000000cf000000a6",
            INIT_0D => X"000000ab000000a6000000a7000000b2000000b1000000a60000009e00000077",
            INIT_0E => X"000000a5000000b4000000ba000000b9000000ba000000b2000000b2000000b7",
            INIT_0F => X"000000ba000000e6000000df000000e0000000dd000000dc000000e4000000cf",
            INIT_10 => X"0000008e000000d6000000e1000000e0000000da000000ca000000cb000000a7",
            INIT_11 => X"000000830000007c0000007e0000008100000081000000780000009800000099",
            INIT_12 => X"0000007b0000008d00000088000000880000008a000000820000008400000086",
            INIT_13 => X"000000b9000000e3000000dc000000de000000d9000000da000000e3000000ba",
            INIT_14 => X"000000a5000000d1000000da000000dc000000d9000000cb000000c9000000a4",
            INIT_15 => X"000000ac000000a3000000a0000000b3000000b40000009c000000b5000000c4",
            INIT_16 => X"000000be000000c6000000c0000000bf000000c9000000be000000c1000000bf",
            INIT_17 => X"000000bc000000e8000000e1000000df000000e1000000e1000000e1000000d4",
            INIT_18 => X"00000068000000ac000000d6000000d9000000d9000000c8000000c6000000a4",
            INIT_19 => X"000000a00000009700000090000000a5000000af000000a6000000a50000009e",
            INIT_1A => X"000000b9000000ad000000b7000000aa000000b6000000bd000000ad000000b2",
            INIT_1B => X"000000bc000000e7000000e0000000dd000000e2000000dc000000b2000000a6",
            INIT_1C => X"0000006f00000092000000cb000000da000000d8000000c7000000c9000000a9",
            INIT_1D => X"000000900000008f0000008f0000009b000000900000009d0000009500000086",
            INIT_1E => X"000000b00000008e0000008d0000007f0000008e000000940000008e00000093",
            INIT_1F => X"000000ba000000e4000000dc000000d9000000dc000000d10000009500000089",
            INIT_20 => X"000000c5000000c1000000cd000000db000000d9000000c7000000ce000000b1",
            INIT_21 => X"000000bd000000bb000000ba000000c0000000b8000000bb000000b7000000b8",
            INIT_22 => X"000000c8000000bc000000ba000000b2000000bf000000c2000000c2000000c0",
            INIT_23 => X"000000b9000000e4000000dd000000db000000db000000d6000000c6000000c1",
            INIT_24 => X"000000d2000000dc000000d6000000d7000000d6000000c5000000d4000000ba",
            INIT_25 => X"000000ba000000b9000000b4000000b6000000ba000000b6000000bb000000b9",
            INIT_26 => X"000000c6000000b6000000b6000000b5000000b8000000c3000000c6000000c1",
            INIT_27 => X"000000b7000000e3000000de000000df000000df000000dd000000de000000de",
            INIT_28 => X"000000cc000000d6000000d4000000d7000000d8000000c8000000de000000bc",
            INIT_29 => X"000000bf000000bc000000b8000000b5000000b0000000b6000000b8000000b5",
            INIT_2A => X"000000c9000000ba000000b8000000b6000000b9000000b8000000ba000000bd",
            INIT_2B => X"000000b8000000e3000000dc000000db000000db000000dc000000dd000000df",
            INIT_2C => X"000000de000000d7000000d1000000dc000000e0000000cf000000e2000000bf",
            INIT_2D => X"000000df000000df000000db000000d9000000d7000000d6000000d7000000d9",
            INIT_2E => X"000000db000000d9000000d6000000d8000000da000000db000000dd000000df",
            INIT_2F => X"000000ba000000e3000000db000000d7000000d6000000d9000000db000000db",
            INIT_30 => X"000000d9000000ac00000099000000b5000000ce000000d4000000dc000000bc",
            INIT_31 => X"000000e2000000e1000000df000000de000000dc000000dd000000e1000000e2",
            INIT_32 => X"000000da000000dc000000db000000d9000000da000000dc000000dd000000e1",
            INIT_33 => X"000000bb000000e6000000e0000000e0000000e0000000de000000dc000000d9",
            INIT_34 => X"00000073000000630000007e0000009d000000c1000000d6000000df000000bd",
            INIT_35 => X"000000e2000000df000000dc000000da000000dd000000dd000000c60000009d",
            INIT_36 => X"000000e0000000e0000000dd000000dc000000df000000e1000000e0000000e2",
            INIT_37 => X"000000b7000000e2000000dd000000dd000000de000000de000000de000000df",
            INIT_38 => X"0000005a00000092000000c4000000dc000000e9000000de000000e2000000bd",
            INIT_39 => X"000000e4000000e3000000e0000000da000000ca000000a10000007100000054",
            INIT_3A => X"000000d9000000d8000000d7000000d7000000dc000000e0000000e1000000e2",
            INIT_3B => X"000000b6000000e1000000da000000d7000000d8000000d8000000d8000000d8",
            INIT_3C => X"000000b3000000da000000e1000000e1000000ea000000e0000000e5000000bb",
            INIT_3D => X"000000e1000000e4000000dd000000c0000000910000006a0000005800000073",
            INIT_3E => X"000000db000000d9000000d6000000d6000000d9000000da000000db000000df",
            INIT_3F => X"000000b7000000e2000000dc000000d9000000da000000dc000000dd000000db",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000e1000000e0000000e2000000e4000000e9000000de000000e9000000be",
            INIT_41 => X"000000d9000000c0000000920000006a0000005b0000005000000062000000b5",
            INIT_42 => X"000000d9000000da000000da000000d9000000da000000dd000000e1000000e0",
            INIT_43 => X"000000bc000000e3000000dc000000dd000000dd000000dd000000dd000000da",
            INIT_44 => X"000000dd000000e2000000e3000000e7000000e9000000dd000000ea000000bf",
            INIT_45 => X"0000008800000064000000500000004b0000004f0000004900000082000000d5",
            INIT_46 => X"000000de000000df000000d9000000d9000000dc000000d7000000c8000000ad",
            INIT_47 => X"000000bd000000e3000000db000000da000000db000000db000000dd000000dd",
            INIT_48 => X"000000dc000000e2000000e1000000e3000000e4000000d9000000e8000000bd",
            INIT_49 => X"0000004c0000004e0000004c0000004a000000500000004a00000090000000dd",
            INIT_4A => X"000000e2000000e1000000c9000000b0000000a1000000810000006400000053",
            INIT_4B => X"000000bb000000e1000000d9000000d7000000d7000000d9000000dc000000df",
            INIT_4C => X"000000e2000000e3000000e1000000e0000000e1000000d7000000e8000000bb",
            INIT_4D => X"000000520000004d000000450000003b000000380000003200000077000000d5",
            INIT_4E => X"000000a2000000850000005b000000410000003f000000420000004800000050",
            INIT_4F => X"000000bc000000e3000000dd000000dd000000df000000da000000cc000000b8",
            INIT_50 => X"000000e1000000e4000000e6000000df000000df000000de000000e7000000b7",
            INIT_51 => X"0000004e000000440000004300000035000000270000003c00000062000000a2",
            INIT_52 => X"000000430000003f000000310000003900000048000000530000005200000051",
            INIT_53 => X"000000c3000000df000000d7000000c6000000a80000008b0000006d0000004b",
            INIT_54 => X"000000d4000000e2000000e2000000de000000de000000e2000000e2000000b0",
            INIT_55 => X"0000005e0000003300000039000000350000006a000000960000008b0000009b",
            INIT_56 => X"000000430000005a00000072000000630000004900000082000000a10000009a",
            INIT_57 => X"000000be000000d0000000c5000000b7000000a9000000ab0000008600000045",
            INIT_58 => X"000000de000000de000000de000000df000000df000000e1000000e1000000af",
            INIT_59 => X"000000b3000000a00000009f0000009f000000cc000000e4000000e0000000de",
            INIT_5A => X"000000ad000000c0000000c1000000b2000000a9000000cf000000dc000000d6",
            INIT_5B => X"000000bd000000d2000000d1000000d8000000d6000000d2000000c3000000ab",
            INIT_5C => X"000000c7000000c9000000cc000000ce000000d1000000d7000000d4000000a6",
            INIT_5D => X"000000c4000000c2000000c1000000c0000000c2000000c5000000c3000000c7",
            INIT_5E => X"000000cd000000c8000000c4000000c8000000ca000000c4000000c2000000c4",
            INIT_5F => X"000000b5000000c9000000c5000000c5000000bf000000c0000000c5000000ce",
            INIT_60 => X"0000006a0000006b000000700000007600000078000000820000007800000065",
            INIT_61 => X"000000800000006c000000650000006200000063000000660000006200000065",
            INIT_62 => X"0000009e00000098000000960000009400000093000000920000009200000090",
            INIT_63 => X"00000092000000a7000000a5000000a8000000a8000000a8000000a6000000a4",
            INIT_64 => X"0000008800000089000000880000008a0000008600000086000000820000006f",
            INIT_65 => X"0000008300000083000000800000007f0000007e000000830000008600000084",
            INIT_66 => X"0000007e0000007c0000008000000081000000810000007f000000860000008a",
            INIT_67 => X"0000006000000073000000730000007700000084000000840000008200000081",
            INIT_68 => X"000000640000006c000000760000007a00000078000000780000007100000068",
            INIT_69 => X"0000005600000057000000550000005800000059000000550000005b00000060",
            INIT_6A => X"0000003c0000003f000000410000004200000043000000460000004f00000056",
            INIT_6B => X"0000004b0000003f00000032000000360000003b0000003c0000003c0000003b",
            INIT_6C => X"000000360000003b0000003f0000003a000000390000003d000000370000003d",
            INIT_6D => X"000000320000003100000032000000300000002f0000002f0000003300000038",
            INIT_6E => X"00000037000000320000002e0000002d0000002f000000350000003700000033",
            INIT_6F => X"00000068000000680000003a0000003000000034000000340000003400000036",
            INIT_70 => X"00000039000000370000003d0000003e0000003c000000410000003d00000044",
            INIT_71 => X"0000003600000038000000380000003b0000003a00000037000000380000003d",
            INIT_72 => X"0000003400000034000000330000003300000034000000370000003b00000039",
            INIT_73 => X"0000004b00000078000000710000004b00000039000000370000003500000033",
            INIT_74 => X"00000036000000340000003900000039000000350000003b000000340000003e",
            INIT_75 => X"0000003500000034000000380000003900000032000000300000003200000036",
            INIT_76 => X"0000003000000035000000370000003600000033000000340000003600000039",
            INIT_77 => X"000000320000003e000000650000007c0000005f0000003d0000003400000032",
            INIT_78 => X"0000003c0000003c0000003d0000003b000000370000003a000000350000003e",
            INIT_79 => X"0000004500000044000000480000004c0000004b0000003a0000003700000039",
            INIT_7A => X"00000035000000370000003a00000046000000490000004b0000004a0000004b",
            INIT_7B => X"00000033000000360000003a0000005b0000007f0000006b0000004500000033",
            INIT_7C => X"000000350000003900000038000000330000002e000000330000003300000040",
            INIT_7D => X"000000390000003c0000003e000000400000003e000000320000003300000034",
            INIT_7E => X"0000003700000034000000350000004000000040000000400000003e0000003c",
            INIT_7F => X"0000003200000034000000320000003500000048000000690000006700000046",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY11;


    MEM_IFMAP_LAYER0_ENTITY12 : if BRAM_NAME = "ifmap_layer0_entity12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d0000002c00000028000000170000001e000000300000004600000041",
            INIT_01 => X"0000003000000033000000350000002c0000000f0000000a000000280000002d",
            INIT_02 => X"000000370000003c000000510000005f0000005b0000005d0000005a00000041",
            INIT_03 => X"0000004300000036000000330000004d00000044000000290000006f00000070",
            INIT_04 => X"000000310000003100000041000000290000001e0000003c0000004f00000045",
            INIT_05 => X"0000003100000037000000450000004100000019000000070000002300000031",
            INIT_06 => X"0000003b0000003700000051000000570000005000000053000000550000004d",
            INIT_07 => X"0000003d0000004100000036000000380000002f0000001f0000007900000083",
            INIT_08 => X"00000036000000320000004a0000004000000029000000480000005400000049",
            INIT_09 => X"000000270000002f000000430000003c000000240000000b0000002000000036",
            INIT_0A => X"0000003f0000003000000055000000530000003e0000003b0000004d0000004b",
            INIT_0B => X"00000030000000490000004e000000460000002900000017000000800000008b",
            INIT_0C => X"0000003f00000037000000440000005000000036000000500000004b00000058",
            INIT_0D => X"0000002700000028000000330000002b00000025000000110000001c0000003a",
            INIT_0E => X"00000044000000320000005400000056000000460000004b0000006200000055",
            INIT_0F => X"00000026000000410000005d000000640000004b0000002f000000890000008e",
            INIT_10 => X"000000440000003d0000003d00000051000000420000006f000000590000005f",
            INIT_11 => X"0000003f00000033000000230000001f000000160000000f000000160000003e",
            INIT_12 => X"0000004e00000033000000530000004d00000047000000480000004b00000048",
            INIT_13 => X"000000580000004b0000005f0000006300000057000000570000009c00000095",
            INIT_14 => X"00000039000000400000003a000000470000004d000000520000005300000052",
            INIT_15 => X"00000047000000470000003d000000320000001c00000011000000140000003b",
            INIT_16 => X"0000004e00000046000000530000002900000038000000440000004300000045",
            INIT_17 => X"00000063000000700000006f0000005e0000005900000062000000ac0000009c",
            INIT_18 => X"00000031000000490000004a000000480000003b000000200000004000000045",
            INIT_19 => X"0000003f0000005600000055000000520000003e0000001d0000001200000031",
            INIT_1A => X"0000004e000000550000005e000000190000002b0000005f0000003400000022",
            INIT_1B => X"0000002f00000056000000830000006c0000006b0000006d000000b4000000a6",
            INIT_1C => X"0000003d000000500000004e000000510000004600000019000000350000003b",
            INIT_1D => X"000000190000004b00000058000000570000005e000000350000000a00000028",
            INIT_1E => X"00000062000000590000006500000032000000390000005c0000002d0000000d",
            INIT_1F => X"0000001800000034000000800000007c0000007c00000078000000b300000090",
            INIT_20 => X"0000004f0000003f000000590000007700000066000000310000002f00000044",
            INIT_21 => X"0000000e000000290000005a0000005900000060000000510000002200000042",
            INIT_22 => X"000000730000006e000000710000006f00000047000000430000005c00000034",
            INIT_23 => X"000000160000001f000000730000007c0000007f000000790000009c00000088",
            INIT_24 => X"00000037000000410000007b000000800000007200000037000000350000004d",
            INIT_25 => X"0000002500000014000000450000006a0000006e0000006f000000520000004f",
            INIT_26 => X"0000005c0000007300000078000000760000006100000053000000690000005c",
            INIT_27 => X"000000170000000e0000005f000000770000007f0000007d0000009300000090",
            INIT_28 => X"0000003100000064000000840000008100000070000000360000003a00000055",
            INIT_29 => X"000000530000003f0000005d0000007d0000006d000000680000005400000027",
            INIT_2A => X"00000039000000550000007f0000006d0000006e000000680000005e00000061",
            INIT_2B => X"000000150000000c0000005d000000720000007c0000007b0000009600000098",
            INIT_2C => X"0000004b00000080000000830000007e0000006b00000032000000350000006c",
            INIT_2D => X"00000093000000810000006e0000008a0000006b000000550000005b00000033",
            INIT_2E => X"0000005d0000005a000000730000007500000077000000710000007800000084",
            INIT_2F => X"000000090000000e00000065000000790000007d000000710000008d000000a0",
            INIT_30 => X"0000007700000082000000800000006a0000005c0000002b0000002a00000060",
            INIT_31 => X"00000084000000690000006e0000009400000089000000720000007b00000078",
            INIT_32 => X"000000770000007e000000780000008c00000086000000800000008700000092",
            INIT_33 => X"000000280000001200000063000000820000006a000000630000009100000098",
            INIT_34 => X"00000088000000850000006f00000064000000590000003b0000004200000061",
            INIT_35 => X"0000007f00000083000000880000008e00000091000000960000008c00000093",
            INIT_36 => X"000000880000009c0000008e0000009700000093000000880000007b0000007d",
            INIT_37 => X"00000053000000320000005c00000082000000700000006d0000009000000092",
            INIT_38 => X"00000085000000850000005e000000680000005f0000004b0000004800000069",
            INIT_39 => X"00000098000000a000000096000000930000008500000080000000870000008f",
            INIT_3A => X"000000a5000000a20000008a0000008a00000087000000840000009000000091",
            INIT_3B => X"0000004d0000003b0000005f00000076000000770000007e0000007f000000a3",
            INIT_3C => X"000000830000007b00000062000000650000005b00000044000000440000005e",
            INIT_3D => X"000000a200000093000000930000007c0000004f0000008a000000c100000093",
            INIT_3E => X"000000b30000009400000079000000900000009000000098000000ab000000b4",
            INIT_3F => X"000000540000001a0000003f000000700000007b00000080000000a0000000b4",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008100000078000000780000006e000000590000004a0000004f00000058",
            INIT_41 => X"000000a6000000a40000009c0000007200000057000000c0000000b800000078",
            INIT_42 => X"0000008f00000094000000ad000000bb000000b6000000b7000000a10000009a",
            INIT_43 => X"00000076000000290000002c0000006b0000007c0000008e000000c3000000b5",
            INIT_44 => X"0000006a0000006f00000064000000740000006000000067000000590000005b",
            INIT_45 => X"000000ac000000ac000000990000008c000000a8000000bb0000008000000072",
            INIT_46 => X"0000009c000000ab000000a5000000a1000000a30000009d000000a4000000a7",
            INIT_47 => X"0000005e0000002a0000004a0000006a00000072000000a700000091000000a1",
            INIT_48 => X"0000005b0000005f0000004e000000720000007a000000780000006100000065",
            INIT_49 => X"00000099000000a000000089000000a7000000cc000000810000006e00000073",
            INIT_4A => X"000000a5000000a20000009c000000b3000000b2000000aa000000ba000000b3",
            INIT_4B => X"0000007200000046000000590000005400000048000000680000008c0000009c",
            INIT_4C => X"00000064000000480000004c0000005a000000600000007a0000006b0000006e",
            INIT_4D => X"000000b4000000a60000009f000000bd0000008c000000570000007f0000006d",
            INIT_4E => X"000000a1000000a200000099000000a2000000bc000000be000000ad000000ae",
            INIT_4F => X"0000008a000000700000003e000000420000004a0000004b0000009500000099",
            INIT_50 => X"000000670000003c00000047000000590000004e000000590000006a00000077",
            INIT_51 => X"000000be000000ae000000b50000007f00000042000000720000005f0000004b",
            INIT_52 => X"000000a5000000ab000000a0000000a4000000c1000000b8000000ab000000ba",
            INIT_53 => X"00000073000000700000005e0000004d0000005c000000680000008b00000092",
            INIT_54 => X"0000005f000000480000004c0000006a000000670000003a0000005e0000007e",
            INIT_55 => X"000000bc000000c4000000a10000005b0000006300000078000000410000005e",
            INIT_56 => X"000000a10000009a000000a0000000aa000000a7000000a7000000c1000000b6",
            INIT_57 => X"000000640000006d0000008800000069000000510000006e0000008a00000091",
            INIT_58 => X"00000054000000450000005e000000710000006800000046000000520000006f",
            INIT_59 => X"000000c8000000ba0000009b0000007f0000007d000000550000006d00000074",
            INIT_5A => X"000000a6000000a4000000a2000000940000009d000000b1000000bb000000bb",
            INIT_5B => X"00000061000000610000007300000078000000610000007900000095000000a2",
            INIT_5C => X"0000004c000000550000007b00000097000000b40000008c0000005c00000065",
            INIT_5D => X"000000c8000000ad000000af00000092000000540000005a0000007c00000067",
            INIT_5E => X"000000ad000000a3000000ac0000009f0000009f000000ad000000ad000000bc",
            INIT_5F => X"00000060000000640000005f0000007000000083000000830000008b000000a4",
            INIT_60 => X"0000006c0000007f0000009d000000c2000000d1000000c00000009000000077",
            INIT_61 => X"000000c5000000b0000000af0000007c0000006f0000006a0000005e0000006a",
            INIT_62 => X"000000a3000000af000000c50000009c000000a5000000b0000000aa000000b8",
            INIT_63 => X"000000660000006b0000006000000064000000650000007a0000008300000093",
            INIT_64 => X"00000088000000a0000000c4000000c5000000a90000008a000000740000006e",
            INIT_65 => X"000000a9000000b40000009f000000920000008a0000005c0000006300000081",
            INIT_66 => X"00000097000000b3000000bc000000a6000000b2000000af0000008d0000008e",
            INIT_67 => X"0000004900000066000000650000005b0000003a000000700000009a0000008f",
            INIT_68 => X"000000a3000000bf000000b9000000a50000006b0000004a000000570000005b",
            INIT_69 => X"00000074000000920000008400000076000000660000006a0000008000000086",
            INIT_6A => X"000000a7000000ad0000009f000000b7000000b6000000a1000000630000004d",
            INIT_6B => X"0000004d000000440000005c0000005b0000002b0000005e000000870000009c",
            INIT_6C => X"000000bb000000a6000000940000005f0000002c000000320000005f00000051",
            INIT_6D => X"0000006b000000770000007200000068000000720000007e00000090000000ae",
            INIT_6E => X"00000096000000a9000000b2000000a9000000b60000009d0000005200000051",
            INIT_6F => X"000000560000005000000045000000610000003f0000002c0000006c00000098",
            INIT_70 => X"000000b0000000920000006d0000001c00000015000000340000005f0000005a",
            INIT_71 => X"000000820000007200000077000000780000007f0000008e000000b5000000ca",
            INIT_72 => X"00000098000000b4000000ad0000009f000000a9000000900000007600000081",
            INIT_73 => X"0000006a000000a70000007200000033000000550000002c0000004400000077",
            INIT_74 => X"0000009c00000077000000310000001800000034000000390000005b0000005f",
            INIT_75 => X"0000007500000074000000850000008d0000009b000000ba000000cb000000bb",
            INIT_76 => X"0000007d0000009c000000a70000009f000000990000008b000000770000006d",
            INIT_77 => X"0000007a000000aa000000900000003700000040000000440000004100000065",
            INIT_78 => X"0000007300000036000000210000002e00000049000000200000004b0000005e",
            INIT_79 => X"00000092000000880000009b000000b1000000c2000000c3000000b000000096",
            INIT_7A => X"00000069000000600000005f00000065000000770000005e000000650000008b",
            INIT_7B => X"0000006a0000009a0000008f000000800000006d0000006b0000007600000083",
            INIT_7C => X"0000003b0000001b00000028000000410000004c00000018000000230000004e",
            INIT_7D => X"000000ba000000a5000000b7000000c0000000b0000000960000008800000078",
            INIT_7E => X"0000008c000000700000005500000042000000560000006b000000aa000000cf",
            INIT_7F => X"000000800000009a0000008f00000096000000890000008900000095000000a9",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY12;


    MEM_IFMAP_LAYER0_ENTITY13 : if BRAM_NAME = "ifmap_layer0_entity13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000500000004b00000039000000210000002e000000400000005100000044",
            INIT_01 => X"00000042000000460000004b0000004700000022000000140000004600000053",
            INIT_02 => X"00000052000000540000006c0000007e000000790000007c0000007800000057",
            INIT_03 => X"000000570000004c00000043000000600000005b0000003b0000008100000088",
            INIT_04 => X"00000054000000540000005c000000380000002f0000004a0000006600000050",
            INIT_05 => X"000000490000004d0000005c0000005d00000030000000120000003e00000058",
            INIT_06 => X"000000530000004d0000006c000000750000006a0000006f000000750000006b",
            INIT_07 => X"000000510000005a0000004200000047000000410000002d0000008b00000097",
            INIT_08 => X"0000005a00000056000000690000005400000038000000580000006d0000005f",
            INIT_09 => X"0000003c0000004200000058000000590000003c00000014000000350000005c",
            INIT_0A => X"00000056000000420000007200000072000000540000004e0000006600000067",
            INIT_0B => X"0000003b00000062000000620000005400000037000000230000008f0000009e",
            INIT_0C => X"0000006000000058000000660000006d00000049000000640000006400000074",
            INIT_0D => X"00000037000000360000004300000041000000380000001a0000002d0000005e",
            INIT_0E => X"0000005b0000004500000072000000760000006200000061000000750000006a",
            INIT_0F => X"000000320000005e0000007e000000780000005d0000004000000096000000a0",
            INIT_10 => X"0000005e0000005a0000005e000000720000005d000000800000006800000078",
            INIT_11 => X"0000005600000049000000370000002f000000240000001a000000270000005d",
            INIT_12 => X"000000670000004a0000006d00000067000000650000006b0000007100000069",
            INIT_13 => X"0000006c0000006700000084000000810000007400000070000000ac000000a2",
            INIT_14 => X"0000004e0000005b000000590000005f00000062000000620000006600000069",
            INIT_15 => X"0000006c0000006a0000005d0000004d0000002b0000001b0000002300000058",
            INIT_16 => X"00000066000000620000006e000000390000004e000000640000006500000067",
            INIT_17 => X"000000780000008400000090000000810000007f00000082000000ba000000a7",
            INIT_18 => X"0000003f0000005d000000640000005a0000004f00000030000000600000005e",
            INIT_19 => X"0000006300000082000000810000007e0000005a000000260000001d0000004a",
            INIT_1A => X"0000006a000000710000007b000000250000003900000073000000470000003a",
            INIT_1B => X"0000003b00000065000000a0000000890000008c0000008d000000c1000000b7",
            INIT_1C => X"000000470000005e0000006100000067000000690000002f0000005400000056",
            INIT_1D => X"00000029000000720000008c0000008a0000008b000000490000001400000038",
            INIT_1E => X"0000008c000000780000007d0000003b0000004f00000073000000410000001a",
            INIT_1F => X"000000180000003f0000009b000000900000009400000096000000c3000000b0",
            INIT_20 => X"0000005c0000005000000072000000950000008c0000004a0000004e00000062",
            INIT_21 => X"000000170000003f000000860000008800000090000000710000002c00000047",
            INIT_22 => X"000000a50000009b0000008b00000070000000560000005e0000007c00000045",
            INIT_23 => X"00000016000000290000008e000000920000009600000096000000b1000000aa",
            INIT_24 => X"00000045000000540000009b000000a3000000940000004e0000005100000074",
            INIT_25 => X"00000038000000210000005d0000008a0000008e000000890000005a00000051",
            INIT_26 => X"000000810000009c0000009c0000009700000080000000730000008f0000007c",
            INIT_27 => X"000000180000001600000079000000940000009a00000098000000ad000000a7",
            INIT_28 => X"000000410000007f000000a6000000a500000091000000490000004f00000078",
            INIT_29 => X"0000006c000000470000005d0000007e0000007f0000008e0000007200000036",
            INIT_2A => X"0000005700000075000000a50000009c000000a1000000920000008500000087",
            INIT_2B => X"000000170000001300000074000000910000009c00000097000000af000000a9",
            INIT_2C => X"0000005f000000a5000000a8000000a10000008a00000042000000450000007b",
            INIT_2D => X"000000a200000088000000660000006d000000700000008a0000008c0000004b",
            INIT_2E => X"0000008800000076000000850000007c00000087000000970000009a00000099",
            INIT_2F => X"0000000b0000001400000077000000940000009d00000092000000aa000000bd",
            INIT_30 => X"00000098000000ad000000a400000087000000790000003c000000390000006a",
            INIT_31 => X"0000008b000000660000005c00000073000000760000007f0000009300000090",
            INIT_32 => X"00000088000000770000006b0000007800000074000000850000008a0000008d",
            INIT_33 => X"0000002b0000001a00000072000000a10000009100000087000000ae000000b0",
            INIT_34 => X"000000ab000000ac0000008c0000007f000000740000004e0000005500000074",
            INIT_35 => X"0000006e00000071000000760000007700000078000000820000007c00000099",
            INIT_36 => X"00000075000000810000007a000000830000007d000000770000006c00000069",
            INIT_37 => X"0000005f0000004100000070000000a60000009a0000008d000000a200000090",
            INIT_38 => X"000000a8000000a5000000720000008200000078000000630000006000000084",
            INIT_39 => X"000000840000008e000000810000007c00000070000000680000006b0000008b",
            INIT_3A => X"000000900000008d00000076000000730000006f0000006b000000770000007a",
            INIT_3B => X"0000005e00000048000000700000009d0000009f000000920000007b0000008e",
            INIT_3C => X"000000a6000000970000007c0000007f000000760000005d0000005a00000079",
            INIT_3D => X"0000008b0000007b0000007c0000006b0000004500000079000000ab00000099",
            INIT_3E => X"000000a700000083000000670000007a0000007700000080000000900000009b",
            INIT_3F => X"00000068000000220000004b00000095000000a0000000800000008c0000009f",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a300000095000000980000008d0000007e000000640000006400000070",
            INIT_41 => X"0000008d0000008b000000850000006400000047000000a6000000a30000008a",
            INIT_42 => X"0000007e0000007d00000097000000a30000009e000000a00000008800000081",
            INIT_43 => X"0000008b000000330000003d0000008f0000008f0000007a000000b1000000a9",
            INIT_44 => X"00000089000000900000007c0000009300000081000000830000007000000070",
            INIT_45 => X"00000093000000920000007f0000007a00000099000000a8000000790000008f",
            INIT_46 => X"00000086000000990000008f000000860000008a000000840000008b0000008d",
            INIT_47 => X"0000006f0000003a00000064000000860000007a000000920000008200000091",
            INIT_48 => X"000000760000007b000000610000008d0000008e000000950000007600000079",
            INIT_49 => X"00000082000000880000006e00000091000000bb000000790000007e0000008f",
            INIT_4A => X"000000910000009600000086000000970000009a00000094000000a10000009a",
            INIT_4B => X"0000008600000061000000770000006700000057000000610000007b00000086",
            INIT_4C => X"0000007d0000005d000000650000007a0000006f000000970000008700000088",
            INIT_4D => X"000000a00000009200000088000000a90000007d000000600000009900000086",
            INIT_4E => X"0000009100000090000000800000008d000000a7000000a60000009400000096",
            INIT_4F => X"000000a90000009500000057000000530000005e0000004b0000008200000084",
            INIT_50 => X"000000820000005400000068000000790000005e000000700000008c00000094",
            INIT_51 => X"000000aa0000009b000000a3000000760000004a0000008d0000007400000066",
            INIT_52 => X"00000091000000930000008900000092000000a70000009d00000095000000a5",
            INIT_53 => X"000000a10000009c0000007700000060000000710000006d0000007c0000007f",
            INIT_54 => X"000000790000006300000065000000810000007d000000480000007700000098",
            INIT_55 => X"000000a9000000b5000000960000005d0000007d0000009a0000005b00000078",
            INIT_56 => X"0000008b00000081000000870000008f0000008f00000091000000ad000000a2",
            INIT_57 => X"000000990000009a000000ab000000810000006600000075000000780000007d",
            INIT_58 => X"000000730000006200000076000000880000007b000000520000006800000088",
            INIT_59 => X"000000b3000000ad000000950000008100000094000000750000008d00000096",
            INIT_5A => X"0000008d0000008c0000008b0000007e0000008f0000009f000000a8000000a5",
            INIT_5B => X"0000009500000096000000a4000000980000006d0000007a0000008500000088",
            INIT_5C => X"0000006f000000790000009e000000ac000000bf000000960000006f0000007d",
            INIT_5D => X"000000ac0000009a000000a10000009400000069000000730000009900000091",
            INIT_5E => X"0000008f0000008800000093000000890000008d0000009c0000009b000000a1",
            INIT_5F => X"000000950000009e000000950000009c000000860000007b0000008c00000089",
            INIT_60 => X"00000093000000aa000000bd000000d1000000dc000000c8000000a200000095",
            INIT_61 => X"000000a4000000960000009f0000008b000000880000007d0000007a00000091",
            INIT_62 => X"0000008800000093000000a9000000850000008e0000009f0000009b0000009b",
            INIT_63 => X"0000009c000000a00000008f0000009a000000720000006b0000007e0000007f",
            INIT_64 => X"000000b0000000bf000000d7000000d5000000be0000009d000000890000008b",
            INIT_65 => X"0000008f0000009a00000097000000ad000000a30000007500000084000000a9",
            INIT_66 => X"0000007c00000095000000a3000000910000009800000099000000810000007c",
            INIT_67 => X"000000780000009700000095000000910000004a000000600000008300000077",
            INIT_68 => X"000000c1000000d3000000cf000000bf00000086000000610000006f00000073",
            INIT_69 => X"00000068000000860000008f000000900000007f00000091000000ad000000b1",
            INIT_6A => X"0000008e000000940000008a000000a10000009b0000008b0000005c00000049",
            INIT_6B => X"0000006d0000006f00000091000000920000003c000000550000007500000083",
            INIT_6C => X"000000d5000000c3000000b2000000780000004000000041000000720000006a",
            INIT_6D => X"0000007d0000008d000000960000008e00000099000000ad000000b9000000ca",
            INIT_6E => X"0000007f00000095000000a1000000900000009a0000008e000000600000006c",
            INIT_6F => X"00000075000000760000006c0000009300000061000000310000006200000083",
            INIT_70 => X"000000c7000000b40000008700000029000000260000003e0000007000000074",
            INIT_71 => X"000000a10000009e000000a4000000ab000000b2000000b7000000cc000000d4",
            INIT_72 => X"0000007e0000009c00000099000000870000008d000000870000008b0000009d",
            INIT_73 => X"00000083000000c500000088000000540000007c0000003b0000004200000067",
            INIT_74 => X"000000bf0000009500000042000000250000004e0000004f0000007b0000007f",
            INIT_75 => X"0000009f000000a5000000b4000000b8000000c2000000d6000000db000000d0",
            INIT_76 => X"0000007200000087000000930000008a000000830000007b0000007d00000087",
            INIT_77 => X"0000008f000000c9000000ac0000004e0000005b000000550000004f0000006c",
            INIT_78 => X"000000970000004e00000030000000430000006b00000034000000680000007d",
            INIT_79 => X"000000b6000000b4000000c3000000cd000000da000000d9000000cb000000bd",
            INIT_7A => X"0000006f0000005900000059000000610000007a0000005e00000074000000a5",
            INIT_7B => X"00000081000000bc000000b50000009f00000086000000820000008a00000096",
            INIT_7C => X"0000004e000000290000003a0000006000000073000000280000003300000066",
            INIT_7D => X"000000ce000000c4000000d2000000da000000cf000000b9000000b5000000a0",
            INIT_7E => X"000000a0000000840000006600000056000000710000007c000000b4000000d6",
            INIT_7F => X"0000009c000000b9000000b3000000b4000000a7000000a7000000a7000000ba",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY13;


    MEM_IFMAP_LAYER0_ENTITY14 : if BRAM_NAME = "ifmap_layer0_entity14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000390000003700000024000000160000001e0000002e0000004000000032",
            INIT_01 => X"00000032000000310000002c0000002b000000120000000c000000360000003b",
            INIT_02 => X"00000039000000380000004e000000530000004d000000510000004d0000003a",
            INIT_03 => X"000000420000003500000029000000410000003a0000001f0000005d00000061",
            INIT_04 => X"0000003c0000003b0000003d000000230000001d00000039000000510000003a",
            INIT_05 => X"0000002f0000003b0000003e000000380000001b000000070000002f00000040",
            INIT_06 => X"0000003c00000033000000510000004e000000440000004a0000004a00000044",
            INIT_07 => X"00000042000000450000002c0000002d0000002700000015000000600000006f",
            INIT_08 => X"000000410000003c000000480000003500000023000000460000005700000048",
            INIT_09 => X"0000002100000030000000410000003400000023000000070000002600000045",
            INIT_0A => X"0000003e0000002d000000520000004d00000037000000320000004200000043",
            INIT_0B => X"000000330000004d0000004b0000003f00000026000000100000006300000074",
            INIT_0C => X"0000004a0000004100000048000000470000002f000000500000004c0000005e",
            INIT_0D => X"0000001e000000230000003400000028000000220000000c0000001e00000048",
            INIT_0E => X"000000430000002e0000004d000000510000004500000044000000570000004b",
            INIT_0F => X"0000002200000044000000600000005f000000490000002a0000006b00000077",
            INIT_10 => X"0000004c00000048000000440000004b0000003c0000006a0000004f00000061",
            INIT_11 => X"0000003b00000033000000250000001c000000110000000c0000001800000049",
            INIT_12 => X"0000004d0000002d0000004900000047000000470000004b0000004f00000048",
            INIT_13 => X"0000005000000049000000610000005e00000055000000520000008100000080",
            INIT_14 => X"0000003d0000004d000000450000003d000000430000004b0000004d00000052",
            INIT_15 => X"00000049000000470000003b0000002c000000160000000d0000001300000043",
            INIT_16 => X"0000004d0000003e000000490000002200000035000000490000004800000048",
            INIT_17 => X"0000005c000000680000006e0000005c0000005b000000600000009300000088",
            INIT_18 => X"000000320000004f0000004f0000003e00000033000000190000004600000048",
            INIT_19 => X"0000003e0000004d0000004b0000004900000036000000180000000f00000038",
            INIT_1A => X"0000004a0000004800000058000000160000002a000000600000003300000022",
            INIT_1B => X"0000002b00000051000000830000006b0000006c00000068000000a100000095",
            INIT_1C => X"0000003a0000004b000000480000004d00000046000000150000003b0000003f",
            INIT_1D => X"000000120000003e0000004b0000004b000000510000002f0000000800000029",
            INIT_1E => X"00000053000000480000005e0000002a00000040000000590000002700000006",
            INIT_1F => X"000000150000003400000085000000760000007800000072000000a200000083",
            INIT_20 => X"0000004600000039000000580000007900000068000000310000003500000049",
            INIT_21 => X"00000007000000220000004f0000004e00000053000000470000001700000033",
            INIT_22 => X"0000005d0000005b00000063000000500000003e0000003c0000005100000028",
            INIT_23 => X"00000014000000210000007c0000007900000079000000780000008d00000073",
            INIT_24 => X"00000033000000400000007f0000008300000076000000380000003a00000056",
            INIT_25 => X"0000001c0000000d0000003a0000005e0000006300000061000000400000003b",
            INIT_26 => X"0000004a0000005f000000690000006200000050000000490000005d00000053",
            INIT_27 => X"000000170000000d000000650000007f0000007e000000770000008400000074",
            INIT_28 => X"0000003000000067000000870000008400000074000000350000003b0000005b",
            INIT_29 => X"00000049000000320000004a0000006600000061000000600000004b00000020",
            INIT_2A => X"00000031000000470000006c000000620000006100000059000000520000005a",
            INIT_2B => X"000000140000000a0000005b0000007b0000008a000000770000007c00000077",
            INIT_2C => X"000000480000008700000087000000810000006e0000002f0000003300000065",
            INIT_2D => X"0000008700000075000000560000005e0000004f00000052000000540000002e",
            INIT_2E => X"000000580000004a000000580000005c0000005e0000005d0000006600000078",
            INIT_2F => X"000000070000000b0000005b000000770000008d000000760000007300000084",
            INIT_30 => X"000000770000008b000000830000006b00000060000000280000002800000058",
            INIT_31 => X"0000006c000000510000004a0000005f0000005900000057000000660000006b",
            INIT_32 => X"0000005f0000005700000055000000660000005d000000640000006e00000076",
            INIT_33 => X"000000200000000f000000590000007b0000007100000065000000780000007c",
            INIT_34 => X"000000890000008b0000006e000000640000005c000000370000003f0000005f",
            INIT_35 => X"0000005600000056000000580000005a0000005c00000065000000610000007b",
            INIT_36 => X"0000005f0000006e0000006c000000720000006c000000640000005800000055",
            INIT_37 => X"0000004c000000310000005800000080000000730000006b000000750000006d",
            INIT_38 => X"000000870000008600000056000000680000006000000047000000450000006a",
            INIT_39 => X"0000006a0000006e000000600000006000000058000000510000005700000074",
            INIT_3A => X"000000800000007f0000006b000000610000005c000000570000005f00000062",
            INIT_3B => X"00000046000000350000005c0000007a00000077000000740000005e0000007a",
            INIT_3C => X"00000085000000790000005f000000670000005c000000400000004000000060",
            INIT_3D => X"0000007100000062000000650000005800000033000000640000009600000081",
            INIT_3E => X"000000980000007100000053000000600000005f000000650000007700000083",
            INIT_3F => X"000000480000000d00000039000000760000007c000000620000007800000094",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000082000000780000007c000000730000005a000000470000004c00000057",
            INIT_41 => X"000000780000007700000074000000540000003a000000960000008e0000006e",
            INIT_42 => X"0000006e000000670000007e000000890000008600000085000000710000006c",
            INIT_43 => X"0000006b000000210000002a000000750000007200000063000000a30000009f",
            INIT_44 => X"000000690000007500000063000000750000005d000000640000005800000056",
            INIT_45 => X"00000081000000810000006f0000006b0000008b0000009b000000660000006e",
            INIT_46 => X"000000710000007c0000007600000071000000760000006d000000770000007c",
            INIT_47 => X"0000005700000027000000480000006900000063000000830000007500000083",
            INIT_48 => X"0000005600000063000000470000006d0000007300000078000000600000005f",
            INIT_49 => X"000000750000007b0000005e00000082000000b00000006a000000630000006c",
            INIT_4A => X"00000079000000780000006f0000008300000088000000810000008d00000089",
            INIT_4B => X"0000006e00000043000000510000004800000043000000500000006b00000075",
            INIT_4C => X"0000005e000000470000004800000058000000570000007d000000700000006d",
            INIT_4D => X"0000009400000087000000760000009800000073000000490000007900000064",
            INIT_4E => X"0000007a00000079000000710000007d00000095000000940000008200000085",
            INIT_4F => X"0000008a00000073000000380000003d0000004e0000003a0000007100000072",
            INIT_50 => X"000000660000003c000000480000005800000043000000590000007400000077",
            INIT_51 => X"0000009c0000008d0000009200000065000000370000006d0000005700000048",
            INIT_52 => X"0000007c0000007f0000007b00000086000000980000008c0000008800000098",
            INIT_53 => X"000000770000007a000000620000004d000000620000005d000000690000006d",
            INIT_54 => X"000000600000004b00000046000000600000005d00000032000000610000007e",
            INIT_55 => X"00000097000000a2000000830000004900000061000000760000003b0000005a",
            INIT_56 => X"000000750000006e000000760000007d0000007f00000084000000a300000096",
            INIT_57 => X"0000006a000000700000008e0000006b0000004f0000005e0000006600000069",
            INIT_58 => X"00000059000000450000004e0000005c00000059000000370000005100000070",
            INIT_59 => X"0000009c000000970000007d0000006b00000076000000530000006b00000077",
            INIT_5A => X"00000075000000780000007b0000006c0000007e000000940000009b00000094",
            INIT_5B => X"0000006900000063000000790000008100000056000000540000006600000072",
            INIT_5C => X"0000004e000000450000005f000000770000009a000000780000005600000062",
            INIT_5D => X"00000096000000840000008b0000007d0000004e000000570000007e00000073",
            INIT_5E => X"0000007b0000007600000084000000790000007e000000920000008e0000008d",
            INIT_5F => X"000000670000006a00000065000000790000006f000000520000005800000073",
            INIT_60 => X"0000005c00000060000000770000009f000000b6000000a70000008800000074",
            INIT_61 => X"0000008f0000008300000088000000700000006f000000660000005a00000066",
            INIT_62 => X"00000077000000840000009c0000007500000080000000960000008e00000086",
            INIT_63 => X"0000006c00000071000000600000006a000000530000004e0000005900000066",
            INIT_64 => X"000000690000007b0000009e000000a600000092000000710000006d0000006c",
            INIT_65 => X"0000007b000000860000007e000000910000008c000000550000005200000066",
            INIT_66 => X"0000006a0000008a0000009600000083000000890000008a0000007300000068",
            INIT_67 => X"0000004b0000006900000065000000600000002d0000004a0000006f00000061",
            INIT_68 => X"0000007e00000097000000970000008b00000056000000370000005500000058",
            INIT_69 => X"000000520000006e0000006e0000006f00000057000000570000006800000068",
            INIT_6A => X"0000007a0000008100000078000000910000008c000000790000004b00000035",
            INIT_6B => X"00000040000000410000006200000061000000200000003e0000006200000074",
            INIT_6C => X"0000009c00000086000000750000004b00000020000000220000005c00000052",
            INIT_6D => X"0000005f0000005b0000005a0000005200000057000000620000006d0000008d",
            INIT_6E => X"0000006b000000800000008f000000810000008b000000790000004600000052",
            INIT_6F => X"000000420000004700000047000000630000003f0000001d0000004e00000071",
            INIT_70 => X"00000094000000720000004e0000000f0000000d00000023000000560000005a",
            INIT_71 => X"00000071000000560000005b00000061000000620000006f0000008b000000a2",
            INIT_72 => X"0000006a0000008700000087000000760000007e000000730000006a00000078",
            INIT_73 => X"0000005300000099000000600000002c0000005b000000260000002a0000004f",
            INIT_74 => X"0000007a000000570000001f0000000d000000250000002d000000560000005c",
            INIT_75 => X"0000005c0000005d00000072000000750000007a0000009e000000ad00000096",
            INIT_76 => X"0000005b00000073000000850000007e0000007100000067000000550000004d",
            INIT_77 => X"00000062000000860000006c0000002a0000003c0000003b000000320000004e",
            INIT_78 => X"0000005400000023000000170000002400000038000000180000004700000052",
            INIT_79 => X"000000790000006f0000008200000096000000a5000000a50000009200000076",
            INIT_7A => X"0000005600000046000000450000004e000000620000003f000000420000006c",
            INIT_7B => X"000000590000007b000000740000007800000062000000600000006c00000075",
            INIT_7C => X"000000250000000f0000001d0000003400000040000000110000001b00000041",
            INIT_7D => X"0000009c0000008800000098000000aa00000096000000740000006400000059",
            INIT_7E => X"0000007f00000066000000470000002f0000004a0000004500000079000000a6",
            INIT_7F => X"0000007500000092000000880000009300000082000000830000008b0000009c",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY14;


    MEM_IFMAP_LAYER0_ENTITY15 : if BRAM_NAME = "ifmap_layer0_entity15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000970000009c0000009d0000008d000000580000004d0000008b000000b3",
            INIT_01 => X"0000007600000079000000880000009700000097000000900000009e0000009c",
            INIT_02 => X"000000530000005e000000620000006200000054000000540000006c0000007e",
            INIT_03 => X"0000004d0000004c00000057000000750000006000000054000000560000005a",
            INIT_04 => X"000000a70000009e0000009f0000009f000000920000008000000085000000b8",
            INIT_05 => X"0000007d0000008800000096000000960000009a00000099000000a2000000a5",
            INIT_06 => X"000000580000005e000000620000005d000000520000005a0000006d00000081",
            INIT_07 => X"0000005a0000005b00000062000000760000006a0000005b0000004c0000004e",
            INIT_08 => X"000000a40000009b00000098000000a4000000aa000000b000000098000000b4",
            INIT_09 => X"0000008c00000092000000970000009c0000009f000000a2000000aa000000a2",
            INIT_0A => X"0000006b00000067000000620000005500000047000000580000007c00000092",
            INIT_0B => X"0000005f0000005d000000650000006f0000006f0000006f0000006d00000065",
            INIT_0C => X"000000a3000000a400000098000000a8000000b5000000b8000000ae000000af",
            INIT_0D => X"000000a40000009f000000a2000000ae000000a8000000a7000000b3000000a6",
            INIT_0E => X"0000006b000000630000005a000000480000003a000000590000008900000097",
            INIT_0F => X"0000006f0000006d0000006100000069000000790000007d0000008000000075",
            INIT_10 => X"000000af000000b0000000a1000000a2000000ac000000a7000000ae000000af",
            INIT_11 => X"000000a4000000a0000000a8000000b0000000b4000000b3000000b2000000b2",
            INIT_12 => X"0000005e000000630000005a0000004200000045000000780000009c000000ad",
            INIT_13 => X"000000740000007100000068000000700000007b0000007f0000007c00000069",
            INIT_14 => X"000000b3000000b0000000a6000000a9000000aa00000090000000ae000000b5",
            INIT_15 => X"000000960000009f000000ae000000b0000000b5000000b4000000b4000000b4",
            INIT_16 => X"00000070000000830000007d00000060000000740000009b000000af000000b5",
            INIT_17 => X"0000007c000000760000007800000079000000790000007a0000007800000075",
            INIT_18 => X"000000af000000b0000000ae000000af000000b20000008a0000009c000000c0",
            INIT_19 => X"00000099000000ad000000bb000000bb000000b8000000ba000000b4000000b8",
            INIT_1A => X"00000079000000940000009500000096000000a7000000ad000000ad000000a6",
            INIT_1B => X"000000800000007b0000007a000000780000006f0000006d0000007500000073",
            INIT_1C => X"000000b8000000af000000af000000ad000000ab0000009c0000007d000000b9",
            INIT_1D => X"000000a6000000b8000000b9000000bd000000c2000000c1000000b7000000bc",
            INIT_1E => X"0000007a0000008f00000089000000aa000000b0000000b1000000ac000000a4",
            INIT_1F => X"0000007d0000007b000000760000007500000067000000600000006e0000006b",
            INIT_20 => X"000000b4000000b2000000ad000000ac000000a00000009f000000950000009b",
            INIT_21 => X"000000a0000000ac000000af000000bb000000bf000000ba000000ba000000bb",
            INIT_22 => X"00000085000000a60000009b000000b7000000b0000000a6000000970000009a",
            INIT_23 => X"0000007d0000007a0000007a0000007600000077000000700000006800000068",
            INIT_24 => X"000000aa000000b7000000b2000000b2000000a900000093000000980000009a",
            INIT_25 => X"000000a9000000a5000000a7000000ae000000c1000000c6000000bc000000b0",
            INIT_26 => X"0000008d000000ab000000a0000000b3000000a9000000920000008c0000009d",
            INIT_27 => X"0000007d000000760000007b000000740000007700000075000000680000005f",
            INIT_28 => X"000000ba000000b8000000b8000000ae000000b10000009f0000007000000086",
            INIT_29 => X"000000bb000000a70000009e0000009b000000b0000000bf000000c2000000ba",
            INIT_2A => X"0000007c0000009b0000009c000000a0000000970000008600000093000000ae",
            INIT_2B => X"0000007f0000007b000000750000006b0000006600000069000000660000004a",
            INIT_2C => X"000000be000000bf000000b1000000930000009d000000ae0000005b00000041",
            INIT_2D => X"000000a300000094000000ae000000b8000000b0000000ac000000b0000000bc",
            INIT_2E => X"0000005000000083000000950000009800000095000000850000009a000000b0",
            INIT_2F => X"0000007d00000078000000710000006700000066000000670000006100000042",
            INIT_30 => X"000000b6000000bd000000ca000000bc000000b1000000bf0000005c00000015",
            INIT_31 => X"0000007200000098000000ae000000c8000000bc000000a50000009c000000b3",
            INIT_32 => X"0000004e00000072000000880000009700000089000000780000007f0000005f",
            INIT_33 => X"0000007600000075000000710000006200000062000000590000004900000040",
            INIT_34 => X"000000bb000000bc000000c3000000c8000000ad000000a8000000630000002c",
            INIT_35 => X"0000009a000000a8000000a8000000b9000000c2000000b400000095000000a5",
            INIT_36 => X"00000048000000640000007f0000009c0000008a00000091000000920000006b",
            INIT_37 => X"0000006f0000006c0000006a0000006200000060000000530000004000000039",
            INIT_38 => X"000000bb000000b4000000be000000c40000009f000000750000007600000069",
            INIT_39 => X"000000bc000000b4000000a5000000ab000000c1000000c6000000ad000000ad",
            INIT_3A => X"000000480000006900000080000000a0000000b3000000ad000000bb000000ae",
            INIT_3B => X"000000660000006100000064000000630000006c000000570000004500000043",
            INIT_3C => X"000000a8000000b4000000c4000000c60000009d00000068000000710000008a",
            INIT_3D => X"000000c8000000c4000000bf000000d2000000cd000000cb000000bf000000b4",
            INIT_3E => X"000000500000007100000099000000a8000000be000000bc000000bb000000c0",
            INIT_3F => X"000000620000005a0000005a0000007800000087000000600000004000000046",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000096000000b0000000bb000000be00000093000000730000008a00000096",
            INIT_41 => X"000000cb000000be000000c2000000d3000000c6000000d3000000c7000000ab",
            INIT_42 => X"0000004600000064000000a6000000be000000bd000000b8000000ba000000bf",
            INIT_43 => X"0000005e0000004a0000005c000000950000008f0000006a000000380000002f",
            INIT_44 => X"00000091000000bf000000c0000000bd000000a5000000920000009b0000009b",
            INIT_45 => X"000000a8000000b2000000c2000000c000000095000000a9000000d20000009c",
            INIT_46 => X"0000002b00000043000000750000009a000000a7000000aa000000b5000000a9",
            INIT_47 => X"000000500000003f0000006a0000009c0000008f000000680000003100000022",
            INIT_48 => X"00000089000000ba000000be000000c4000000a60000008a000000a2000000a5",
            INIT_49 => X"0000008f00000080000000b6000000d2000000a90000009d000000c900000074",
            INIT_4A => X"000000330000002f0000003800000052000000610000007f000000930000007c",
            INIT_4B => X"00000041000000390000007b0000009d0000009d00000069000000400000002b",
            INIT_4C => X"00000098000000be000000be000000be0000009e0000007800000096000000a9",
            INIT_4D => X"000000ce00000090000000a5000000c3000000b9000000bc000000990000003c",
            INIT_4E => X"000000500000004700000033000000370000003d0000006500000089000000b1",
            INIT_4F => X"00000032000000360000008e000000b0000000a00000006e0000004a00000037",
            INIT_50 => X"0000009a000000ba000000bc000000ba000000a600000096000000a0000000aa",
            INIT_51 => X"000000c00000008c0000008c0000009b000000920000007e0000003100000020",
            INIT_52 => X"000000570000005200000049000000490000003e000000610000009c000000cc",
            INIT_53 => X"0000003300000048000000a7000000bc000000a60000006b0000003e0000003a",
            INIT_54 => X"0000007c000000a3000000b2000000b50000009c00000097000000ab000000b2",
            INIT_55 => X"0000008200000065000000630000004e00000037000000280000001d00000024",
            INIT_56 => X"000000550000003c0000003300000034000000370000005f0000007b00000090",
            INIT_57 => X"0000003700000059000000b1000000bb00000099000000660000004d0000004e",
            INIT_58 => X"0000006900000095000000a7000000a90000009800000092000000ab000000b5",
            INIT_59 => X"000000780000005c000000470000002f0000002e000000420000005e0000004f",
            INIT_5A => X"000000370000001e00000022000000230000002900000038000000370000005a",
            INIT_5B => X"0000003c0000006a000000ae000000ad00000077000000610000005600000052",
            INIT_5C => X"0000008900000094000000a00000009c000000a30000009e0000009c000000b1",
            INIT_5D => X"000000670000007d0000006d0000006e0000006b00000066000000760000008f",
            INIT_5E => X"000000130000000e0000001c000000180000001300000010000000110000002f",
            INIT_5F => X"0000004300000085000000ad0000008c0000006300000060000000410000002b",
            INIT_60 => X"000000c0000000ab0000008c00000097000000b6000000a70000008b0000009e",
            INIT_61 => X"000000650000007f0000008d00000092000000880000008500000074000000ac",
            INIT_62 => X"0000000f0000000a000000110000001800000019000000200000002500000041",
            INIT_63 => X"000000690000009c00000094000000620000004e000000610000004200000014",
            INIT_64 => X"000000b100000094000000880000009e000000ab000000ae000000a4000000a0",
            INIT_65 => X"0000007d0000008e0000008b0000007f00000097000000a900000093000000b8",
            INIT_66 => X"0000001a0000001100000018000000210000002b0000003f0000004d00000067",
            INIT_67 => X"00000088000000780000005a0000004800000032000000480000003e0000001f",
            INIT_68 => X"000000780000008c000000a8000000b1000000a7000000a7000000a3000000a0",
            INIT_69 => X"00000091000000a60000009c0000007b00000082000000760000008f000000ab",
            INIT_6A => X"0000004300000038000000420000004c0000004e0000005b000000690000007c",
            INIT_6B => X"0000006a000000510000007b0000006400000049000000410000004100000046",
            INIT_6C => X"0000007b00000099000000aa000000b4000000930000008c0000009f0000009c",
            INIT_6D => X"000000a2000000a80000009e000000830000007e000000730000009c0000008b",
            INIT_6E => X"00000077000000690000006800000070000000780000007b000000770000007f",
            INIT_6F => X"000000680000005c000000860000007a0000006d000000680000006900000074",
            INIT_70 => X"0000008c0000008d0000009c000000ad0000008b0000007b0000009e000000a4",
            INIT_71 => X"000000a8000000a60000009d00000097000000a100000082000000790000008d",
            INIT_72 => X"000000940000008a0000008500000081000000840000008f0000008a00000090",
            INIT_73 => X"000000930000007300000064000000780000008400000086000000890000008f",
            INIT_74 => X"0000009e0000009e000000a1000000a7000000a800000090000000950000008e",
            INIT_75 => X"000000a20000009e000000a0000000a1000000a90000009700000090000000a5",
            INIT_76 => X"0000009e00000096000000950000008d0000007f000000890000009100000099",
            INIT_77 => X"0000009f0000008b000000770000007b0000008f00000094000000960000009f",
            INIT_78 => X"000000a8000000aa000000a7000000a7000000b9000000b3000000a600000098",
            INIT_79 => X"00000085000000890000009d000000a9000000b2000000ad000000a4000000a7",
            INIT_7A => X"0000009d00000098000000970000008c000000880000008c0000008f00000092",
            INIT_7B => X"0000009900000090000000830000008500000090000000990000009c000000a6",
            INIT_7C => X"0000009f000000910000007d0000008b000000ab000000b7000000b20000009f",
            INIT_7D => X"0000007300000083000000980000009e0000009c000000950000008b000000a2",
            INIT_7E => X"000000a10000009c0000009d000000900000008f000000940000008e00000084",
            INIT_7F => X"0000009800000099000000960000009c0000009c000000940000009f000000a7",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY15;


    MEM_IFMAP_LAYER0_ENTITY16 : if BRAM_NAME = "ifmap_layer0_entity16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000053000000540000005f000000600000003b000000310000006000000076",
            INIT_01 => X"0000004f0000004b000000520000005c0000005a00000053000000610000005f",
            INIT_02 => X"00000033000000380000003800000037000000320000003b000000500000005b",
            INIT_03 => X"0000002f0000002f000000350000004c0000003a00000033000000380000003c",
            INIT_04 => X"000000680000005d000000600000006c00000069000000590000005800000082",
            INIT_05 => X"000000480000004f00000057000000540000005b0000005a0000006200000065",
            INIT_06 => X"00000033000000370000003800000037000000320000003d0000004800000052",
            INIT_07 => X"000000390000003a0000003d0000004b0000004100000035000000280000002b",
            INIT_08 => X"0000006a0000005f000000590000006c0000007a000000810000006800000084",
            INIT_09 => X"0000004c0000004f00000050000000550000005e000000620000006900000062",
            INIT_0A => X"000000420000003f0000003a000000330000002a000000360000004c00000055",
            INIT_0B => X"00000039000000380000003e000000430000004200000043000000420000003c",
            INIT_0C => X"00000069000000680000005a0000007000000084000000880000007f00000081",
            INIT_0D => X"0000005d000000570000005a0000006700000066000000650000007100000065",
            INIT_0E => X"0000003e00000039000000330000002a0000001f000000330000004e0000004f",
            INIT_0F => X"0000004500000043000000370000003c0000004a0000004b0000004d00000046",
            INIT_10 => X"0000007200000072000000630000006d0000007f000000790000007f00000080",
            INIT_11 => X"0000005c00000059000000630000006c00000071000000700000006f0000006f",
            INIT_12 => X"0000002e0000003800000034000000270000002c0000004e000000590000005e",
            INIT_13 => X"00000047000000450000003b0000004200000049000000470000004300000035",
            INIT_14 => X"00000074000000710000006a000000760000007f000000680000008300000089",
            INIT_15 => X"000000540000005a000000690000006d00000071000000740000007500000073",
            INIT_16 => X"0000003d000000520000004d0000003a0000004f00000067000000680000006a",
            INIT_17 => X"0000004b00000046000000480000004900000046000000430000003f0000003e",
            INIT_18 => X"0000006f00000073000000750000007a00000087000000660000007700000098",
            INIT_19 => X"0000005c000000660000007100000073000000700000007c0000007b00000079",
            INIT_1A => X"000000430000005b000000570000005c0000006e0000006d0000006500000064",
            INIT_1B => X"0000004e0000004a00000048000000450000003b00000038000000400000003e",
            INIT_1C => X"000000790000007200000076000000780000007e000000780000005900000093",
            INIT_1D => X"000000640000006c0000006d00000073000000730000007c0000007a00000080",
            INIT_1E => X"00000048000000570000004b000000660000006a0000006d0000006800000065",
            INIT_1F => X"0000004b000000490000004400000042000000350000002e0000003c0000003b",
            INIT_20 => X"0000007700000075000000740000007700000072000000780000006f00000076",
            INIT_21 => X"0000005e0000006100000067000000730000006d0000006f0000007a00000080",
            INIT_22 => X"00000059000000720000005f0000006d0000006400000061000000590000005e",
            INIT_23 => X"0000004b00000048000000480000004600000047000000400000003a0000003e",
            INIT_24 => X"0000006f0000007b0000007a0000007c00000078000000690000007100000077",
            INIT_25 => X"0000006f000000650000006d00000076000000790000007d0000007b00000076",
            INIT_26 => X"000000670000007a000000640000006a00000060000000520000005500000069",
            INIT_27 => X"0000004b000000440000004b0000004700000049000000470000003e0000003d",
            INIT_28 => X"0000007e0000007c0000007f000000780000007e000000720000004800000064",
            INIT_29 => X"000000900000007800000077000000790000007b00000080000000810000007f",
            INIT_2A => X"0000005b0000006c000000610000005f000000580000004f0000006300000083",
            INIT_2B => X"0000004c0000004900000046000000400000003b0000003d0000003e0000002e",
            INIT_2C => X"00000083000000840000007a0000005d000000690000007f0000003400000022",
            INIT_2D => X"000000850000007400000097000000a60000008c000000780000007300000081",
            INIT_2E => X"00000031000000560000005c0000006000000061000000560000006e0000008d",
            INIT_2F => X"0000004a00000045000000420000003e0000003c0000003e0000003c0000002a",
            INIT_30 => X"000000840000008c0000009a0000008c0000007d0000008e0000004000000004",
            INIT_31 => X"000000530000007700000093000000b20000009c0000007b0000006b0000007f",
            INIT_32 => X"000000310000004d0000005c0000006f00000064000000530000005b00000040",
            INIT_33 => X"0000004400000042000000430000003b00000039000000370000002f00000029",
            INIT_34 => X"0000008d0000008f000000960000009c0000007b0000007a0000004800000018",
            INIT_35 => X"00000077000000800000008100000097000000a00000008f0000006a00000077",
            INIT_36 => X"0000002d000000440000005a0000007b0000006d00000073000000740000004d",
            INIT_37 => X"0000003e0000003a0000003e0000003b00000037000000330000002b00000023",
            INIT_38 => X"0000008f000000860000009100000096000000700000004a0000005200000045",
            INIT_39 => X"0000009700000085000000720000007d0000009c000000a10000008400000083",
            INIT_3A => X"0000002f0000004b0000005d000000810000009800000092000000a000000091",
            INIT_3B => X"00000039000000360000003c0000003c0000004400000038000000300000002f",
            INIT_3C => X"0000007d000000860000009600000098000000700000003b0000004100000057",
            INIT_3D => X"000000a00000008f000000840000009b000000a5000000a70000009b0000008f",
            INIT_3E => X"00000039000000540000007800000089000000a10000009f0000009e000000a2",
            INIT_3F => X"000000390000003600000037000000510000005f000000400000002b00000033",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006c000000810000008d0000009000000066000000400000004e00000058",
            INIT_41 => X"0000009f00000086000000860000009e0000009d000000af000000a50000008b",
            INIT_42 => X"0000003100000049000000870000009a0000009800000093000000940000009a",
            INIT_43 => X"000000390000002c0000003d0000006f000000670000004b000000230000001e",
            INIT_44 => X"0000006900000091000000930000008f00000074000000570000005700000056",
            INIT_45 => X"000000790000007a0000008b000000910000006c00000085000000b300000080",
            INIT_46 => X"000000180000002a0000005800000072000000790000007c000000870000007d",
            INIT_47 => X"0000002e00000027000000500000007500000066000000490000001d00000013",
            INIT_48 => X"0000006200000091000000990000009c000000760000004d0000005c0000005c",
            INIT_49 => X"000000620000004b00000083000000a50000007a00000074000000aa0000005c",
            INIT_4A => X"0000001b000000110000001b000000360000004000000055000000610000004c",
            INIT_4B => X"0000002800000024000000640000007f0000007500000045000000280000001a",
            INIT_4C => X"000000730000009b000000a30000009c0000006e0000003c000000540000005e",
            INIT_4D => X"0000009c00000057000000710000009500000089000000940000007c00000027",
            INIT_4E => X"0000002e000000220000001800000027000000270000003d0000005000000078",
            INIT_4F => X"00000020000000220000007b0000009900000078000000450000002d0000001f",
            INIT_50 => X"0000007500000098000000a20000009600000072000000590000005d00000061",
            INIT_51 => X"0000007c00000049000000560000007300000074000000640000001d0000000d",
            INIT_52 => X"000000320000003100000032000000310000001b0000002f0000005b00000086",
            INIT_53 => X"000000200000003800000096000000a20000007d000000420000001e00000019",
            INIT_54 => X"0000005700000081000000960000008d0000006300000057000000680000006a",
            INIT_55 => X"0000003e00000029000000390000003600000025000000160000000b0000000f",
            INIT_56 => X"000000330000002200000023000000200000001a000000360000004800000053",
            INIT_57 => X"0000001f0000004a0000009e0000009b000000700000003e0000002b00000028",
            INIT_58 => X"0000004200000073000000890000007b0000005a0000004f0000006800000070",
            INIT_59 => X"000000450000002c000000260000001b0000001700000028000000420000002f",
            INIT_5A => X"0000001f0000000f00000016000000190000001d000000260000001f00000036",
            INIT_5B => X"0000001f0000005700000094000000860000004e0000003a0000003300000031",
            INIT_5C => X"0000005e0000007300000081000000690000006000000059000000580000006d",
            INIT_5D => X"0000003c0000004b0000003e000000420000003c000000360000004700000061",
            INIT_5E => X"0000000c0000000b00000013000000110000000e000000090000000a0000001a",
            INIT_5F => X"0000002300000069000000880000005e0000003b0000003a0000001f00000017",
            INIT_60 => X"000000930000008900000068000000600000007000000060000000460000005b",
            INIT_61 => X"000000350000003f000000450000004a00000043000000450000003a00000075",
            INIT_62 => X"000000120000000d000000090000000c0000000d000000130000001900000029",
            INIT_63 => X"00000047000000790000006800000034000000270000003e000000240000000c",
            INIT_64 => X"0000008600000069000000560000006100000062000000620000005c0000005b",
            INIT_65 => X"000000490000004e0000004900000044000000610000007c0000006b0000008e",
            INIT_66 => X"000000140000000b0000000e000000160000001c000000260000002b0000003e",
            INIT_67 => X"0000006400000058000000380000002500000014000000300000002a00000014",
            INIT_68 => X"0000004c0000005b0000006f0000007100000062000000610000005e0000005b",
            INIT_69 => X"00000054000000630000005f0000004700000051000000500000006e00000084",
            INIT_6A => X"0000002b000000200000002b0000003500000033000000380000003d00000048",
            INIT_6B => X"00000042000000300000005a000000400000002800000025000000280000002e",
            INIT_6C => X"00000048000000620000006d0000007100000052000000500000006000000057",
            INIT_6D => X"00000058000000600000005e0000004a0000004600000045000000730000005c",
            INIT_6E => X"0000004b0000003d0000003c000000420000004a0000004c0000004700000045",
            INIT_6F => X"0000003a000000360000005e0000004c000000410000003f0000004000000049",
            INIT_70 => X"000000500000004e0000005a000000690000004c000000430000006100000060",
            INIT_71 => X"0000005a0000005d0000005c00000057000000620000004c0000004800000057",
            INIT_72 => X"000000570000004d00000048000000420000004600000055000000540000004f",
            INIT_73 => X"0000005e0000004600000035000000430000004f000000500000005200000053",
            INIT_74 => X"0000005b000000580000005b0000006100000065000000510000005400000049",
            INIT_75 => X"0000005a0000005d0000005d00000059000000630000005b0000005900000069",
            INIT_76 => X"0000005b0000005400000052000000490000003c000000490000005500000058",
            INIT_77 => X"000000640000005700000044000000430000005500000057000000560000005d",
            INIT_78 => X"0000005f000000600000005f00000060000000710000006a0000006000000053",
            INIT_79 => X"0000004a000000520000005a0000005b000000680000006d0000006900000066",
            INIT_7A => X"0000005c00000057000000550000004d0000004a0000004d0000004e00000052",
            INIT_7B => X"0000005a000000570000004d0000004e000000540000005a0000005900000064",
            INIT_7C => X"0000005c0000004d000000420000005200000068000000710000006b0000005c",
            INIT_7D => X"0000003d0000004d0000005b000000580000005a0000005b000000510000005f",
            INIT_7E => X"000000600000005b0000005c0000005300000052000000560000004d00000046",
            INIT_7F => X"000000570000005b0000005a0000005c0000005b000000570000005c00000065",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY16;


    MEM_IFMAP_LAYER0_ENTITY17 : if BRAM_NAME = "ifmap_layer0_entity17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000360000003a0000004300000041000000240000001a0000003d00000053",
            INIT_01 => X"000000340000002e000000350000003e0000003b00000034000000410000003f",
            INIT_02 => X"000000260000002d0000002f0000002f000000270000002b0000004100000047",
            INIT_03 => X"00000029000000290000002e00000045000000320000002a0000002d0000002f",
            INIT_04 => X"0000004d000000440000004300000046000000460000003a0000003500000061",
            INIT_05 => X"0000002e00000032000000390000003400000039000000380000004100000044",
            INIT_06 => X"000000280000002c0000002f0000002f000000260000002b000000340000003c",
            INIT_07 => X"00000031000000330000003500000043000000380000002b0000001e00000020",
            INIT_08 => X"0000004e000000440000003900000044000000510000005c0000004700000064",
            INIT_09 => X"000000300000003100000030000000340000003b0000003f0000004700000040",
            INIT_0A => X"0000003800000035000000300000002b0000001e00000021000000320000003b",
            INIT_0B => X"000000310000002f000000350000003900000038000000390000003800000033",
            INIT_0C => X"0000004800000049000000370000004900000059000000610000005f00000060",
            INIT_0D => X"0000003f00000036000000370000004300000042000000420000004e00000041",
            INIT_0E => X"000000350000002f0000002900000022000000120000001a0000002e0000002f",
            INIT_0F => X"0000003c0000003a0000002d000000300000003e00000040000000440000003d",
            INIT_10 => X"0000004b0000004c0000003f000000490000005700000054000000610000005c",
            INIT_11 => X"0000003b000000350000003b000000430000004b0000004b0000004a0000004a",
            INIT_12 => X"000000270000002e000000290000001f0000001e00000033000000340000003b",
            INIT_13 => X"0000003c0000003a00000030000000340000003d0000003d0000003b0000002e",
            INIT_14 => X"0000004c0000004c000000460000005100000059000000470000006600000065",
            INIT_15 => X"00000031000000350000004300000044000000470000004e000000510000004c",
            INIT_16 => X"00000032000000420000003e0000002b00000039000000480000004100000043",
            INIT_17 => X"000000410000003c0000003d0000003c0000003a000000380000003600000038",
            INIT_18 => X"0000004b00000051000000500000005300000063000000490000005900000078",
            INIT_19 => X"00000035000000430000004f0000004c00000042000000550000005700000051",
            INIT_1A => X"0000002f0000004100000040000000410000004d0000004a000000400000003c",
            INIT_1B => X"000000420000003f0000003d0000003a000000300000002d0000003600000035",
            INIT_1C => X"000000540000004f00000051000000510000005b0000005b0000003b00000075",
            INIT_1D => X"0000003f0000004a0000004c0000004d00000048000000560000005600000057",
            INIT_1E => X"0000002f000000380000002f00000047000000490000004c0000004900000042",
            INIT_1F => X"000000400000003e00000039000000370000002a00000023000000310000002c",
            INIT_20 => X"00000050000000500000004f00000053000000510000005b000000540000005c",
            INIT_21 => X"0000003d00000043000000480000005100000046000000490000005300000058",
            INIT_22 => X"0000003c0000004f000000400000004f00000046000000460000004100000043",
            INIT_23 => X"000000400000003d0000003d0000003a0000003b000000340000002d0000002c",
            INIT_24 => X"0000004700000053000000560000005b0000005a0000004c0000005800000061",
            INIT_25 => X"000000550000004d00000053000000580000005300000054000000520000004f",
            INIT_26 => X"0000004b00000059000000480000005000000046000000390000003e00000051",
            INIT_27 => X"00000040000000390000003f0000003a0000003c0000003a000000310000002b",
            INIT_28 => X"00000054000000520000005b0000005900000062000000560000003000000051",
            INIT_29 => X"0000007e00000067000000650000005e0000005000000050000000540000005b",
            INIT_2A => X"00000044000000510000004c0000004b0000004300000037000000490000006b",
            INIT_2B => X"000000410000003e0000003a000000330000002d0000002f0000003100000020",
            INIT_2C => X"0000005a0000005a00000056000000400000004d000000630000001f00000014",
            INIT_2D => X"0000007900000067000000880000008f0000005f00000045000000450000005f",
            INIT_2E => X"00000021000000420000004d00000052000000500000003f0000005200000076",
            INIT_2F => X"0000003f0000003b00000036000000300000002e000000300000003000000021",
            INIT_30 => X"00000062000000690000007a0000006e0000005c000000700000003200000000",
            INIT_31 => X"000000490000005f0000007d0000009d00000077000000540000004800000060",
            INIT_32 => X"0000002a000000410000004f0000006000000054000000410000004700000034",
            INIT_33 => X"0000003a00000039000000380000002d00000029000000290000002500000025",
            INIT_34 => X"0000006f00000070000000780000007d0000005c000000610000003c00000014",
            INIT_35 => X"0000006c00000062000000640000007f000000800000006e0000004c00000059",
            INIT_36 => X"000000290000003a0000004c0000006a0000005b000000620000006300000044",
            INIT_37 => X"0000003500000032000000340000002e00000026000000250000002300000021",
            INIT_38 => X"000000730000006a000000750000007b000000580000003a000000460000003b",
            INIT_39 => X"0000008900000066000000500000005f0000007d000000820000006700000066",
            INIT_3A => X"0000002a000000400000004e0000006f000000840000007e0000008c00000083",
            INIT_3B => X"000000310000002e000000320000002f000000320000002a000000280000002b",
            INIT_3C => X"000000620000006c0000007c0000007e0000005e000000320000003500000049",
            INIT_3D => X"0000008c00000071000000620000007b000000880000008a0000007d00000072",
            INIT_3E => X"000000330000004900000069000000750000008c0000008a000000890000008f",
            INIT_3F => X"000000320000002d0000002d000000430000004d00000032000000230000002f",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000053000000690000007500000077000000560000003a0000004100000048",
            INIT_41 => X"000000870000006d0000006b000000820000008200000093000000890000006e",
            INIT_42 => X"0000002a0000003d0000007700000087000000830000007e0000007f00000084",
            INIT_43 => X"00000033000000240000003300000061000000550000003c0000001b0000001a",
            INIT_44 => X"000000500000007a0000007c0000007800000066000000510000004800000047",
            INIT_45 => X"0000005c00000065000000790000007c000000540000006a0000009700000063",
            INIT_46 => X"000000110000001f000000480000005e00000065000000680000007300000063",
            INIT_47 => X"000000290000001f0000004600000068000000550000003a000000150000000e",
            INIT_48 => X"0000004b0000007d000000880000008600000064000000440000004e0000004f",
            INIT_49 => X"0000004800000037000000710000008e000000610000005b0000009300000047",
            INIT_4A => X"000000160000000d000000140000002a00000032000000450000004f00000035",
            INIT_4B => X"000000230000001e0000005b0000006f00000060000000370000002300000014",
            INIT_4C => X"0000005d0000008a000000990000008700000058000000320000004800000051",
            INIT_4D => X"0000008d000000470000005c0000007c000000710000007f0000006f0000001f",
            INIT_4E => X"0000002c00000024000000190000002400000021000000330000004100000067",
            INIT_4F => X"0000001a0000001e000000730000008900000060000000360000002b0000001a",
            INIT_50 => X"000000620000008600000096000000820000005f0000004f0000005200000053",
            INIT_51 => X"00000074000000420000004c000000650000006300000056000000170000000a",
            INIT_52 => X"0000002e0000002f0000002f0000002e00000017000000270000004e0000007a",
            INIT_53 => X"000000190000002f000000890000009200000067000000340000001b00000014",
            INIT_54 => X"000000460000006e000000870000007b000000530000004e0000005c0000005c",
            INIT_55 => X"0000003800000025000000340000002f0000001d00000010000000080000000c",
            INIT_56 => X"0000002c0000001d0000001c00000019000000120000002b0000003900000046",
            INIT_57 => X"000000180000003d0000008d0000008c0000005e000000310000002600000021",
            INIT_58 => X"0000003000000060000000760000006b0000004e000000460000005d00000061",
            INIT_59 => X"0000003b000000260000001f0000001300000013000000220000003a00000025",
            INIT_5A => X"000000180000000a0000001100000011000000120000001b0000001300000027",
            INIT_5B => X"0000001800000046000000800000007800000040000000300000002c0000002a",
            INIT_5C => X"0000004b0000005f0000006b0000005b00000058000000520000004d0000005e",
            INIT_5D => X"0000003300000043000000350000003a0000003900000030000000370000004a",
            INIT_5E => X"0000000600000007000000130000000e00000008000000030000000400000010",
            INIT_5F => X"0000001b0000005700000073000000510000002f000000300000001700000011",
            INIT_60 => X"0000007e00000075000000520000005300000069000000570000003b0000004b",
            INIT_61 => X"0000002e000000390000003d000000420000003e000000390000002200000055",
            INIT_62 => X"0000000e0000000c0000000e0000000f0000000d000000120000001700000024",
            INIT_63 => X"0000003e0000006800000055000000280000001e000000360000001c00000007",
            INIT_64 => X"0000007000000057000000450000005500000056000000510000004d0000004d",
            INIT_65 => X"0000003a00000045000000430000003b0000004f000000640000004f0000006f",
            INIT_66 => X"0000000e000000060000000c0000001100000015000000200000002600000033",
            INIT_67 => X"0000005a0000004c0000002e0000001f0000000f00000029000000220000000f",
            INIT_68 => X"000000390000004a00000060000000650000005500000052000000510000004f",
            INIT_69 => X"000000440000005a000000580000003d0000003e0000003a000000570000006d",
            INIT_6A => X"0000002300000018000000230000002c0000002a0000002f000000350000003b",
            INIT_6B => X"000000380000002700000052000000390000001f0000001b0000001d00000026",
            INIT_6C => X"00000039000000530000005f000000660000004a0000004a000000570000004c",
            INIT_6D => X"0000004d00000057000000540000003f0000003a00000037000000630000004d",
            INIT_6E => X"0000003f00000031000000310000003b00000044000000430000003c00000039",
            INIT_6F => X"0000002f0000002d000000540000003f0000003300000030000000310000003c",
            INIT_70 => X"00000044000000410000004e0000005e00000045000000400000005a00000055",
            INIT_71 => X"00000051000000530000004e0000004a0000005a000000420000003c0000004c",
            INIT_72 => X"000000480000003e000000390000003b000000400000004c0000004700000043",
            INIT_73 => X"000000530000003d00000029000000320000003e000000400000004200000044",
            INIT_74 => X"000000500000004e00000051000000570000005c000000490000004b0000003d",
            INIT_75 => X"000000500000004e0000004c0000004a00000059000000500000004c0000005d",
            INIT_76 => X"0000004b000000440000004200000040000000350000003e000000450000004a",
            INIT_77 => X"000000590000004e00000038000000320000004400000048000000480000004d",
            INIT_78 => X"00000055000000570000005500000056000000640000005a0000005100000046",
            INIT_79 => X"0000003c0000003f000000460000004a0000005a0000005d0000005700000056",
            INIT_7A => X"0000004c0000004700000046000000410000003e0000003e0000003c00000042",
            INIT_7B => X"0000004f0000004d000000410000003e000000470000004e0000004d00000055",
            INIT_7C => X"00000051000000460000003900000046000000590000005f0000005d0000004f",
            INIT_7D => X"0000002f0000003d0000004c0000004a00000047000000470000004000000053",
            INIT_7E => X"000000500000004b0000004c0000004500000046000000480000003f00000038",
            INIT_7F => X"000000490000004f0000004c0000004f0000004e000000490000004f00000056",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY17;


    MEM_IFMAP_LAYER0_ENTITY18 : if BRAM_NAME = "ifmap_layer0_entity18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000f6000000f9000000f6000000e6000000d9000000d1000000b9000000a0",
            INIT_01 => X"000000c7000000d8000000dd000000da000000dd000000e6000000f3000000f8",
            INIT_02 => X"0000008b0000007900000090000000a6000000b4000000b8000000bb000000bc",
            INIT_03 => X"0000005e0000005b000000650000005e0000004f00000066000000660000006a",
            INIT_04 => X"000000eb000000f3000000f5000000e8000000e6000000f2000000ef000000e1",
            INIT_05 => X"000000ba000000c8000000cb000000c9000000cd000000d8000000e6000000ed",
            INIT_06 => X"000000870000007a0000008d0000008e0000007f000000a1000000ab000000af",
            INIT_07 => X"00000064000000610000006b0000005f00000034000000250000005200000076",
            INIT_08 => X"000000d6000000df000000e2000000d9000000dc000000f1000000f9000000fc",
            INIT_09 => X"000000a7000000b3000000b6000000b3000000b8000000c3000000cf000000d5",
            INIT_0A => X"00000072000000800000008c000000800000008100000094000000980000009f",
            INIT_0B => X"0000006900000069000000730000006300000026000000040000002800000057",
            INIT_0C => X"000000c0000000c8000000cb000000d3000000d3000000de000000e1000000e9",
            INIT_0D => X"00000099000000a0000000a5000000a0000000a4000000ae000000b7000000bb",
            INIT_0E => X"000000690000007f0000007d0000007d0000008a0000008c0000008d00000091",
            INIT_0F => X"0000006d000000700000007800000070000000370000001a000000250000003b",
            INIT_10 => X"000000ab000000b3000000b4000000be000000c9000000cf000000c3000000cf",
            INIT_11 => X"0000008d00000093000000970000009100000092000000990000009f000000a3",
            INIT_12 => X"0000005a000000840000007a0000008100000087000000830000008800000087",
            INIT_13 => X"0000006d00000072000000780000007500000056000000300000003d0000003a",
            INIT_14 => X"000000970000009f0000009c00000099000000a2000000aa000000ab000000b6",
            INIT_15 => X"0000008a0000008a0000008d0000008b0000008a0000008c0000008d00000090",
            INIT_16 => X"0000004500000066000000890000008c0000008a000000860000008c00000087",
            INIT_17 => X"0000006e00000070000000800000008100000074000000430000003e0000004b",
            INIT_18 => X"000000850000008c00000086000000880000008600000088000000880000008d",
            INIT_19 => X"000000910000008e000000920000008f0000008d0000008b0000008900000087",
            INIT_1A => X"000000210000002f0000006b0000008e0000008f0000008a0000009100000091",
            INIT_1B => X"000000700000006f00000084000000840000007f0000006c0000004b00000048",
            INIT_1C => X"000000840000008a000000830000008800000081000000800000007d00000076",
            INIT_1D => X"000000990000009a0000009e0000009600000093000000900000008c00000088",
            INIT_1E => X"000000110000000d000000420000008000000094000000930000009500000092",
            INIT_1F => X"0000007000000072000000800000007b0000007a000000800000007500000050",
            INIT_20 => X"000000890000008f000000870000008b00000085000000840000007e00000073",
            INIT_21 => X"000000aa000000a30000009a000000940000009800000095000000910000008b",
            INIT_22 => X"0000001e0000000e0000002c00000073000000940000009d000000a20000009e",
            INIT_23 => X"0000006f000000740000007a000000770000007e000000880000008b00000069",
            INIT_24 => X"0000008d00000091000000880000008d00000088000000880000008000000076",
            INIT_25 => X"000000a7000000a20000009a0000009d000000a50000009a000000930000008d",
            INIT_26 => X"000000370000002e00000038000000630000008a00000091000000930000009b",
            INIT_27 => X"0000006e0000007500000074000000730000007e0000007a0000007c0000006d",
            INIT_28 => X"0000008c00000090000000880000008e000000890000008b000000840000007d",
            INIT_29 => X"00000098000000900000008b000000830000009900000096000000900000008b",
            INIT_2A => X"0000002a000000450000005c00000080000000d6000000d3000000ba000000a6",
            INIT_2B => X"0000006b000000710000006f0000007000000073000000630000005f00000055",
            INIT_2C => X"0000008a0000008e000000880000008d0000008a0000008e0000008900000085",
            INIT_2D => X"000000cb000000c9000000b60000008e00000084000000880000008f00000089",
            INIT_2E => X"0000002a00000092000000bd000000a2000000c0000000cf000000ce000000d2",
            INIT_2F => X"000000680000006c0000006a0000006d0000007200000067000000280000001b",
            INIT_30 => X"000000890000008a0000008c0000008f0000008b0000008f0000008b0000008c",
            INIT_31 => X"0000007300000089000000a0000000ab000000a4000000900000008500000087",
            INIT_32 => X"0000005f000000c9000000dc0000006f0000003b0000004b0000005d0000006a",
            INIT_33 => X"00000064000000690000006500000063000000740000003e000000070000000d",
            INIT_34 => X"000000870000008200000092000000920000008c0000008f0000008a00000090",
            INIT_35 => X"00000013000000310000005c0000005e0000006e0000008c0000009100000082",
            INIT_36 => X"0000009d000000d2000000d1000000780000001200000019000000320000001d",
            INIT_37 => X"0000005f00000063000000520000004500000044000000130000000600000026",
            INIT_38 => X"00000080000000790000008e000000900000008e000000920000008b00000091",
            INIT_39 => X"000000160000002e000000520000005600000044000000540000007f00000085",
            INIT_3A => X"000000cb000000cd000000c9000000af000000410000001e0000003200000013",
            INIT_3B => X"000000580000004f000000380000002300000016000000120000001000000066",
            INIT_3C => X"000000830000008b000000840000008a00000090000000940000008b0000008f",
            INIT_3D => X"00000022000000280000004e0000006a00000056000000480000004200000075",
            INIT_3E => X"000000c3000000cd000000c5000000cb000000b6000000730000004600000024",
            INIT_3F => X"00000053000000640000004f0000001800000012000000250000003d0000006c",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007900000084000000720000008500000090000000930000008b0000008e",
            INIT_41 => X"0000009b000000530000004400000055000000450000003c0000005900000051",
            INIT_42 => X"00000072000000d3000000d7000000d7000000eb000000ed000000db000000c0",
            INIT_43 => X"000000540000008f0000008b0000004100000014000000350000005d00000030",
            INIT_44 => X"000000430000003a0000004500000074000000890000008e0000008d0000008f",
            INIT_45 => X"000000f20000008c00000019000000240000001c0000001d0000004b00000051",
            INIT_46 => X"0000003a00000095000000df000000db000000dc000000e3000000eb000000ec",
            INIT_47 => X"0000005b000000a7000000a1000000850000004e0000004e0000005400000039",
            INIT_48 => X"000000340000002d000000470000008d00000086000000880000008c0000008f",
            INIT_49 => X"000000d90000009b000000290000002f00000016000000170000002100000043",
            INIT_4A => X"00000067000000ad000000df000000dc000000d0000000bf000000be000000c7",
            INIT_4B => X"00000059000000a500000094000000980000009500000087000000730000005d",
            INIT_4C => X"0000002b000000210000004c000000bd000000b50000007e0000008c0000008f",
            INIT_4D => X"000000c20000009e000000420000003900000017000000100000001500000039",
            INIT_4E => X"000000b3000000de000000ce000000c2000000c9000000c4000000b3000000b6",
            INIT_4F => X"0000004200000088000000920000009600000097000000950000009c00000097",
            INIT_50 => X"0000002a000000260000005a000000b5000000ea0000009a000000850000008c",
            INIT_51 => X"000000ba000000a000000031000000140000000b0000000b0000000b00000034",
            INIT_52 => X"000000c4000000a10000005a0000004500000073000000b9000000b9000000b0",
            INIT_53 => X"000000260000004d000000880000009300000099000000a0000000aa000000b7",
            INIT_54 => X"0000002e0000002d0000006a0000008b000000a3000000a30000008000000082",
            INIT_55 => X"000000b4000000a2000000360000001e0000000f00000009000000030000001c",
            INIT_56 => X"000000950000003000000015000000140000001500000071000000be000000ac",
            INIT_57 => X"00000027000000150000004300000080000000850000008e000000ab000000bb",
            INIT_58 => X"00000030000000340000006c000000480000001a00000067000000840000007c",
            INIT_59 => X"000000b0000000a5000000630000005a0000003b0000000b0000000700000012",
            INIT_5A => X"000000460000000e000000260000002f0000001d0000002a000000a9000000b1",
            INIT_5B => X"00000030000000150000000e0000003c00000075000000750000008800000095",
            INIT_5C => X"0000001f00000044000000720000003b0000001e000000490000007c00000079",
            INIT_5D => X"000000bb000000bb0000006c0000004f00000048000000180000000e0000000d",
            INIT_5E => X"0000001b0000001c0000001b0000001e0000002b0000001b0000008b000000bf",
            INIT_5F => X"0000003b0000002a0000001500000016000000590000007b000000840000006c",
            INIT_60 => X"0000001c0000004d000000710000003c0000003f00000047000000660000006d",
            INIT_61 => X"000000b3000000bd000000880000004600000047000000300000001f00000010",
            INIT_62 => X"0000000e0000001b0000002900000035000000360000001f00000074000000b4",
            INIT_63 => X"0000003b0000003200000022000000120000003c0000007c0000008500000048",
            INIT_64 => X"000000150000004b000000690000003a0000003c0000003d0000005100000057",
            INIT_65 => X"000000a3000000a40000009100000061000000600000004c0000002e00000014",
            INIT_66 => X"00000011000000250000003100000047000000390000002000000071000000aa",
            INIT_67 => X"00000032000000280000001d0000000c00000021000000600000006c00000029",
            INIT_68 => X"0000002f000000570000005f000000390000003c000000400000004900000049",
            INIT_69 => X"000000b6000000b7000000b0000000a9000000a500000089000000620000003d",
            INIT_6A => X"0000001b000000330000005c0000006000000036000000220000007c000000b6",
            INIT_6B => X"000000280000001d00000012000000060000000c0000003b0000004600000011",
            INIT_6C => X"0000002f0000004500000059000000410000004e000000450000004900000049",
            INIT_6D => X"0000006000000062000000600000005b000000560000004a0000003c00000034",
            INIT_6E => X"000000140000001d0000003e0000003b0000003c000000200000005300000062",
            INIT_6F => X"00000021000000110000000a00000007000000030000000a0000001100000004",
            INIT_70 => X"000000040000000f000000270000002d0000003600000048000000530000004b",
            INIT_71 => X"0000000b0000000a000000080000000700000007000000050000000200000003",
            INIT_72 => X"0000000f000000380000002f0000004300000042000000080000000d0000000b",
            INIT_73 => X"000000200000000f0000000a0000000600000003000000010000000200000002",
            INIT_74 => X"00000019000000100000000a000000150000002f000000510000005900000050",
            INIT_75 => X"0000000c0000000e0000000e0000000e0000000e0000000e0000000a0000000e",
            INIT_76 => X"000000070000002a000000480000003e0000001700000006000000090000000a",
            INIT_77 => X"00000021000000150000000b0000000700000005000000050000000400000003",
            INIT_78 => X"0000003a0000003b0000002f0000002e00000037000000490000004f00000049",
            INIT_79 => X"0000001c0000001d000000200000001f0000001c00000019000000110000001a",
            INIT_7A => X"000000060000000800000016000000140000000c000000100000001500000018",
            INIT_7B => X"0000001f0000001b0000000f0000000b00000008000000080000000700000008",
            INIT_7C => X"000000380000004800000053000000580000004e0000004c0000004800000045",
            INIT_7D => X"0000003100000032000000330000002f0000002a0000002b0000002600000020",
            INIT_7E => X"0000000c0000001300000022000000220000001c0000001e000000260000002c",
            INIT_7F => X"0000001d0000001e0000001a000000120000000d0000000f000000100000000e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY18;


    MEM_IFMAP_LAYER0_ENTITY19 : if BRAM_NAME = "ifmap_layer0_entity19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000051000000500000004e000000420000003a000000390000003100000025",
            INIT_01 => X"0000003800000043000000430000004100000042000000490000005200000056",
            INIT_02 => X"0000002700000032000000380000003400000073000000400000003200000032",
            INIT_03 => X"0000001300000015000000120000001d000000240000002e0000002200000016",
            INIT_04 => X"00000042000000480000004a00000043000000440000004d0000004800000043",
            INIT_05 => X"0000002e00000037000000360000003200000034000000390000004000000044",
            INIT_06 => X"000000210000001e000000230000002800000029000000270000002a00000029",
            INIT_07 => X"0000001200000016000000150000001c0000001b0000001e0000002e00000022",
            INIT_08 => X"00000031000000380000003d0000003a0000003e000000480000004400000048",
            INIT_09 => X"000000260000002b0000002a00000026000000280000002b0000002d00000030",
            INIT_0A => X"000000220000001f00000021000000230000001c0000001e0000002300000022",
            INIT_0B => X"000000110000001300000014000000150000000e0000000d0000002200000030",
            INIT_0C => X"000000240000002b000000300000003e0000003c0000003d0000003600000038",
            INIT_0D => X"0000002000000022000000210000001f00000020000000220000002300000023",
            INIT_0E => X"000000250000001d0000001c000000200000001d0000001b0000001e0000001d",
            INIT_0F => X"000000110000001000000013000000160000000f0000000b000000120000002a",
            INIT_10 => X"0000001b0000002000000024000000340000003b000000420000003900000039",
            INIT_11 => X"0000001e0000001c0000001a0000001a0000001a0000001c0000001d0000001c",
            INIT_12 => X"0000002a00000043000000300000001c0000001c0000001c0000001c0000001c",
            INIT_13 => X"00000011000000130000001f0000001b000000190000000d0000001200000019",
            INIT_14 => X"00000016000000190000001a0000001a000000210000002f0000003a0000003b",
            INIT_15 => X"0000001f0000001b0000001800000018000000190000001a0000001900000017",
            INIT_16 => X"0000003c0000005e0000005d000000210000001e000000210000001e0000001d",
            INIT_17 => X"00000013000000180000002d0000002b0000002c0000001e0000001b00000029",
            INIT_18 => X"0000001500000016000000170000001600000014000000170000001c00000022",
            INIT_19 => X"000000230000001d00000019000000180000001a000000190000001600000016",
            INIT_1A => X"000000250000003700000059000000330000001e000000230000001f00000020",
            INIT_1B => X"00000015000000170000001e000000240000002d0000002b0000002800000038",
            INIT_1C => X"0000001600000016000000170000001600000012000000100000001100000011",
            INIT_1D => X"000000270000001d0000001b000000190000001b0000001a0000001700000018",
            INIT_1E => X"0000000b00000012000000400000004100000030000000330000002d00000028",
            INIT_1F => X"00000015000000160000001600000019000000200000001f0000002500000022",
            INIT_20 => X"0000001700000017000000160000001500000012000000120000001200000011",
            INIT_21 => X"0000003b0000003300000038000000250000001e0000001c0000001800000019",
            INIT_22 => X"0000001000000011000000280000003d00000036000000370000003a0000003b",
            INIT_23 => X"0000001400000015000000170000001a0000001b00000018000000190000001a",
            INIT_24 => X"0000001800000016000000140000001500000012000000120000001200000013",
            INIT_25 => X"00000034000000390000004c0000003e00000031000000200000001900000018",
            INIT_26 => X"0000002c0000003000000031000000380000003a000000320000002e00000031",
            INIT_27 => X"0000001400000014000000180000001900000019000000190000002300000029",
            INIT_28 => X"0000001700000015000000150000001500000012000000130000001200000014",
            INIT_29 => X"0000004a0000003e000000420000003100000035000000240000001900000019",
            INIT_2A => X"000000210000004b000000680000007c000000b8000000a60000008900000068",
            INIT_2B => X"0000001300000012000000190000001800000019000000260000003d00000038",
            INIT_2C => X"0000001800000016000000180000001800000013000000140000001200000015",
            INIT_2D => X"000000be000000b20000009700000055000000300000001f0000001d00000019",
            INIT_2E => X"0000001600000098000000d0000000b2000000c5000000ca000000cd000000cd",
            INIT_2F => X"0000001100000011000000160000001500000028000000460000002500000018",
            INIT_30 => X"0000001a00000019000000180000001800000015000000160000001400000014",
            INIT_31 => X"000000750000008c0000009b0000009000000070000000420000002000000019",
            INIT_32 => X"0000004e000000d5000000e8000000750000003d000000470000005800000064",
            INIT_33 => X"0000001000000011000000150000001a00000046000000320000000a0000000f",
            INIT_34 => X"0000001a00000019000000170000001700000016000000190000001600000014",
            INIT_35 => X"000000120000003400000056000000500000005b00000067000000480000001a",
            INIT_36 => X"0000009b000000e0000000dd0000007c000000100000000f0000002200000011",
            INIT_37 => X"000000100000001200000013000000210000003b000000160000000700000024",
            INIT_38 => X"00000015000000130000001900000018000000160000001b0000001700000018",
            INIT_39 => X"00000018000000320000004e0000003d000000290000003a0000005500000037",
            INIT_3A => X"000000cd000000d1000000d8000000bf000000490000001e0000002b0000000b",
            INIT_3B => X"0000001200000014000000160000001b00000017000000100000000e00000067",
            INIT_3C => X"000000340000003c0000002500000019000000170000001a000000160000001a",
            INIT_3D => X"000000260000002e0000004d000000500000003b00000038000000340000004c",
            INIT_3E => X"000000d2000000d9000000d8000000df000000c40000007c0000004900000023",
            INIT_3F => X"000000110000003e000000470000001f0000000e000000150000003900000076",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005c00000060000000350000002100000017000000190000001400000019",
            INIT_41 => X"000000a20000005a0000004700000051000000420000003e0000005d00000049",
            INIT_42 => X"00000079000000de000000e4000000e3000000f5000000f5000000df000000c4",
            INIT_43 => X"00000013000000750000008c0000004800000009000000110000003b00000025",
            INIT_44 => X"00000045000000350000002c000000280000001a000000180000001500000019",
            INIT_45 => X"000000fb00000094000000200000003100000029000000250000005200000058",
            INIT_46 => X"0000001f0000008b000000e2000000e1000000e2000000e9000000f2000000f6",
            INIT_47 => X"0000002200000097000000a2000000850000004300000028000000190000000b",
            INIT_48 => X"000000360000002e000000460000005d00000026000000160000001300000016",
            INIT_49 => X"000000e3000000a300000031000000380000001b00000018000000260000004b",
            INIT_4A => X"0000004a000000a3000000e4000000e5000000da000000cb000000cd000000d6",
            INIT_4B => X"00000033000000a0000000960000009700000095000000800000005a00000039",
            INIT_4C => X"0000002a000000240000005a000000af0000007c000000260000000f00000013",
            INIT_4D => X"000000d0000000aa0000004f00000040000000150000000b000000170000003f",
            INIT_4E => X"000000b1000000e3000000d9000000ce000000d6000000d3000000c5000000c7",
            INIT_4F => X"0000002a00000088000000970000009a000000a2000000a7000000a800000098",
            INIT_50 => X"0000002e0000002f0000006f000000be000000dc000000650000000a00000012",
            INIT_51 => X"000000cc000000b1000000420000001f0000000e000000090000000a00000039",
            INIT_52 => X"000000d3000000ac000000660000004f0000007c000000c6000000ca000000c2",
            INIT_53 => X"000000110000004a0000008c0000009c000000a9000000b1000000b8000000c8",
            INIT_54 => X"00000034000000370000008000000096000000a500000084000000140000000e",
            INIT_55 => X"000000c6000000b4000000480000002d000000160000000a000000030000001e",
            INIT_56 => X"000000a3000000380000001e0000001a000000190000007b000000cd000000be",
            INIT_57 => X"000000110000000d0000004400000088000000930000009e000000b8000000ca",
            INIT_58 => X"000000350000003e00000082000000530000002100000053000000230000000a",
            INIT_59 => X"000000c2000000b7000000750000006c00000048000000100000000700000013",
            INIT_5A => X"0000004f000000140000002b000000310000001e0000002f000000b7000000c3",
            INIT_5B => X"00000018000000090000000a00000040000000810000008400000094000000a1",
            INIT_5C => X"000000240000004e00000088000000460000002300000037000000210000000a",
            INIT_5D => X"000000cd000000cd0000007e000000610000005800000022000000110000000f",
            INIT_5E => X"0000001f000000200000001f000000200000002b0000002000000098000000d0",
            INIT_5F => X"00000021000000190000000c00000017000000630000008a0000009100000075",
            INIT_60 => X"000000210000005700000088000000470000004100000036000000150000000a",
            INIT_61 => X"000000c5000000cf0000009a00000056000000570000003f0000002700000015",
            INIT_62 => X"0000000f0000001c0000002c00000037000000380000002500000081000000c6",
            INIT_63 => X"0000001f0000001c000000140000000e000000430000008b000000930000004d",
            INIT_64 => X"0000001c0000005600000080000000450000003e0000002f0000000e00000007",
            INIT_65 => X"000000b4000000b6000000a20000006f0000006f0000005e0000003c0000001e",
            INIT_66 => X"0000000f00000023000000350000004b0000003c000000290000007f000000bc",
            INIT_67 => X"00000016000000100000000d00000007000000260000006f0000007a0000002c",
            INIT_68 => X"0000003d0000006800000075000000460000003b00000027000000110000000b",
            INIT_69 => X"000000c7000000c9000000c3000000b9000000b70000009f0000007900000051",
            INIT_6A => X"0000001c0000003400000062000000660000003c0000002a00000088000000c6",
            INIT_6B => X"000000160000000c000000070000000300000010000000450000004f00000015",
            INIT_6C => X"0000003c000000550000006700000049000000430000001d0000001400000013",
            INIT_6D => X"0000006d000000710000007100000068000000640000005b0000005000000045",
            INIT_6E => X"000000170000001f00000042000000400000004100000025000000590000006d",
            INIT_6F => X"000000180000000b0000000600000006000000050000000e0000001400000008",
            INIT_70 => X"00000007000000160000002c0000002c000000250000001d0000001c00000017",
            INIT_71 => X"0000001000000011000000100000000d0000000c0000000c0000000a0000000a",
            INIT_72 => X"0000001000000038000000300000004400000043000000090000000f0000000f",
            INIT_73 => X"000000190000000e000000090000000600000004000000030000000300000004",
            INIT_74 => X"0000002000000019000000120000001700000020000000270000002500000021",
            INIT_75 => X"0000000f00000013000000150000001700000017000000170000001500000017",
            INIT_76 => X"0000000800000029000000470000003e00000018000000070000000a0000000b",
            INIT_77 => X"0000001d000000180000000e0000000900000006000000050000000500000004",
            INIT_78 => X"0000004d00000051000000430000003c00000032000000290000002500000023",
            INIT_79 => X"00000023000000270000002c00000031000000300000002d000000240000002c",
            INIT_7A => X"000000090000000a000000190000001700000010000000150000001b0000001d",
            INIT_7B => X"0000001e0000001f000000140000000e0000000b0000000a000000090000000b",
            INIT_7C => X"00000052000000660000006f0000006d000000570000003b0000002a0000002a",
            INIT_7D => X"0000004300000046000000480000004a00000047000000450000003e00000037",
            INIT_7E => X"00000012000000180000002c0000002f000000290000002b000000330000003b",
            INIT_7F => X"0000001e000000200000001c0000001600000013000000150000001600000014",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY19;


    MEM_IFMAP_LAYER0_ENTITY20 : if BRAM_NAME = "ifmap_layer0_entity20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000002000000050000000a000000090000000a0000000e0000000b0000000d",
            INIT_01 => X"0000000000000005000000060000000400000002000000010000000300000003",
            INIT_02 => X"000000080000001d000000170000001600000056000000230000000000000001",
            INIT_03 => X"000000050000000600000008000000130000001d000000270000001b0000000d",
            INIT_04 => X"00000000000000030000000800000007000000040000000a0000000c0000000d",
            INIT_05 => X"0000000100000004000000040000000200000001000000010000000200000004",
            INIT_06 => X"0000000700000006000000060000000700000013000000100000000100000001",
            INIT_07 => X"0000000600000004000000080000001300000016000000170000002e00000021",
            INIT_08 => X"0000000000000001000000040000000400000000000000030000000400000007",
            INIT_09 => X"0000000300000005000000060000000400000004000000040000000400000004",
            INIT_0A => X"0000000a000000060000000700000004000000090000000c0000000300000004",
            INIT_0B => X"0000000600000003000000060000000f0000000c0000000d0000002300000028",
            INIT_0C => X"000000030000000300000004000000120000000b000000080000000300000001",
            INIT_0D => X"0000000600000006000000090000000800000007000000080000000600000005",
            INIT_0E => X"00000017000000100000000a00000004000000090000000a0000000500000007",
            INIT_0F => X"0000000800000005000000060000000f0000000e00000011000000160000001e",
            INIT_10 => X"000000080000000700000006000000170000001a0000001d000000130000000c",
            INIT_11 => X"00000008000000070000000a0000000900000008000000090000000800000007",
            INIT_12 => X"0000002700000040000000250000000800000007000000080000000700000009",
            INIT_13 => X"000000090000000d0000000f0000000e000000150000000e0000001000000010",
            INIT_14 => X"000000080000000900000006000000090000000c000000160000001e00000018",
            INIT_15 => X"00000009000000070000000a0000000b0000000a000000090000000500000005",
            INIT_16 => X"0000003b0000005d0000005500000014000000070000000b0000000b0000000a",
            INIT_17 => X"00000009000000100000001b0000001700000020000000130000000e00000022",
            INIT_18 => X"000000070000000a0000000800000008000000070000000a0000000b0000000c",
            INIT_19 => X"0000000c0000000a0000000c0000000d0000000e0000000a0000000500000006",
            INIT_1A => X"000000280000003c0000005600000025000000070000000e0000000e00000009",
            INIT_1B => X"000000070000000600000010000000140000001c0000001c0000001c00000035",
            INIT_1C => X"000000090000000c0000000a0000000b00000007000000060000000600000003",
            INIT_1D => X"0000001300000010000000120000000e0000000e0000000c0000000800000009",
            INIT_1E => X"0000000a000000140000003e00000031000000160000001a0000001500000010",
            INIT_1F => X"000000070000000400000008000000090000000d000000100000001a0000001e",
            INIT_20 => X"0000000b0000000e0000000a0000000b00000008000000090000000a00000007",
            INIT_21 => X"000000280000002200000024000000130000000f0000000e0000000c0000000d",
            INIT_22 => X"000000090000000f0000002b0000003300000022000000220000002000000024",
            INIT_23 => X"000000080000000800000008000000080000000a000000090000000c00000014",
            INIT_24 => X"0000000d0000000e0000000a0000000c000000080000000b0000000c0000000c",
            INIT_25 => X"0000002600000028000000310000002700000022000000140000000e0000000e",
            INIT_26 => X"00000026000000340000003b0000003600000032000000270000001b00000020",
            INIT_27 => X"0000000a0000000b00000009000000060000000c0000000b0000001500000023",
            INIT_28 => X"0000000d0000000d0000000a0000000c000000090000000b0000000b0000000c",
            INIT_29 => X"0000003f000000320000003200000020000000280000001b000000100000000d",
            INIT_2A => X"00000022000000540000007100000079000000b4000000a10000007700000058",
            INIT_2B => X"0000000a0000000c0000000a00000009000000110000001d0000003100000032",
            INIT_2C => X"0000000c0000000d0000000c0000000e0000000b0000000e0000000a00000009",
            INIT_2D => X"000000ba000000af000000930000004d0000002700000018000000120000000c",
            INIT_2E => X"0000001c0000009e000000d5000000b1000000ca000000d2000000c8000000c8",
            INIT_2F => X"000000090000000b000000090000000a00000025000000460000002200000013",
            INIT_30 => X"0000000e0000000d0000000e000000100000000d0000000f0000000a00000008",
            INIT_31 => X"0000007d00000093000000a20000008e0000006c0000003e000000180000000c",
            INIT_32 => X"00000054000000d7000000f10000007e0000004a000000540000005e0000006e",
            INIT_33 => X"00000008000000090000000d000000190000004900000034000000090000000c",
            INIT_34 => X"0000000e0000000c00000010000000110000000e0000000f0000000b0000000b",
            INIT_35 => X"000000190000003d0000005f000000560000005d000000670000004400000014",
            INIT_36 => X"000000a7000000eb000000eb0000008900000017000000110000002300000016",
            INIT_37 => X"000000070000000900000011000000280000004200000017000000070000002a",
            INIT_38 => X"000000120000000b00000012000000100000000e000000120000000d0000000f",
            INIT_39 => X"0000001b0000003700000053000000440000002e0000003b0000005300000036",
            INIT_3A => X"000000e0000000e7000000e8000000c80000004c0000001c000000270000000c",
            INIT_3B => X"000000080000000d000000160000001f0000001a000000130000001600000073",
            INIT_3C => X"00000037000000390000001e0000000e0000000e000000130000000d00000010",
            INIT_3D => X"00000029000000320000004e000000520000003c00000039000000350000004f",
            INIT_3E => X"000000dd000000ec000000e6000000e7000000c80000007c0000004700000023",
            INIT_3F => X"000000090000003f00000049000000200000000e0000001a000000440000007e",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005c0000005d0000002f0000001800000011000000130000000e00000011",
            INIT_41 => X"000000a60000005e000000470000004c0000003d0000003c000000620000004f",
            INIT_42 => X"0000007c000000e7000000f0000000ed000000fc000000fa000000e2000000c6",
            INIT_43 => X"000000110000007e000000950000004c0000000c0000001c0000004a0000002a",
            INIT_44 => X"00000048000000380000002a0000002400000015000000120000001000000012",
            INIT_45 => X"000001000000009a000000220000002d00000024000000240000005800000060",
            INIT_46 => X"0000002700000096000000ee000000ed000000ed000000f4000000f9000000fa",
            INIT_47 => X"00000026000000a3000000ae0000008e0000004d0000003b0000002e00000015",
            INIT_48 => X"000000420000003c000000490000005c00000022000000100000001000000011",
            INIT_49 => X"000000f0000000ae000000370000003e000000210000001c0000002c00000054",
            INIT_4A => X"00000056000000b1000000ee000000ef000000e7000000d9000000d9000000e1",
            INIT_4B => X"00000037000000a9000000a1000000a4000000a4000000920000006a00000045",
            INIT_4C => X"000000380000003500000062000000b40000007d000000200000000a0000000d",
            INIT_4D => X"000000e0000000b900000059000000490000001b0000000e0000001c00000048",
            INIT_4E => X"000000c0000000f2000000e1000000d7000000e3000000e4000000d5000000d5",
            INIT_4F => X"0000002a0000008d0000009f000000a6000000b0000000b5000000b4000000a5",
            INIT_50 => X"000000390000003e0000007b000000c9000000e500000065000000070000000c",
            INIT_51 => X"000000da000000bf0000004f000000260000000f000000090000000f00000041",
            INIT_52 => X"000000e4000000b80000006d000000580000008a000000d8000000db000000d0",
            INIT_53 => X"0000000e0000004d00000093000000a6000000b5000000bf000000c9000000da",
            INIT_54 => X"0000003d000000450000008d000000a2000000b30000008b000000180000000d",
            INIT_55 => X"000000d4000000c200000056000000360000001b0000000b0000000400000023",
            INIT_56 => X"000000b10000004000000022000000200000002400000088000000db000000cc",
            INIT_57 => X"0000000d0000000f00000049000000900000009f000000ad000000cc000000dd",
            INIT_58 => X"0000003e0000004c0000008f00000060000000310000005b0000002700000009",
            INIT_59 => X"000000d0000000c5000000830000007900000051000000150000000700000015",
            INIT_5A => X"00000059000000190000002e000000370000002600000038000000c1000000d1",
            INIT_5B => X"00000014000000080000000e000000480000008d00000095000000a9000000b2",
            INIT_5C => X"0000002d0000005c0000009500000053000000300000003b0000002200000005",
            INIT_5D => X"000000db000000db0000008c0000006f000000640000002a000000130000000f",
            INIT_5E => X"000000270000002400000023000000250000003300000026000000a0000000de",
            INIT_5F => X"0000001e000000160000000c0000001d0000006e0000009b000000a400000082",
            INIT_60 => X"0000002a0000006500000094000000540000004d0000003a0000001700000007",
            INIT_61 => X"000000d3000000dd000000a800000064000000650000004a0000002b00000016",
            INIT_62 => X"0000001500000023000000340000003f000000400000002b00000089000000d4",
            INIT_63 => X"0000001c0000001800000012000000130000004e0000009a000000a200000056",
            INIT_64 => X"00000025000000650000008c000000520000004c000000370000001500000009",
            INIT_65 => X"000000c2000000c3000000b00000007e0000007f0000006c0000004300000021",
            INIT_66 => X"000000150000002e0000004100000056000000460000003000000087000000c9",
            INIT_67 => X"000000140000000b0000000a0000000b000000310000007b0000008300000032",
            INIT_68 => X"0000004b0000007800000084000000570000004900000031000000170000000b",
            INIT_69 => X"000000d5000000d4000000cf000000c8000000c8000000b1000000860000005d",
            INIT_6A => X"00000022000000400000006e00000071000000480000003500000094000000d6",
            INIT_6B => X"000000160000000d0000000900000007000000160000004c0000005500000018",
            INIT_6C => X"000000480000006000000073000000570000004e00000025000000160000000f",
            INIT_6D => X"0000007b0000007e0000007d0000007700000072000000690000005d00000052",
            INIT_6E => X"0000001b000000290000004e0000004b0000004c00000030000000660000007c",
            INIT_6F => X"000000190000000f0000000a0000000800000006000000100000001800000009",
            INIT_70 => X"0000000c0000001900000030000000320000002b000000230000001f00000015",
            INIT_71 => X"000000190000001a000000180000001400000011000000110000000e0000000e",
            INIT_72 => X"00000012000000410000003b0000004e0000004a0000000d0000001400000018",
            INIT_73 => X"0000001a0000000d000000090000000500000003000000040000000500000003",
            INIT_74 => X"000000250000001e000000170000001e000000250000002c0000002800000021",
            INIT_75 => X"0000001300000017000000180000001b0000001c0000001c000000190000001c",
            INIT_76 => X"000000080000002f00000053000000470000001c00000006000000090000000f",
            INIT_77 => X"0000001c000000150000000b0000000600000004000000050000000500000002",
            INIT_78 => X"000000590000005c0000004f000000490000003b000000300000002900000025",
            INIT_79 => X"000000280000002b00000030000000390000003b000000380000002f00000038",
            INIT_7A => X"0000000800000010000000250000002100000015000000150000001b00000023",
            INIT_7B => X"0000001c0000001d000000120000000d0000000a0000000a0000000900000008",
            INIT_7C => X"000000630000007600000080000000800000006500000046000000310000002c",
            INIT_7D => X"0000004f00000051000000530000005700000055000000540000004e00000047",
            INIT_7E => X"0000001300000020000000380000003a00000031000000310000003c00000047",
            INIT_7F => X"0000001c000000220000001f0000001900000015000000180000001800000013",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY20;


    MEM_IFMAP_LAYER0_ENTITY21 : if BRAM_NAME = "ifmap_layer0_entity21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005c0000005b00000055000000510000004d000000510000005200000053",
            INIT_01 => X"0000004c0000005000000052000000570000005c000000650000005f0000005c",
            INIT_02 => X"0000002f00000034000000380000003c0000003e0000003f0000004100000044",
            INIT_03 => X"00000015000000190000001d000000240000002200000023000000250000002a",
            INIT_04 => X"0000005d0000005a00000054000000500000004d000000530000005300000054",
            INIT_05 => X"0000004c0000004e0000005200000058000000610000005f000000580000005a",
            INIT_06 => X"0000002e00000034000000360000003d00000042000000400000004400000047",
            INIT_07 => X"0000001f0000001d0000001e000000240000002300000024000000260000002a",
            INIT_08 => X"0000004c00000058000000540000004b0000004b000000500000005100000052",
            INIT_09 => X"0000004c0000004d000000580000006500000063000000570000005600000052",
            INIT_0A => X"0000002d00000034000000370000003a00000040000000400000004400000049",
            INIT_0B => X"000000350000003100000030000000310000002c00000029000000280000002b",
            INIT_0C => X"0000003200000050000000570000004a0000004e000000500000005100000053",
            INIT_0D => X"000000500000005800000066000000680000005b000000570000006100000055",
            INIT_0E => X"0000003a00000039000000380000003b0000003f0000003f0000004000000049",
            INIT_0F => X"0000004500000045000000470000004900000047000000440000003f0000003d",
            INIT_10 => X"000000370000004c000000530000004a0000004f0000004f0000004f0000004f",
            INIT_11 => X"000000570000005a000000590000004e0000004b0000004b0000005400000053",
            INIT_12 => X"0000005700000054000000500000004e00000046000000430000004200000053",
            INIT_13 => X"000000490000004f000000540000005800000059000000590000005600000057",
            INIT_14 => X"000000460000004600000049000000490000004d0000004b0000004a0000004c",
            INIT_15 => X"000000510000004e0000004e0000004b00000049000000470000004500000046",
            INIT_16 => X"000000680000006600000068000000640000006200000060000000590000005a",
            INIT_17 => X"000000420000004900000050000000570000005e000000610000005f00000063",
            INIT_18 => X"000000330000002b0000003e0000004a0000004900000047000000480000004a",
            INIT_19 => X"0000005e000000510000004a0000004b00000047000000440000004000000044",
            INIT_1A => X"0000006d000000680000006400000066000000720000006e0000006200000060",
            INIT_1B => X"0000004300000046000000490000004c00000050000000550000005b00000063",
            INIT_1C => X"000000290000002a0000003a0000004700000048000000470000004800000047",
            INIT_1D => X"000000600000005200000047000000410000003f0000003a0000003600000039",
            INIT_1E => X"000000610000006c0000006a00000067000000670000005d0000005e00000069",
            INIT_1F => X"0000004d0000004f000000500000005000000050000000540000005b0000005d",
            INIT_20 => X"0000002e000000570000006700000058000000520000004b0000004900000049",
            INIT_21 => X"000000570000005a000000570000005100000052000000450000003800000038",
            INIT_22 => X"000000660000006a00000066000000610000005b0000005e0000006300000062",
            INIT_23 => X"0000005f0000005b00000059000000590000005c00000061000000630000005e",
            INIT_24 => X"000000330000006800000099000000880000007b0000006d0000005f00000056",
            INIT_25 => X"0000005a000000660000006c0000006500000061000000490000003b0000003c",
            INIT_26 => X"0000006e00000069000000630000005d0000005d00000061000000610000005f",
            INIT_27 => X"0000006e0000006e0000006e0000006d0000006c0000006c0000006900000067",
            INIT_28 => X"0000003200000057000000a2000000a00000009d000000960000008b0000007f",
            INIT_29 => X"0000005a0000006b000000700000006500000058000000350000003800000043",
            INIT_2A => X"00000065000000600000005f00000060000000600000005e000000600000005e",
            INIT_2B => X"0000007000000074000000770000007b0000007e0000007d0000007100000068",
            INIT_2C => X"0000002c0000005a0000009f000000a0000000a20000009f0000009d00000098",
            INIT_2D => X"0000005c000000610000005a00000067000000560000003a0000004500000048",
            INIT_2E => X"0000005c0000005700000062000000630000005e0000005f000000600000005a",
            INIT_2F => X"0000006c00000074000000790000007f00000083000000830000007000000061",
            INIT_30 => X"000000300000007200000094000000980000009d000000a00000009e0000009b",
            INIT_31 => X"0000005d000000580000006000000073000000670000005e0000005800000044",
            INIT_32 => X"000000550000005400000065000000630000005e000000620000006500000059",
            INIT_33 => X"0000005f0000006b000000760000007f000000840000007d0000006e00000069",
            INIT_34 => X"00000050000000880000008e0000009000000092000000950000009400000094",
            INIT_35 => X"0000005e0000005c0000007100000072000000680000005e000000480000002f",
            INIT_36 => X"000000520000005500000061000000600000005d00000061000000670000005d",
            INIT_37 => X"0000004d000000570000006400000070000000790000006f0000006b0000006b",
            INIT_38 => X"0000008900000097000000930000008e0000008c0000008a0000008700000086",
            INIT_39 => X"000000620000005a0000005e000000590000003e00000032000000490000005d",
            INIT_3A => X"00000053000000560000005e0000005e00000061000000670000006900000066",
            INIT_3B => X"0000004b0000004a000000520000005f000000660000005c000000650000005f",
            INIT_3C => X"000000980000009a0000009f00000098000000900000008b0000008600000083",
            INIT_3D => X"000000660000005f00000064000000670000003900000035000000760000009e",
            INIT_3E => X"00000055000000570000005b000000610000006a0000006f000000740000006e",
            INIT_3F => X"0000005f0000005a000000550000005300000053000000550000006200000054",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007300000089000000a1000000a4000000a0000000980000009000000087",
            INIT_41 => X"00000067000000680000007a0000007b0000006e00000080000000910000009d",
            INIT_42 => X"00000057000000580000005a00000061000000680000006c0000006d00000069",
            INIT_43 => X"0000005e00000069000000690000006500000055000000570000005c0000004f",
            INIT_44 => X"0000007f000000b0000000b3000000aa000000a40000009f0000009a00000094",
            INIT_45 => X"00000067000000800000009100000071000000980000009d000000c5000000b0",
            INIT_46 => X"000000590000005b0000005f0000006100000066000000680000006500000067",
            INIT_47 => X"0000004600000056000000680000006d0000005b0000005b000000560000004f",
            INIT_48 => X"000000c4000000f8000000ee000000dd000000c5000000b2000000a40000009b",
            INIT_49 => X"0000006a000000890000008e0000006c000000b8000000b0000000c80000009c",
            INIT_4A => X"000000590000005f000000630000006500000065000000640000006300000064",
            INIT_4B => X"00000047000000490000005200000058000000530000005c0000005100000050",
            INIT_4C => X"000000f4000000fb000000f6000000fd000000f9000000eb000000d6000000bf",
            INIT_4D => X"0000006e0000008b0000007200000071000000c3000000ac0000009e000000a0",
            INIT_4E => X"0000005c00000066000000680000006700000063000000610000006200000062",
            INIT_4F => X"000000480000004a000000500000004b00000049000000550000004e00000053",
            INIT_50 => X"000000c9000000ba000000bb000000f3000000fe000000fd000000fc000000f5",
            INIT_51 => X"00000072000000800000006a000000740000009c000000970000008000000091",
            INIT_52 => X"0000005c000000690000006e0000006c00000067000000650000006700000068",
            INIT_53 => X"000000490000004d000000530000004e00000055000000540000004c00000052",
            INIT_54 => X"000000720000006b0000007e000000e900000100000000fc000000fc000000fb",
            INIT_55 => X"000000670000006800000063000000630000006e000000780000007300000069",
            INIT_56 => X"00000056000000600000006e000000700000006b0000006b0000006e0000006d",
            INIT_57 => X"0000004f00000052000000520000005b000000680000005a0000004c0000004e",
            INIT_58 => X"00000076000000720000007c000000c8000000eb000000f6000000f8000000f8",
            INIT_59 => X"000000440000004b00000056000000500000004f00000053000000570000005d",
            INIT_5A => X"000000610000006100000061000000620000006100000062000000640000005f",
            INIT_5B => X"0000005200000052000000550000006e0000006f0000005b000000570000005b",
            INIT_5C => X"0000008400000085000000880000008a00000096000000b5000000d6000000eb",
            INIT_5D => X"0000003a0000006000000059000000430000003c000000390000003d00000064",
            INIT_5E => X"0000006500000068000000650000005e00000050000000470000004500000033",
            INIT_5F => X"000000510000005100000062000000770000006d0000005e000000570000005d",
            INIT_60 => X"000000670000006f0000007a0000007c000000780000007a0000008200000099",
            INIT_61 => X"000000530000006a000000660000004500000034000000390000005a0000006a",
            INIT_62 => X"0000006d000000660000006700000064000000550000004d0000004700000040",
            INIT_63 => X"000000500000005c0000007300000071000000630000005d000000570000006a",
            INIT_64 => X"0000006d0000006600000061000000650000006d000000720000006f0000006d",
            INIT_65 => X"000000590000005f000000650000005d00000055000000670000007800000075",
            INIT_66 => X"000000660000006900000077000000720000005a000000520000004b0000004a",
            INIT_67 => X"0000004f0000006b0000007500000065000000620000005e0000006b0000006f",
            INIT_68 => X"000000710000006f0000006a000000630000005b0000005d0000006200000069",
            INIT_69 => X"0000005c000000540000004c000000500000005f000000610000006800000070",
            INIT_6A => X"0000005e000000690000007b00000075000000590000004f0000004800000051",
            INIT_6B => X"0000005a0000006f000000690000006000000065000000670000006700000060",
            INIT_6C => X"000000640000006b0000006e0000006c000000650000005e0000005700000057",
            INIT_6D => X"0000005c0000004c000000490000005d0000006800000056000000510000005b",
            INIT_6E => X"000000560000005d000000640000005b0000004f0000004f0000004d00000058",
            INIT_6F => X"0000006500000066000000600000006000000060000000610000005c00000057",
            INIT_70 => X"00000050000000560000005f000000650000006900000067000000600000005a",
            INIT_71 => X"0000005d0000006000000055000000620000006a000000600000005500000051",
            INIT_72 => X"0000005b000000540000004c000000470000004c0000004f0000005100000058",
            INIT_73 => X"000000600000005b00000060000000620000005a00000053000000560000005c",
            INIT_74 => X"0000004f0000004f0000004f00000050000000560000005f0000006300000064",
            INIT_75 => X"000000590000006100000060000000630000006c000000620000005300000052",
            INIT_76 => X"00000059000000520000004a0000004c000000510000004f000000540000005c",
            INIT_77 => X"00000053000000530000005c0000005d0000005600000052000000550000005a",
            INIT_78 => X"0000005300000059000000570000004d00000047000000490000004e00000057",
            INIT_79 => X"0000005c0000005900000067000000640000006a000000610000004f00000051",
            INIT_7A => X"00000053000000540000004f0000005200000059000000580000005700000060",
            INIT_7B => X"000000490000004f000000560000005600000053000000560000005a00000056",
            INIT_7C => X"0000005100000053000000560000005400000049000000460000003f0000003e",
            INIT_7D => X"000000580000005b000000680000005f0000006b0000005e0000004a0000004e",
            INIT_7E => X"000000530000005500000050000000550000005900000058000000580000005b",
            INIT_7F => X"000000480000004c0000004d0000004c00000050000000560000005900000054",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY21;


    MEM_IFMAP_LAYER0_ENTITY22 : if BRAM_NAME = "ifmap_layer0_entity22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000060000000600000005a0000005a000000590000005d0000005e0000005e",
            INIT_01 => X"0000005200000055000000580000005e000000650000006e0000006600000061",
            INIT_02 => X"000000380000003d000000410000004500000048000000490000004b0000004e",
            INIT_03 => X"000000190000001d000000220000002800000027000000290000002e00000033",
            INIT_04 => X"000000620000005f0000005900000059000000590000005f0000005f00000060",
            INIT_05 => X"000000520000005500000059000000600000006b0000006a0000006000000061",
            INIT_06 => X"000000350000003b0000003d0000004400000049000000470000004b0000004f",
            INIT_07 => X"0000001f0000001f000000200000002600000025000000270000002c00000031",
            INIT_08 => X"000000510000005d0000005a00000054000000570000005c0000005c0000005e",
            INIT_09 => X"000000540000005600000062000000700000006e000000630000006000000059",
            INIT_0A => X"00000030000000360000003a0000003f0000004600000044000000490000004f",
            INIT_0B => X"00000031000000300000002e0000002f0000002b000000290000002b0000002e",
            INIT_0C => X"00000039000000560000005d000000530000005a0000005c0000005d0000005f",
            INIT_0D => X"0000005a00000065000000720000007400000068000000630000006b0000005d",
            INIT_0E => X"0000003900000038000000380000003e0000004200000042000000430000004e",
            INIT_0F => X"0000003d0000003f000000410000004300000042000000410000003e0000003c",
            INIT_10 => X"0000003e0000005200000059000000530000005b0000005b0000005b0000005c",
            INIT_11 => X"0000006400000069000000680000005c00000058000000580000005f0000005c",
            INIT_12 => X"00000053000000500000004d000000500000004800000045000000460000005b",
            INIT_13 => X"0000003f000000460000004b0000004f00000050000000510000005100000053",
            INIT_14 => X"0000004d0000004c0000004f0000005200000059000000570000005600000058",
            INIT_15 => X"0000005f0000005e0000005e0000005a00000057000000550000005200000050",
            INIT_16 => X"0000006200000060000000640000006400000063000000620000005e00000063",
            INIT_17 => X"000000370000003e000000450000004c0000005300000058000000580000005d",
            INIT_18 => X"000000370000002a0000003d0000005100000054000000520000005400000055",
            INIT_19 => X"000000650000005d000000570000005b00000059000000580000005700000053",
            INIT_1A => X"0000006700000067000000670000006900000073000000700000006400000062",
            INIT_1B => X"00000036000000390000003f000000440000004a0000004e000000500000005b",
            INIT_1C => X"0000002c00000026000000370000004c00000054000000520000005300000052",
            INIT_1D => X"000000630000005b00000053000000500000005100000052000000550000004c",
            INIT_1E => X"0000005e00000071000000720000006d0000006c000000610000006000000067",
            INIT_1F => X"0000003b0000004000000044000000470000004b0000004d0000004d00000052",
            INIT_20 => X"0000003100000055000000680000005e0000005b000000540000005200000051",
            INIT_21 => X"0000005e000000650000006400000061000000630000005b0000005400000049",
            INIT_22 => X"00000067000000720000006f0000006a00000062000000650000006800000065",
            INIT_23 => X"0000004800000047000000460000004a0000004e000000520000005500000057",
            INIT_24 => X"00000036000000680000009d0000008e0000008000000073000000650000005c",
            INIT_25 => X"00000065000000750000007c00000075000000710000005d000000540000004b",
            INIT_26 => X"00000076000000740000006e00000068000000670000006b0000006a00000067",
            INIT_27 => X"0000005200000055000000550000005500000054000000550000005a00000064",
            INIT_28 => X"0000003500000059000000aa000000a6000000a0000000990000008e00000082",
            INIT_29 => X"0000006b0000007f000000820000007700000068000000460000004d00000050",
            INIT_2A => X"000000720000006e000000690000006a0000006a000000690000006c0000006a",
            INIT_2B => X"00000055000000590000005b0000005e00000060000000620000006200000069",
            INIT_2C => X"0000002e0000005d000000a9000000a7000000a4000000a20000009f0000009a",
            INIT_2D => X"000000720000007a000000700000007b000000670000004a0000005600000051",
            INIT_2E => X"0000006e00000067000000690000006b000000670000006a0000006d0000006a",
            INIT_2F => X"000000550000005a0000005e0000006000000063000000650000006100000066",
            INIT_30 => X"00000030000000750000009f0000009e0000009e000000a10000009f0000009d",
            INIT_31 => X"00000075000000740000007800000087000000780000006c0000006500000049",
            INIT_32 => X"00000069000000640000006a00000069000000660000006c000000730000006b",
            INIT_33 => X"0000004c000000550000005d0000006200000065000000600000006000000070",
            INIT_34 => X"0000004c00000087000000930000009300000093000000970000009800000099",
            INIT_35 => X"000000710000007300000085000000830000007500000067000000490000002c",
            INIT_36 => X"00000064000000650000006a0000006a0000006b00000071000000770000006c",
            INIT_37 => X"000000400000004a000000550000005d000000620000005d0000006900000075",
            INIT_38 => X"0000008300000095000000940000008f0000008e0000008e0000008e0000008f",
            INIT_39 => X"0000006d000000680000006b0000006300000046000000350000004100000054",
            INIT_3A => X"00000062000000650000006c0000006e000000750000007d0000007c00000072",
            INIT_3B => X"0000003f0000004100000048000000550000005a000000580000006f0000006c",
            INIT_3C => X"0000009300000099000000a000000099000000910000008e0000008d0000008c",
            INIT_3D => X"0000006e00000065000000680000006a0000003a000000340000006f00000097",
            INIT_3E => X"00000065000000680000006c000000730000008000000087000000890000007b",
            INIT_3F => X"0000004d0000004a000000480000004a0000004e000000590000006f00000063",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007200000088000000a0000000a40000009f0000009b000000950000008f",
            INIT_41 => X"0000006c000000660000007700000076000000680000007a0000008f0000009b",
            INIT_42 => X"0000006a0000006b0000006d0000007500000080000000850000008400000078",
            INIT_43 => X"000000440000004f000000540000005a00000056000000620000006c00000061",
            INIT_44 => X"00000081000000b0000000b1000000a7000000a10000009f0000009d0000009a",
            INIT_45 => X"0000006c0000007b00000089000000680000008e00000097000000c7000000b3",
            INIT_46 => X"0000006e00000070000000730000007700000080000000830000007e00000079",
            INIT_47 => X"00000027000000340000004a0000005c0000005e0000006a0000006900000063",
            INIT_48 => X"000000c7000000f7000000ec000000da000000c1000000b0000000a40000009d",
            INIT_49 => X"00000071000000860000008800000065000000b1000000ad000000ce000000a3",
            INIT_4A => X"00000071000000760000007a0000007d00000081000000820000007e00000077",
            INIT_4B => X"00000027000000250000002c0000003e000000500000006a0000006700000068",
            INIT_4C => X"000000f7000000fa000000f2000000fa000000f6000000e8000000d4000000c0",
            INIT_4D => X"000000780000008b000000700000006e000000c1000000ae000000aa000000a9",
            INIT_4E => X"000000740000007e0000007f0000008000000080000000800000007e00000076",
            INIT_4F => X"0000002b00000027000000250000002a0000003e00000060000000660000006c",
            INIT_50 => X"000000d2000000be000000ba000000f1000000fb000000fa000000fb000000f5",
            INIT_51 => X"0000007a00000087000000730000007d000000a00000009c00000092000000a1",
            INIT_52 => X"000000740000007d0000007f0000007f00000080000000810000007f00000078",
            INIT_53 => X"00000029000000290000002a0000002d0000004200000057000000620000006a",
            INIT_54 => X"000000820000007400000083000000ea000000fe000000fb000000fb000000fb",
            INIT_55 => X"0000006b00000072000000770000007a0000007c000000820000008a0000007f",
            INIT_56 => X"0000006c0000006f000000770000007d0000007f000000820000008000000076",
            INIT_57 => X"000000290000002c0000002f0000003d00000050000000520000005a00000063",
            INIT_58 => X"000000830000007b00000080000000cb000000ef000000f9000000fc000000fc",
            INIT_59 => X"0000004400000051000000690000006a00000067000000660000006c0000006f",
            INIT_5A => X"00000073000000700000006b0000006e00000074000000780000007500000066",
            INIT_5B => X"0000002d0000002d0000003400000051000000540000004b0000005900000068",
            INIT_5C => X"0000008a000000890000008900000090000000a0000000bf000000df000000f5",
            INIT_5D => X"0000003a00000063000000660000005a00000057000000510000004b0000006d",
            INIT_5E => X"000000740000007a000000740000006d000000650000005f000000560000003a",
            INIT_5F => X"0000002f0000002f000000420000005900000050000000460000004d00000061",
            INIT_60 => X"00000069000000700000007b0000008200000084000000860000008d000000a5",
            INIT_61 => X"000000560000006f0000006e00000053000000470000004a0000005e0000006b",
            INIT_62 => X"0000007c0000007b0000007b000000760000006c000000660000005a00000048",
            INIT_63 => X"000000300000003d00000054000000520000004400000042000000490000006c",
            INIT_64 => X"0000006a00000065000000610000006a000000750000007a0000007800000075",
            INIT_65 => X"0000006100000068000000680000005c000000570000006a0000007300000070",
            INIT_66 => X"0000007a000000820000008e00000086000000720000006c0000005f00000054",
            INIT_67 => X"000000320000004f000000570000004500000040000000450000006400000077",
            INIT_68 => X"0000006b0000006e0000006b000000650000005e00000060000000660000006c",
            INIT_69 => X"000000680000005d000000480000004200000051000000560000005d00000067",
            INIT_6A => X"0000007a000000850000009400000089000000710000006b0000005f0000005e",
            INIT_6B => X"0000003f000000550000004b0000004000000042000000510000006b00000072",
            INIT_6C => X"00000057000000650000006c0000006b000000630000005d0000005700000058",
            INIT_6D => X"0000005e0000004e0000003f0000004a00000053000000410000003c00000049",
            INIT_6E => X"000000720000007a0000007b000000690000005d0000005f0000005700000059",
            INIT_6F => X"0000004b0000004a0000003f0000003c0000003b0000004e000000680000006d",
            INIT_70 => X"0000003800000045000000540000005b0000005f000000610000005f0000005d",
            INIT_71 => X"0000004800000055000000490000005300000055000000420000003100000032",
            INIT_72 => X"0000006800000064000000580000004500000044000000430000003e0000003e",
            INIT_73 => X"000000450000003a000000360000003500000033000000400000005a00000065",
            INIT_74 => X"0000003000000034000000370000003b00000044000000510000005b00000060",
            INIT_75 => X"000000390000004d0000004f0000005200000052000000400000002e0000002f",
            INIT_76 => X"0000004a000000470000003f0000003a0000003a000000340000003200000035",
            INIT_77 => X"000000360000003000000031000000300000002e000000340000004100000048",
            INIT_78 => X"0000003000000034000000300000002c0000002b000000310000003c00000049",
            INIT_79 => X"000000350000003e0000004f0000004b000000490000003a0000002c00000030",
            INIT_7A => X"0000002f000000330000002f0000003400000039000000340000002e00000032",
            INIT_7B => X"0000002a0000002b0000002d0000002b0000002a0000002e000000310000002f",
            INIT_7C => X"0000002d00000029000000290000002a00000025000000270000002500000029",
            INIT_7D => X"0000002e0000003b0000004c0000004300000047000000360000002b0000002f",
            INIT_7E => X"0000002d000000310000002d0000002f000000300000002d0000002a0000002b",
            INIT_7F => X"00000026000000280000002800000025000000270000002a0000002d0000002b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY22;


    MEM_IFMAP_LAYER0_ENTITY23 : if BRAM_NAME = "ifmap_layer0_entity23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005f0000005d00000052000000500000004f000000530000005400000055",
            INIT_01 => X"0000004f000000540000004e0000004b000000480000004f000000550000005a",
            INIT_02 => X"00000033000000380000003b0000003c0000003d0000003c0000003e00000044",
            INIT_03 => X"00000015000000190000001e000000240000002300000025000000290000002e",
            INIT_04 => X"0000005d0000005a000000500000004e0000004f000000550000005500000056",
            INIT_05 => X"0000004800000047000000450000004400000047000000460000004900000054",
            INIT_06 => X"0000002e0000003400000035000000380000003e0000003e0000004300000046",
            INIT_07 => X"0000001b0000001a0000001b0000002100000020000000220000002500000029",
            INIT_08 => X"000000480000005600000050000000490000004e000000520000005300000054",
            INIT_09 => X"0000003c000000360000003f0000004800000043000000380000004100000046",
            INIT_0A => X"000000260000002d0000002f000000300000003a0000003d0000004100000042",
            INIT_0B => X"0000002c0000002a000000290000002a00000025000000220000002100000024",
            INIT_0C => X"0000002b0000004d000000520000004800000050000000520000005300000055",
            INIT_0D => X"0000002f000000320000003f0000004100000034000000320000004500000043",
            INIT_0E => X"0000002c0000002b0000002b0000002d00000036000000390000003400000032",
            INIT_0F => X"00000037000000380000003b0000003c0000003b00000038000000320000002f",
            INIT_10 => X"0000002c000000460000004c0000004800000051000000510000005100000052",
            INIT_11 => X"0000002300000026000000270000001f0000001d00000022000000330000003d",
            INIT_12 => X"00000044000000410000003d0000003d0000003b000000390000002b00000029",
            INIT_13 => X"000000380000003e000000430000004700000048000000470000004200000044",
            INIT_14 => X"000000380000003e00000042000000470000004f0000004c0000004c0000004d",
            INIT_15 => X"0000000e0000000f0000001400000016000000170000001a000000210000002c",
            INIT_16 => X"000000500000004e0000005200000053000000540000004f000000350000001f",
            INIT_17 => X"0000002e000000350000003c000000440000004b0000004d000000480000004c",
            INIT_18 => X"0000002000000020000000370000004700000048000000460000004700000049",
            INIT_19 => X"000000150000000e0000000b0000001200000013000000140000001800000026",
            INIT_1A => X"000000520000004f000000500000005600000059000000460000002900000018",
            INIT_1B => X"0000002a0000002d000000340000003b0000004300000048000000480000004b",
            INIT_1C => X"000000110000001c000000330000004300000045000000440000004500000044",
            INIT_1D => X"00000018000000110000000b000000090000000b0000000a0000000c00000017",
            INIT_1E => X"000000400000004d0000004f0000004d0000003f00000021000000160000001c",
            INIT_1F => X"0000002b0000002f000000360000003c00000042000000480000004900000041",
            INIT_20 => X"00000013000000460000005d000000520000004e000000470000004500000044",
            INIT_21 => X"0000001400000021000000210000002000000025000000190000000c00000012",
            INIT_22 => X"0000003b0000003c000000380000003100000021000000190000001800000016",
            INIT_23 => X"000000350000003400000034000000390000003f000000490000004b0000003b",
            INIT_24 => X"00000016000000550000008d0000008000000075000000670000005900000050",
            INIT_25 => X"0000001c000000350000003d0000003900000038000000210000000f00000015",
            INIT_26 => X"0000003a0000002d000000230000001800000014000000160000001600000015",
            INIT_27 => X"0000003d0000003f00000040000000410000004100000046000000480000003d",
            INIT_28 => X"00000018000000470000009800000098000000950000008e0000008300000077",
            INIT_29 => X"000000210000003f000000440000003c0000003100000015000000110000001e",
            INIT_2A => X"0000002b0000001c000000140000000f00000011000000150000001b00000019",
            INIT_2B => X"000000410000004400000047000000490000004a0000004d0000004600000037",
            INIT_2C => X"000000170000004f00000099000000990000009900000096000000940000008f",
            INIT_2D => X"0000002700000037000000300000003d0000002e000000190000002200000028",
            INIT_2E => X"0000001f000000120000001500000013000000150000001f000000240000001d",
            INIT_2F => X"000000450000004a0000004c0000004d0000004d0000004c0000003b0000002a",
            INIT_30 => X"000000200000006b000000920000009200000094000000970000009500000092",
            INIT_31 => X"000000290000002c00000034000000470000003b00000034000000370000002b",
            INIT_32 => X"00000019000000120000001c0000001a0000001e0000002c0000003200000022",
            INIT_33 => X"00000042000000490000004f000000510000005100000045000000320000002e",
            INIT_34 => X"000000400000007e000000890000008a0000008b0000008f0000008f00000090",
            INIT_35 => X"00000024000000280000004000000046000000410000003d0000002e0000001a",
            INIT_36 => X"00000013000000120000001d0000002100000028000000330000003600000024",
            INIT_37 => X"00000037000000400000004a0000004f0000004e0000003c000000330000002f",
            INIT_38 => X"0000007700000089000000880000008600000086000000860000008400000085",
            INIT_39 => X"00000022000000200000002a0000002e000000210000001b0000003100000047",
            INIT_3A => X"00000011000000110000001c00000027000000320000003d0000003900000028",
            INIT_3B => X"00000032000000360000003e0000004600000041000000300000003300000024",
            INIT_3C => X"0000008100000088000000910000008c00000085000000810000007f0000007d",
            INIT_3D => X"000000270000002700000033000000400000001e0000001e0000005a00000084",
            INIT_3E => X"00000013000000140000001c0000002c0000003d000000450000004500000031",
            INIT_3F => X"0000003d0000003c00000039000000350000002d000000290000003000000019",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005a000000750000009100000095000000910000008b000000840000007d",
            INIT_41 => X"00000028000000310000004d0000005700000050000000620000007200000080",
            INIT_42 => X"00000017000000190000001f0000002d0000003c000000440000003f0000002e",
            INIT_43 => X"000000320000003e00000042000000400000002d0000002b0000002a00000015",
            INIT_44 => X"000000680000009e000000a40000009a00000093000000900000008c00000088",
            INIT_45 => X"000000290000004b0000006700000050000000770000007a000000a600000095",
            INIT_46 => X"0000001b0000001f00000028000000300000003c00000041000000380000002d",
            INIT_47 => X"00000014000000230000003900000041000000320000002f0000002300000015",
            INIT_48 => X"000000b2000000eb000000e6000000d2000000b6000000a40000009700000090",
            INIT_49 => X"0000002d00000055000000670000004d000000950000008a000000ab00000085",
            INIT_4A => X"0000001d0000002700000030000000350000003c0000003f000000380000002b",
            INIT_4B => X"00000015000000160000001f00000027000000270000002f0000001d00000017",
            INIT_4C => X"000000e6000000f2000000f2000000f8000000f0000000e1000000cd000000b7",
            INIT_4D => X"00000031000000560000004d000000530000009f00000084000000840000008d",
            INIT_4E => X"000000210000002f00000037000000390000003a0000003c000000370000002a",
            INIT_4F => X"0000001b0000001c0000001d000000190000001c000000270000001a00000019",
            INIT_50 => X"000000b5000000ab000000b0000000ec000000f9000000f7000000f8000000f1",
            INIT_51 => X"00000034000000470000003c0000004d00000076000000720000006200000078",
            INIT_52 => X"0000002000000030000000390000003b0000003a00000039000000360000002e",
            INIT_53 => X"0000001a0000001f000000200000001c00000025000000250000001700000018",
            INIT_54 => X"00000055000000530000006a000000e0000000fd000000f9000000f9000000f8",
            INIT_55 => X"00000031000000340000002e0000003000000041000000510000004e00000047",
            INIT_56 => X"0000001b00000024000000330000003d00000039000000360000003700000033",
            INIT_57 => X"0000001c0000001f0000001f0000002800000036000000270000001600000015",
            INIT_58 => X"0000005e000000600000006d000000c2000000eb000000f5000000f8000000f7",
            INIT_59 => X"000000200000002d0000002b0000001c00000019000000230000003500000041",
            INIT_5A => X"000000290000002b0000002d000000300000002f0000002f000000330000002e",
            INIT_5B => X"0000001e0000001d00000021000000390000003a000000240000001e00000022",
            INIT_5C => X"000000740000007a000000810000008800000098000000b6000000d7000000ec",
            INIT_5D => X"00000022000000490000003400000014000000090000000d0000002300000051",
            INIT_5E => X"000000310000003b0000003b0000002f000000200000001a0000001c00000011",
            INIT_5F => X"0000001d0000001c0000002c0000003f00000034000000220000001a00000023",
            INIT_60 => X"0000005c00000068000000760000007b000000780000007a000000820000009a",
            INIT_61 => X"00000034000000450000003d0000001d000000120000001f000000460000005a",
            INIT_62 => X"0000003d00000041000000470000003a00000028000000240000002400000022",
            INIT_63 => X"0000001c000000270000003c00000038000000280000001f0000001700000030",
            INIT_64 => X"0000005d0000005b000000580000005f000000680000006d0000006b00000069",
            INIT_65 => X"000000310000002f00000038000000380000003e000000560000006200000060",
            INIT_66 => X"00000039000000480000005b0000004c000000300000002a0000002500000028",
            INIT_67 => X"0000001d000000370000003d0000002a000000230000001d0000002c00000036",
            INIT_68 => X"000000580000005b00000058000000560000005100000053000000590000005f",
            INIT_69 => X"000000340000002c00000023000000280000003e000000440000004900000053",
            INIT_6A => X"00000032000000470000005f0000005100000031000000270000001e00000028",
            INIT_6B => X"000000280000003a000000300000002200000023000000250000002a00000029",
            INIT_6C => X"000000400000004c0000005300000057000000550000004f000000490000004b",
            INIT_6D => X"000000310000002900000022000000320000003b0000002a0000002700000033",
            INIT_6E => X"0000002d0000003c000000450000003700000027000000240000001e00000026",
            INIT_6F => X"000000330000003000000024000000200000001d000000220000002600000026",
            INIT_70 => X"000000210000002c00000039000000440000004d0000004f0000004e0000004c",
            INIT_71 => X"000000260000003200000029000000370000003d0000002e0000001e0000001d",
            INIT_72 => X"000000300000002e000000250000001d0000001e0000001d0000001a0000001d",
            INIT_73 => X"0000002f00000024000000200000001e0000001800000019000000250000002e",
            INIT_74 => X"0000001b0000001e000000200000002600000032000000400000004a00000050",
            INIT_75 => X"0000001d0000002c0000002f000000350000003c0000002d0000001b0000001b",
            INIT_76 => X"000000250000002000000018000000190000001c00000017000000170000001c",
            INIT_77 => X"000000220000001c0000001e0000001a00000015000000150000001d00000023",
            INIT_78 => X"0000001c000000210000001d0000001a0000001a000000210000002d0000003a",
            INIT_79 => X"0000001c0000002100000032000000310000003300000027000000180000001b",
            INIT_7A => X"000000170000001900000015000000180000001d00000019000000150000001b",
            INIT_7B => X"00000017000000190000001a0000001500000012000000160000001a00000017",
            INIT_7C => X"0000001900000018000000190000001a0000001500000018000000170000001b",
            INIT_7D => X"0000001800000023000000330000002a0000003000000021000000160000001a",
            INIT_7E => X"000000190000001d000000170000001700000018000000150000001400000015",
            INIT_7F => X"0000001600000018000000160000001100000012000000160000001b00000018",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY23;


    MEM_IFMAP_LAYER0_ENTITY24 : if BRAM_NAME = "ifmap_layer0_entity24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b2000000b7000000bc000000a400000041000000150000001300000017",
            INIT_01 => X"000000b7000000b6000000b7000000b8000000ba000000ba000000ac000000aa",
            INIT_02 => X"000000c2000000990000006e0000006b0000005c0000007f000000a4000000b4",
            INIT_03 => X"000000c5000000c7000000c8000000c9000000c6000000c5000000c9000000c3",
            INIT_04 => X"000000b2000000bf000000ca000000990000002e000000150000001300000017",
            INIT_05 => X"000000b2000000b4000000b8000000ba000000b7000000a90000009e000000a4",
            INIT_06 => X"000000ce000000b40000006a0000004a000000560000008a000000ad000000b4",
            INIT_07 => X"000000ca000000cc000000cd000000cf000000ce000000d0000000d5000000cf",
            INIT_08 => X"000000a8000000b9000000c80000007f0000001f000000170000001400000017",
            INIT_09 => X"000000b2000000b3000000b2000000b2000000a20000009a0000009e0000009f",
            INIT_0A => X"000000d1000000c500000072000000470000007d000000b6000000be000000b5",
            INIT_0B => X"000000ce000000d0000000d3000000d4000000d3000000d5000000d8000000d5",
            INIT_0C => X"000000a0000000af000000bd0000006300000017000000180000001500000017",
            INIT_0D => X"000000c3000000bf000000ba000000aa00000095000000a6000000a8000000a8",
            INIT_0E => X"000000d6000000d200000092000000630000008d000000bc000000c8000000c3",
            INIT_0F => X"000000d6000000d7000000d9000000d9000000d5000000d4000000d4000000d5",
            INIT_10 => X"00000097000000a5000000aa0000004800000015000000170000001700000019",
            INIT_11 => X"000000bc000000a90000009d000000920000009b000000b9000000b7000000af",
            INIT_12 => X"000000db000000d3000000ac000000790000008d000000b2000000c4000000c5",
            INIT_13 => X"000000ce000000d1000000d4000000d6000000d9000000d9000000d9000000dd",
            INIT_14 => X"0000009a000000a40000008f00000031000000170000001a0000001b0000001a",
            INIT_15 => X"00000097000000800000007d00000082000000a6000000c8000000c2000000a9",
            INIT_16 => X"000000c9000000bc000000b6000000930000008f00000094000000a5000000a5",
            INIT_17 => X"000000d3000000d7000000d7000000dc000000db000000d5000000d9000000d4",
            INIT_18 => X"000000ab000000b40000007d00000025000000190000001b0000001a0000001e",
            INIT_19 => X"000000820000007a000000710000008b000000b3000000ca000000c5000000a9",
            INIT_1A => X"000000c9000000bf000000cb000000b90000008c0000007a0000008500000077",
            INIT_1B => X"000000e0000000dc000000da000000dc000000db000000d7000000da000000d7",
            INIT_1C => X"000000a8000000c1000000af00000064000000240000001f000000300000005e",
            INIT_1D => X"000000840000008e00000091000000ae000000c3000000c6000000c0000000a3",
            INIT_1E => X"000000d5000000bd000000d1000000c00000008b0000007a000000790000006a",
            INIT_1F => X"000000e5000000de000000d5000000d0000000e8000000ef000000ed000000f2",
            INIT_20 => X"000000a0000000be000000be000000b10000007a000000720000009e000000b4",
            INIT_21 => X"00000092000000a7000000b9000000c2000000c8000000c5000000ad00000085",
            INIT_22 => X"000000dc000000bd000000c9000000b10000008d000000850000008100000081",
            INIT_23 => X"000000ea000000e1000000c7000000bd000000d5000000e8000000eb000000f1",
            INIT_24 => X"0000009d000000c5000000c3000000c1000000ba000000b2000000c0000000c5",
            INIT_25 => X"00000097000000b2000000c3000000c1000000bf000000b9000000a300000080",
            INIT_26 => X"000000ea000000d0000000c2000000aa00000086000000830000008100000072",
            INIT_27 => X"000000eb000000d0000000bb000000b9000000c9000000eb000000f0000000ec",
            INIT_28 => X"00000097000000c5000000cd000000c8000000c0000000bb000000c4000000ca",
            INIT_29 => X"00000088000000a8000000bb000000c1000000bd000000b8000000af00000095",
            INIT_2A => X"000000f0000000cd000000b5000000a700000081000000800000008000000075",
            INIT_2B => X"000000dd000000c1000000bb000000ba000000ce000000ee000000f3000000f3",
            INIT_2C => X"000000a0000000c2000000d0000000cb000000c0000000c5000000cd000000cd",
            INIT_2D => X"0000007700000092000000ac000000c1000000bf000000c1000000bf000000a8",
            INIT_2E => X"000000ea000000bf000000b0000000a700000087000000850000008e0000007c",
            INIT_2F => X"000000c4000000b9000000b8000000ba000000d7000000ec000000f1000000f3",
            INIT_30 => X"000000b4000000bf000000c7000000c5000000c1000000c8000000cc000000ce",
            INIT_31 => X"0000008300000098000000ae000000ae000000ad000000b7000000b3000000ac",
            INIT_32 => X"000000e6000000bf000000ac000000a90000009a0000008e000000a60000008d",
            INIT_33 => X"000000c0000000b8000000ba000000c8000000e4000000ef000000f1000000f0",
            INIT_34 => X"000000ca000000b1000000b4000000c9000000bf000000c6000000ca000000d2",
            INIT_35 => X"0000009c00000093000000a8000000a80000008e0000008e0000009a000000ab",
            INIT_36 => X"000000e6000000c5000000a00000009e000000a400000096000000a9000000af",
            INIT_37 => X"000000d7000000c3000000bf000000e2000000f2000000f4000000f1000000f1",
            INIT_38 => X"000000d7000000a1000000aa000000cf000000c0000000c7000000c9000000d3",
            INIT_39 => X"0000007f00000089000000b1000000be000000ac000000ad000000ba000000bd",
            INIT_3A => X"000000ec000000c1000000b0000000af000000a000000096000000ae000000b4",
            INIT_3B => X"000000e1000000d4000000c9000000ef000000fb000000f3000000f2000000f5",
            INIT_3C => X"000000d90000009a000000b5000000d1000000c1000000c5000000c4000000d3",
            INIT_3D => X"00000098000000a6000000ad000000aa000000b9000000c3000000c5000000ce",
            INIT_3E => X"000000cc000000af000000b5000000c000000098000000a6000000b8000000a3",
            INIT_3F => X"000000e2000000e2000000d5000000df000000f7000000f4000000f3000000ee",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000c60000009b000000c4000000c5000000b5000000b4000000c2000000d6",
            INIT_41 => X"000000b2000000ae000000a1000000ad000000b7000000ae000000c0000000d6",
            INIT_42 => X"000000760000009c000000b4000000a700000093000000bd000000a400000080",
            INIT_43 => X"000000e4000000ea000000d6000000ce000000eb000000ef000000d70000009d",
            INIT_44 => X"000000b9000000be000000ca000000b4000000a3000000a6000000c6000000d7",
            INIT_45 => X"000000ad000000b0000000ae000000c1000000d6000000cd000000d2000000cf",
            INIT_46 => X"00000087000000ab000000c8000000a300000099000000bf0000008900000081",
            INIT_47 => X"000000eb000000ef000000d2000000bb000000c1000000b80000009000000074",
            INIT_48 => X"000000c2000000d2000000cb000000b9000000a4000000ae000000cd000000d8",
            INIT_49 => X"000000b3000000be000000cb000000e1000000e2000000da000000d3000000bf",
            INIT_4A => X"000000ac000000aa000000c2000000a70000009e000000a80000007900000097",
            INIT_4B => X"000000ec000000de000000b8000000a2000000a900000099000000830000009a",
            INIT_4C => X"000000d2000000d1000000ca000000c5000000b4000000c0000000d0000000d8",
            INIT_4D => X"000000b5000000cf000000d5000000d1000000cc000000c5000000bd000000ba",
            INIT_4E => X"000000ab0000009c000000ae000000b7000000af0000009200000095000000b2",
            INIT_4F => X"000000cc000000ac000000a0000000a6000000b4000000a900000094000000a3",
            INIT_50 => X"000000ca000000c9000000cb000000bf000000b6000000ca000000d5000000da",
            INIT_51 => X"000000c7000000cf000000c6000000b2000000c0000000c1000000c3000000ca",
            INIT_52 => X"000000a6000000930000009b000000b1000000bb000000a6000000cb000000d3",
            INIT_53 => X"000000a70000009f0000009c0000009c000000af000000b6000000ab000000a7",
            INIT_54 => X"000000c8000000d0000000c8000000b3000000ba000000d1000000d7000000d9",
            INIT_55 => X"000000c2000000c4000000b6000000a1000000ba000000d2000000d7000000d1",
            INIT_56 => X"000000a60000009b0000008e0000009b000000b9000000be000000cf000000cb",
            INIT_57 => X"0000008f0000009e0000009e000000960000009f000000ad000000b3000000ac",
            INIT_58 => X"000000d9000000da000000c5000000a9000000c0000000d6000000d5000000d6",
            INIT_59 => X"000000bf000000c3000000b3000000aa000000c3000000d4000000d9000000d7",
            INIT_5A => X"000000aa000000a70000008e00000084000000aa000000c0000000c0000000be",
            INIT_5B => X"0000007d00000086000000930000009d0000009d000000ad000000b3000000aa",
            INIT_5C => X"000000de000000d8000000c1000000a8000000ca000000d3000000d1000000d5",
            INIT_5D => X"000000c6000000c9000000c2000000c2000000cd000000d3000000de000000df",
            INIT_5E => X"000000a7000000ab0000009b0000008600000099000000bc000000c4000000c6",
            INIT_5F => X"00000089000000850000008e000000a3000000a5000000b2000000bd000000a6",
            INIT_60 => X"000000d5000000d3000000bf000000af000000ca000000ce000000ce000000d3",
            INIT_61 => X"000000c9000000c9000000ce000000c2000000ab000000c6000000d8000000d6",
            INIT_62 => X"0000009d000000a70000009e0000009000000096000000b1000000c5000000c8",
            INIT_63 => X"00000090000000950000009600000098000000a8000000b0000000b50000009f",
            INIT_64 => X"000000d2000000d0000000bc000000b5000000c1000000c9000000cc000000d2",
            INIT_65 => X"000000c2000000c6000000d0000000b10000007a000000a0000000ce000000cd",
            INIT_66 => X"00000099000000a00000009c0000008b00000096000000a6000000b8000000c1",
            INIT_67 => X"000000830000008c00000098000000980000009b0000009f000000a00000009b",
            INIT_68 => X"000000d6000000cd000000b2000000ae000000bb000000c6000000ca000000d2",
            INIT_69 => X"000000b6000000bb000000ca000000b400000083000000a4000000cb000000d1",
            INIT_6A => X"000000900000009a00000099000000860000008b0000009d000000a9000000b6",
            INIT_6B => X"00000093000000960000009b0000009d0000008d000000830000008d00000097",
            INIT_6C => X"000000d7000000c4000000a8000000a8000000b5000000c2000000c8000000d2",
            INIT_6D => X"000000ac000000ad000000b9000000cb000000b8000000bd000000c7000000d4",
            INIT_6E => X"0000008d00000091000000940000008300000076000000930000009b000000a3",
            INIT_6F => X"0000009c000000a2000000a300000095000000850000007f0000008400000090",
            INIT_70 => X"000000d3000000bd0000009e000000a2000000b4000000bd000000c2000000d0",
            INIT_71 => X"000000a4000000a3000000ac000000bf000000c7000000c2000000c5000000d3",
            INIT_72 => X"000000910000009000000090000000890000006d00000082000000930000009e",
            INIT_73 => X"000000930000009f000000a200000097000000860000007c0000008400000090",
            INIT_74 => X"000000cd000000b30000008f0000009f000000b5000000b0000000b1000000c2",
            INIT_75 => X"000000a10000009c000000a5000000b5000000be000000c2000000c7000000d0",
            INIT_76 => X"000000920000008a000000850000008900000072000000700000008800000095",
            INIT_77 => X"0000008d00000094000000950000009600000090000000830000008300000092",
            INIT_78 => X"000000c70000009c00000085000000a7000000b2000000a50000009d000000ac",
            INIT_79 => X"0000008b0000008400000085000000a0000000c2000000c7000000c7000000ce",
            INIT_7A => X"000000950000008a00000081000000820000007e0000006b0000007e0000008c",
            INIT_7B => X"00000098000000950000008c000000880000008e000000910000008c0000008d",
            INIT_7C => X"000000b7000000820000007d0000009e0000009b000000900000008600000097",
            INIT_7D => X"000000690000005e0000006700000080000000a5000000b7000000bf000000c5",
            INIT_7E => X"0000008f0000008b0000007d000000790000007c000000750000007000000077",
            INIT_7F => X"000000960000009b00000095000000840000007d000000810000008c0000008b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY24;


    MEM_IFMAP_LAYER0_ENTITY25 : if BRAM_NAME = "ifmap_layer0_entity25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008e0000009300000093000000830000002f000000100000001500000013",
            INIT_01 => X"0000008f0000008c0000008c0000008d0000008e000000900000008900000087",
            INIT_02 => X"000000a4000000820000005d0000005f00000049000000600000007e0000008c",
            INIT_03 => X"00000097000000980000009b0000009e0000009d0000009b0000009c0000009b",
            INIT_04 => X"000000920000009b000000a10000007a0000001f000000110000001400000014",
            INIT_05 => X"00000097000000920000009600000098000000950000008b000000880000008a",
            INIT_06 => X"000000af0000009c00000058000000410000004900000075000000960000009f",
            INIT_07 => X"000000a3000000a4000000a8000000ac000000ad000000ab000000a9000000a8",
            INIT_08 => X"0000008c00000097000000a20000006600000015000000140000001400000014",
            INIT_09 => X"0000009f00000098000000990000009a0000008b00000088000000950000008d",
            INIT_0A => X"000000b7000000b1000000610000003a0000006d000000a1000000ab000000a6",
            INIT_0B => X"000000a6000000a9000000ad000000b1000000b2000000b1000000b2000000b3",
            INIT_0C => X"000000820000008c000000990000004f00000011000000150000001400000014",
            INIT_0D => X"000000b0000000a9000000a600000099000000870000009d000000a400000097",
            INIT_0E => X"000000c3000000c4000000850000005200000076000000a1000000af000000b0",
            INIT_0F => X"000000ab000000ad000000b1000000b3000000b3000000b4000000b7000000bd",
            INIT_10 => X"0000007700000082000000890000003800000013000000150000001400000015",
            INIT_11 => X"000000a7000000940000008b0000008400000092000000b3000000b20000009c",
            INIT_12 => X"000000d2000000ce000000a70000006d0000007800000098000000a9000000af",
            INIT_13 => X"000000ac000000b1000000b6000000ba000000bf000000c3000000c9000000d1",
            INIT_14 => X"0000007800000082000000730000002600000016000000170000001600000016",
            INIT_15 => X"000000840000006b0000006c000000760000009e000000c3000000b900000092",
            INIT_16 => X"000000c7000000be000000b70000008f00000084000000810000008f00000092",
            INIT_17 => X"000000c2000000c7000000ca000000d1000000d1000000cc000000d1000000cf",
            INIT_18 => X"00000094000000a1000000710000001e00000014000000150000001300000018",
            INIT_19 => X"00000071000000690000006200000080000000aa000000c2000000ba00000097",
            INIT_1A => X"000000c5000000c0000000ca000000b2000000800000006b0000007400000068",
            INIT_1B => X"000000da000000d7000000d6000000d8000000d7000000d1000000cf000000ce",
            INIT_1C => X"0000009c000000ba000000ae000000600000001d000000180000002900000058",
            INIT_1D => X"000000760000008100000084000000a4000000ba000000bd000000b500000095",
            INIT_1E => X"000000ce000000bb000000cc000000b40000007c0000006c0000006b0000005c",
            INIT_1F => X"000000e2000000dc000000d3000000cd000000e4000000e7000000e0000000e6",
            INIT_20 => X"00000093000000b7000000bd000000af000000750000006d00000099000000b1",
            INIT_21 => X"000000830000009a000000ad000000b8000000c0000000bc000000a100000078",
            INIT_22 => X"000000d8000000bc000000c5000000a60000007f000000770000007300000073",
            INIT_23 => X"000000e8000000e0000000c6000000bc000000d3000000e3000000e2000000e9",
            INIT_24 => X"00000090000000be000000c2000000bf000000b6000000af000000bc000000c2",
            INIT_25 => X"0000008a000000a4000000b6000000b7000000b6000000b10000009800000073",
            INIT_26 => X"000000e9000000d0000000bd000000a00000007b000000770000007600000066",
            INIT_27 => X"000000eb000000d1000000bd000000bb000000cb000000ea000000eb000000e8",
            INIT_28 => X"0000008a000000bf000000cd000000c6000000bb000000b7000000c0000000c7",
            INIT_29 => X"0000007c0000009a000000af000000b8000000b5000000b0000000a500000088",
            INIT_2A => X"000000f0000000cd000000b00000009e0000007800000077000000760000006b",
            INIT_2B => X"000000e0000000c6000000c0000000c0000000d4000000f2000000f4000000f3",
            INIT_2C => X"00000092000000bc000000d1000000c9000000bb000000c1000000c9000000c9",
            INIT_2D => X"0000006b000000840000009f000000b7000000b7000000b9000000b60000009b",
            INIT_2E => X"000000eb000000bd000000aa0000009e0000007e0000007c0000008500000073",
            INIT_2F => X"000000ca000000c0000000c0000000c2000000de000000f2000000f6000000f6",
            INIT_30 => X"000000a5000000b7000000c6000000c4000000bd000000c5000000c9000000cb",
            INIT_31 => X"000000780000008a000000a2000000a4000000a5000000b0000000aa0000009f",
            INIT_32 => X"000000e7000000bd000000a5000000a100000092000000870000009f00000085",
            INIT_33 => X"000000c7000000c1000000c3000000d0000000ea000000f7000000f8000000f4",
            INIT_34 => X"000000b90000009c000000a7000000c1000000b9000000c4000000ca000000d0",
            INIT_35 => X"0000008f000000890000009e000000a1000000870000008700000091000000a1",
            INIT_36 => X"000000e4000000c30000009d00000099000000a200000095000000a4000000a4",
            INIT_37 => X"000000de000000cc000000c7000000e8000000f5000000f9000000f7000000f2",
            INIT_38 => X"000000c10000007d0000008e000000bf000000b6000000c5000000cc000000d2",
            INIT_39 => X"0000007200000082000000aa000000b8000000a7000000a6000000b1000000b5",
            INIT_3A => X"000000e7000000bd000000ae000000ab0000009e00000098000000aa000000a5",
            INIT_3B => X"000000e9000000dd000000cf000000f2000000fb000000f5000000f4000000f2",
            INIT_3C => X"000000c00000007000000091000000bd000000b9000000c5000000c8000000d4",
            INIT_3D => X"00000089000000a0000000a7000000a4000000b4000000bd000000be000000c7",
            INIT_3E => X"000000c3000000a8000000b1000000b800000091000000a2000000b000000092",
            INIT_3F => X"000000eb000000ec000000dd000000e4000000f9000000f5000000f1000000e8",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ad0000006e0000009b000000b0000000ae000000b6000000c7000000d8",
            INIT_41 => X"000000a4000000a70000009b000000a8000000b2000000a8000000ba000000d0",
            INIT_42 => X"0000006800000090000000ab0000009a00000086000000b1000000960000006e",
            INIT_43 => X"000000ed000000f3000000dd000000d2000000ed000000ee000000d100000091",
            INIT_44 => X"000000a200000095000000a7000000a30000009e000000a9000000ce000000db",
            INIT_45 => X"000000a1000000aa000000a8000000bc000000d1000000c8000000cd000000ca",
            INIT_46 => X"000000730000009b000000ba0000009300000087000000ad0000007800000070",
            INIT_47 => X"000000ef000000f3000000d4000000b9000000bc000000b20000008400000062",
            INIT_48 => X"000000b1000000b3000000b5000000af000000a1000000b3000000d6000000dd",
            INIT_49 => X"000000ab000000b8000000c5000000dc000000dd000000d4000000cf000000bd",
            INIT_4A => X"0000009300000094000000b1000000970000008c00000095000000670000008b",
            INIT_4B => X"000000ea000000d9000000b1000000970000009c0000008a0000007000000083",
            INIT_4C => X"000000c8000000be000000c2000000c2000000b2000000c6000000da000000df",
            INIT_4D => X"000000b1000000c8000000d0000000cb000000c7000000bf000000b8000000ba",
            INIT_4E => X"0000008f000000830000009b000000a80000009e0000007f00000087000000ab",
            INIT_4F => X"000000c50000009e00000090000000930000009f000000940000007e00000089",
            INIT_50 => X"000000c2000000be000000c7000000bf000000b7000000d0000000dd000000e1",
            INIT_51 => X"000000bf000000c6000000c1000000ab000000ba000000be000000bc000000c6",
            INIT_52 => X"0000008d0000007b00000087000000a0000000a900000094000000bf000000cf",
            INIT_53 => X"0000009a0000008c0000008800000087000000980000009f000000950000008e",
            INIT_54 => X"000000be000000c8000000c3000000b3000000be000000d6000000dd000000de",
            INIT_55 => X"000000b5000000b6000000b300000097000000b2000000d1000000cd000000c6",
            INIT_56 => X"00000093000000890000007c00000086000000a5000000ae000000c4000000c5",
            INIT_57 => X"0000007d0000008b0000008b000000830000008b00000099000000a100000099",
            INIT_58 => X"000000cf000000d2000000bf000000aa000000c6000000db000000da000000db",
            INIT_59 => X"000000b0000000b4000000ae0000009c000000b4000000cf000000ce000000cb",
            INIT_5A => X"00000098000000960000007d0000006f00000096000000b0000000b5000000b6",
            INIT_5B => X"0000006a00000073000000800000008a0000008a0000009a000000a100000098",
            INIT_5C => X"000000d5000000d2000000bc000000aa000000cf000000d9000000d6000000da",
            INIT_5D => X"000000b5000000ba000000ba000000ae000000b6000000c7000000d3000000d4",
            INIT_5E => X"000000950000009a000000890000007200000085000000ab000000b6000000ba",
            INIT_5F => X"00000076000000730000007b00000090000000920000009f000000ab00000094",
            INIT_60 => X"000000cd000000cf000000bd000000b3000000d1000000d4000000d4000000d8",
            INIT_61 => X"000000b6000000bb000000c3000000a70000008a000000b1000000cd000000cd",
            INIT_62 => X"0000008c000000960000008d0000007d000000820000009e000000b5000000b9",
            INIT_63 => X"0000007c000000820000008300000085000000950000009d000000a30000008d",
            INIT_64 => X"000000cc000000ce000000be000000bb000000c8000000d0000000d2000000d7",
            INIT_65 => X"000000ae000000b8000000c2000000910000005000000083000000c4000000c6",
            INIT_66 => X"000000880000008f0000008b000000780000008300000093000000a5000000ae",
            INIT_67 => X"00000070000000790000008500000085000000880000008c0000008e00000089",
            INIT_68 => X"000000d1000000cd000000b7000000b5000000c2000000cd000000d0000000d7",
            INIT_69 => X"000000a1000000ab000000ba0000008e0000005100000081000000c2000000cc",
            INIT_6A => X"0000007e000000890000008700000073000000780000008900000095000000a1",
            INIT_6B => X"0000008000000083000000880000008a0000007a000000700000007b00000085",
            INIT_6C => X"000000d4000000c6000000af000000b0000000bc000000c8000000cd000000d6",
            INIT_6D => X"000000950000009b000000a8000000aa0000008e000000a0000000c0000000d0",
            INIT_6E => X"0000007b000000800000008300000071000000640000007f000000850000008d",
            INIT_6F => X"00000089000000900000009000000082000000720000006c000000720000007e",
            INIT_70 => X"000000d2000000c0000000a6000000a9000000b7000000c0000000c4000000d2",
            INIT_71 => X"0000008c0000008d00000099000000ab000000b4000000b6000000c0000000d1",
            INIT_72 => X"0000007f0000007e0000007e000000780000005c0000006f0000007d00000086",
            INIT_73 => X"000000810000008d00000090000000850000007400000069000000720000007e",
            INIT_74 => X"000000cc000000b500000097000000a6000000b9000000b3000000b3000000c4",
            INIT_75 => X"000000880000008500000092000000a6000000b3000000ba000000c2000000cd",
            INIT_76 => X"00000080000000780000007300000078000000610000005d000000720000007e",
            INIT_77 => X"0000007b0000008200000083000000840000007e000000710000007100000080",
            INIT_78 => X"000000c30000009c0000008c000000ae000000b8000000aa000000a1000000b1",
            INIT_79 => X"000000730000006c0000007100000091000000b6000000bf000000c1000000c9",
            INIT_7A => X"000000830000007800000070000000720000006e000000590000006a00000076",
            INIT_7B => X"00000086000000820000007a000000750000007c0000007f0000007a0000007b",
            INIT_7C => X"000000b10000008000000082000000a6000000a1000000970000008c0000009d",
            INIT_7D => X"000000530000004700000053000000700000009a000000af000000b7000000bf",
            INIT_7E => X"0000007e000000790000006c0000006c0000006e000000650000005e00000063",
            INIT_7F => X"000000840000008900000084000000730000006b0000006f0000007a00000079",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY25;


    MEM_IFMAP_LAYER0_ENTITY26 : if BRAM_NAME = "ifmap_layer0_entity26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000740000006d000000730000007100000028000000130000001c00000017",
            INIT_01 => X"0000006b000000690000006900000069000000690000006a0000006700000071",
            INIT_02 => X"000000890000007200000056000000540000003a0000004c000000630000006a",
            INIT_03 => X"000000780000007a0000007d0000007f0000007d0000007c0000007d0000007c",
            INIT_04 => X"0000007c00000076000000820000006a0000001a000000140000001b00000018",
            INIT_05 => X"00000079000000720000007600000078000000750000006d000000720000007d",
            INIT_06 => X"000000960000008c000000510000003e000000440000006a0000008300000085",
            INIT_07 => X"0000008000000081000000850000008800000088000000890000008c0000008a",
            INIT_08 => X"0000007b00000074000000830000005800000012000000170000001a00000018",
            INIT_09 => X"000000840000007d0000007f0000008100000074000000740000008d0000008b",
            INIT_0A => X"0000009e0000009f000000590000003700000069000000980000009a0000008e",
            INIT_0B => X"00000084000000880000008b0000008e0000008e000000920000009700000097",
            INIT_0C => X"000000730000006a0000007c0000004500000012000000190000001900000018",
            INIT_0D => X"000000970000009500000094000000890000007800000092000000a60000009c",
            INIT_0E => X"000000a9000000b10000007a0000004a0000006d000000940000009c00000096",
            INIT_0F => X"0000008e00000091000000940000009600000095000000980000009d000000a1",
            INIT_10 => X"00000068000000600000006d0000003300000017000000190000001800000019",
            INIT_11 => X"0000009300000086000000800000007c0000008d000000b2000000b8000000a1",
            INIT_12 => X"000000b5000000b700000098000000600000006c000000890000009600000097",
            INIT_13 => X"00000093000000980000009c000000a0000000a4000000a8000000ae000000b3",
            INIT_14 => X"000000660000005f00000059000000230000001c0000001b0000001a0000001a",
            INIT_15 => X"000000760000006200000066000000740000009f000000c7000000c100000096",
            INIT_16 => X"000000aa000000a6000000a7000000840000007a000000770000008300000082",
            INIT_17 => X"000000a9000000af000000b1000000b7000000b7000000b3000000b7000000b2",
            INIT_18 => X"0000007b000000800000005c0000001d0000001a00000019000000160000001a",
            INIT_19 => X"0000006a000000630000005e0000007e000000ab000000c7000000c300000093",
            INIT_1A => X"000000b0000000aa000000c0000000ac0000007a000000650000006d00000060",
            INIT_1B => X"000000c2000000bf000000bf000000c5000000ca000000c5000000c4000000c3",
            INIT_1C => X"0000007e0000009b0000009a000000580000001900000011000000210000004d",
            INIT_1D => X"000000710000007b00000081000000a3000000b9000000c1000000be0000008c",
            INIT_1E => X"000000bd000000a5000000c6000000b100000079000000680000006700000058",
            INIT_1F => X"000000cd000000c4000000bb000000ba000000da000000e0000000db000000e4",
            INIT_20 => X"0000007700000099000000a70000009b00000060000000560000008000000095",
            INIT_21 => X"0000007f00000094000000aa000000b7000000bf000000bf000000a80000006f",
            INIT_22 => X"000000c1000000a2000000bb000000a30000007c000000740000007000000070",
            INIT_23 => X"000000d2000000c4000000a60000009d000000bb000000cf000000d5000000df",
            INIT_24 => X"000000750000009f000000a9000000a70000009b000000920000009e000000a1",
            INIT_25 => X"000000870000009f000000b4000000b6000000b5000000b30000009b00000068",
            INIT_26 => X"000000cc000000b2000000b20000009e00000079000000750000007400000064",
            INIT_27 => X"000000cf000000b00000009600000093000000a7000000cb000000d6000000d8",
            INIT_28 => X"00000070000000a0000000b0000000af000000a50000009e000000a5000000aa",
            INIT_29 => X"0000007900000095000000ac000000b6000000b4000000b1000000a40000007b",
            INIT_2A => X"000000d1000000af000000a60000009c0000007600000075000000740000006a",
            INIT_2B => X"000000ba0000009f0000009300000091000000a9000000cd000000d8000000de",
            INIT_2C => X"0000007a0000009d000000b0000000b0000000a6000000a9000000ae000000ac",
            INIT_2D => X"000000680000007f0000009d000000b6000000b6000000b9000000b10000008d",
            INIT_2E => X"000000ce000000a3000000a40000009f0000007d0000007b0000008400000073",
            INIT_2F => X"0000009c000000930000008e00000092000000b5000000cd000000d9000000e0",
            INIT_30 => X"0000008f00000099000000a4000000a5000000a0000000a5000000a7000000a7",
            INIT_31 => X"00000076000000850000009f000000a3000000a4000000ae000000a300000091",
            INIT_32 => X"000000cd000000a8000000a3000000a300000092000000870000009f00000086",
            INIT_33 => X"000000980000009000000090000000a3000000c7000000d6000000dc000000df",
            INIT_34 => X"000000a40000008300000088000000a30000009b000000a0000000a2000000a9",
            INIT_35 => X"00000092000000870000009e0000009f00000085000000840000008800000092",
            INIT_36 => X"000000cb000000b000000098000000980000009e00000090000000a2000000a7",
            INIT_37 => X"000000b6000000a20000009f000000c5000000da000000dd000000d8000000d7",
            INIT_38 => X"000000b20000006d00000078000000a80000009d000000a2000000a4000000ae",
            INIT_39 => X"0000007800000084000000ab000000b6000000a3000000a1000000a7000000a6",
            INIT_3A => X"000000cc000000aa000000a4000000a6000000950000008c000000a3000000a9",
            INIT_3B => X"000000c7000000bb000000b0000000d6000000e4000000da000000d5000000d3",
            INIT_3C => X"000000b70000006800000084000000aa0000009f000000a1000000a0000000af",
            INIT_3D => X"0000008d000000a3000000a8000000a2000000b0000000b8000000b6000000bc",
            INIT_3E => X"000000a900000096000000a5000000af0000008500000092000000a500000091",
            INIT_3F => X"000000c7000000c7000000ba000000c4000000dd000000d9000000d4000000ca",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a80000006d00000097000000a100000094000000920000009f000000b3",
            INIT_41 => X"000000a6000000aa0000009c000000a5000000ae000000a4000000b5000000c7",
            INIT_42 => X"000000500000007e0000009e0000008f000000770000009f0000008800000069",
            INIT_43 => X"000000c5000000c9000000b7000000af000000cd000000d1000000b700000076",
            INIT_44 => X"0000009f00000097000000a5000000950000008300000085000000a4000000b5",
            INIT_45 => X"000000a2000000ac000000a8000000b9000000cd000000c4000000c7000000c2",
            INIT_46 => X"0000005c00000088000000ad00000086000000770000009b0000006900000068",
            INIT_47 => X"000000c8000000cb000000b0000000980000009e000000980000006f0000004b",
            INIT_48 => X"000000aa000000b1000000b00000009f000000850000008e000000ac000000b7",
            INIT_49 => X"000000aa000000bb000000c6000000d9000000d9000000cf000000c5000000b1",
            INIT_4A => X"0000007e00000082000000a20000008b0000007e000000850000005a00000083",
            INIT_4B => X"000000c7000000b8000000920000007c0000008400000076000000600000006f",
            INIT_4C => X"000000bc000000b6000000b7000000af00000095000000a1000000b0000000b9",
            INIT_4D => X"000000af000000ca000000d0000000c9000000c2000000b9000000aa000000aa",
            INIT_4E => X"0000007b000000710000008c0000009d00000091000000710000007b000000a4",
            INIT_4F => X"000000a600000084000000790000007f0000008e000000860000007000000077",
            INIT_50 => X"000000b2000000b1000000ba000000ab0000009b000000ad000000b7000000bd",
            INIT_51 => X"000000bd000000c3000000bc000000a4000000b1000000b2000000ac000000b4",
            INIT_52 => X"0000007c0000006a00000078000000930000009d00000088000000b6000000c9",
            INIT_53 => X"000000820000007a00000077000000780000008a000000940000008a00000080",
            INIT_54 => X"000000b0000000bb000000b70000009e000000a1000000b7000000bc000000bd",
            INIT_55 => X"000000b1000000ad000000a60000008b000000a4000000c0000000bf000000b8",
            INIT_56 => X"00000085000000790000006b0000007600000096000000a2000000bc000000c0",
            INIT_57 => X"0000006c0000007d0000007c000000750000007d0000008d000000960000008e",
            INIT_58 => X"000000c5000000c7000000b400000094000000a6000000bb000000ba000000ba",
            INIT_59 => X"000000aa000000a90000009f00000091000000a8000000c0000000c3000000c1",
            INIT_5A => X"0000008b000000860000006c0000005d00000086000000a3000000ac000000af",
            INIT_5B => X"0000005b00000065000000720000007c0000007c0000008e000000970000008d",
            INIT_5C => X"000000cf000000c9000000b00000008f000000ac000000b7000000b5000000ba",
            INIT_5D => X"000000ac000000ae000000ab000000a5000000af000000bd000000cb000000ce",
            INIT_5E => X"000000880000008a0000007800000061000000750000009e000000ab000000b2",
            INIT_5F => X"00000068000000640000006d000000820000008400000092000000a10000008a",
            INIT_60 => X"000000ca000000c6000000aa00000092000000a9000000af000000b2000000b8",
            INIT_61 => X"000000aa000000ab000000b4000000a100000088000000ab000000c5000000c8",
            INIT_62 => X"0000007e000000860000007c0000006c0000007300000090000000a8000000ad",
            INIT_63 => X"0000006f00000074000000750000007700000087000000910000009900000082",
            INIT_64 => X"000000c8000000c0000000a2000000930000009d000000a8000000b0000000b8",
            INIT_65 => X"0000009f000000a6000000b30000008d0000005200000081000000b9000000bf",
            INIT_66 => X"0000007a0000007f0000007a000000690000007400000084000000960000009f",
            INIT_67 => X"000000620000006b00000077000000770000007a00000080000000840000007f",
            INIT_68 => X"000000ca000000ba000000920000008600000094000000a3000000ac000000b8",
            INIT_69 => X"0000009000000098000000ac0000008c0000005800000082000000b2000000c0",
            INIT_6A => X"00000070000000790000007700000064000000690000007a0000008400000091",
            INIT_6B => X"00000072000000750000007a0000007c0000006c00000064000000710000007a",
            INIT_6C => X"000000cc000000b2000000840000007e0000008e0000009e000000a9000000b7",
            INIT_6D => X"000000830000008700000098000000a4000000900000009d000000af000000c3",
            INIT_6E => X"0000006d000000710000007300000061000000540000006f000000740000007c",
            INIT_6F => X"0000007b000000820000008200000074000000640000005f0000006600000072",
            INIT_70 => X"000000cc000000b20000007a000000770000008e00000099000000a1000000b1",
            INIT_71 => X"0000007b0000007a000000870000009d000000a8000000aa000000b4000000c5",
            INIT_72 => X"00000071000000700000006f000000680000004b0000005e0000006d00000077",
            INIT_73 => X"000000730000007e0000008200000077000000660000005c0000006400000070",
            INIT_74 => X"000000c8000000a90000006b00000074000000910000008d00000090000000a3",
            INIT_75 => X"00000079000000730000008100000096000000a3000000ac000000b7000000c2",
            INIT_76 => X"000000720000006a0000006500000068000000510000004e0000006400000070",
            INIT_77 => X"0000006e00000074000000750000007600000070000000630000006300000072",
            INIT_78 => X"000000c0000000910000005f0000007c0000008f000000830000007e0000008e",
            INIT_79 => X"000000650000005c0000006200000082000000a8000000b2000000b7000000be",
            INIT_7A => X"000000740000006a00000061000000630000005f0000004b0000005c00000068",
            INIT_7B => X"00000077000000740000006c000000670000006e000000710000006c0000006d",
            INIT_7C => X"000000ae0000007600000057000000740000007800000070000000680000007b",
            INIT_7D => X"000000460000003900000045000000630000008d000000a4000000ae000000b5",
            INIT_7E => X"000000700000006b0000005e0000005d00000060000000580000005100000057",
            INIT_7F => X"000000760000007b00000076000000650000005d000000610000006c0000006b",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY26;


    MEM_IFMAP_LAYER0_ENTITY27 : if BRAM_NAME = "ifmap_layer0_entity27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bd000000cf000000d6000000da000000c7000000cd000000d2000000d9",
            INIT_01 => X"0000008f0000008c0000009a00000096000000a9000000a6000000ae000000bb",
            INIT_02 => X"000000e1000000e2000000d7000000db000000df000000db000000bf000000a7",
            INIT_03 => X"000000a2000000a1000000aa000000c8000000bb000000af000000be000000db",
            INIT_04 => X"000000b3000000d3000000e1000000d8000000d7000000dc000000dd000000de",
            INIT_05 => X"000000db000000d1000000ce000000c7000000bc000000be000000c0000000b4",
            INIT_06 => X"000000e5000000e1000000e2000000e9000000ec000000ec000000eb000000e5",
            INIT_07 => X"000000c8000000ba000000b7000000d8000000cd000000d0000000d4000000e7",
            INIT_08 => X"000000ad000000d9000000ef000000e9000000e8000000e7000000e9000000ea",
            INIT_09 => X"000000e0000000d4000000bc000000be000000b7000000ad000000b4000000a4",
            INIT_0A => X"000000e1000000d6000000df000000e5000000e1000000e3000000eb000000da",
            INIT_0B => X"000000d3000000d0000000ca000000d1000000d8000000e6000000e8000000ea",
            INIT_0C => X"0000009e000000e4000000f3000000f4000000f2000000f4000000f4000000f5",
            INIT_0D => X"0000009f000000a200000088000000910000009f000000830000009d00000092",
            INIT_0E => X"000000e2000000d0000000cb000000d1000000d3000000c3000000cb000000a9",
            INIT_0F => X"000000d4000000e0000000db000000c7000000d5000000e4000000e9000000e6",
            INIT_10 => X"00000075000000cf000000f1000000f5000000f4000000f4000000f3000000f5",
            INIT_11 => X"0000005c000000640000005b000000640000006b000000590000006c00000063",
            INIT_12 => X"000000e9000000ca000000b9000000b6000000950000007c0000007c00000066",
            INIT_13 => X"000000de000000e2000000d5000000c2000000cd000000e3000000e2000000e1",
            INIT_14 => X"0000007e000000d8000000ed000000f5000000f3000000f4000000f4000000f5",
            INIT_15 => X"000000630000006b0000006700000065000000660000005b0000005a00000048",
            INIT_16 => X"000000eb000000d8000000be0000007e0000005d0000005b0000005900000059",
            INIT_17 => X"000000ec000000d9000000bd000000ae000000c4000000d8000000df000000e7",
            INIT_18 => X"0000009e000000d9000000db000000f1000000f4000000f3000000f3000000f5",
            INIT_19 => X"0000008a0000008f000000840000008c00000097000000840000007200000050",
            INIT_1A => X"000000e9000000dd0000009b0000006e00000078000000720000007a00000082",
            INIT_1B => X"000000eb000000cc000000ab000000a7000000c0000000c6000000e0000000eb",
            INIT_1C => X"00000099000000d7000000c7000000e3000000f6000000f3000000f3000000f4",
            INIT_1D => X"00000083000000830000009e000000cf000000ca000000bb0000009200000051",
            INIT_1E => X"000000d70000009f000000840000009f00000084000000830000008d00000081",
            INIT_1F => X"000000dd000000b2000000ab000000c5000000d1000000d4000000d7000000e5",
            INIT_20 => X"00000082000000da000000ce000000e3000000f5000000f4000000f3000000f4",
            INIT_21 => X"0000007d0000007400000091000000b800000081000000800000008200000051",
            INIT_22 => X"000000c60000009000000093000000990000007d0000008e000000890000007c",
            INIT_23 => X"000000c9000000a9000000a4000000b8000000dc000000e9000000db000000d6",
            INIT_24 => X"0000006e000000a8000000be000000e4000000f2000000f4000000f3000000f3",
            INIT_25 => X"0000007800000073000000800000008f0000006e000000770000008600000053",
            INIT_26 => X"000000c40000008c0000009b000000950000007d00000092000000830000007d",
            INIT_27 => X"000000dc000000d7000000c8000000c8000000e9000000f0000000f0000000e9",
            INIT_28 => X"0000005f0000008200000085000000dc000000f5000000f4000000f1000000ef",
            INIT_29 => X"0000006c0000006d0000006b0000006d0000006c00000074000000740000004e",
            INIT_2A => X"000000a70000008f000000960000008800000073000000780000007800000073",
            INIT_2B => X"000000f4000000f5000000f5000000f4000000f3000000f5000000e4000000d0",
            INIT_2C => X"00000059000000a5000000a9000000d8000000f4000000f2000000e9000000de",
            INIT_2D => X"00000060000000620000005f0000005f000000640000005b000000430000003d",
            INIT_2E => X"0000007e000000810000007900000069000000610000005a0000005f00000060",
            INIT_2F => X"000000f4000000f4000000f4000000f4000000f3000000f8000000d80000009b",
            INIT_30 => X"00000064000000b5000000b7000000bf000000e3000000ec000000df000000d0",
            INIT_31 => X"0000005400000056000000630000006f00000065000000580000003800000037",
            INIT_32 => X"0000008100000070000000620000006d000000710000005d0000005400000052",
            INIT_33 => X"000000f4000000f4000000f4000000f4000000f4000000f5000000e2000000ae",
            INIT_34 => X"000000660000009c0000009a000000aa000000c3000000db000000cc000000c8",
            INIT_35 => X"000000550000005e0000007500000073000000660000006c0000006300000068",
            INIT_36 => X"0000007c0000006c00000068000000800000008c0000007a0000006a0000005a",
            INIT_37 => X"000000f4000000f4000000f5000000ef000000d4000000c3000000b300000096",
            INIT_38 => X"0000008a0000009300000094000000a4000000a9000000cf000000d2000000c8",
            INIT_39 => X"0000004d000000540000005d000000590000005d0000006a0000005c00000081",
            INIT_3A => X"000000520000004b0000004a0000004f0000005100000051000000510000004c",
            INIT_3B => X"000000f4000000f4000000f4000000bf0000008f0000008c0000007b00000065",
            INIT_3C => X"000000c0000000ba000000960000007000000077000000c4000000e2000000d2",
            INIT_3D => X"0000003f0000003c0000002f0000002d000000370000004d0000004d0000006c",
            INIT_3E => X"000000400000003d0000003200000031000000360000003b0000003f0000003b",
            INIT_3F => X"000000f4000000f6000000e100000087000000670000005b0000004b00000047",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a1000000c0000000910000005d00000060000000b4000000c1000000c7",
            INIT_41 => X"000000470000004f0000004f00000068000000620000005c0000004900000056",
            INIT_42 => X"0000001c0000001600000032000000340000001b0000001e0000001c00000025",
            INIT_43 => X"000000f3000000f7000000ce00000080000000680000005b0000003500000018",
            INIT_44 => X"000000470000009f0000009d0000007800000071000000c2000000c7000000d3",
            INIT_45 => X"000000660000008000000079000000950000007c000000740000005a00000044",
            INIT_46 => X"000000630000005c00000093000000940000006400000070000000620000004e",
            INIT_47 => X"000000f5000000f2000000b70000009c0000008e000000870000006c0000005e",
            INIT_48 => X"0000001e00000084000000a50000006e00000066000000b7000000ca000000dc",
            INIT_49 => X"00000064000000810000006500000052000000530000006b0000006200000039",
            INIT_4A => X"000000a3000000a2000000a8000000ac0000009f0000009e000000ae00000099",
            INIT_4B => X"000000f7000000e40000008700000072000000770000009c000000af000000a0",
            INIT_4C => X"0000002a0000006f0000008d0000005300000062000000bc000000cf000000db",
            INIT_4D => X"0000005d0000004000000038000000350000003e0000004c000000480000003a",
            INIT_4E => X"00000067000000670000006b00000074000000650000005b0000007c000000a0",
            INIT_4F => X"000000f8000000d90000007600000051000000430000007e0000009b00000063",
            INIT_50 => X"0000003c0000005d000000580000003800000065000000c7000000d2000000d9",
            INIT_51 => X"0000004100000040000000360000003c000000460000003f0000002e00000038",
            INIT_52 => X"000000610000005d000000600000006400000067000000690000007200000063",
            INIT_53 => X"000000f9000000d4000000720000005200000049000000640000006f00000066",
            INIT_54 => X"0000004400000051000000460000005300000075000000ca000000cd000000d1",
            INIT_55 => X"0000003f000000570000004d00000044000000330000002b0000002300000032",
            INIT_56 => X"0000005d0000003e000000430000004000000048000000520000004700000034",
            INIT_57 => X"000000fa000000cc0000006c000000700000006c000000530000003c00000058",
            INIT_58 => X"00000049000000470000006f0000005d00000068000000c5000000ca000000cd",
            INIT_59 => X"0000004f0000008e000000630000004b0000002200000026000000290000003f",
            INIT_5A => X"000000990000006600000072000000630000007600000093000000560000001e",
            INIT_5B => X"000000f6000000c30000005a000000770000008d0000004a0000003f000000b2",
            INIT_5C => X"00000063000000610000006c0000003100000057000000b9000000c2000000c6",
            INIT_5D => X"000000370000005700000032000000280000002400000027000000330000005f",
            INIT_5E => X"0000009c00000074000000880000007a0000007f000000970000004f00000020",
            INIT_5F => X"000000f0000000c20000004e0000003e0000004a00000035000000370000009f",
            INIT_60 => X"000000900000006c0000003b000000250000004d000000a9000000b4000000b6",
            INIT_61 => X"000000210000001e0000001c0000001d000000200000002b0000003c0000006a",
            INIT_62 => X"000000750000007a000000790000006a000000580000003a0000002a00000027",
            INIT_63 => X"000000e1000000ba000000500000003300000032000000330000002f00000043",
            INIT_64 => X"0000008d0000006f000000600000005b0000007d000000a4000000a5000000a8",
            INIT_65 => X"0000001f0000001d0000001e0000001e00000024000000370000004a00000060",
            INIT_66 => X"000000b5000000b3000000cb000000cd000000ae000000400000001800000023",
            INIT_67 => X"000000d3000000ae0000005b00000042000000300000002b0000002600000057",
            INIT_68 => X"0000008d0000006c0000007600000098000000b4000000af000000a3000000a2",
            INIT_69 => X"0000001d000000190000001800000019000000300000004e000000530000005b",
            INIT_6A => X"000000a6000000a9000000b1000000b8000000a4000000470000002600000027",
            INIT_6B => X"000000ce000000a90000005f0000004e000000310000001e0000001e00000051",
            INIT_6C => X"00000092000000670000007500000092000000a6000000b3000000ac0000009a",
            INIT_6D => X"00000025000000210000001e0000002000000036000000520000005500000057",
            INIT_6E => X"000000890000008e000000790000006b00000065000000560000004d00000036",
            INIT_6F => X"000000c7000000a50000005b0000004e00000036000000210000001e0000003c",
            INIT_70 => X"0000007100000067000000850000008f000000940000009e000000a9000000a6",
            INIT_71 => X"0000002c0000002a000000270000002a0000003c0000004b000000510000004f",
            INIT_72 => X"0000008b000000830000006e0000005a0000004d000000410000003600000030",
            INIT_73 => X"000000c4000000a90000005b0000004600000036000000260000001d00000035",
            INIT_74 => X"0000004e0000006b00000085000000890000008d0000009300000097000000a2",
            INIT_75 => X"000000300000002e0000002a000000320000003c000000460000004e00000048",
            INIT_76 => X"0000007100000065000000590000004c000000420000003b0000003300000031",
            INIT_77 => X"000000ba000000ae000000620000003f00000034000000230000001d00000045",
            INIT_78 => X"0000003c0000006a0000008c0000008f0000008c0000008e0000008d00000094",
            INIT_79 => X"0000003a00000036000000340000003900000037000000420000004a00000042",
            INIT_7A => X"0000005d00000057000000500000004900000046000000410000003a0000003a",
            INIT_7B => X"000000b4000000b3000000830000004a0000003700000026000000250000004d",
            INIT_7C => X"0000003d0000007e000000920000009e000000a2000000a00000009500000090",
            INIT_7D => X"00000048000000490000004500000046000000430000003a0000003900000039",
            INIT_7E => X"0000006100000063000000610000005e00000062000000590000004900000044",
            INIT_7F => X"000000ba000000b6000000a40000007700000047000000400000004500000052",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY27;


    MEM_IFMAP_LAYER0_ENTITY28 : if BRAM_NAME = "ifmap_layer0_entity28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b9000000ca000000d1000000d7000000ca000000d0000000d0000000d7",
            INIT_01 => X"0000009d0000009a000000a70000009d000000a000000098000000a8000000b8",
            INIT_02 => X"000000e4000000e5000000db000000de000000e1000000e1000000cb000000b5",
            INIT_03 => X"000000a5000000b0000000b8000000d0000000c4000000b8000000c5000000dd",
            INIT_04 => X"000000ab000000cc000000dd000000d5000000d9000000e1000000e0000000e2",
            INIT_05 => X"000000e0000000d0000000cd000000c4000000b1000000b2000000bd000000b4",
            INIT_06 => X"000000e7000000e4000000e5000000ee000000f3000000f2000000f0000000ec",
            INIT_07 => X"000000c5000000bf000000be000000de000000d2000000d4000000d6000000e7",
            INIT_08 => X"000000a6000000d6000000ef000000ea000000eb000000ea000000ea000000eb",
            INIT_09 => X"000000df000000ce000000b7000000b8000000b1000000a8000000b1000000a6",
            INIT_0A => X"000000e0000000d9000000e4000000eb000000e8000000e3000000ec000000dc",
            INIT_0B => X"000000d2000000d1000000ce000000d9000000dd000000e6000000e9000000e9",
            INIT_0C => X"00000099000000e3000000f4000000f4000000f3000000f4000000f4000000f5",
            INIT_0D => X"000000a0000000a20000008a000000900000009f000000820000009b00000092",
            INIT_0E => X"000000e0000000d3000000d3000000de000000dc000000c2000000cd000000ac",
            INIT_0F => X"000000d4000000e2000000df000000cf000000db000000e5000000e9000000e6",
            INIT_10 => X"00000070000000cd000000f0000000f5000000f4000000f4000000f4000000f5",
            INIT_11 => X"0000005c000000640000005c000000650000006d0000005b0000006d00000062",
            INIT_12 => X"000000e3000000c9000000c2000000c20000009a0000007c0000007d00000068",
            INIT_13 => X"000000e1000000e8000000dc000000cb000000d3000000e3000000de000000dc",
            INIT_14 => X"0000007b000000d4000000eb000000f6000000f3000000f4000000f4000000f5",
            INIT_15 => X"000000660000006e0000006a00000067000000690000005f0000005d00000047",
            INIT_16 => X"000000e6000000d9000000c5000000810000005d0000005b000000590000005b",
            INIT_17 => X"000000ed000000e2000000c5000000b4000000c6000000d6000000da000000dd",
            INIT_18 => X"0000009c000000d5000000d6000000f0000000f4000000f3000000f3000000f5",
            INIT_19 => X"000000960000009b0000008b000000900000009a00000089000000770000004f",
            INIT_1A => X"000000e9000000e1000000a0000000720000007e00000079000000800000008e",
            INIT_1B => X"000000ec000000d4000000b0000000a5000000ba000000c0000000da000000e9",
            INIT_1C => X"00000096000000d3000000c1000000e2000000f7000000f3000000f3000000f4",
            INIT_1D => X"000000900000008d000000a5000000cd000000c8000000bc0000009800000051",
            INIT_1E => X"000000d6000000a30000008c000000a70000008f0000008d000000960000008e",
            INIT_1F => X"000000dc000000af000000ae000000c7000000d2000000d3000000d1000000e0",
            INIT_20 => X"0000007f000000d8000000ca000000e1000000f5000000f4000000f3000000f4",
            INIT_21 => X"000000870000007c00000097000000b900000087000000840000008600000051",
            INIT_22 => X"000000c00000008e0000009e000000a400000088000000960000009100000086",
            INIT_23 => X"000000c40000009c0000009e000000b1000000d7000000e7000000d8000000cf",
            INIT_24 => X"0000006e000000a8000000bd000000e3000000f2000000f4000000f2000000f2",
            INIT_25 => X"000000810000007c000000870000009300000076000000800000008c00000053",
            INIT_26 => X"000000c100000091000000a40000009e00000086000000970000008b00000085",
            INIT_27 => X"000000d7000000cc000000be000000c1000000e6000000ef000000ef000000e5",
            INIT_28 => X"0000005e0000008000000081000000da000000f4000000f3000000ef000000e8",
            INIT_29 => X"00000073000000730000007000000071000000700000007a0000007a0000004f",
            INIT_2A => X"000000aa000000990000009e000000900000007e0000007f000000800000007c",
            INIT_2B => X"000000f4000000f5000000f3000000f3000000f4000000f6000000e3000000ce",
            INIT_2C => X"000000580000009f000000a1000000d3000000f2000000f2000000e3000000cd",
            INIT_2D => X"00000066000000670000006100000062000000660000005e000000450000003c",
            INIT_2E => X"00000080000000890000007f00000071000000670000005f0000006400000068",
            INIT_2F => X"000000f4000000f4000000f4000000f4000000f3000000f8000000d700000099",
            INIT_30 => X"00000063000000ad000000aa000000b4000000dc000000e4000000d5000000bc",
            INIT_31 => X"00000055000000580000006700000072000000660000005a0000003900000037",
            INIT_32 => X"00000086000000760000006500000070000000730000005d0000005500000055",
            INIT_33 => X"000000f4000000f4000000f4000000f4000000f4000000f5000000e1000000b0",
            INIT_34 => X"000000630000008d0000008600000098000000b5000000ca000000bc000000b8",
            INIT_35 => X"00000056000000600000007800000076000000670000006f0000006600000067",
            INIT_36 => X"0000007f0000006e0000006a00000084000000920000007d0000006b0000005c",
            INIT_37 => X"000000f4000000f4000000f5000000ee000000d2000000c3000000b300000098",
            INIT_38 => X"0000007e0000007f0000007b0000009200000098000000bd000000c2000000b6",
            INIT_39 => X"0000004f000000550000005d0000005a0000005e000000690000005d0000007c",
            INIT_3A => X"000000530000004c0000004b000000510000005500000054000000530000004e",
            INIT_3B => X"000000f4000000f4000000f4000000bc0000008a0000008a0000007a00000065",
            INIT_3C => X"000000ae000000a90000007d0000006500000065000000a7000000cc000000bd",
            INIT_3D => X"0000003e0000003b0000002f0000002b000000360000004f0000004d00000067",
            INIT_3E => X"000000400000003d000000300000002f00000034000000390000003e0000003b",
            INIT_3F => X"000000f4000000f6000000df00000080000000610000005a0000004a00000046",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000092000000ac0000007c000000520000005400000097000000a4000000ae",
            INIT_41 => X"000000440000004c0000004b000000640000005a000000570000004900000053",
            INIT_42 => X"00000019000000140000002f00000030000000170000001a0000001700000021",
            INIT_43 => X"000000f3000000f7000000ca0000007800000064000000560000003200000015",
            INIT_44 => X"000000400000008e000000870000006800000068000000b3000000b4000000c0",
            INIT_45 => X"000000620000007d0000007600000095000000780000006c0000005700000041",
            INIT_46 => X"00000060000000590000009000000090000000600000006a0000005900000046",
            INIT_47 => X"000000f4000000f1000000b2000000970000008b00000082000000670000005a",
            INIT_48 => X"0000001c0000007600000092000000620000005e000000ab000000bd000000d1",
            INIT_49 => X"0000005f0000008000000064000000530000004f000000670000005f00000036",
            INIT_4A => X"000000a1000000a0000000a8000000ab0000009e0000009b000000aa00000092",
            INIT_4B => X"000000f7000000e2000000800000006f000000770000009b000000ac0000009e",
            INIT_4C => X"00000028000000640000007f0000004c0000005b000000b0000000c1000000d0",
            INIT_4D => X"000000590000003d000000350000003200000039000000490000004400000035",
            INIT_4E => X"000000640000006300000068000000710000006200000057000000770000009c",
            INIT_4F => X"000000f8000000d6000000700000004d0000003f0000007a0000009800000060",
            INIT_50 => X"00000038000000530000004e000000330000005f000000be000000c3000000ca",
            INIT_51 => X"0000003d0000003b0000003300000039000000440000003c0000002700000033",
            INIT_52 => X"000000600000005c0000005f0000006300000065000000660000006e0000005f",
            INIT_53 => X"000000f9000000d00000006c0000004f00000046000000600000006c00000064",
            INIT_54 => X"0000003f000000490000003e0000004c0000006e000000c0000000c0000000c2",
            INIT_55 => X"0000003b00000053000000480000004100000030000000280000001d0000002e",
            INIT_56 => X"000000580000003b000000400000003c000000430000004d0000004300000030",
            INIT_57 => X"000000f9000000c9000000650000006b000000690000004e0000003600000052",
            INIT_58 => X"0000004300000041000000630000005500000061000000bb000000be000000c3",
            INIT_59 => X"0000004c0000008d00000060000000480000002000000023000000260000003a",
            INIT_5A => X"00000092000000610000006d0000005e000000710000008c0000004f00000019",
            INIT_5B => X"000000f4000000c000000053000000740000008a000000450000003a000000ab",
            INIT_5C => X"0000005e00000059000000630000002c00000052000000b0000000b7000000bd",
            INIT_5D => X"00000034000000550000002f000000260000002100000024000000300000005a",
            INIT_5E => X"000000970000007100000086000000770000007b000000910000004a0000001c",
            INIT_5F => X"000000ee000000c0000000470000003b0000004700000032000000330000009c",
            INIT_60 => X"0000008b00000065000000360000002200000048000000a3000000ad000000ae",
            INIT_61 => X"0000001e0000001a000000190000001a0000001e000000280000003a00000066",
            INIT_62 => X"0000007200000076000000750000006800000056000000350000002600000025",
            INIT_63 => X"000000df000000b80000004b0000002f0000002e000000300000002b0000003e",
            INIT_64 => X"00000088000000670000005900000057000000780000009e000000a0000000a2",
            INIT_65 => X"0000001d0000001b0000001b0000001c0000002200000034000000480000005c",
            INIT_66 => X"000000b4000000b1000000ca000000cf000000af0000003d0000001500000020",
            INIT_67 => X"000000d1000000ab000000570000003e0000002c000000280000002200000054",
            INIT_68 => X"00000088000000660000007000000093000000b0000000a80000009c0000009c",
            INIT_69 => X"0000001a0000001700000016000000160000002d0000004b0000005100000056",
            INIT_6A => X"000000a5000000a9000000b1000000b9000000a4000000450000002200000023",
            INIT_6B => X"000000cc000000a70000005c0000004b0000002d0000001a000000190000004e",
            INIT_6C => X"0000008e00000063000000710000008d000000a1000000ad000000a700000095",
            INIT_6D => X"000000220000001f0000001c0000001d000000330000004f0000005300000053",
            INIT_6E => X"000000850000008a000000740000006600000061000000510000004800000032",
            INIT_6F => X"000000c6000000a4000000590000004c000000320000001d0000001b00000037",
            INIT_70 => X"0000006c00000063000000820000008b000000900000009b000000a6000000a4",
            INIT_71 => X"000000290000002700000024000000260000003800000048000000500000004c",
            INIT_72 => X"000000830000007c0000006700000054000000480000003d000000330000002d",
            INIT_73 => X"000000c3000000a9000000590000004500000032000000210000001a00000031",
            INIT_74 => X"000000490000006600000082000000870000008d0000009200000094000000a0",
            INIT_75 => X"0000002d0000002b000000280000002f00000038000000420000004d00000045",
            INIT_76 => X"0000006a0000005e00000054000000460000003d00000036000000300000002e",
            INIT_77 => X"000000ba000000af000000620000003d000000300000001f0000001a00000040",
            INIT_78 => X"00000039000000680000008b0000008f0000008c0000008e0000008d00000093",
            INIT_79 => X"00000036000000330000003100000037000000340000003f0000004a00000040",
            INIT_7A => X"00000057000000510000004a00000044000000420000003d0000003600000036",
            INIT_7B => X"000000b5000000b6000000840000004800000034000000230000002100000048",
            INIT_7C => X"0000003a0000007c000000910000009d000000a3000000a10000009600000092",
            INIT_7D => X"0000004500000046000000420000004300000041000000390000003800000037",
            INIT_7E => X"0000005e000000600000005f0000005c0000005f000000570000004800000043",
            INIT_7F => X"000000b9000000b6000000a300000076000000460000003e0000004400000051",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY28;


    MEM_IFMAP_LAYER0_ENTITY29 : if BRAM_NAME = "ifmap_layer0_entity29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000af000000c6000000d1000000d1000000b6000000bf000000ca000000d1",
            INIT_01 => X"0000008f0000008d0000009a00000095000000a00000009d000000a5000000ab",
            INIT_02 => X"000000d6000000d9000000ca000000d1000000db000000d6000000bc000000a4",
            INIT_03 => X"00000095000000950000009d000000b7000000ad000000a1000000b1000000d0",
            INIT_04 => X"000000a3000000c8000000db000000cf000000cd000000d2000000d4000000d4",
            INIT_05 => X"000000d7000000cd000000c9000000c2000000b6000000b8000000b6000000a5",
            INIT_06 => X"000000d7000000d3000000d4000000dd000000e4000000e3000000e3000000df",
            INIT_07 => X"000000ba000000ad000000aa000000c6000000bb000000c3000000cd000000df",
            INIT_08 => X"000000a4000000d3000000ec000000e3000000e2000000e3000000e5000000e6",
            INIT_09 => X"000000e0000000cf000000bf000000bc000000b8000000b7000000ad0000009f",
            INIT_0A => X"000000d3000000c8000000d0000000d6000000d6000000e0000000e5000000db",
            INIT_0B => X"000000c6000000c5000000bc000000b9000000c5000000db000000e0000000de",
            INIT_0C => X"000000af000000e3000000f1000000f2000000f1000000f4000000f4000000f5",
            INIT_0D => X"000000b6000000b8000000a0000000ae000000bb000000a1000000b0000000a8",
            INIT_0E => X"000000d4000000c4000000ba000000b9000000ca000000d0000000d5000000b9",
            INIT_0F => X"000000c8000000d4000000c5000000a9000000bb000000d5000000dc000000d7",
            INIT_10 => X"00000084000000cd000000f1000000f5000000f4000000f4000000f3000000f5",
            INIT_11 => X"0000008d0000009b0000008b0000009f000000a70000008a000000a10000008b",
            INIT_12 => X"000000e0000000c4000000a9000000a9000000a400000099000000a60000008e",
            INIT_13 => X"000000d2000000cc000000b8000000a0000000b1000000d4000000d1000000d1",
            INIT_14 => X"00000081000000d7000000ee000000f6000000f3000000f4000000f4000000f5",
            INIT_15 => X"000000a7000000b1000000aa000000aa000000aa000000a00000009c00000071",
            INIT_16 => X"000000e4000000cd000000b3000000940000008f000000980000009d0000009d",
            INIT_17 => X"000000df000000c0000000a000000093000000aa000000c1000000ce000000da",
            INIT_18 => X"000000b4000000dd000000dd000000f1000000f4000000f3000000f3000000f5",
            INIT_19 => X"000000d3000000d9000000cb000000c8000000cf000000c4000000b400000083",
            INIT_1A => X"000000e1000000cd000000a6000000a3000000bf000000c0000000c3000000cc",
            INIT_1B => X"000000da000000b20000009200000091000000a9000000b1000000d5000000e3",
            INIT_1C => X"000000c0000000d9000000ca000000e6000000f7000000f2000000f2000000f4",
            INIT_1D => X"000000d1000000ce000000d7000000ea000000e8000000e0000000c200000086",
            INIT_1E => X"000000cc0000009a000000b4000000e0000000cf000000ca000000d0000000cf",
            INIT_1F => X"000000c70000009a00000092000000ab000000bc000000c4000000c9000000dc",
            INIT_20 => X"000000ae000000df000000d1000000e3000000f5000000f3000000f3000000f5",
            INIT_21 => X"000000c9000000c1000000cc000000dd000000c1000000c1000000ba00000087",
            INIT_22 => X"000000bc000000a3000000d0000000dc000000c6000000cd000000cd000000ca",
            INIT_23 => X"000000b2000000940000008b000000a1000000cb000000df000000d1000000cb",
            INIT_24 => X"000000a4000000c2000000cd000000e5000000f2000000f3000000f1000000f2",
            INIT_25 => X"000000c4000000c0000000c4000000ca000000b8000000bd000000c10000008c",
            INIT_26 => X"000000c8000000bc000000e0000000d7000000c6000000d0000000ca000000c7",
            INIT_27 => X"000000d3000000ca000000ba000000bc000000e3000000ed000000ee000000e6",
            INIT_28 => X"0000009c000000a9000000a0000000df000000f4000000f3000000ee000000ea",
            INIT_29 => X"000000b7000000b4000000ae000000ae000000ac000000b3000000b100000086",
            INIT_2A => X"000000c4000000d0000000dc000000cd000000be000000bc000000be000000bb",
            INIT_2B => X"000000f4000000f4000000f4000000f4000000f4000000f6000000e6000000d9",
            INIT_2C => X"00000097000000be000000b6000000d8000000f2000000f2000000e6000000d3",
            INIT_2D => X"000000aa000000a60000009f0000009e000000a0000000930000006e0000006a",
            INIT_2E => X"000000af000000c6000000bd000000ad000000a60000009e000000a3000000a9",
            INIT_2F => X"000000f4000000f4000000f4000000f4000000f3000000f8000000e0000000b7",
            INIT_30 => X"0000009f000000c3000000b4000000bd000000e1000000e9000000da000000c4",
            INIT_31 => X"0000008c0000008f000000a8000000ba000000a00000008d0000005c0000005d",
            INIT_32 => X"000000960000008f0000008300000098000000a700000092000000890000008b",
            INIT_33 => X"000000f4000000f4000000f4000000f4000000f4000000f3000000e3000000bc",
            INIT_34 => X"00000089000000a200000095000000a4000000c1000000d3000000c7000000c3",
            INIT_35 => X"00000092000000a6000000cd000000bd000000a6000000b2000000aa00000096",
            INIT_36 => X"0000008a0000008000000080000000af000000d3000000c0000000ac00000099",
            INIT_37 => X"000000f3000000f3000000f5000000ef000000d3000000bf000000b1000000a0",
            INIT_38 => X"000000890000008e000000880000009c000000a2000000c8000000cf000000c2",
            INIT_39 => X"0000008b00000095000000a3000000960000009f000000b1000000b2000000a2",
            INIT_3A => X"000000850000007f0000007c000000860000009300000092000000920000008d",
            INIT_3B => X"000000f4000000f3000000f5000000cc000000a6000000ad000000a300000095",
            INIT_3C => X"000000b9000000b40000008b000000710000006e000000ad000000d0000000c3",
            INIT_3D => X"0000005f000000590000004c00000049000000570000007f0000009a00000085",
            INIT_3E => X"00000067000000630000005600000056000000580000005e000000600000005c",
            INIT_3F => X"000000f5000000f5000000e8000000af0000009b0000008f000000740000006d",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a1000000b5000000880000006000000065000000a1000000aa000000b7",
            INIT_41 => X"0000006a0000007d0000007d0000008c00000087000000810000008400000080",
            INIT_42 => X"0000002800000023000000470000004d000000270000002c0000002b00000035",
            INIT_43 => X"000000f3000000f6000000db000000a700000097000000910000005000000020",
            INIT_44 => X"000000490000009900000092000000780000007c000000c2000000c1000000ca",
            INIT_45 => X"00000083000000a90000009f000000b800000094000000830000008700000069",
            INIT_46 => X"000000730000006f000000aa000000af0000007a000000840000007600000066",
            INIT_47 => X"000000f4000000f2000000c5000000bb000000b5000000b2000000910000006f",
            INIT_48 => X"00000024000000820000009d0000007300000072000000b8000000c8000000d8",
            INIT_49 => X"000000840000009d000000810000006f0000006300000081000000950000004f",
            INIT_4A => X"000000bd000000ba000000c1000000c8000000b9000000b7000000c1000000b1",
            INIT_4B => X"000000f6000000e8000000a20000009400000097000000b6000000c7000000b5",
            INIT_4C => X"0000003d000000710000008b0000006000000071000000bb000000cc000000d9",
            INIT_4D => X"0000007d0000005e00000053000000550000005d00000073000000700000004e",
            INIT_4E => X"0000008f0000008c00000095000000a00000008a0000007f0000009f000000bf",
            INIT_4F => X"000000f7000000e20000009a00000073000000630000009f000000bd0000008a",
            INIT_50 => X"00000054000000630000005c0000004900000075000000c7000000d0000000d5",
            INIT_51 => X"0000005f00000067000000570000005f0000006900000061000000410000004b",
            INIT_52 => X"0000008f0000008900000090000000960000009700000099000000a200000086",
            INIT_53 => X"000000f7000000de00000092000000730000006f0000008f0000009900000093",
            INIT_54 => X"0000005a0000005c000000510000006500000083000000cc000000ce000000cc",
            INIT_55 => X"000000570000007d0000006f0000006200000045000000390000002d00000046",
            INIT_56 => X"0000007d0000005e00000065000000620000006700000070000000660000004a",
            INIT_57 => X"000000f8000000d4000000890000009a00000095000000710000005200000073",
            INIT_58 => X"0000005e000000560000007a0000006900000075000000ce000000d0000000d1",
            INIT_59 => X"00000063000000ad00000083000000660000002f000000330000003600000056",
            INIT_5A => X"000000ab0000007c0000008a00000079000000820000009e000000640000002d",
            INIT_5B => X"000000fa000000cf0000007500000098000000ab0000005f0000004b000000bb",
            INIT_5C => X"0000008000000072000000740000003b00000068000000cc000000d6000000dd",
            INIT_5D => X"0000004b0000006c00000046000000380000003000000034000000410000007c",
            INIT_5E => X"000000af0000008f000000a7000000910000008f000000a60000005f00000030",
            INIT_5F => X"000000fb000000d6000000680000005400000062000000480000004a000000af",
            INIT_60 => X"000000b000000080000000440000002f00000063000000c9000000d4000000d7",
            INIT_61 => X"0000002f0000002b00000027000000280000002d000000380000005000000087",
            INIT_62 => X"0000008b00000090000000930000007d0000006e000000500000003c00000037",
            INIT_63 => X"000000fb000000d90000006d000000450000004300000046000000430000005c",
            INIT_64 => X"000000aa0000008500000075000000730000009d000000cb000000cf000000cf",
            INIT_65 => X"0000002d0000002900000029000000280000003000000048000000650000007e",
            INIT_66 => X"000000c9000000c7000000dc000000da000000c0000000530000002700000032",
            INIT_67 => X"000000f7000000d20000007e0000005a0000003f00000038000000340000006b",
            INIT_68 => X"000000a1000000860000009a000000bf000000d8000000ce000000c0000000bc",
            INIT_69 => X"000000290000002300000022000000210000003e000000680000007300000079",
            INIT_6A => X"000000bb000000be000000c0000000c7000000b3000000550000003100000033",
            INIT_6B => X"000000f5000000d1000000850000006f00000042000000260000002700000060",
            INIT_6C => X"000000a0000000840000009e000000b5000000c6000000cd000000c6000000bf",
            INIT_6D => X"000000310000002c0000002600000027000000460000006f0000007600000072",
            INIT_6E => X"000000a6000000ad00000096000000870000007e000000690000005d00000044",
            INIT_6F => X"000000f2000000cf0000008200000071000000470000002a0000002800000048",
            INIT_70 => X"0000008500000082000000a3000000ab000000b8000000c6000000d1000000ce",
            INIT_71 => X"00000039000000350000002f000000320000004d000000680000006f0000006b",
            INIT_72 => X"000000b0000000a800000091000000780000006800000057000000480000003f",
            INIT_73 => X"000000ee000000d40000007e0000006600000047000000300000002800000045",
            INIT_74 => X"0000006500000086000000a6000000b2000000bd000000c2000000c2000000c7",
            INIT_75 => X"0000003e0000003b000000360000003e0000004f000000600000006900000063",
            INIT_76 => X"0000008f000000810000007400000064000000570000004e0000004500000041",
            INIT_77 => X"000000e8000000df0000008500000059000000470000002c0000002700000057",
            INIT_78 => X"0000005000000090000000bc000000bd000000bc000000be000000bc000000c1",
            INIT_79 => X"0000004e0000004a00000045000000490000004600000058000000630000005a",
            INIT_7A => X"000000720000006d00000066000000610000005d000000560000004e0000004e",
            INIT_7B => X"000000e7000000e8000000ad000000640000004a00000030000000300000005e",
            INIT_7C => X"00000055000000a5000000bb000000c8000000cd000000d0000000c7000000c4",
            INIT_7D => X"00000063000000620000005900000054000000540000004e0000004c0000004c",
            INIT_7E => X"0000007f00000080000000810000007d0000007c00000072000000630000005e",
            INIT_7F => X"000000df000000e1000000cc0000009400000060000000540000005b00000070",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY29;


    MEM_GOLD_LAYER0_ENTITY0 : if BRAM_NAME = "gold_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000101000000bc00000051000001040000004000000012000000a0",
            INIT_01 => X"00000000000000ba00000000000000000000001c000000000000004700000000",
            INIT_02 => X"0000000000000092000000000000000000000031000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000200000000000000000000010400000000000000000000000000000000",
            INIT_05 => X"0000003800000000000000a80000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000037000000530000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000000000000000000000000000000f0000000000000000",
            INIT_0A => X"000000b7000000820000011300000037000001340000017a000000a800000000",
            INIT_0B => X"000000620000014d00000000000000790000002d000000000000000000000035",
            INIT_0C => X"00000035000000100000007e0000000000000000000000000000000000000000",
            INIT_0D => X"00000000000000000000000000000000000000d1000000000000006a00000000",
            INIT_0E => X"00000081000000d20000007700000033000000a000000000000000b0000000b0",
            INIT_0F => X"000000650000000000000057000000a9000000080000000000000000000000c6",
            INIT_10 => X"000000000000007a00000058000000000000003c000000a100000000000000c8",
            INIT_11 => X"0000000000000000000000000000005c00000000000000060000000000000000",
            INIT_12 => X"000000ff00000000000000480000007700000000000000e60000002c00000000",
            INIT_13 => X"0000000000000000000000360000000000000019000000000000000000000024",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000aa0000006c000000b50000004d0000005d0000000000000000",
            INIT_17 => X"000000300000001b000000000000003f00000000000000000000000000000000",
            INIT_18 => X"0000001200000000000000b30000011900000000000000000000000000000015",
            INIT_19 => X"000000000000000000000026000000b6000000bd00000000000000aa00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000028",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001700000068000000d00000014f0000014400000124000000c000000000",
            INIT_1D => X"0000000000000016000000570000000900000000000000000000004000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000005d000000cf",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"000000b800000001000000a80000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000063000000150000009000000096000000280000001e",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000009e0000011b000000000000000000000000000000000000000000000000",
            INIT_24 => X"00000079000000000000000000000000000000000000006c0000000000000000",
            INIT_25 => X"00000000000000110000001200000067000000ff0000000400000043000000f8",
            INIT_26 => X"0000004e00000086000000000000004100000069000000000000001c00000000",
            INIT_27 => X"0000002600000017000000510000006c00000091000000000000000000000031",
            INIT_28 => X"000000000000007800000000000000e0000000fd000000b00000000000000046",
            INIT_29 => X"000000ab00000059000000000000000000000000000000000000000000000010",
            INIT_2A => X"000000530000003b000000db0000008f0000006a000000ef000000fb000000c1",
            INIT_2B => X"00000062000000ab000000460000007b00000000000000000000001000000014",
            INIT_2C => X"00000051000001230000007a0000008c0000006d000000a20000013c0000005a",
            INIT_2D => X"000000000000003c00000000000000000000000000000000000000a100000097",
            INIT_2E => X"0000010400000000000000000000000000000000000000000000000000000007",
            INIT_2F => X"0000012f000000a20000004f0000001e00000000000000000000000000000000",
            INIT_30 => X"000000a100000083000001610000013a0000015b00000000000000000000008c",
            INIT_31 => X"000000dc00000070000000880000000000000000000000120000013800000072",
            INIT_32 => X"000000000000000000000000000000ae000000cd0000013e000000ad000000e0",
            INIT_33 => X"0000001f000000c8000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001e00000000000000260000001b0000004e0000004b00000046000000bf",
            INIT_35 => X"000000a5000000aa000000060000001e000000360000009f0000013b00000073",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000010100000076000000430000006a00000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000007c00000066",
            INIT_3C => X"0000005900000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000003d00000000000000000000000000000000000000310000000000000069",
            INIT_3E => X"0000000000000000000000ed0000007200000031000000100000000000000000",
            INIT_3F => X"0000012c00000070000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000003200000000000000000000000000000000000000d00000017f",
            INIT_41 => X"00000076000000440000006d000000de00000021000000390000000800000067",
            INIT_42 => X"0000000000000000000000000000000000000000000000eb0000014100000084",
            INIT_43 => X"0000003f0000006e00000078000000b200000000000000000000000000000000",
            INIT_44 => X"0000001c0000000000000000000000000000000000000000000000920000007f",
            INIT_45 => X"00000000000000000000014800000087000000340000001e0000000000000191",
            INIT_46 => X"0000004a00000058000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000c5000000d7000000f30000000000000000000000000000000000000046",
            INIT_48 => X"0000006b00000118000000000000000000000000000000000000000000000000",
            INIT_49 => X"000001a4000000710000003a000000fe00000000000000310000000000000000",
            INIT_4A => X"000000000000000000000000000000000000000000000000000000b600000130",
            INIT_4B => X"0000000000000000000000000000000000000000000000f300000000000000e3",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000c70000004d000001690000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000520000007800000100000000000000002a000000aa000000f5",
            INIT_4F => X"000000000000000000000000000001c000000076000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000007d000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000007400000000000000000000000000000000000000110000000000000000",
            INIT_53 => X"000000000000000000000000000000b90000000600000139000000c800000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000005c00000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"000000c300000000000000000000004500000000000000000000000000000000",
            INIT_59 => X"00000149000001db000001b4000000d4000001d5000001a10000016c000000eb",
            INIT_5A => X"00000000000000000000005c000000830000007c000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"00000255000002030000004d000000d4000000a0000000d10000017600000079",
            INIT_5E => X"00000000000000630000000000000129000001b6000002700000022a00000218",
            INIT_5F => X"0000000000000000000000000000000000000059000000000000000000000000",
            INIT_60 => X"00000000000000000000000000000000000000da0000003d0000000000000000",
            INIT_61 => X"0000000000000022000001d6000001480000005f000000dd0000004a000000a8",
            INIT_62 => X"0000018a000000900000000e0000000000000000000000af0000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000013d000001370000004200000090000000d4000000f90000000000000000",
            INIT_66 => X"000000000000000000000000000000000000000000000016000000b700000138",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"000000b80000019b000001450000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000002c00000000000001060000014f00000115",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000029f000000000000019d0000016d000000b9000000000000000000000000",
            INIT_6C => X"00000121000000fb000000000000000000000000000000000000000000000000",
            INIT_6D => X"00000000000000000000000000000000000000000000000000000000000000fa",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"00000000000000000000009f00000083000000d00000000000000000000000d3",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000003d00000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"000000000000000000000000000000000000000000000000000000000000000f",
            INIT_73 => X"0000000000000000000000380000006f00000000000000000000000000000000",
            INIT_74 => X"0000007a00000079000000000000008b00000000000000000000003400000034",
            INIT_75 => X"0000000000000000000000000000000000000054000000a0000001430000018e",
            INIT_76 => X"00000000000000c2000000a40000009a00000124000000e40000009000000000",
            INIT_77 => X"000000000000000000000000000000000000000800000000000000a600000028",
            INIT_78 => X"0000009d0000016e000000ec000000db000000e4000000000000000b0000006f",
            INIT_79 => X"000000000000000000000000000000000000000000000000000001d90000005f",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000001f0000008b000000000000000000000000000000000000000000000000",
            INIT_7C => X"000000000000000000000000000000330000000000000000000000000000001c",
            INIT_7D => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_7E => X"000000000000011b000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000c100000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY0;


    MEM_GOLD_LAYER0_ENTITY1 : if BRAM_NAME = "gold_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000000000000000000930000009f",
            INIT_01 => X"0000000000000000000000000000000000000000000000dc00000000000000f5",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000006f000000f5000000c50000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000210000000000000000000000d60000003c0000009e",
            INIT_05 => X"0000018f000000d3000001610000026000000048000000000000000000000000",
            INIT_06 => X"0000002f000001a40000008f00000079000000d1000001a3000000c100000002",
            INIT_07 => X"000000b2000000710000005b0000005200000000000000000000000000000000",
            INIT_08 => X"00000000000000dc000000e900000096000000b7000000620000002d00000000",
            INIT_09 => X"000001db000001ed000001c5000000b00000006f000000470000000800000105",
            INIT_0A => X"0000000000000000000000000000000000000000000001dc000002dc000001b6",
            INIT_0B => X"0000000000000000000000000000000000000053000000c0000000fd00000000",
            INIT_0C => X"0000000000000000000000000000003700000000000000000000000000000000",
            INIT_0D => X"000000c7000001a7000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000000000007000000000000000000000010400000061000000b3000000c0",
            INIT_0F => X"000000d2000000e300000111000001ac000001c100000167000000c700000045",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_11 => X"000000ec0000000000000000000000000000004a0000009f000000fe00000000",
            INIT_12 => X"00000000000000000000000000000000000000000000000000000025000000b3",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000002b00000000000000840000000000000000000000000000000000000000",
            INIT_16 => X"000000e100000131000000740000009d000000c20000008b00000104000000c2",
            INIT_17 => X"000000000000010c000000f7000000f1000000000000000000000000000000b9",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000006100000027000000000000008900000000000000000000000000000000",
            INIT_1C => X"0000006b00000072000000000000000000000000000000000000000700000000",
            INIT_1D => X"0000000700000000000000000000000000000000000000000000000000000090",
            INIT_1E => X"0000003000000000000000000000001f00000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000018b00000000000000000000000000000000000000000000004300000003",
            INIT_21 => X"0000009d0000010d0000011300000053000000a00000003800000179000000de",
            INIT_22 => X"0000000000000025000000d7000000170000004e000000000000000000000000",
            INIT_23 => X"00000000000000000000000000000000000000000000000000000000000000dc",
            INIT_24 => X"0000000000000000000000000000000d0000002a000000140000000000000000",
            INIT_25 => X"000000df000000a00000007c000000e500000099000000000000000000000000",
            INIT_26 => X"00000023000000000000001500000023000000a000000073000000c6000000a6",
            INIT_27 => X"0000000000000000000000000000001a00000018000000000000000000000000",
            INIT_28 => X"0000005700000073000000820000000000000036000000000000000000000000",
            INIT_29 => X"000000000000008c0000009c000000660000001e000000450000001800000158",
            INIT_2A => X"00000000000000510000001c0000000000000067000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000009000000000000000000000000000000000000000000000000",
            INIT_2D => X"000000d5000000c500000000000000d0000000cf000001810000000000000000",
            INIT_2E => X"000000000000000000000000000000000000000000000062000000cf000000b1",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"00000029000000b4000000a20000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000000000006a0000006c0000009400000053000000580000009f",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000c0000000000000006300000000000000000000007e0000002c00000050",
            INIT_34 => X"0000000000000000000000000000000000000085000000000000000000000000",
            INIT_35 => X"0000001200000018000000b00000006700000000000000000000000000000022",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000003000000049",
            INIT_37 => X"0000000000000000000000000000002800000038000000590000001d00000000",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000000000001c",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000001100000000000000100000000b000000000000007100000077000000d6",
            INIT_3B => X"0000001f00000008000000000000000000000000000000000000000900000000",
            INIT_3C => X"000000eb000000900000000000000083000000a2000000530000009200000000",
            INIT_3D => X"000000000000000000000000000000000000000b00000000000000cc00000054",
            INIT_3E => X"00000032000000a9000000b7000000b700000090000000db0000009300000000",
            INIT_3F => X"000000000000000000000000000000000000001b0000000c000000200000004d",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000011e0000012300000150000000090000008400000010",
            INIT_41 => X"0000001800000000000000000000000000000089000000bb0000006c00000030",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000004a00000000",
            INIT_43 => X"000000a7000000a0000000000000000000000000000000000000000000000000",
            INIT_44 => X"000000000000009c000000a90000002800000000000000670000001200000051",
            INIT_45 => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000048",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000000000000bc000000710000000000000000000000000000000000000000",
            INIT_4C => X"000000000000000000000000000000250000005d00000000000000c9000000a5",
            INIT_4D => X"000001970000004900000031000000750000000000000000000000000000002f",
            INIT_4E => X"00000000000000420000001f0000007f000000470000005b0000013c00000091",
            INIT_4F => X"0000006d000000ae000000000000000e0000013c0000004e0000000000000041",
            INIT_50 => X"0000003e0000000000000001000000a10000011600000000000000b40000007d",
            INIT_51 => X"00000182000000bb000000fa000000d90000007d000000fc0000000e00000000",
            INIT_52 => X"00000000000000000000000000000000000000000000014d0000010500000102",
            INIT_53 => X"000000000000000000000000000000000000000a0000004f0000003e00000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"000000fc0000019f0000000000000000000000000000005c0000001a00000000",
            INIT_56 => X"000000eb0000007a000000b2000001060000008000000094000000e1000000c2",
            INIT_57 => X"000000740000008e000000f5000000000000008e000000a50000001100000107",
            INIT_58 => X"0000014c000000a8000000000000000000000000000000000000002600000037",
            INIT_59 => X"0000002c00000212000003050000000000000000000000000000000000000088",
            INIT_5A => X"000000a900000101000000000000007500000000000000000000006d00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000054000000c90000001200000000000000000000000000000000",
            INIT_5D => X"00000000000000000000006a0000000000000000000000000000000000000000",
            INIT_5E => X"00000000000000000000006100000054000000000000016a000001aa000000a0",
            INIT_5F => X"000000000000000000000000000000a800000000000000000000000000000002",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"00000000000000000000001b00000026000000e1000000000000000000000000",
            INIT_63 => X"0000008300000000000000000000002c0000000000000044000000b400000097",
            INIT_64 => X"0000000000000000000000240000004a00000056000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"000000000000000a0000000000000000000000130000005f0000000000000000",
            INIT_67 => X"0000000000000000000000a300000048000000000000000a0000009100000044",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000007",
            INIT_69 => X"000001ba00000155000000bd000000ac00000167000000a90000000000000000",
            INIT_6A => X"000000a200000000000000020000001400000083000000790000009a0000000c",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000017",
            INIT_6C => X"0000000a000000800000000e0000000000000000000000000000000000000000",
            INIT_6D => X"000000f900000009000000ca00000107000000450000006e0000000000000027",
            INIT_6E => X"000000b5000000000000004d000000770000035e000002bc00000266000000cd",
            INIT_6F => X"000000000000002500000000000000000000000000000000000001190000005f",
            INIT_70 => X"0000000000000000000000c50000011700000006000000000000000000000000",
            INIT_71 => X"00000000000001250000013c0000008f000000000000005f0000008800000000",
            INIT_72 => X"000000b80000008a000000ff0000001f00000000000000420000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"000000000000000000000000000000000000006b000000a40000000000000000",
            INIT_75 => X"0000002800000034000000d90000009a000000600000009f0000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000001780000016400000168",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"000001150000011b000000c90000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000230000000c0000007e000001730000007700000040",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000028e0000021c00000137000000000000000000000000000000a2000000be",
            INIT_7C => X"0000007300000000000000000000000000000000000000490000003e00000000",
            INIT_7D => X"000000000000000000000000000000ff000000530000005a000000930000008a",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000005b0000004300000181000000a700000081000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY1;


    MEM_GOLD_LAYER0_ENTITY2 : if BRAM_NAME = "gold_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000000000000000000000000009c",
            INIT_01 => X"000000710000000f000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000000000000000000002d0000000000000000000000000000000000000000",
            INIT_03 => X"000000c7000000320000004f0000007200000000000000000000002b0000000a",
            INIT_04 => X"0000012800000176000001db000000000000000000000053000000000000003a",
            INIT_05 => X"000000000000008c000001040000003f0000002c0000009e000000cc00000083",
            INIT_06 => X"0000007e0000008a000000000000007b00000000000000640000012900000000",
            INIT_07 => X"0000005100000000000000430000000000000000000000000000000a0000005c",
            INIT_08 => X"0000017800000000000000000000002b00000021000000000000000000000000",
            INIT_09 => X"000000600000005800000042000000790000008d0000002400000001000000f1",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000004400000003000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000800000010000000000000002b00000096000000000000000e",
            INIT_0D => X"00000000000000000000000000000000000000000000001f0000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000062000000f80000005a0000005000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000e20000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000ae00000087000000510000000000000000000000000000000000000000",
            INIT_14 => X"00000000000000000000010d000000e30000011a000000cf0000009000000000",
            INIT_15 => X"000000ae00000138000000520000000000000000000000910000000000000000",
            INIT_16 => X"000000f90000007f0000006a0000007c00000197000000000000005000000047",
            INIT_17 => X"00000098000000000000000000000000000000ef00000101000000bc0000002b",
            INIT_18 => X"000000330000010a0000017b00000000000000210000003d00000000000000e3",
            INIT_19 => X"00000030000000e70000013b00000059000000890000013b00000162000001c3",
            INIT_1A => X"00000000000000000000000000000000000000000000017f0000011300000115",
            INIT_1B => X"00000000000000000000000000000000000001320000009b0000006300000000",
            INIT_1C => X"00000000000000ca000001aa00000008000000270000000f00000000000000a5",
            INIT_1D => X"0000016400000138000000000000000000000000000000000000000000000162",
            INIT_1E => X"00000042000001540000002d0000003200000192000000950000000000000158",
            INIT_1F => X"0000026d000002120000012e000000da0000015e000000490000007c00000114",
            INIT_20 => X"000000760000000000000000000000000000001400000000000000000000003f",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000004900000036000000000000005500000009000000000000000b00000000",
            INIT_23 => X"00000000000000000000000000000000000000000000009c0000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000010d000000aa0000000000000000000000000000001c0000002b",
            INIT_26 => X"00000000000000000000004e000000b10000010e00000074000000cf000000e0",
            INIT_27 => X"0000000000000071000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000000320000017c0000006e0000000000000059000000610000003400000000",
            INIT_2B => X"000000e80000009c000000ee000001d3000000a0000000c50000010000000000",
            INIT_2C => X"000000e6000000fc000000ff00000069000000ed000000750000014e00000190",
            INIT_2D => X"000000840000012600000065000000d400000000000000de000000550000002e",
            INIT_2E => X"0000000000000000000000000000000000000000000000520000007b00000094",
            INIT_2F => X"0000000000000054000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000830000000800000000000000000000003e000000000000000000000000",
            INIT_31 => X"0000000000000000000000730000004c0000000000000000000000030000004f",
            INIT_32 => X"0000000000000032000000800000008300000000000000000000001600000000",
            INIT_33 => X"00000078000000ad000000bf00000077000000f5000000000000006900000000",
            INIT_34 => X"00000076000000a90000000000000011000000fb00000000000000790000005a",
            INIT_35 => X"0000000000000000000000000000001a00000000000000000000000000000037",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_37 => X"0000000000000007000000080000002a0000005a000000000000000000000000",
            INIT_38 => X"0000008d0000004400000000000000000000001b00000000000000000000001a",
            INIT_39 => X"0000000000000000000000600000000000000000000000000000003e00000000",
            INIT_3A => X"0000004800000010000000660000001b0000001f000000000000000000000010",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000086000000be0000014a000000590000003d000000370000009700000000",
            INIT_3D => X"0000001c0000000000000000000000000000000000000000000000e100000073",
            INIT_3E => X"00000000000000000000000000000000000000000000002e0000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000890000002a0000002c0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000f80000000100000039000000810000003700000048",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"000000000000000000000030000000000000003e000000000000000000000037",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001b000000ec000000d900000152000000b2000000d1000000ee00000000",
            INIT_46 => X"0000004200000000000000680000006f000000de000000a60000009b0000008e",
            INIT_47 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000000000000000000000d30000003b00000000000000be",
            INIT_49 => X"0000015c00000151000000dd0000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000009c00000115000000a9000000e600000156",
            INIT_4B => X"0000010e00000012000000000000000000000042000000000000000000000000",
            INIT_4C => X"0000002b00000008000000af00000000000000000000010f0000007800000052",
            INIT_4D => X"0000005500000000000000170000000000000000000000000000000000000007",
            INIT_4E => X"00000039000000000000004700000000000000000000003700000000000000b8",
            INIT_4F => X"00000000000000000000003f0000000e00000000000000000000000000000054",
            INIT_50 => X"0000000000000000000000000000000000000000000000190000000000000000",
            INIT_51 => X"00000075000000ad000000000000004700000039000000000000000000000000",
            INIT_52 => X"00000000000000000000000000000000000000f00000003f0000000c00000000",
            INIT_53 => X"0000010e000000f4000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000d10000000000000166000001a200000000000000000000015300000191",
            INIT_55 => X"00000039000000150000000400000000000000000000003b0000001700000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000029",
            INIT_5A => X"0000008500000000000000000000006600000000000000000000000000000000",
            INIT_5B => X"00000000000000450000000000000000000000a300000005000000000000003f",
            INIT_5C => X"000000050000002800000000000000000000003c000000600000000000000000",
            INIT_5D => X"000000000000006d000000000000000000000092000000000000000000000000",
            INIT_5E => X"00000000000000a20000004a000000000000003e000000950000002200000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"000000ce00000016000000ab0000003c00000000000001110000000000000000",
            INIT_61 => X"00000043000000a5000000960000002b0000007f000000c70000000000000000",
            INIT_62 => X"0000003f000000d7000000ab0000015b000000260000001e000000dd000000ba",
            INIT_63 => X"000000f2000001390000015a0000016100000000000000da000000f400000000",
            INIT_64 => X"000000000000000000000000000001140000007b000001900000011b000000b2",
            INIT_65 => X"0000000000000000000000000000004400000000000000000000000000000098",
            INIT_66 => X"0000000000000000000000a60000002300000000000000370000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000089000000de000000e000000000000000c60000010e000000a500000070",
            INIT_69 => X"000000000000005400000051000000a000000078000000860000001900000083",
            INIT_6A => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000002d000000cd00000118000000e400000000000000000000000000000000",
            INIT_6D => X"00000000000000000000007d00000096000000910000003b00000000000000c4",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000002600000076",
            INIT_6F => X"000000000000002c000000000000003d000000d4000000000000000000000056",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000970000005d000000be0000008a000000480000000000000000",
            INIT_73 => X"000000dd00000001000000000000005c000000030000004d0000004e00000056",
            INIT_74 => X"00000000000000550000000000000000000000200000002a000000000000001a",
            INIT_75 => X"0000000000000041000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000002b0000002f000000be0000000000000000",
            INIT_77 => X"000000000000000000000000000000000000000000000000000000000000001c",
            INIT_78 => X"00000000000000b0000000490000000000000055000000000000002600000000",
            INIT_79 => X"00000025000000930000003e000000220000001e000000000000000000000000",
            INIT_7A => X"000000290000000000000000000000be0000004c0000003d0000005400000034",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000006d00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"000000df00000000000000000000002b00000000000000000000000000000000",
            INIT_7E => X"0000006d0000000000000086000000cf000000000000005a0000000000000000",
            INIT_7F => X"000000000000000000000000000000000000003200000000000000000000001e",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY2;


    MEM_GOLD_LAYER0_ENTITY3 : if BRAM_NAME = "gold_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000010e000000ea000000440000002d000000820000000000000041",
            INIT_02 => X"000000000000000000000000000000000000002f000000270000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"000000c3000000bf000000c2000000de000000a400000087000000cf00000000",
            INIT_05 => X"000000000000000300000000000000000000000000000000000000e4000000cc",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000070000000820000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000001000000073000000ae000000000000009d000000e4",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000054000000000000001b00000000000000000000000000000000",
            INIT_0C => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000d3000000000000000000000109000000720000007e000000ed0000007d",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000023",
            INIT_0F => X"00000000000000a60000009e000000b8000000ca000000000000000000000000",
            INIT_10 => X"0000004e000000830000008f000000920000004e00000000000000660000003a",
            INIT_11 => X"00000000000000000000000000000136000000b5000000db0000007c00000006",
            INIT_12 => X"00000000000000000000004d0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000040000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000000000031000000e400000015000000f8000000bc",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000a500000049000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000340000005c000000000000000000000000000000000000000000000065",
            INIT_19 => X"0000000000000070000000690000002d000000000000000000000000000000c4",
            INIT_1A => X"0000000000000000000000000000006f00000084000000b50000006400000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"000000780000002a000000ae000000bc00000000000000c30000005c00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000000000000000000000000004b",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000b9000000ae0000006e0000009400000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000000000077000000bc0000006e0000012c00000077",
            INIT_24 => X"0000000000000019000000000000000000000047000000000000000000000000",
            INIT_25 => X"00000000000000e3000000aa00000082000000700000007e000000820000005d",
            INIT_26 => X"0000007000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000011600000145000000fe000000e0000000ae000001150000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000f50000011c00000059",
            INIT_2B => X"000000bc00000034000000570000005a00000000000000000000000000000000",
            INIT_2C => X"00000000000000000000003200000034000000660000006400000096000000ac",
            INIT_2D => X"0000000b0000005e000000a7000000800000004e000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000060000000400000000000000000000000c1000000000000000000000025",
            INIT_30 => X"00000057000000d3000000e2000000090000012000000108000000400000004b",
            INIT_31 => X"000000000000000000000000000001b900000004000002150000016d00000169",
            INIT_32 => X"000000000000004100000073000000000000000000000000000001da000001b7",
            INIT_33 => X"000000000000000000000000000000000000000000000000000000af0000008f",
            INIT_34 => X"0000014900000120000002790000037c00000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000160000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000004b00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000003b000000eb000001bf0000013b0000009e000000080000000000000000",
            INIT_3B => X"000001340000000000000000000000000000000000000000000000be00000000",
            INIT_3C => X"000000000000000000000000000000000000000000000000000001420000001e",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"000000d100000069000000000000000000000000000000e30000000000000000",
            INIT_3F => X"00000000000000000000000000000000000000000000000e000000eb000000fe",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b4000000ca000000d00000016c000000cc000001630000000000000000",
            INIT_41 => X"0000015600000094000000260000006500000000000000000000000000000073",
            INIT_42 => X"00000000000000000000008600000000000000000000006c0000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000262000000db000000420000022f000001ec000000000000000000000000",
            INIT_46 => X"00000027000000310000017a000000c6000000000000008c0000009e0000005f",
            INIT_47 => X"00000000000001b700000011000000000000006a00000000000000000000000d",
            INIT_48 => X"0000008c00000051000000000000000000000000000000000000012000000170",
            INIT_49 => X"000000000000013900000097000000a1000000a4000000c40000008200000148",
            INIT_4A => X"0000000000000000000000000000010000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"000001090000011c000000e60000002900000062000000000000000000000000",
            INIT_4D => X"000000000000000000000000000000000000000000000000000000000000009f",
            INIT_4E => X"0000000000000000000000000000000000000000000002360000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"00000033000000aa000000840000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000f50000004600000000000000000000000000000040",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000008a000001f90000019400000000000000c8",
            INIT_54 => X"00000000000001270000000000000356000001d20000016a0000026b0000028f",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000026",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000002a00000135000000d8000002000000008e",
            INIT_58 => X"00000000000000fb000000000000000000000000000000000000000800000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000000000001100000000000001240000003f000001cf0000008700000000",
            INIT_5B => X"0000000000000059000000000000012d0000000000000112000000f400000000",
            INIT_5C => X"000000c70000000000000000000000bc0000000000000084000000880000004f",
            INIT_5D => X"0000004600000000000000000000009a000001bf00000082000001c900000115",
            INIT_5E => X"0000000000000089000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000002800000000000000000000000000000000000000000000000000000179",
            INIT_60 => X"000000b300000374000001a8000002a2000000a60000019b000001ba000000d7",
            INIT_61 => X"000000530000007a0000005e00000064000002310000027b00000026000001c7",
            INIT_62 => X"0000000000000000000000000000000000000000000000ca000000d70000005a",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000009c0000001a000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000009d000000b10000000000000051000000780000002b0000000000000000",
            INIT_66 => X"00000000000000000000000000000000000000000000000000000000000000bb",
            INIT_67 => X"0000007800000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000170000012700000059000000ce00000000000000000000000000000000",
            INIT_6B => X"000000000000000000000000000000370000000000000000000000b300000000",
            INIT_6C => X"0000007f00000224000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000000000019800000168000001750000000000000072000000f300000040",
            INIT_6E => X"000000000000010300000045000000000000011e000000000000000000000011",
            INIT_6F => X"000000780000000000000000000000b500000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"00000182000002670000012c00000134000001de000002c80000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000001650000013800000154",
            INIT_73 => X"00000010000000000000000000000000000000ad000000000000000000000000",
            INIT_74 => X"0000000000000000000000c30000000000000000000000590000000000000000",
            INIT_75 => X"000001530000001a000000100000000000000000000000c10000000000000000",
            INIT_76 => X"000001a500000000000000000000000000000000000000000000002000000000",
            INIT_77 => X"0000000000000134000000af0000000400000096000001a000000089000001d1",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"000000000000006f000000000000000000000075000000330000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"00000155000001b50000017e0000002a00000029000000000000001e00000000",
            INIT_7E => X"0000006f00000000000001e80000018f00000081000001ea00000168000000bd",
            INIT_7F => X"000000000000003d000000d3000000f100000091000000160000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY3;


    MEM_GOLD_LAYER0_ENTITY4 : if BRAM_NAME = "gold_layer0_entity4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000e300000000000001140000010c0000000000000000000000e700000000",
            INIT_03 => X"0000014300000182000000f600000092000000f2000000fe00000000000000b9",
            INIT_04 => X"0000000000000000000000cb00000001000000000000013a0000010400000081",
            INIT_05 => X"0000006400000069000000360000001a0000002100000000000000000000005c",
            INIT_06 => X"00000000000000000000000000000036000000b30000012e0000000000000093",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000500000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000000000011900000000000000b500000166000000380000000000000066",
            INIT_0B => X"0000000000000090000001340000001c00000072000000be0000004f00000000",
            INIT_0C => X"0000000000000001000000000000000000000011000000240000004e00000089",
            INIT_0D => X"00000000000000000000008a0000000f000000000000002e000000940000000c",
            INIT_0E => X"0000009f00000000000000600000005e0000000000000000000000a400000000",
            INIT_0F => X"000000000000000000000000000000ae00000000000000000000008100000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000001000000000000000000000002b00000000000000000000000000000000",
            INIT_12 => X"00000000000000000000006000000000000000290000013d000000cd00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000001f0000000000000000000000b100000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000002e00000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000016",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000000000005e000000a30000000000000000000000000000000000000000",
            INIT_19 => X"000000000000000000000000000000c300000063000000000000009800000096",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000870000000000000000000000000000001800000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"000000000000010b00000089000000d600000146000000db000000cd00000000",
            INIT_1E => X"0000000000000071000000000000000000000000000000410000010400000072",
            INIT_1F => X"00000130000000500000000900000075000000a20000001b000000d2000000a7",
            INIT_20 => X"00000000000000000000000000000000000000940000011500000000000000c5",
            INIT_21 => X"0000004500000000000000820000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000000d0000000000000046000000fd",
            INIT_23 => X"000001450000000000000000000000000000001900000000000000000000003c",
            INIT_24 => X"0000000000000039000001720000000e00000066000001e60000002000000088",
            INIT_25 => X"00000000000000000000014c000000240000000000000069000000e600000021",
            INIT_26 => X"0000000000000062000000000000000000000000000000000000000000000122",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000008b00000000",
            INIT_28 => X"0000000700000000000000000000000000000031000000050000000000000000",
            INIT_29 => X"00000055000000b5000000500000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000b0000000000000000000000d100000000",
            INIT_2B => X"0000011700000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"000000700000000d0000000000000000000000e8000000ad0000000000000105",
            INIT_2D => X"000000000000002f0000007b000000000000000e000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000a10000001400000000000000bc0000007c000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000001400000000000000000000007b00000000000000000000000000000000",
            INIT_33 => X"0000008100000076000000000000000c00000000000000160000000000000021",
            INIT_34 => X"00000000000000000000000000000000000000000000000d0000000000000000",
            INIT_35 => X"0000006200000000000000440000006a00000000000000000000000000000000",
            INIT_36 => X"0000006100000084000000000000005b0000003d00000000000000000000007d",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000120000001b00000124000000000000002d000000d1000000a700000000",
            INIT_39 => X"0000007d0000004b0000006b0000008f0000005d000000570000002500000112",
            INIT_3A => X"000000b900000000000001b10000019c000000000000008400000057000001ad",
            INIT_3B => X"0000007f00000079000000b6000000ae000001d2000000eb00000091000001f5",
            INIT_3C => X"0000003f000000000000000000000093000000fd000000950000005800000139",
            INIT_3D => X"000000dd0000001600000000000000000000000000000010000000000000004b",
            INIT_3E => X"000000000000003e0000000000000000000000a900000000000000000000006a",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000049000000af0000004500000047000000a200000035000000a900000140",
            INIT_41 => X"0000000000000033000000000000000000000000000000000000000000000092",
            INIT_42 => X"0000001d0000000000000000000000aa00000000000000000000000000000062",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"000000000000000000000000000000500000002e000000000000000000000000",
            INIT_46 => X"0000003300000000000000000000001c00000034000000250000000000000000",
            INIT_47 => X"00000000000000b9000000160000004900000012000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"00000000000000780000001b000000bc000000f50000009d000000cf00000000",
            INIT_4B => X"000000ec000000db000001010000010c000000b100000177000000640000003c",
            INIT_4C => X"000000a0000000e8000001310000007a0000013700000056000000b8000000aa",
            INIT_4D => X"0000000f00000000000000a700000020000000720000000e000000fd00000000",
            INIT_4E => X"000000000000000000000000000000880000001500000000000000000000005c",
            INIT_4F => X"0000001a0000014b000000000000000000000000000000000000000000000000",
            INIT_50 => X"000000180000004d000000000000000000000000000000000000000000000045",
            INIT_51 => X"0000000900000041000000330000008600000012000000000000000000000000",
            INIT_52 => X"0000003e00000000000000000000000000000000000000050000000000000000",
            INIT_53 => X"00000000000000000000001c00000039000000f1000000180000002200000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000065000000000000000000000030000000450000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_58 => X"0000004600000032000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000006000000000000000000000000000000024000000170000000000000000",
            INIT_5A => X"00000008000000aa000000230000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000006900000001000000bb0000010d000001730000011a0000014e00000000",
            INIT_5D => X"000000490000000b0000004b0000004800000000000000000000011e0000007b",
            INIT_5E => X"0000000000000000000000000000000000000000000000a40000015000000126",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"000000210000000b000000120000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000a9000000ab000000350000006d000000a4000000dd",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000000000000000000000000000000000000000000000000000000000001c",
            INIT_64 => X"0000000000000000000000000000000000000000000000650000000000000000",
            INIT_65 => X"0000010800000000000000ca000000e9000000640000002f0000001000000007",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000008a000000c0",
            INIT_67 => X"00000081000000cc000000ab000000820000004e000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000081000000b80000006d00000053",
            INIT_69 => X"000000e60000003a000001d10000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000000000000071000000500000008a",
            INIT_6B => X"0000000000000000000000000000001600000000000000000000004100000000",
            INIT_6C => X"0000000000000045000000000000000000000084000000000000000000000000",
            INIT_6D => X"00000033000000ce000000870000006800000092000000890000000000000000",
            INIT_6E => X"0000006700000036000000460000005600000000000000b30000002100000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000014",
            INIT_70 => X"0000000000000000000000000000000000000047000000000000000000000000",
            INIT_71 => X"0000010e000001130000010b000000f600000000000000000000000000000002",
            INIT_72 => X"00000000000000000000000000000048000000060000009f000000000000004c",
            INIT_73 => X"00000000000000c6000000000000000000000000000000000000000000000000",
            INIT_74 => X"000000dc0000000000000000000000770000002700000000000000a200000026",
            INIT_75 => X"000000690000000f000000490000000000000018000000000000019f000000b5",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000190000005400000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000300000038000000000000003c00000055",
            INIT_7C => X"0000000000000000000000000000001000000000000000020000006200000095",
            INIT_7D => X"000000980000004c000000000000000000000035000000000000000000000000",
            INIT_7E => X"000000000000001b00000000000000b50000000000000000000000190000000b",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY4;


    MEM_GOLD_LAYER0_ENTITY5 : if BRAM_NAME = "gold_layer0_entity5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000012000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000006f0000008000000000000000f200000088000000900000001d00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000f5000000ef000000aa",
            INIT_03 => X"000000a9000000000000000e0000000000000001000000000000000000000022",
            INIT_04 => X"00000000000000b800000000000000d6000000a20000008a000000970000004b",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_06 => X"0000000000000000000000000000004800000053000000000000000000000058",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000010a0000004e000000000000000e0000019b000000000000000000000141",
            INIT_09 => X"0000000000000122000001560000013a000000000000004d0000003200000075",
            INIT_0A => X"000000000000000000000000000000000000000000000000000001d400000172",
            INIT_0B => X"0000000000000000000000000000000000000000000000ce0000000600000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000c8000000aa000000000000000000000000000000000000000000000000",
            INIT_0E => X"000000440000016000000000000000000000000000000000000000bb00000000",
            INIT_0F => X"00000000000000620000002c0000000000000000000000000000011c00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000600000000000000000000000e50000000000000000000000b300000000",
            INIT_13 => X"0000002e0000000000000000000001740000000000000000000000ec00000058",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000005700000000",
            INIT_16 => X"000000000000000c0000000000000000000000000000002e0000000000000000",
            INIT_17 => X"00000000000000000000000000000009000000000000006b0000000000000012",
            INIT_18 => X"0000005f00000000000000820000006e00000029000000210000006c00000000",
            INIT_19 => X"0000000000000053000000bb000001910000017400000179000000920000008a",
            INIT_1A => X"000000000000000000000000000000000000000000000000000000410000004b",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000048000000580000003f0000000000000000000000000000000000000000",
            INIT_1D => X"000001f800000000000000000000017300000000000000000000000000000000",
            INIT_1E => X"00000000000000690000003c00000000000000830000009a00000000000001ce",
            INIT_1F => X"000000000000002c000000000000000000000000000000000000000000000062",
            INIT_20 => X"0000006f00000054000000ac000000b800000000000000890000001500000000",
            INIT_21 => X"000000190000008100000122000000c6000001d90000015a000000de00000000",
            INIT_22 => X"0000014400000000000000000000009f00000022000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"000000fb00000000000000000000009200000000000000000000000000000000",
            INIT_25 => X"00000000000000070000018c000000cb00000056000001690000000000000000",
            INIT_26 => X"00000000000000000000000000000000000000000000003c00000044000000d9",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000077000000f9000001100000000000000000000000000000000000000000",
            INIT_29 => X"00000000000000000000000000000000000000d700000000000000430000016a",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000a9000000fb00000000000001340000004200000000000000000000009f",
            INIT_2C => X"000000000000004c000000190000004b00000000000000000000005400000000",
            INIT_2D => X"0000006300000000000000000000000000000029000000650000000000000058",
            INIT_2E => X"00000000000000000000003c0000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000038000000f2000000770000006400000081000000040000002b",
            INIT_30 => X"000000000000000000000000000000000000000000000000000000d700000000",
            INIT_31 => X"0000007c00000053000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000400000016100000000000000540000001a0000007b0000000000000000",
            INIT_33 => X"0000001700000000000000850000000000000000000000420000017400000000",
            INIT_34 => X"0000000000000000000000ea0000004d000000000000002e0000004a00000018",
            INIT_35 => X"00000000000000000000000000000098000000000000001a000000000000000f",
            INIT_36 => X"000000000000015200000035000000000000000b000000000000008e00000000",
            INIT_37 => X"0000000000000000000000d20000000000000000000000b90000012400000000",
            INIT_38 => X"0000009e000001d10000005c0000000b00000052000000740000000000000098",
            INIT_39 => X"000000000000000000000000000000270000010b000001110000004000000131",
            INIT_3A => X"0000000000000000000000000000000000000000000001570000001500000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000005500000000",
            INIT_3D => X"0000004a0000005d000000c70000000000000000000000000000010d00000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000000000000c2000000210000000000000000000000000000000000000008",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004e000000b900000000000000000000000000000000000000430000004f",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000017000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000069000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000004d000000000000000000000000000000000000010a000000db00000000",
            INIT_45 => X"000000000000014400000069000000000000004800000022000000be00000000",
            INIT_46 => X"000000550000011e00000000000000ef0000002600000000000000c400000000",
            INIT_47 => X"0000007f000000580000004e0000008700000000000000000000012700000000",
            INIT_48 => X"0000000000000022000000d3000000aa00000000000000cf000000000000001f",
            INIT_49 => X"000001410000017c00000129000000ca000001a8000000e40000000000000056",
            INIT_4A => X"00000000000000000000000000000000000000000000018400000169000000c0",
            INIT_4B => X"0000006f00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000003700000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000008200000000000000000000005e00000102000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000dc0000000000000064",
            INIT_4F => X"000000a4000000ac0000000000000184000001ba0000000000000000000000f9",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY5;



end a1;