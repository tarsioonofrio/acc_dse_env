LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE ifmap_package is
		type padroes is array(0 to 4000000) of integer;

		constant input_map: padroes := ( 

			0, 25, 35, 
			66, 0, 3, 
			209, 0, 0, 
			

			145, 0, 0, 
			0, 0, 0, 
			0, 0, 131, 
			

			0, 0, 0, 
			0, 0, 56, 
			54, 60, 201, 
			

			57, 86, 10, 
			0, 45, 0, 
			0, 0, 0, 
			

			61, 93, 194, 
			150, 32, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 130, 
			0, 94, 95, 
			16, 0, 100, 
			

			0, 33, 31, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 62, 20, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 8, 78, 
			

			43, 52, 0, 
			71, 0, 0, 
			0, 0, 0, 
			

			0, 0, 126, 
			0, 71, 8, 
			259, 122, 234, 
			

			44, 53, 0, 
			0, 0, 0, 
			0, 154, 269, 
			

			0, 0, 0, 
			0, 0, 57, 
			0, 0, 50, 
			

			61, 7, 0, 
			0, 0, 0, 
			0, 0, 48, 
			

			0, 0, 0, 
			0, 0, 0, 
			40, 8, 29, 
			

			92, 335, 246, 
			184, 58, 30, 
			41, 0, 4, 
			

			4, 104, 56, 
			0, 0, 0, 
			0, 0, 14, 
			

			43, 144, 131, 
			188, 171, 144, 
			169, 35, 0, 
			

			0, 0, 0, 
			0, 42, 24, 
			0, 0, 0, 
			

			0, 40, 0, 
			201, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 40, 0, 
			45, 0, 123, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 184, 16, 
			82, 0, 0, 
			2, 129, 43, 
			

			0, 59, 28, 
			1, 50, 134, 
			77, 0, 3, 
			

			0, 0, 0, 
			0, 21, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 117, 59, 
			0, 0, 0, 
			0, 0, 72, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 208, 
			0, 0, 95, 
			125, 0, 16, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 50, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 5, 0, 
			0, 14, 0, 
			

			32, 0, 16, 
			251, 0, 0, 
			67, 53, 28, 
			

			40, 86, 115, 
			87, 61, 22, 
			0, 0, 0, 
			

			87, 0, 140, 
			168, 188, 115, 
			156, 0, 0, 
			

			128, 0, 85, 
			41, 0, 18, 
			0, 0, 0, 
			

			23, 36, 43, 
			0, 55, 0, 
			0, 0, 0, 
			

			0, 0, 66, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			94, 58, 0, 
			191, 0, 18, 
			0, 102, 93, 
			

			29, 61, 65, 
			25, 0, 0, 
			0, 0, 0, 
			

			0, 0, 68, 
			0, 0, 46, 
			101, 0, 35, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			19, 0, 0, 
			0, 95, 198, 
			338, 245, 176, 
			

			0, 0, 0, 
			0, 106, 23, 
			214, 563, 506, 
			

			99, 55, 86, 
			58, 181, 46, 
			0, 0, 0, 
			

			10, 0, 0, 
			0, 24, 55, 
			66, 55, 19, 
			

			44, 0, 0, 
			86, 103, 120, 
			53, 112, 46, 
			

			0, 0, 60, 
			0, 150, 68, 
			27, 0, 0, 
			

			0, 0, 0, 
			53, 0, 0, 
			0, 0, 0, 
			

			33, 106, 0, 
			0, 0, 0, 
			0, 0, 21, 
			

			0, 0, 43, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			58, 0, 0, 
			

			75, 0, 53, 
			41, 0, 2, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			

			0, 0, 0, 
			0, 0, 138, 
			0, 0, 0, 
			

			0, 0, 0, 
			22, 83, 0, 
			0, 0, 0, 
			

			72, 21, 0, 
			0, 59, 0, 
			0, 0, 0, 
			

			16, 0, 0, 
			0, 0, 0, 
			0, 0, 51, 
			

			0, 0, 0, 
			0, 0, 0, 
			0, 0, 0, 
			
		others=>0 );
END ifmap_package;
