-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity ifmap_18k_layer2_entity0 is
    generic (
        DEVICE: string := "7SERIES"
        );
  
    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic_vector(2-1 downto 0);;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(10-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
  end ifmap_18k_layer2_entity0;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "18Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_03 => X"00000000000000000060006c003700210038000c004c00000000000000170000",
       INIT_04 => X"000f002a00000000001500070000002b005f0061001100130000000000000029",
       INIT_05 => X"0000005d007300000043004600b8005a000000000000001700d6002300000000",
       INIT_06 => X"00000000000500000000001c003a001f0027013a000e0000001d00c200240038",
       INIT_07 => X"0080006f0000001701cf00220000000000160000006000f2000000000000017a",
       INIT_08 => X"009200000000000a00000000009d00ce0000000d00000000007b0000007c000c",
       INIT_09 => X"00000003000000000000000f0000000000000000000000000000000000110000",
       INIT_0A => X"0000000000000000000000360000000000000000003800000000000000000000",
       INIT_0B => X"00000000004b0000000000770000009d000000000000002d0000001500000000",
       INIT_0C => X"00000013000000210000000600000000000000000000000000000000000d0000",
       INIT_0D => X"000000790000006e000000000000006a00000000000600000000000000cb0000",
       INIT_0E => X"00000000003c0039001b003700000000000000000000000600000000003200b6",
       INIT_0F => X"000000080000000a0000003900670000000c00200011002e0000002a00000015",
       INIT_10 => X"0036000900170000000000000009000b00190006000000170000000d00290009",
       INIT_11 => X"00000008000000000000000000000000000000000000000000170000000d0009",
       INIT_12 => X"000000160026001a001300000000000000000000000000000000000000000000",
       INIT_13 => X"0000000000000000000500000001000200000000000000000000001b0000000e",
       INIT_14 => X"00110000000000000000000000000000000000000000000f0000000000000000",
       INIT_15 => X"003b00020000000100060018001500000000000000000000000b000000050000",
       INIT_16 => X"000000110006001c004000010000001f000c00050017002d0008002100120008",
       INIT_17 => X"00130022003000000000003800310000002e001a000000080000000000000000",
       INIT_18 => X"00000000000000000000000000000000002200000000004a004a002a00320000",
       INIT_19 => X"00090009000a00000011003200000000000000050000003e00040019001f0000",
       INIT_1A => X"005b0000004e00000000000000160000005d005b0000000d00000083005f0000",
       INIT_1B => X"000000000000005b001c00000000000000000000000000000000000000000000",
       INIT_1C => X"0000000000000029000000190000000000000000003c00000017000000360000",
       INIT_1D => X"00000010000000000000001f000000080017000e000000000000000000aa003b",
       INIT_1E => X"00560027002f0000002700870056004d004c00720068006100510094002d0000",
       INIT_1F => X"004d00000038002500000018000c000a0000009b002d0000000e001c00000000",
       INIT_20 => X"00000074003900390036001b0000000000130000004b001d0002004d00500092",
       INIT_21 => X"00500000000000000024009e000000000000001200150032004b001c00000000",
       INIT_22 => X"000000000000000000000000004e0000000000000037002c0000002500000000",
       INIT_23 => X"0000000000640000003f000000110013000000000000000000000000005f0002",
       INIT_24 => X"0000000700000014000b00040053000400180032002e00170000000000000000",
       INIT_25 => X"0000000000000000000000000000000d000d0000000000000000000000000000",
       INIT_26 => X"0000000d00000000000000160000000e001e0000000000060000000000010021",
       INIT_27 => X"00000000000000000012001b000000000000003900380041002e000000000000",
       INIT_28 => X"0000000000000000000000000000000000000022000000000000000000000000",
       INIT_29 => X"00000000000000000000000000000000002300000017007c00030000001a0000",
       INIT_2A => X"0000001a0000001500060018001700000000000c001e00240035004000810092",
       INIT_2B => X"0027006c00190000003300000000000000000000000000000000007000000000",
       INIT_2C => X"00000005000000000000001c004f003800380000003600000000000000000000",
       INIT_2D => X"0000000000000000000000000000000000000013000000000000000000000000",
       INIT_2E => X"000000000000000000000000000000000000001c004200650026006600000000",
       INIT_2F => X"0062004e00590056007700190000004d00600035004700b70074000c00280025",
       INIT_30 => X"001800390085007800390050006e0084008a009a008b00a90092009c00ab00bb",
       INIT_31 => X"00000000000a00a600b500a90067005000460097004d00000000001c002d0011",
       INIT_32 => X"001c0000000000210000001d0068001d000000000000000000000000002b002f",
       INIT_33 => X"00370034006a0040002400d10067005600730042001700610000000000000000",
       INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_35 => X"0000000f00000000000000000000000000000000000000000000000000000006",
       INIT_36 => X"00000000002100000068000000b3009b007d009c007c00c1007d00a0009800a9",
       INIT_37 => X"00c200b00006001c000000000000000000000000001100000000000000000000",
       INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INIT_3A => X"00000000000000620061004b0051005000490041006100880053005b005e005a",
       INIT_3B => X"002a0068005a00600076005f0073003c0076006d004e007b00460041005d005c",
       INIT_3C => X"00970046003b004f001000150023002e002f00000000000000000000000d0000",
       INIT_3D => X"000000000000000000630073007b00570056004b004800450070004300400005",
       INIT_3E => X"00120044002b00320022001e00000024003c0007005d00000009000000210021",
       INIT_3F => X"000000060000001500190017002b000000000000000000000000000000000000",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
