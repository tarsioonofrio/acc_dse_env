library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    -12555, 5187, 421, -594, 6712, -7672, 9532, 3569, -7946, 2656,

    -- weights
    -- filter=0 channel=0
    -2, -4, -11, -10, -7, -4, -9, -2, -5, -5, -4, -4, -9, -10, -8, -4, -11, -6, -10, -10, -7, -4, -11, -4, -9, -10, -5, -5, -2, -9, -5, -7, -1, -1, -4, -1, -5, -7, -1, -2, -5, -7, -8, -2, -1, -4, -9, -3, -9, -5, -10, -3, -8, -10, -1, -5, -8, -3, -3, -8, -6, -8, -7, -7, -5, -3, -5, -9, -5, -1, -7, -9, -8, -8, -7, -3, 0, -6, 0, -7, -1, -7, -8, -8, -8, -6, -1, 0, 0, -8, -2, -7, -7, -7, -9, 0, -6, -7, -5, -8, -3, -2, -7, -3, -9, -9, -10, -5, -1, -5, -8, -4, -9, -5, -4, -8, -9, -6, -7, -1, -7, -1, -2, -5, -3, -8, -8, -3, -4, -6, -2, -1, -8, -9, -4, -5, -5, -4, -4, -5, -1, -1, -1, -7, -1, -1, -9, -2, -5, 0, 0, 0, -5, -5, -3, -5, -4, -1, -2, 0, -3, 0, -8, 0, -2, -7, -6, -6, -4, -3, -4, -3, -3, -3, 0, -5, -3, -5, -9, -3, -2, 0, -6, -3, -6, -5, -6, -2, 0, -7, 0, -3, -5, -2, 0, -7, -5, -2, 0, -4, -1, -6, -7, 0, 0, -4, -2, -4, -4, -3, -1, -6, -6, -1, -6, -7, 0, -1, -8, -4, -4, -5, -6, -2, 0, -4, 0, -4, -1, -3, 0, 0, 0, 0, -6, -8, -6, -6, -2, -6, -10, -10, -3, -3, -3, -2, -6, -4, -6, -2, 0, -1, -9, -2, -1, 0, 1, -4, -3, -1, 0, -2, -6, -3, 0, -3, -5, -1, -6, -4, -8, -9, -7, -6, -10, -5, -6, -4, -10, -7, -1, -1, -4, 0, -1, -5, -4, 1, -3, -2, -4, -7, -3, -3, -4, -3, 1, -5, -3, -4, -6, -8, -5, -3, -12, -6, -3, -7, -9, -10, -7, -8, -7, -9, -7, -5, -8, -2, -3, 2, -2, -1, -3, -7, -6, 0, -7, -5, -7, -5, -7, -3, -11, -4, -4, -10, -5, -4, -9, -3, -9, -6, -1, -8, -2, -4, -6, -4, -7, -4, -2, -1, -5, -3, 0, -4, -4, -7, -8, -8, -2, -8, -3, -8, -7, -6, -6, -7, -13, -4, -5, -9, -4, -3, -8, -5, -2, -7, -3, -9, -10, -4, 0, 0, 3, 1, -3, -4, -8, -7, -10, -9, -9, -6, -9, -12, -10, -9, -14, -14, -13, -10, -10, -11, -5, -3, -8, -4, -9, -9, -2, -2, -6, -3, -5, 3, 0, -4, -2, -2, 1, -4, -5, -7, -4, -4, -13, -14, -9, -14, -17, -13, -13, -15, -12, -7, -4, -6, -5, -2, -8, -3, -2, -1, -2, 0, -4, 1, 0, -2, -1, -3, -2, -7, -3, -7, -9, -10, -9, -9, -14, -12, -12, -17, -11, -9, -14, -11, -13, -6, -10, -9, -7, -3, -2, -3, -3, 0, -3, 1, -3, -2, -2, -2, 0, -4, -1, -6, -9, -11, -11, -14, -15, -11, -13, -14, -15, -12, -15, -5, -6, -9, -5, -7, -9, -10, -8, 1, 0, -5, 2, 0, 0, 2, 1, -3, -5, -1, -5, -3, -11, -10, -7, -6, -8, -10, -15, -16, -17, -17, -16, -8, -10, -6, -8, -5, -12, -7, -5, 1, 3, -4, 0, 0, 0, 1, -1, 2, -1, -4, -7, -3, -8, -6, -11, -11, -16, -14, -20, -14, -17, -21, -15, -11, -9, -5, -8, -10, -6, -8, -1, 0, -4, -3, 1, -6, 0, -4, -2, 3, 1, 0, -4, -2, -4, -12, -7, -9, -11, -12, -16, -16, -18, -23, -16, -11, -11, -11, -12, -11, -8, -2, 0, 2, -5, -5, 1, 1, -5, -2, -2, 3, 0, 1, -5, 0, -5, -10, -12, -16, -17, -17, -14, -14, -19, -15, -18, -11, -9, -4, -10, -4, -9, 0, 1, 0, -6, -1, -4, -3, -4, 3, -1, 0, -3, -1, 1, -1, -8, -12, -11, -7, -8, -12, -13, -17, -14, -21, -10, -13, -6, -5, -3, -1, -7, -6, -4, -3, -3, 1, -5, 0, -6, 0, 0, -3, 3, 4, -3, -5, -2, -8, -10, -11, -5, -9, -13, -12, -12, -18, -12, -8, -8, -12, -3, -7, 1, 1, -1, -2, -2, -3, -7, -7, -3, -5, -3, -2, 2, 0, -4, -3, 0, -7, -5, -3, -5, -11, -7, -8, -9, -12, -8, -4, -7, -4, -3, -6, -4, -3, 1, 0, 0, -5, -5, -4, -2, 0, -2, 3, -3, 0, 1, -1, 0, -7, -7, -5, -10, -7, -9, -8, -4, -3, -7, -7, -7, -4, -6, -6, -4, -5, 3, 0, 2, -5, -3, 0, -2, -7, 1, 0, -2, 0, 1, -1, -5, 0, -6, -2, -7, -9, -3, -7, -5, 0, -5, -2, 0, -5, -4, 0, -3, 1, -4, 3, -2, 1, -2, -6, -2, -3, 0, 1, -1, -5, -2, -4, 3, -4, 1, 0, -7, -7, -6, -1, -6, -5, 0, -2, 0, 1, -6, 1, 0, 2, -4, -4, 0, -4, -1, -5, -5, 0, 0, -5, 0, -5, -4, 3, 1, 1, -1, -3, -5, -4, -3, -4, -1, 1, -3, -3, -2, -2, -6, -1, 2, 1, 0, 0, -3, 1, 0, -6, -2, -7, -4, 0, 0, -5, 0, 0, 1, -3, 2, 0, -1, -4, -1, -6, -4, -2, -4, -1, 0, 0, -3, 0, 1, 0, -3, -4, -1, -1, -6, 0, -7, -8, 0, 1, 1, 0, 3, 0, -1, 0, 2, -2, 0, 0, 2, 1, -2, 5, -2, 3, -5, -3, 1, -6, 0, -4, -2, -1, -1, -3, -6, -6, -8, -4, -4, -4, -5, 0, 2, -3, -2, -3, 0, 0, -3, -1, 0, 1, 2, 0, -3, -2, -1, 0, -1, -4, 1, -4, 0, 0, -4, -8, -9, -8, -4, 0, -4, 0, -5, -1, 1, 0, 0, -3, 2, 1, 2, 0, 0, 2, 3, 0, -4, -2, -2, 0, -5, 0, -2, -2, -3, 0, -7, -3, -1, 0, -9, -6, -7, -5, -5, -6, -8, 0, -6, -5, -8, 0, -5, -5, -1, -1, 0, 0, -1, -2, -6, -6, -7, -3, -6, -1, -2, -2, -4, -9, -2, -9, -2, -1, -9, -7, -4, -5, -1, -1, -4, -6, -3, -1, -4, -4, -8, -4, -6, -4, -6, -10, -4, -8, -4, -1, -6, -6, -6, -8, -7, -9, -4, -7, -1, -1, -7, -3, 0, -6, -1, -4, -8, -8, -8, -5, 1, -2, -3, -1, -3, -2, -1, -1, -1, 0, -3, -8, -3, -8, -8, -1, -6, -6, -3, 0, -3, -7, -9, -3, -7, -1, -3, -1, -6, -1, -7, -2, -1, -4, -5, 1, -3, 0, 0, -6, 0, 1, 2, 0, -3, 0, 0, -1, -8, -2, -2, 0, -6, -5, -8, -7, -8, 0, -3, 0, -3, -6, -2, -6, -4, -4, -5, 1, 1, 0, 0, 0, -3, -5, -3, 0, -4, -2, 0, -5, -8, -6, -6, 0, -6, 1, 0, -4, -9, -1, 0, -2, -5, 2, -2, -2, 0, 0, 0, -3, -2, 2, -1, 2, -2, 1, -4, -4, -5, -1, -2, 0, -4, -6, -5, -1, -1, -7, 0, 1, -7, -1, -2, -1, -5, -5, 2, -2, 5, 1, -3, -1, -4, 0, -1, 3, 4, 0, -5, -2, -5, 0, 0, -2, -5, 0, 1, -3, -2, -6, 0, 0, -3, 0, -1, 4, -1, -2, 2, -1, 5, 1, -1, 2, 4, -3, 3, 3, 4, 4, 1, 0, 4, -2, -4, -5, 0, -2, -6, 0, -4, -6, -1, -5, -5, -4, 0, 0, 4, 3, -4, 4, 2, 0, 4, 4, -4, 3, -1, 4, 2, 3, -1, 0, -3, 0, 2, -2, 1, -4, -3, 0, -3, -4, -6, -2, -2, -3, 2, 0, 1, 0, -3, -2, 0, 0, 1, 0, 1, 4, 2, 3, -1, -2, -3, -3, 0, 2, 0, 0, -7, -5, 0, 1, -5, 1, -2, 0, -2, 0, 1, -1, 2, 0, 3, -1, 3, -1, -2, 0, 0, 4, -3, -1, 4, 0, -4, 1, -3, 0, -1, -7, -1, 0, 1, 2, -4, 2, -1, -5, -7, -7, -4, -1, -3, 0, 3, 4, -2, 1, 0, 0, -2, -3, 5, -1, 4, 3, -2, -1, 0, -3, -5, -3, -6, -5, -3, -1, -2, -3, 0, -6, -4, -2, -5, -4, -2, 4, 1, -1, 0, -3, 0, -4, -2, 2, 0, -1, 0, 0, 3, 1, 2, -4, -2, -3, -9, -3, 0, 2, -2, -2, -3, -4, -1, -7, -7, 0, -3, 0, 1, -4, -7, 0, -6, -1, -7, 0, 0, -3, 0, 2, 1, -1, -2, -7, -5, -6, -5, -7, -3, 2, 4, -2, -3, -4, -1, -5, -3, -1, -3, -1, -2, 0, -6, -3, 0, -4, 0, 0, -4, -1, 1, -6, -3, 0, -1, -5, -6, -8, -5, -2, 4, -1, 0, -2, 3, 0, -2, -6, 0, -2, -8, 1, -2, -7, -4, -1, -1, 0, -5, 1, 2, 0, -1, -4, 3, 1, -4, -4, -5, -3, -7, 0, -5, -2, 0, 4, 0, 1, -3, -6, -1, 0, -6, -2, 0, -3, -7, -4, -4, -7, -5, -10, -1, -4, 1, -3, -3, -3, -3, 1, -2, 0, -6, -1, -5, -4, -2, 3, 3, 0, 1, -4, -6, 0, -3, 2, -3, -3, -3, -10, -4, -4, -11, -11, 0, -1, 0, -1, 0, -2, -3, -4, -3, -1, 3, -1, 0, 2, 3, -2, -1, 4, 0, 1, 2, 3, -5, -5, -2, -5, -5, -4, -8, -6, -10, -8, -8, -8, 0, 0, 0, 0, -4, -3, 3, -1, 2, 2, -3, 1, -4, -2, 0, 2, -1, 4, 2, -1, -3, -4, 0, -4, 0, -9, -8, -8, -6, -14, -7, -3, -6, 0, 0, -3, -2, 0, 0, 5, 4, 2, -5, -4, -2, -2, -2, 2, 2, 7, 3, 1, -4, -4, -1, -7, -5, -2, -7, -13, -9, -7, -6, -2, -4, -3, 2, 2, 1, 0, 0, 2, 6, 1, -2, -5, -4, 3, 2, 2, 5, 1, 7, 5, -2, 3, 0, -3, -5, -7, -7, -11, -9, -5, -9, -6, -4, -4, 0, -1, 5, 3, 8, 5, 1, -1, 2, 0, 0, 0, 6, 6, 6, 5, 4, 1, -1, 0, 0, -1, 0, -3, -5, -6, -3, -3, -2, 0, 1, 4, 5, 3, 1, 8, 10, 9, 4, -1, 0, -6, -1, -1, -1, 7, 8, 2, 2, 5, 5, 1, 1, 0, 3, -1, 1, -3, -3, -2, 0, -3, 0, 0, 2, 0, 1, 0, 6, 2, 8, 5, -4, -5, -2, -1, 4, -1, 0, 1, 2, 3, 0, 4, 4, 5, 3, 0, 6, 3, 3, -3, -2, 0, -2, -1, 0, 7, 6, 7, 1, 1, 4, 0, -2, -3, -3, 0, -3, -3, 1, -1, 7, -1, 2, 4, 3, 2, 1, 4, 3, 4, 1, 2, 5, -1, 3, 1, 1, 5, 7, 3, 0, 2, 0, 1, -3, -3, -2, -8, -1, 1, 0, 2, 4, 0, 3, 3, 6, 5, 1, -1, 4, 0, 5, 7, 2, 2, 0, 0, 0, 0, 5, 2, 2, -2, 2, -2, -4, -5, -7, -7, -1, 0, -2, -5, 0, 6, 2, 0, 0, 5, 1, -2, 4, 3, 3, 2, 3, 5, 4, 2, 5, 3, 4, -2, 0, 2, 3, -3, -1, -4, -6, -3, -5, -6, 0, -4, 5, 0, 6, 1, 2, 1, 0, 5, 3, 4, 4, 0, 7, 0, 1, 0, 0, -1, -1, -4, -3, -1, 0, -3, -4, -11, -3, -7, -5, -6, -1, 1, -1, -1, 3, 3, 1, 2, 7, 6, 0, 1, 2, 7, 7, 0, 2, 0, 1, 2, -1, -3, -3, -6, -6, -8, -11, -7, -12, -5, -9, -5, -2, -5, 0, 1, 1, 4, -1, 4, 1, 3, -1, 0, 5, -1, 1, -3, 0, -1, -4, -3, -3, 0, -4, -1, -7, -3, -3, -4, -10, -4, -5, -7, -5, -4, 0, -2, 0, -1, -6, 1, 0, 3, 4, -2, 4, 1, 2, -4, -1, 0, 0, -2, 1, -3, -7, -10, -6, -6, -12, -11, -8, -3, -11, -5, -6, -7, -8, -4, -6, -3, -7, -3, -6, 0, -7, 0, -2, -6, -4, -7, -5, -3, -2, 0, -6, -3, -9, -6, -3, -7, -6, -10, 7, 4, 8, 8, 6, 3, 5, 8, 2, 3, 7, 5, 6, 8, 8, 6, 6, 4, 7, 6, 4, 1, 0, 3, 1, 5, 0, 4, 5, 3, 2, 7, 6, 9, 6, 9, 2, 7, 5, 4, 3, 8, 11, 9, 4, 4, 10, 7, 6, 10, 8, 4, 2, 5, 3, 2, 4, 2, 11, 4, 1, 2, 6, 9, 5, 6, 3, 6, 8, 9, 6, 8, 4, 7, 3, 6, 5, 4, 10, 7, 5, 4, 7, 4, 3, 5, 12, 9, 9, 8, 10, 11, 3, 9, 10, 8, 8, 8, 2, 7, 3, 11, 5, 8, 13, 12, 9, 6, 7, 11, 10, 9, 5, 7, 12, 9, 12, 12, 13, 7, 12, 8, 11, 10, 10, 10, 4, 4, 6, 4, 2, 4, 4, 3, 5, 5, 11, 10, 5, 5, 5, 12, 11, 10, 8, 12, 5, 11, 5, 8, 13, 10, 5, 5, 5, 4, 10, 5, 8, 5, 9, 3, 10, 10, 10, 10, 8, 11, 7, 13, 8, 10, 8, 9, 8, 8, 13, 7, 6, 9, 15, 13, 11, 12, 7, 7, 7, 10, 7, 7, 11, 14, 13, 6, 7, 7, 9, 6, 9, 14, 6, 15, 6, 9, 11, 15, 9, 9, 12, 13, 9, 11, 9, 10, 9, 11, 8, 11, 5, 11, 4, 7, 11, 10, 14, 13, 11, 6, 5, 6, 8, 11, 12, 10, 12, 11, 8, 13, 6, 13, 7, 11, 13, 8, 13, 12, 5, 7, 12, 7, 7, 12, 8, 5, 15, 13, 8, 5, 9, 7, 1, 5, 8, 6, 12, 12, 11, 11, 8, 11, 12, 12, 9, 13, 13, 9, 10, 12, 6, 10, 7, 12, 10, 9, 5, 6, 15, 9, 7, 7, 10, 2, 6, 6, 11, 5, 11, 9, 9, 6, 11, 13, 10, 14, 10, 11, 7, 6, 11, 6, 9, 10, 5, 12, 3, 6, 10, 8, 11, 16, 6, 6, 2, 4, 7, 8, 3, 9, 12, 8, 4, 9, 9, 5, 8, 6, 9, 14, 12, 13, 10, 12, 9, 12, 4, 5, 9, 3, 4, 4, 15, 10, 14, 8, 6, 2, 7, 0, 6, 9, 12, 10, 7, 7, 2, 8, 3, 6, 5, 8, 6, 11, 7, 8, 5, 11, 7, 2, 7, 0, 4, 3, 6, 17, 10, 7, 8, 8, 5, 6, 5, 8, 5, 6, 5, 3, 4, 7, 6, 2, 0, 7, 0, 6, 5, 5, 1, 5, 5, 6, 0, 7, 1, 10, 11, 15, 11, 12, 6, 9, 2, 4, 5, 7, 2, 1, 1, 3, 2, 2, 2, 0, 0, 0, 3, 1, 3, -1, 4, 9, 6, 3, -2, 7, 5, 8, 9, 13, 11, 11, 13, 3, 3, 4, 1, 6, 1, 2, 4, 3, 2, -3, -3, 2, -3, 3, -1, 5, 5, 1, 4, 1, 3, 2, -2, 3, 4, 9, 9, 14, 16, 13, 11, 7, 7, 0, 3, 6, -1, 0, 2, -4, -5, 0, -6, -6, -5, -5, -5, 2, -1, 6, 1, 5, -1, 5, 5, 6, 1, 6, 8, 15, 8, 11, 9, 4, 8, 2, 7, 4, 5, 3, 6, -1, 0, -1, -8, -6, -7, -7, 0, 0, 0, 3, 5, -1, 1, 4, 7, 7, 5, 13, 7, 12, 10, 8, 12, 5, 5, 9, 2, 3, 6, 4, -1, 0, -3, -10, -3, -8, -5, -9, -7, 0, -3, 6, 3, 3, 3, 3, 10, 5, 5, 13, 11, 6, 9, 13, 10, 13, 7, 8, 5, 12, 1, 4, -2, 3, -1, -3, -7, -5, -5, -3, -3, -1, 5, 3, 2, 10, 6, 12, 13, 10, 12, 8, 10, 8, 11, 6, 8, 12, 13, 8, 8, 8, 4, 0, 5, 2, -2, 0, -5, -5, -4, -6, -7, 4, 5, 5, 4, 9, 7, 7, 8, 11, 14, 7, 5, 13, 11, 9, 13, 12, 11, 9, 13, 7, 4, 7, 8, 6, 5, -3, 1, -8, -3, -5, 0, 3, 4, 4, 7, 11, 14, 9, 11, 11, 10, 11, 11, 3, 3, 11, 15, 9, 13, 13, 15, 8, 9, 4, 6, 2, 10, 2, 3, 2, 1, 0, -1, 8, 6, 11, 9, 9, 18, 13, 18, 19, 17, 12, 4, 3, 6, 8, 9, 16, 13, 16, 15, 10, 8, 14, 11, 7, 3, 11, 5, 4, 0, 8, 7, 9, 10, 10, 9, 9, 12, 14, 19, 18, 14, 9, 11, 2, 2, 4, 7, 10, 14, 11, 9, 9, 13, 13, 15, 10, 11, 7, 10, 13, 5, 9, 6, 8, 13, 11, 8, 12, 17, 19, 16, 16, 10, 10, 11, 2, 7, 10, 7, 14, 8, 11, 16, 8, 10, 14, 10, 7, 9, 7, 7, 14, 8, 11, 9, 13, 13, 10, 16, 9, 16, 14, 14, 16, 7, 9, 3, 6, 6, 9, 8, 11, 11, 12, 9, 9, 10, 15, 11, 9, 7, 12, 9, 11, 11, 17, 13, 10, 15, 14, 9, 13, 14, 7, 10, 7, 14, 3, 8, 6, 4, 5, 1, 8, 8, 7, 8, 12, 11, 17, 13, 14, 15, 8, 12, 16, 8, 12, 13, 11, 12, 12, 11, 15, 10, 13, 14, 8, 13, 7, 2, 6, -2, 4, 3, 2, 6, 13, 7, 13, 17, 7, 8, 10, 16, 11, 8, 8, 12, 11, 15, 16, 11, 15, 11, 11, 12, 6, 10, 10, 7, 8, 2, 5, -3, 0, 6, 2, 6, 6, 8, 8, 8, 8, 11, 11, 14, 9, 13, 9, 13, 11, 12, 12, 12, 9, 7, 9, 10, 5, 8, 3, 7, 3, 4, 2, 0, 5, 0, 4, 10, 9, 10, 7, 13, 9, 6, 15, 8, 12, 13, 14, 16, 11, 8, 14, 5, 6, 4, 8, 7, 6, 1, 2, 3, -2, -1, -1, 1, -4, 3, 2, 8, 8, 4, 9, 7, 10, 11, 8, 9, 8, 11, 12, 10, 6, 13, 10, 10, 9, 3, 11, 10, 5, 5, 6, 0, -1, -1, -2, -3, -3, 1, 1, 0, 3, 0, 5, 7, 3, 3, 2, 8, 4, 3, 9, 3, 4, 5, 0, 8, 7, 3, 6, 0, 1, -1, 0, 2, -1, -1, 1,
    -- filter=0 channel=1
    0, 1, 6, 4, 1, 8, 1, 7, 6, 6, 4, 5, 9, 6, 7, 3, 8, 8, 8, 8, 4, 5, 6, 8, 4, 7, 9, 4, 3, 8, 4, 6, 0, 5, 8, 3, 6, 3, 2, 5, 2, 3, 3, 10, 6, 3, 6, 1, 1, 6, 5, 5, 2, 7, 7, 3, 2, 2, 3, 8, 8, 6, 4, -2, -2, 2, 1, 7, 7, 7, 1, 7, 7, 5, 10, 8, 5, 0, 7, 7, 5, 2, 0, 5, 3, 9, 1, 3, 1, 8, 8, 5, 5, 6, 7, 0, -5, 1, 3, 1, -2, 5, 3, 3, 4, 5, 7, 6, 2, 1, 3, 2, 4, 6, 0, 2, 3, 7, 1, 8, 0, 1, 3, 5, 5, -1, 4, -1, 1, 5, 1, 3, -1, 6, 6, 1, 4, 4, 3, 0, 4, 0, 2, 5, 0, -2, 0, 7, 4, 2, 6, 4, 4, 2, 1, 2, 7, 6, 2, 0, -1, -1, 2, 3, -1, -1, -2, -2, 0, 3, 0, 5, -3, 0, 0, -5, 1, -1, -3, 4, 2, -2, 5, 0, 5, 0, -2, -2, 2, -1, 0, 0, 5, -1, 6, 0, 3, -1, 1, -4, 3, 0, -3, -2, -5, -4, -1, -8, -5, -4, -7, -5, -4, -3, -3, 0, -3, 2, 2, 0, 3, -1, 0, 1, 1, 6, 3, 2, 4, -2, 3, -4, 0, -1, -7, -8, -2, -7, -8, -3, -5, -6, -10, -7, -9, -6, 0, 0, -1, 0, 2, -2, 2, -2, 4, 2, 4, 5, 5, 5, -1, -4, -6, 0, -7, -6, -6, -13, -10, -13, -12, -10, -7, -13, -7, -9, -11, -7, -10, -2, -2, 0, -6, 4, 1, 5, 0, 3, -1, 0, 9, 8, 1, 2, -2, 0, -2, -8, -8, -9, -8, -16, -16, -17, -16, -15, -9, -7, -7, -6, -9, -3, -6, -6, -1, -1, 7, 2, 2, 2, 0, 0, 9, 2, 0, -3, 1, -5, -4, -7, -5, -11, -7, -11, -16, -13, -10, -9, -14, -13, -6, -8, -3, -1, 0, -2, 0, 2, 9, 5, 3, -2, 3, 7, 9, 2, 4, 0, 1, 1, -2, -4, -7, -3, -7, -12, -10, -7, -3, -7, -3, -2, -8, -3, -3, -2, 4, 0, 2, 8, 6, 2, 6, 0, 6, 2, 10, 3, 9, 5, 6, 9, 5, 2, 2, -1, -6, -2, -4, -6, -1, 0, -1, -4, 0, -3, -2, 1, 3, 11, 11, 10, 11, 10, 7, 3, 6, 1, 8, 7, 4, 6, 13, 9, 10, 7, 7, 2, 1, 3, 4, 0, 6, 4, 4, 4, 5, 5, 2, 4, 4, 7, 5, 8, 5, 8, 7, 1, 0, 3, 2, 10, 7, 13, 16, 9, 11, 9, 12, 13, 4, 5, 9, 12, 5, 9, 8, 4, 9, 11, 8, 10, 13, 7, 9, 5, 5, 10, 3, 4, 2, 6, 0, 5, 6, 12, 12, 14, 13, 16, 12, 6, 7, 11, 10, 7, 14, 14, 11, 6, 9, 9, 12, 12, 7, 11, 13, 8, 4, 3, 9, 3, 6, 5, 4, 9, 8, 13, 5, 15, 15, 10, 7, 7, 11, 13, 12, 10, 8, 5, 8, 9, 9, 6, 5, 4, 4, 8, 7, 4, 3, 0, 3, 7, 2, 4, 3, 5, 1, 0, 2, 7, 8, 11, 5, 3, 9, 11, 7, 3, 6, 7, 4, 9, 5, 6, 5, 0, 3, 3, 1, 2, 5, 4, 1, 4, 11, 1, 5, 0, -4, 2, -3, -1, 1, 4, 5, 8, 2, 6, 4, 0, 5, 2, -1, 2, 0, 0, -2, 4, 4, 0, -1, 0, -2, 1, 1, 2, 6, 2, 4, 0, -7, -5, 1, 2, -4, 2, 0, 1, 3, 5, -1, -2, -2, 4, 1, 5, 3, 2, 3, 1, 0, -5, -4, -4, -4, 4, 8, 4, 13, 10, -1, 1, -1, -5, -3, -3, 0, -3, -2, 1, 2, 2, -2, -1, 0, -5, -4, -4, -4, -3, -7, -3, -7, -10, -8, -2, -5, -3, 5, 12, 15, 5, 1, -1, -1, -2, -1, -7, -6, -6, -3, 0, 0, -6, -9, -6, 0, -7, -7, -1, 0, -7, -7, -7, -3, -11, -11, -7, -6, -1, 7, 13, 9, 11, 1, 0, -9, -7, -5, -7, -7, -5, -3, -8, 0, 0, -7, -4, -5, -5, -1, 0, -7, -9, -7, -9, -12, -8, -4, -10, 0, 5, 2, 10, 17, 3, 0, 1, -8, -6, -2, -9, -8, -6, -12, -4, -5, -2, -12, -11, -4, -6, -10, -7, -3, -10, -8, -13, -12, -9, -5, -7, -4, 2, 4, 11, 14, 6, 0, 0, -7, -11, -12, -9, -11, -8, -9, -10, -5, -13, -5, -5, -13, -11, -9, -12, -14, -14, -16, -13, -7, -14, -5, -7, -4, 0, 8, 10, 18, 8, 6, -1, -2, -5, -3, -7, -14, -8, -6, -12, -14, -14, -13, -14, -11, -8, -15, -14, -10, -16, -12, -8, -12, -7, -6, -8, 0, 4, 11, 13, 12, 7, 3, -6, -9, -6, -7, -12, -6, -6, -11, -12, -11, -14, -14, -13, -11, -14, -16, -11, -16, -13, -8, -4, -4, -8, -7, -6, -1, 2, 4, 12, 16, 12, 5, 3, -4, -6, -2, -8, -4, -6, -9, -8, -16, -18, -10, -12, -14, -16, -16, -12, -9, -6, -3, -2, -4, -8, -7, -6, 1, 0, 10, 12, 7, 7, 3, 3, 1, -5, -3, -2, -3, -5, -5, -6, -11, -11, -10, -13, -16, -8, -6, -5, -9, -7, -1, 0, -2, 1, 0, 1, 6, 7, 10, 15, 11, 12, 11, 8, 3, 1, 2, 2, -4, -5, -1, -7, -7, -5, -5, -6, -7, -6, -5, -8, -8, 2, 3, -1, 0, 5, -1, 5, 3, 13, 10, 14, 12, 6, 8, 10, 2, 8, 5, 3, 6, 2, 0, -1, -2, 1, -3, 1, -1, -3, -1, 0, 4, 3, 4, 2, 8, 2, 10, 9, 9, 14, 10, 16, 12, 13, 7, 5, 11, 11, 2, 3, 8, 6, 6, 6, 0, 3, 2, -2, -1, 3, 0, 2, 5, 3, 6, 8, 2, 11, 7, 13, 11, 5, 14, 6, -6, 0, -2, 0, -4, 0, -5, 2, -1, 0, -1, 0, 1, -1, 1, 0, -4, -2, -1, -1, -2, 0, 0, -2, -1, 0, 2, -4, -1, -2, -1, 0, -2, 0, -4, 1, -3, -3, 3, 0, 2, -3, -1, 5, 1, 0, 0, -3, 1, -6, 0, -4, 1, 2, 0, -1, 3, -1, 2, 0, -4, -4, 0, -2, -7, -6, 1, 1, -2, -5, -6, -5, -3, 5, 4, -2, 3, -2, -3, 1, -3, -2, 0, -4, -2, -1, 0, 3, -5, 3, -1, -1, -5, -2, 1, -7, -4, -1, 0, -1, 0, -4, -6, 1, -3, 2, 4, -1, -2, -3, -1, 0, 0, 0, 3, -1, -4, 1, 1, 0, -6, -2, -2, -1, 1, -1, 0, -5, -2, -2, -6, 1, -6, -3, -5, -2, 0, 2, 0, -2, 2, -5, -4, 1, 1, -3, -2, -2, 3, -4, 2, 0, -1, 0, 1, -7, 0, -5, -2, -8, -9, 0, -6, 1, -5, -2, -7, -6, -6, 0, 0, -5, 0, -3, 0, 2, -1, 3, -5, 1, 0, 0, -1, 0, 2, -2, -6, -3, -2, 0, -7, -1, -6, -2, 2, -4, 2, -1, -1, -2, 0, -6, -3, -4, -4, -1, 0, -1, 1, -5, -1, -5, -3, -5, -4, -4, 0, -1, -7, -4, 0, -7, -5, 0, -6, -3, 0, 2, -4, -2, -5, 0, -5, -7, -5, -3, -4, -5, -4, 0, -6, -1, -3, -4, -4, -3, -5, 1, -3, -6, -9, -4, 0, 0, 0, -8, -4, -5, 3, 3, -2, -2, -4, -7, -8, -3, -3, -5, -2, -5, -7, -3, -7, -4, -9, -2, -8, 0, -7, -7, -8, -1, -6, -2, -3, -5, 0, -7, -4, 2, 0, 4, -2, -5, 0, -5, -4, -4, -8, -9, -1, -7, -9, -5, -8, -2, -1, -8, -7, -4, -6, -3, -5, 0, -1, -3, -3, 3, -4, -4, -4, -1, 4, 0, 1, 0, 1, -4, 0, -5, -5, -2, -5, -9, -1, -8, 0, -1, 1, -4, -4, -4, -6, -5, -5, 3, -1, 1, 2, 1, -1, -8, -2, 1, -1, 2, 0, -4, -3, -4, 0, 1, -6, 1, -3, 0, 1, -3, 2, -4, 3, -3, 0, 3, 2, 0, 0, 0, 6, 0, 0, 3, 0, -5, 0, -1, 4, 2, 1, 1, 1, 7, 4, -2, 5, 3, 2, 2, 5, 0, -1, 1, 6, 2, 3, 2, 2, 7, 3, 3, 2, 6, 4, 0, 2, -1, -6, -6, -4, 2, 1, 3, 2, 9, 8, 7, 7, 7, 8, 10, 7, 5, 11, 4, 4, 3, 10, 10, 4, 10, 9, 3, 3, 6, 3, 3, 0, 1, 1, -6, -1, 2, 1, 2, 6, 10, 3, 9, 4, 11, 5, 11, 10, 6, 11, 12, 8, 4, 4, 11, 3, 1, 3, 2, 4, 3, 0, 3, 0, 0, 1, 1, 0, 3, 1, 7, 1, 10, 7, 10, 4, 8, 11, 5, 8, 14, 8, 14, 5, 12, 12, 1, 9, 0, 5, 2, 4, 0, 0, 4, -5, -2, 2, 3, 1, 0, 2, 5, 6, 2, 8, 0, 2, 1, 8, 9, 7, 4, 6, 5, 4, 6, 8, 1, 4, -2, -2, -1, 0, -3, -3, 2, 0, 0, 0, 1, 2, 0, 0, -7, -4, 0, 1, 3, 2, 6, -1, 6, 1, 4, 5, 1, -2, 0, -2, -2, -6, -2, -5, -3, -1, -4, -7, 0, 0, 0, 2, 5, 0, -4, -8, -8, -5, -8, -3, -4, 0, -3, 4, 0, 0, -1, -4, -2, 0, 0, 1, -6, 0, 0, -7, -8, -6, -10, -3, -5, 0, 0, 5, 0, 1, -7, -12, -12, -10, -6, -11, -7, -6, -7, -5, -6, -1, -1, -5, -5, -1, -4, -5, -5, -10, -7, -7, -6, -12, -12, -5, -1, 0, 8, 4, 1, 1, -7, -8, -12, -10, -6, -8, -12, -7, -7, -10, -11, -8, -10, -10, -11, -4, -4, -6, -7, -11, -11, -11, -11, -6, -11, -4, -2, 2, 9, 10, 0, -3, -4, -8, -12, -13, -13, -11, -12, -10, -8, -6, -11, -8, -8, -11, -6, -8, -3, -3, -3, -7, -8, -9, -15, -10, -4, -9, -5, 2, 9, 8, 0, 2, -6, -3, -9, -5, -6, -7, -10, -10, -5, -12, -11, -8, -8, -11, -8, -5, -5, -2, -11, -7, -13, -6, -11, -8, -5, -10, 0, 2, 9, 10, 1, -1, -8, -6, -7, -7, -5, -13, -12, -12, -12, -7, -4, -12, -12, -7, -7, -8, -5, -9, -13, -11, -8, -9, -8, -7, -11, -7, -1, 1, 3, 6, 2, 2, -2, -8, -11, -11, -13, -14, -7, -14, -13, -11, -9, -9, -11, -10, -9, -11, -9, -14, -13, -17, -15, -14, -14, -7, -10, -7, 4, 9, 9, 7, 5, 4, -4, -10, -6, -10, -6, -9, -9, -7, -9, -15, -10, -12, -12, -11, -12, -11, -12, -15, -13, -14, -9, -9, -10, -6, -10, -7, 3, 1, 14, 6, 11, 5, -2, -8, -9, -8, -9, -6, -11, -6, -6, -14, -16, -11, -11, -17, -12, -14, -17, -17, -13, -12, -6, -4, -4, -3, -2, -3, 4, 7, 9, 9, 10, 2, -6, -7, -11, -4, -11, -9, -6, -11, -12, -12, -9, -10, -15, -11, -18, -11, -9, -8, -10, -5, -7, -2, -5, -7, 1, -3, 0, 8, 6, 6, 8, 6, 2, -2, 0, -1, -7, -7, -8, -10, -8, -14, -11, -15, -8, -10, -13, -8, -10, -3, -2, -1, 1, 2, -4, -4, 3, 0, 5, 6, 13, 12, 9, 8, 5, -3, 3, 1, 0, -5, -3, -2, -1, -4, -5, -4, -5, -10, -7, -7, -1, -1, -2, 1, 0, 5, 2, 0, 1, 4, 8, 10, 6, 11, 5, 9, 1, 0, 4, 0, 4, -1, 3, 3, 0, -2, 0, -4, -5, -6, 0, 0, 0, 3, -2, 0, 4, 4, 4, 10, 4, 8, 10, 5, 13, 8, 5, 3, 10, 5, 5, 1, 7, 0, 2, 0, 6, 7, 0, 6, 4, 5, 0, -1, 0, 3, 7, 1, 5, 1, 6, 9, 10, 3, 12, 7, 6, -9, -5, -10, -3, -5, -3, -9, -5, -10, -2, -3, 0, -2, -5, -3, -8, -6, -2, -3, -8, -8, -1, -6, -1, -7, -1, -3, -8, -2, -10, -6, -10, -9, -6, -8, -5, -5, -6, -2, -2, -5, -9, -1, -5, -7, -7, -1, -6, -2, -8, -10, -4, -8, -3, -5, -7, -2, -4, -2, -4, -4, -10, -7, -8, -6, -12, -11, -3, -3, -9, -7, -6, -7, -6, -6, -7, -8, -2, -10, -3, -5, -5, -11, -6, -3, -8, -8, -2, -8, -7, -5, -9, -7, -2, -7, -10, -7, -7, -6, -9, -5, -10, -4, -6, -1, -1, -3, -3, -2, -1, -5, -7, -1, -4, -9, -2, -10, -8, -9, -5, -2, -8, -10, -6, -4, -8, -6, -8, -8, -9, -5, -9, -5, -11, -3, -7, -6, -7, -2, -5, -3, -5, -6, -6, -5, -5, -2, -2, 0, -7, -1, -4, -4, -7, -6, -10, -8, -11, -10, -10, -8, -11, -3, -9, -4, -10, -6, -1, -8, -5, -1, -4, -5, -6, -2, 1, -1, 0, 1, -5, -6, -6, -4, 0, -4, -6, -3, -10, -4, -8, -7, -13, -8, -9, -6, -1, -5, -6, -3, -3, -3, -6, -5, -5, 0, -2, 1, 0, -1, 0, 0, -5, 1, -6, -6, -3, -4, -6, -10, -1, -11, -12, -10, -4, -6, -11, -4, -8, -5, -6, -7, -3, -5, -3, -5, 2, 1, -3, -3, 5, 0, 0, 3, -2, 2, 1, -2, 0, -7, -10, -9, -3, -6, -7, -10, -5, -7, -1, -8, 0, -7, -2, 0, -5, -8, -5, 2, 3, -1, 0, 5, 0, -1, 6, 1, 4, 3, 2, -5, -5, -5, -3, -1, -6, -2, -5, -4, -10, -8, 0, -4, -4, -2, -6, 2, 0, -3, -6, 1, 0, -1, 3, 2, 5, 5, 2, 3, 1, 0, 6, 5, 1, 3, 0, 2, 2, 0, -2, 0, -7, -3, 0, -2, 0, 0, 1, 0, 4, -1, 0, 2, 5, 6, 9, 3, 8, 7, 8, 8, 7, 3, 2, 3, 2, 6, 2, 3, 6, 1, 0, -2, -6, -6, -5, -2, -3, -1, 0, 0, 4, 4, 1, 5, 11, 11, 11, 11, 7, 14, 8, 9, 9, 11, 14, 4, 6, 4, 3, 6, 2, 3, -2, -5, -9, -8, -2, 0, 1, 1, 7, 9, 12, 7, 9, 13, 16, 15, 17, 15, 18, 13, 15, 17, 16, 13, 15, 14, 11, 11, 11, 13, 7, 9, 0, 1, -9, -5, -1, 2, 2, 5, 9, 9, 15, 13, 19, 15, 18, 16, 23, 23, 22, 25, 18, 20, 19, 21, 18, 17, 12, 12, 19, 17, 10, 6, -1, 2, -8, -7, -1, -2, 6, 8, 13, 13, 19, 13, 17, 21, 22, 26, 27, 22, 29, 24, 22, 21, 22, 23, 21, 16, 19, 20, 12, 11, 9, 11, 0, 3, -7, -2, -3, 1, 7, 10, 11, 10, 16, 14, 14, 17, 16, 20, 25, 26, 23, 21, 23, 21, 22, 21, 15, 17, 13, 14, 10, 16, 12, 7, 8, -1, -5, -4, 2, 4, 5, 2, 6, 15, 17, 12, 18, 21, 20, 15, 20, 17, 19, 24, 23, 26, 19, 22, 14, 15, 15, 7, 12, 13, 7, 4, 8, 0, 0, 4, 0, 3, 2, 8, 3, 8, 7, 11, 10, 14, 13, 14, 19, 13, 12, 14, 17, 15, 15, 12, 14, 11, 4, 6, 11, 2, 3, 9, 7, 0, -1, 0, 3, 3, 4, 5, 0, 5, 2, 6, 9, 9, 7, 8, 14, 16, 13, 12, 12, 10, 13, 10, 5, 4, 7, 4, 0, 1, 2, 4, 5, 3, 6, 5, 8, 6, 4, -4, 2, 2, 0, 1, 3, 5, 4, 8, 9, 12, 4, 6, 3, 6, 8, 6, 5, 6, 6, 3, 0, -3, 2, 0, 6, 6, 1, 4, 1, 0, 2, 0, 0, 5, -1, 3, 2, 0, 6, 0, 3, 1, 1, 0, 2, 2, 4, 0, 2, 0, 2, 0, -4, 0, 0, -3, 0, 10, 7, 9, 1, 2, 0, 0, 0, 2, 1, 3, 3, 4, 5, 5, 0, -4, -2, 2, 6, 1, 4, 1, 0, 4, 1, 0, -3, -4, -3, -3, 0, 4, 8, 13, 3, 4, -4, -5, 2, 1, 0, 1, 0, -4, -3, -1, -3, 1, -5, -2, 0, 1, -1, 0, 0, -6, -1, -2, -1, -5, -1, 0, 1, 10, 6, 12, 7, 6, 0, 0, -5, -2, -4, -3, 0, -2, -5, -3, 2, 0, -4, 0, -1, -1, -1, -2, -4, -2, -1, -6, -9, -3, 1, -6, 0, 7, 14, 9, 6, 2, -1, -4, -3, -1, -7, -2, -3, -7, -5, -7, -1, -5, -4, 1, 0, -5, -2, 0, -8, -4, -7, -4, -6, -8, -6, -3, 2, 11, 15, 12, 4, 5, -3, 0, -6, -6, -4, -10, -6, -6, -7, -6, -4, -2, -7, -7, -8, -3, -9, -9, -6, -10, -6, -1, -2, -1, 0, 0, 6, 9, 8, 15, 10, 2, -1, 0, -7, -6, 0, -1, -2, -6, -5, -10, -6, -8, -7, -6, -9, -12, -9, -4, -2, -7, -5, -7, -2, -6, -3, 4, 2, 8, 9, 12, 6, 5, 1, -2, 0, -5, -5, -4, -5, -7, -8, -6, -9, -7, -10, -4, -8, -13, -5, -3, -4, -2, -1, 2, 2, 0, -3, -1, 3, 11, 15, 15, 13, 3, 0, 1, 0, 0, -1, 0, -2, -4, -1, -8, -10, -10, -10, -3, -4, -6, -3, -3, 1, 0, 1, 0, 2, 4, 7, 3, 11, 11, 15, 12, 9, 4, 8, 1, 0, 4, 3, 6, -2, -1, 0, 1, -7, -7, -2, -6, -3, -4, -2, -3, 0, 3, 3, 8, 2, 8, 2, 8, 7, 11, 15, 6, 6, 8, 9, 4, 7, 10, 8, 6, 7, 5, 1, 1, 2, 4, -1, 5, 0, 3, 5, 8, 4, 9, 3, 11, 6, 12, 7, 6, 9, 9, 15, 9, 9, 11, 8, 11, 5, 12, 9, 7, 9, 3, 3, 3, 2, 5, 6, 2, 2, 1, 4, 7, 12, 5, 12, 5, 13, 6, 11, 13, 8, 11, 9,
    -- filter=0 channel=2
    3, 0, 0, 4, 4, 0, -1, 0, 3, 0, 3, -1, -2, 0, 2, -4, -1, 0, 0, 0, -3, 3, 1, 1, 4, -2, -1, 0, 0, -2, 1, 0, -1, -1, 1, -3, 0, -2, 3, 0, -2, 1, 2, -4, 0, 0, -2, -1, 0, 3, 0, -3, -3, 0, -3, -4, 2, -2, -1, 0, 0, 0, -3, 3, 4, 3, 1, -3, 0, -1, -2, 1, -1, 3, -2, 0, -3, 3, -3, -4, 1, 3, 3, 4, 3, -2, -1, 0, 0, -1, 1, 0, 3, 3, 1, 1, 0, 2, 4, 1, -2, 1, 0, 4, 1, -2, -2, 1, 1, 0, 3, -3, 3, -1, 1, 0, -1, 3, 0, 0, -3, -4, 0, 0, -3, 4, -1, -1, 4, -2, 3, 4, 1, 0, 1, 2, 2, 3, -1, -1, 0, 0, 4, 0, 2, 3, -1, -4, 0, 2, 0, 2, 0, 0, -2, 0, 1, 2, 2, -2, -2, 4, -3, -3, -1, 0, 4, 0, -3, -2, -1, 0, 0, -4, 0, -3, -1, 3, 4, 0, -3, -2, -3, 0, 1, -4, 0, -1, 1, 1, 0, -1, 0, -1, 2, -3, -3, 3, 4, 0, 0, 0, 4, -3, -3, 1, 3, -2, 0, 4, 3, -1, 0, 3, 2, 3, 2, -1, -3, 0, -2, 1, 0, -1, 0, -1, 0, 1, 0, -1, 1, 0, -2, 0, -3, 0, 3, 0, -1, 2, 4, 4, -2, 1, -2, 3, -4, -3, -4, 4, -3, 3, 5, 5, -1, 2, 0, 1, 1, 3, -3, -3, 1, 2, -1, -4, 1, 3, -1, -2, -2, -2, 3, -4, 3, -3, -1, 3, -4, 2, 0, 2, -2, -3, -2, -1, 0, 3, -1, 3, 1, 0, 4, 5, 0, 1, 3, 1, -2, -3, -4, 0, -1, 0, 0, -2, -1, 3, 0, 0, 4, -3, 0, -1, 0, 4, 0, 0, 0, 4, -2, -2, 0, -2, 0, -1, -3, 1, 4, -1, -3, -2, -2, -2, 0, -2, 2, 3, 3, 0, -3, 0, -1, 4, 0, 3, -2, -3, -3, 0, -1, 0, 4, -2, 4, 5, -3, 2, 0, 4, -4, 2, -1, 0, -1, -5, -5, 0, 3, 3, 0, 0, -5, -2, -3, 0, -3, -3, -3, 3, 5, 1, 0, 0, -2, 4, -3, 1, 2, 0, -3, -3, -2, 1, 3, 0, -4, -3, -2, 1, -3, 0, -4, -4, 2, 0, -2, 0, 3, 3, -2, -3, 4, -1, -1, -3, 1, 5, 4, 0, 1, 2, 4, 3, 2, -5, 0, -2, 2, -2, 0, -6, -6, -5, 0, 0, -1, 0, 0, -1, -1, -3, -4, -3, -1, 3, 1, -2, 1, -2, -3, 0, -2, 0, -2, -1, -2, -3, -1, 0, -5, -3, -2, 1, -5, -5, -3, 1, 0, -5, 2, 0, -3, -1, 3, 0, -1, -2, 2, 0, 0, 3, 2, -3, 4, 0, 0, -1, 0, -4, -5, -6, -2, -4, -5, -1, -2, 1, -4, -4, 1, 1, 0, 0, 0, 3, 0, 4, 0, 4, -1, 4, 1, 1, 2, -3, 0, -1, -1, -2, 2, -1, 2, -3, 0, -6, -1, -4, -2, 0, 0, 0, -1, -1, 2, -4, 2, 2, 2, 0, 1, -3, -1, 2, 3, 0, -2, -2, -1, -2, -3, -2, 0, 0, -4, -4, 0, 0, -2, -3, 0, -4, -5, 0, -5, -3, -3, -2, 2, 0, 1, 0, 3, -1, 0, 0, 1, 4, -2, 2, 5, 0, 3, 1, -2, 1, 2, 2, -5, -3, -7, -5, 0, -5, 0, 2, 0, -4, -1, -4, 0, -4, -1, 0, 3, -2, -3, 1, -2, 4, 5, 0, -2, 0, -2, -4, -3, -4, -2, -5, 0, -5, 0, -5, 0, 0, 0, -6, -6, -3, -2, 2, -3, 3, 4, 4, 0, 0, -1, -3, 3, -2, 4, 3, 1, 4, 1, 0, 1, 1, 3, -1, 2, -1, -5, 1, -5, 1, -4, 0, -4, -4, 0, 1, -3, -1, -2, -1, -3, 3, -2, 0, -1, 0, -1, -2, -1, -3, 0, 1, -4, 0, -1, -5, -4, -1, 1, -5, -1, 2, 0, 1, 2, 0, 3, 0, 0, -2, 0, 0, 4, 4, 4, 4, 3, 0, 3, 1, -3, -2, 0, 0, 2, 2, 0, 0, -5, 1, 1, -6, -3, 0, -1, 2, -1, 3, 2, -2, -1, 1, 0, -3, 2, -2, -2, -2, -4, 0, 2, 1, 0, 3, -3, 1, -4, 4, 4, -5, 1, -3, 0, 2, 0, -4, -4, 0, 2, 1, 1, 1, 2, -3, -1, 3, -1, 1, 3, 2, 0, 1, 1, -1, 4, -3, 2, 1, 4, 2, -2, -4, 1, -2, 4, -3, -3, -2, 1, 1, -3, 0, 1, 4, 0, 0, -3, 0, 3, -2, -2, 1, 1, 0, 3, 1, -1, 0, -3, -3, 1, 2, 3, 2, 0, 3, 0, -4, 0, 2, -1, 2, 2, 0, 2, 3, -2, 3, 2, 0, -2, 0, -1, 3, -3, -1, -2, 0, 1, -2, 3, 0, -2, 2, 2, -2, 1, 3, 0, 0, 4, -1, -1, 0, 2, -3, 2, 0, 1, 3, 2, 1, 0, -1, -4, 1, 3, 0, 3, 3, -1, 4, 2, 1, 0, 3, 3, -2, 3, 3, 2, 0, 2, 3, 3, 0, 0, 1, -4, 0, -2, -3, 0, 1, 1, -3, 1, 2, -2, 2, -2, 1, 3, 1, 2, -1, -2, 4, -1, 4, 4, 0, 2, -2, 3, -1, 1, -2, 1, 3, 4, -2, -3, 0, -3, -4, 0, -1, 2, -1, 1, 2, -1, -3, -2, 0, 3, -3, -1, -2, 0, 4, 0, -2, 3, -3, -1, -3, 3, -2, -2, 0, 2, -1, -1, -2, 4, -1, 3, 0, 0, 3, -3, 0, 1, -3, -4, -4, -1, -1, -2, -3, -4, -4, 2, 1, -3, 0, 0, 0, 1, -1, 2, 3, -4, -4, -3, 0, 0, 0, 0, -1, 0, 0, 0, -5, -4, -4, 0, 0, 3, -4, -5, -2, -1, -1, 3, 2, 1, 3, -3, -4, 0, 0, 0, -2, -4, 0, -3, -4, -5, 2, 3, -3, 1, 0, -3, -2, -3, 3, 4, 0, 0, -1, 3, -1, 1, 2, 2, -1, -3, 3, -3, -3, 2, -3, -3, 4, -1, 3, -3, 3, 0, 3, 0, -2, -1, 3, 0, 1, 1, -1, 2, 1, 3, -1, -2, -1, -3, -2, 0, -2, 3, 1, 0, 2, -1, 1, -2, -1, -2, 2, -1, 1, 4, 4, 4, 4, 0, -1, 0, -2, 1, 3, -2, 0, 0, 1, -2, 3, 2, 2, 3, 2, -1, -1, -2, 2, 0, 4, 2, 1, 2, -1, 1, -2, 0, -1, 1, 0, 2, -2, 1, 4, 2, 0, -1, 0, -3, 3, 3, 1, -3, 2, -1, 0, 2, 0, 1, -1, 0, -3, 4, -2, 2, 0, 1, 1, 0, 3, 1, 2, -2, -1, 1, 1, 0, 1, 3, 0, 0, 4, -2, -3, 1, 1, 0, 3, -1, -2, 2, -3, -2, -1, 1, 1, 2, 0, -1, 4, 2, -1, 0, 3, 4, 0, -3, -3, -1, 0, 1, -2, 2, 2, -1, 4, -2, -1, 0, -3, 0, 1, 1, 2, -3, -1, 1, -1, 0, -4, -1, 3, 0, -1, 0, -3, 3, 0, 0, 4, -2, 3, 2, 4, 1, -3, 4, 1, 3, 0, 3, 0, -1, -4, 1, -3, 4, -2, -1, 0, -2, 3, -1, 3, 3, 5, 4, 0, 3, -2, -2, 4, -1, 2, -3, 1, 0, 4, -1, 3, 0, -1, 4, 0, 0, 0, 0, -3, -3, 0, 3, 2, 4, 2, 4, -1, 4, 0, 1, 3, 2, 1, 5, 5, 2, 4, 0, 4, 5, -1, 0, -1, -1, -2, 4, -2, 4, 2, 0, 4, 0, -3, 3, 3, 3, 0, 0, -3, -2, 5, 2, -2, 0, 0, 5, 3, -1, 2, 5, 0, 3, 0, 0, 3, 5, 1, 1, 1, 3, 0, -2, 2, 2, 2, -1, 0, 3, 0, 3, 3, 2, -1, -1, -2, 0, 3, 3, 5, 6, 0, -1, 2, -1, -1, 0, -1, 0, 2, 2, -1, 3, -1, -4, -1, -1, -3, -1, 2, 2, -1, -1, -1, 0, 2, 1, 0, -3, 1, 0, -1, -1, 5, -2, 3, -2, 0, 3, -3, -3, -1, -1, -2, -5, -3, 2, -2, 0, 2, 2, 2, -2, -2, 3, 1, -3, 1, 3, -2, 1, -2, 2, 0, 5, 0, 4, 5, 4, -3, -1, -2, 1, 3, 1, -4, 2, 0, -1, -2, -4, 1, -3, 2, 3, 2, 5, -1, 1, 0, 3, 2, 2, 2, -2, 3, 1, -1, 3, 0, 0, -3, 2, 3, -1, 2, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -3, 4, -1, 0, -1, 1, 1, 2, 3, 3, -1, 0, 5, 4, 4, -1, 5, 3, 5, -2, -3, 0, -4, -4, -4, 0, -3, -6, 0, 0, 3, -3, 0, 2, 3, -1, 0, 5, 6, -2, 3, 5, 4, 3, 0, -1, 2, 2, -1, -2, 5, 1, 3, -1, 0, 2, 0, -4, -6, 2, 0, -4, -2, 0, 2, 2, 4, 2, 5, 1, 3, 2, 1, 0, 5, -1, 0, 1, 1, 0, 0, 0, 2, -1, 1, -5, 0, -2, 2, 2, -3, -4, -2, -4, -4, -2, 4, -2, 4, 1, -2, 5, 1, 1, 1, 5, 3, -2, -2, 0, 0, 5, -1, 0, -3, 0, 3, -1, -2, -2, 2, -5, -2, -4, 0, 0, 2, -2, 2, 0, 0, -3, 3, 3, 2, 0, 3, 3, 5, 4, 0, 1, 5, 0, -1, 4, 0, 2, -2, 1, -5, 0, -1, -4, -2, -4, -4, -4, -3, 2, -2, 3, -3, -1, -2, 3, 4, 2, 2, 0, -1, 3, 1, 6, 2, 4, 4, 2, 3, 0, 3, 0, -2, -3, 2, -5, 0, 0, 1, -1, -3, 1, -2, 1, 5, 4, 4, 0, 0, 4, 2, -2, -3, -3, -2, 2, -1, 2, 1, 1, 2, 3, -3, 2, 1, -2, -1, -5, 0, -2, -4, 3, 1, -3, 0, -2, -2, 0, 0, -2, -2, 1, 0, 4, 1, 3, -2, 2, 3, 1, 4, -2, 5, 1, 0, 0, 3, -1, 2, -4, 2, -1, -3, -1, 0, 0, 4, -3, 5, 2, -3, -2, 4, 0, 4, 1, 1, 0, -1, 4, 0, 1, 0, -1, 1, 0, -1, 2, -3, -3, 0, 0, -3, 1, 3, 0, -1, 0, 2, 4, 0, 2, -2, 4, 5, 3, 0, 2, 0, 0, 4, 2, 4, 2, 3, 0, 2, 0, -3, -1, 1, 1, 0, 3, 0, -3, 4, 0, 3, 3, 2, 0, 0, 2, 2, 0, -2, 4, 0, 4, 1, 2, -2, -3, 5, 1, -2, 4, 1, -2, 2, 4, 0, 2, -4, -2, 0, 0, 0, -1, -1, 0, -2, 0, -1, -1, -2, 5, 4, 4, 0, 2, 4, -2, -2, -2, 1, 3, 0, 0, 0, 0, 4, -2, 0, -2, 3, 0, 1, -1, 1, -1, 2, 1, 0, 0, 0, 1, 3, 3, 0, -2, 4, -3, 0, -1, 2, 0, -3, 5, -1, 0, 2, -3, 0, -4, -2, -1, 2, -3, 3, 1, 3, 1, 1, -1, 4, 1, 1, -1, -3, 3, -2, 3, -2, 4, 4, 0, -3, 0, 1, 2, -3, 3, -2, 0, 2, 4, 0, 2, 4, 3, 3, -3, 1, 3, -3, 1, 2, -3, -2, 0, -2, -3, 4, -3, -1, -1, 0, 3, 0, 2, -1, 3, -3, 3, 4, -3, 2, -1, -3, -3, 0, 1, -1, -3, -1, -1, 3, 0, 2, 0, -2, 0, -3, -4, 0, 4, 2, 1, -1, 3, -4, -1, 0, -2, 3, 2, 0, 1, -2, 2, -3, -2, -4, 2, 0, -4, -3, 2, -2, -1, 0, -3, -4, 2, -3, -4, 0, 1, 0, -1, -1, -1, 0, -1, 2, 2, 0, 0, 0, 4, -2, -1, 3, 3, 1, 2, -1, -1, -2, -4, -1, 3, 3, -3, -1, 2, 3, -1, 1, 1, -3, -3, -1, -1, 0, -1, -4, -2, 0, -3, 3, 3, 3, 0, 3, -1, -4, 0, 2, -3, 1, 3, -1, 0, 0, -2, -5, -4, -1, -1, 1, -1, 0, -1, -3, -3, -2, -3, 0, -5, -4, 1, 0, -4, 0, -3, -6, -6, 0, -6, -4, -3, 0, 0, 0, 0, -3, -3, -1, -6, -2, 0, -3, -2, -2, 1, -3, 0, -1, -3, -3, 0, -3, 0, -3, -1, -5, -1, 0, 1, 0, 0, 0, 2, -4, -2, -1, -4, -3, -5, -2, -4, -6, 0, -2, -5, 1, 0, 0, -4, -6, -5, -3, -3, -1, 0, 0, 1, -2, -1, -5, -2, 0, -4, -3, -5, -3, -4, -4, -5, 1, -1, -1, -1, -5, -6, -2, 0, -6, 0, -5, -1, -5, -3, 2, 2, 1, 2, -3, 1, 0, 2, -3, -2, -2, 0, -5, 1, 0, -2, -4, 0, -6, 0, -4, -4, 0, -3, 0, 1, -3, 0, -1, 1, -2, 0, -1, 1, 1, -3, 0, -2, 0, -4, 0, 0, -3, 0, -2, 1, 0, 0, -1, -4, -4, -1, -5, -5, 2, 0, 2, -5, 1, -2, -5, -4, 0, -3, -1, -4, -1, -3, -4, -3, 3, 2, 2, 0, 1, 0, -5, 0, -3, -4, 0, 0, -5, -4, 2, 0, 0, 0, -4, -1, 1, 3, 2, -2, 0, -3, 0, 3, -4, 0, 0, -1, -5, -2, -3, 0, -5, 0, -3, 0, -4, -4, -2, 2, -3, 1, -4, -2, -2, -3, -5, -2, 0, 1, 0, 3, 0, -2, -4, 1, 3, 1, -1, -2, 3, -2, -1, -1, -2, 1, -4, 0, 0, 1, -3, 3, 3, 0, 0, 2, 3, -4, 2, -1, 3, 1, -4, 0, 0, -2, -4, 2, 1, -3, -1, -3, 0, 1, -3, 2, 3, -1, -4, -4, 0, 1, -3, -2, 0, 0, 2, 0, -5, 0, 0, 0, -3, 2, -1, 0, 2, 1, 0, 3, 3, 0, 4, 0, 0, -1, 1, 1, 3, -1, 3, 2, -1, 1, -3, 3, -3, -1, -2, 2, 1, 1, 1, 0, -1, -4, -4, 3, 1, -4, 2, -2, 0, -3, -2, -2, 1, 0, -3, 0, 0, -3, 2, -4, 3, -2, -2, 3, 0, -4, -2, -1, 0, -3, 2, -3, -2, -3, -1, -4, 0, 0, 4, 1, -1, -2, -2, 1, 0, -4, 3, 1, -1, -2, 0, -3, 0, -2, -3, -4, 2, -2, 4, -4, -2, -2, 0, -4, -2, 2, -3, 2, -1, 1, 0, 4, -1, -2, -1, 1, 3, 2, 3, -4, -5, 1, -2, -4, 1, 0, 3, 3, -2, -1, 2, -3, 3, 0, 0, 3, 4, -1, -3, -3, 3, 0, 0, -3, 3, -3, -3, 0, 0, -2, 2, -2, 2, 0, 0, -4, -2, -2, -3, 2, -3, 2, 4, -2, 4, -2, 4, 0, 1, 3, 0, 2, -1, 3, 0, 3, -4, 4, -3, 1, 3, 1, 3, -3, -4, -5, -3, -3, 0, -3, -4, -2, 2, -2, 0, 3, 3, -4, 0, 0, -2, -4, -2, -3, -3, -2, 1, -1, 0, 2, -1, 0, 3, 1, -3, 3, 1, -4, -3, 2, 0, 1, -3, -5, -1, -4, -3, -2, 4, -3, 3, -1, 3, 0, 1, 1, -2, 1, -3, 0, -2, -2, -2, 0, 1, -5, 2, -1, -5, -1, 0, -3, -3, 2, -1, 3, 0, -3, -1, -2, 2, 0, -1, 2, 2, 2, -2, -1, -1, -4, 4, 2, -2, 2, 2, 0, -1, 2, -1, 1, -3, 1, -3, -4, 2, -2, 0, 0, -2, 2, 1, 4, -1, -2, -4, 3, 0, 2, 1, 3, -2, 0, 0, 2, 0, 0, -4, 1, -1, -1, 0, -2, 1, -5, 0, -2, -4, 0, -2, 2, -2, 0, 0, 3, 2, 4, 3, 2, -2, -3, 1, 0, 1, 2, -2, 1, -4, 3, -1, 2, -2, -3, 2, 0, 1, -1, -3, 1, -5, 0, -3, -4, 0, -1, 0, 1, -1, 3, -3, 0, 0, -4, 1, 2, -3, 0, -1, 1, 4, -1, -2, 0, -4, 0, 1, 0, 1, 0, 2, -2, -1, -5, -2, -1, -3, 0, 1, -2, 0, 4, 3, 0, 2, 0, -4, -2, 0, -3, 0, -1, -1, 3, -3, -3, 0, 0, -1, -4, -4, 0, -4, -4, 3, 2, -1, 4, -3, -3, -1, -3, 4, 4, -2, 0, 3, -4, -2, 4, -3, 3, 2, 0, 0, -3, -2, 4, 0, -3, -4, 2, 3, -2, 1, -3, 3, 0, -1, -1, -2, -1, -1, -1, 1, -3, 2, 4, 0, -3, -2, -3, -2, 0, -1, -2, 3, 0, 1, -3, -1, 4, 0, -4, -4, 0, 3, 3, -3, 0, 2, 1, 2, 1, -2, 0, 3, -3, -4, -1, -3, 1, -2, -2, 3, -2, -3, 0, -3, 0, -2, 1, -2, 0, -4, 3, 0, -1, -2, 3, -2, 4, 0, -3, -2, 3, 0, 0, -3, 0, 2, -4, 3, 0, -3, 0, -4, -2, 2, 3, 3, 0, -3, 0, 2, -3, 0, 0, -2, -2, 1, 0, 1, -2, 0, -2, -4, 0, 0, 2, -2, 1, 0, -2, -4, 1, -1, 0, 0, -2, -2, 3, 4, -2, 1, 1, 0, -3, 0, -1, 3, -2, -1, -4, 4, 0, 3, 3, 1, 0, -4, -2, -2, 0, 4, -5, -4, -3, 2, 1, 0, 1, -1, 3, 2, 2, 0, 0, 0, -4, -3, 0, 0, -2, 0, 1, 0, 3, -2, -3, -3, -2, -2, 1, 3, -2, -4, -4, -1, 0, -2, -4, -3, 0, 0, 1, 0, 0, -4, -1, 1, -3, -2, -1, 3, 0, 0, 3, 1, -3, -1, 2, -4, -2, 2, 2, 0, 3, -5, -3, 3, 2, -4, 0, -4, 0, 0, 2, -1, 3, 2, -3, 0, 2, 0, 0, -2, 2, -3, 1, -2, 1, 0, 3, -1, -2, 0, 2, -5, 0, -2, 1, -4, 0, 2, -3, 1, 0, -5, 2, 1, -2, 0, 1, 0, 2, -4, 1, 0, 0, -2, 1, 1, 2, 2, -4, -1, -4, -3, 1, 3, -2, -3, 2, -4, -3, 1, -3, -5, -2, 0, 2, -4, 1, 1, 0, -1, -4, -1, 0, 1, 0, -4, 0, -3, -1, 0, -1, -1, -5, 1, 0, 0, -4, -1, 0, -4, 1,
    -- filter=0 channel=3
    0, 0, 4, 5, 3, 0, 2, 4, 4, 4, 2, 0, 1, 4, 0, 1, 4, -3, 1, 3, -1, 0, 4, 0, 0, 4, 0, 0, 2, 1, 3, -2, 5, 4, -1, 0, 5, 5, 3, 1, -2, 3, -3, 2, 4, 1, 1, 0, 1, -3, -3, 5, 1, -2, -1, -1, 1, 1, 6, 4, 2, 1, -1, 3, 0, 2, 3, 2, 1, 4, 2, 4, 5, -1, -2, 2, 2, 0, 0, 1, -3, -1, -3, -2, 1, -2, 1, 4, 5, 5, 3, 7, 3, 1, 0, 4, -2, -1, 2, -1, 6, 6, 5, 4, 4, 0, 3, 0, -3, 0, 2, -2, 2, -4, 1, 1, -3, 3, 2, 0, 1, 0, 4, 2, 2, 1, -1, 4, 0, 6, 1, 5, 2, 5, 0, 0, -1, -2, 0, 0, -3, -1, -3, -2, -1, -5, -3, 0, -3, 3, 4, 1, 2, 3, 0, 2, 2, 0, 7, 3, 1, 7, 0, 4, 4, -1, 5, 1, 2, -1, 3, -2, -2, 0, -2, -5, -2, -1, -6, 0, 0, 0, -1, -2, 0, 1, 8, 0, 2, 2, 0, 6, 4, 5, 6, 3, 3, 5, 0, 4, 0, 2, -4, 1, 0, -6, -2, -2, 0, -4, -1, 0, 0, 0, 0, -2, 3, 1, 7, 1, 0, 2, 7, 2, 0, 6, 0, 2, 0, 2, 4, 3, 2, 0, 0, 3, 0, 0, -6, -4, -3, 0, 0, -2, -3, -5, 1, 0, 0, 6, 0, 7, -1, 1, 0, 6, 0, 5, 0, 2, 0, 0, 3, -1, 2, 1, 2, 2, 1, -5, -3, -5, 1, 0, 0, -5, -3, 0, 1, -2, -1, 0, 5, 2, 1, 1, 1, 3, 6, 3, 3, 0, 0, 5, 5, -1, -2, 2, 0, -2, -6, -1, -3, -3, -6, -6, -5, 0, -4, 2, 0, 3, 2, 0, 1, 4, 7, -1, 7, 4, 7, 4, 5, 1, 6, 0, 1, -2, 1, 0, -4, 0, 1, -2, -4, 0, -4, -5, 0, 0, 2, -5, -1, 0, 0, -2, 4, 2, 0, 2, 0, 5, 5, 1, 0, -1, 4, 2, 0, 0, 1, 0, 0, 2, 0, -1, -1, -4, -4, -2, -3, -4, -1, 0, 2, -3, 0, 3, 2, 6, 0, 0, 2, 2, 3, 4, 6, 0, 0, 2, 2, -1, 0, -1, -1, -5, 2, -4, -2, -3, -6, -5, -2, -4, -3, 0, 1, -2, 1, 0, 3, 2, 6, 6, 1, 6, 3, 0, 2, 0, 3, 1, -1, -4, -4, 2, 2, -5, -3, 0, 0, -4, -2, 0, -4, 2, 0, 2, 1, 2, 1, 4, 1, 4, 4, 3, 0, 0, 3, 4, -1, 0, -3, -3, 3, 2, -4, -5, -5, -4, 2, 0, 0, -1, -4, 2, -3, 1, 2, 3, -3, 0, -4, 3, 0, 0, 4, 0, 3, 3, 4, 1, 5, 4, -4, 0, -3, -2, 1, 0, 1, 1, 0, -3, 2, -2, 1, -3, -4, 1, -4, -2, 1, 0, 1, -2, 1, 2, -1, 5, 0, 3, 1, 0, 0, 1, 0, -2, 0, 0, 1, 3, -1, 0, 0, -3, -3, -1, 0, 2, 0, -1, 0, 2, -1, 2, 3, 1, -1, 5, 2, 1, 4, 2, -2, -2, 4, 0, 2, 0, 0, -2, 0, -4, 1, 0, -1, 1, 3, 0, 3, 1, 0, -4, -3, 0, -3, 1, 1, 0, -1, 0, 2, 6, -1, -3, 0, 1, 1, 0, -2, 3, 0, -1, 0, 1, -4, 0, 0, -3, 0, 1, 3, -4, -1, 3, -2, 0, 0, 2, -1, 0, 5, -2, 0, 0, 0, 0, 0, -3, 2, 1, 4, 3, 3, 1, -1, -3, 2, 0, 0, 2, 0, 0, -1, 4, 4, -1, 2, 0, -3, 4, 0, 0, 5, 1, 4, 4, 4, -3, 3, 4, -2, -3, 3, 1, 0, 0, 4, 1, -3, 0, 1, 2, 0, 6, 2, 0, 3, 0, 0, -3, -2, 4, -3, 0, 3, -2, 2, 5, -1, -3, 2, -2, -3, -2, 0, -3, 2, 1, -1, 2, 4, 2, 0, -1, -1, 0, 2, -2, 1, 2, 0, 0, -3, 3, -1, -1, 0, 1, -2, 0, -1, 1, -3, 4, 4, -2, 2, 2, 4, 4, -3, 5, -2, 2, 2, -2, 4, 5, 5, 3, 4, 3, 0, 0, -2, -2, 2, 5, 4, 1, -1, 4, 2, -1, 4, -1, 0, 0, 2, 1, 3, 0, 4, 5, 1, 0, 5, 4, -1, 0, 6, 7, 4, 2, -2, 2, -3, -1, 4, 1, 0, 2, 2, 0, 0, -3, 1, 1, 1, -1, 3, -2, 1, 0, 3, -1, 4, 4, -1, 4, 5, 2, 5, 0, 5, 3, 2, 4, 3, 6, 2, 5, -1, 0, 3, 1, 5, -2, 2, 1, -2, -3, 4, 0, 4, 6, 5, 0, 3, 4, 0, 5, 2, 4, 8, 2, 0, 1, -1, 0, -1, -2, 6, 0, 0, 1, 2, 2, -1, 2, 2, 3, 2, 0, 2, 3, -1, -2, 5, 4, -1, 2, 7, 6, 4, 3, 0, 4, 4, 6, 7, 1, -1, 4, -2, -2, 1, 0, -2, 3, -3, 0, 0, 3, 1, 5, -2, 4, 5, 2, 5, 0, -2, 4, 3, 1, 2, 5, 8, 4, 4, 7, 3, 6, 1, 2, 3, -1, -1, 1, 5, 5, 0, 0, 4, 3, -3, 4, -1, 5, 0, 6, 6, 1, 6, 2, 0, 6, 6, 7, 5, 6, 2, 3, 1, 3, -1, 3, 4, 0, 4, 1, 3, -2, 2, 0, 0, 3, -3, 4, 0, -2, 1, 6, 0, 6, 2, 0, 0, 2, 7, 2, 2, 3, 0, 4, 1, 1, 0, 0, 0, 3, 0, -2, 5, -1, 2, 2, 3, 1, 0, -1, 3, 1, 4, -1, 1, 0, -1, 2, 0, -1, 2, 4, 6, 3, 2, 6, -1, 0, 0, 1, 3, 0, -2, -1, -1, -3, -3, 0, 0, 0, -4, 3, 4, -2, 0, -1, 5, 1, 0, 2, 0, -1, 0, 4, 0, 4, 0, 5, 4, 5, 5, 0, -2, 1, 1, -1, -1, 2, 2, 0, -3, -3, 2, 3, -5, -1, 1, -4, 1, 0, -4, -3, -5, -4, 0, 0, -1, -3, -3, 0, -4, -1, -6, -5, -1, 2, -2, -2, -2, 0, -2, 0, 1, 2, -3, 0, -1, 3, -1, 0, -1, -5, -1, -3, 1, -1, -1, -6, -2, -6, 1, -1, 2, 1, 1, -5, 0, -2, 0, 0, 0, -2, 1, -3, 2, -4, -2, 0, 3, 2, 2, 0, 1, -1, -2, -5, -5, -7, -4, -5, 0, -1, -5, -6, 0, -2, -3, -3, 1, 0, -1, -1, 0, 1, 1, -4, 3, -4, -2, 0, 2, 0, -2, -2, 2, -2, -3, -1, -2, -6, -6, -6, -2, 0, 0, 0, -4, -1, 0, -4, 1, 3, 2, 0, 3, -2, -3, -3, 0, 1, 1, 2, 1, 1, 2, -5, -3, 0, -2, 0, -3, -5, -4, 0, -7, -5, -4, -6, -7, 0, -2, -1, -2, 2, 2, -3, 2, 1, 1, -1, 3, 1, 0, -1, -3, 2, 0, 3, 1, 0, -7, -4, -7, -8, -7, -6, -2, -1, -1, -1, -7, -7, -3, 1, -2, 0, 0, -2, -2, 0, 0, 0, 4, 1, 0, 2, 0, -1, 0, 3, -4, 1, 0, -6, -4, 0, -2, -4, -8, -1, -8, -5, -6, -5, -4, -2, 2, 2, 3, -1, -3, 1, 0, 2, 2, -1, -3, 2, -3, -2, 1, 0, -4, -6, -5, -7, -8, -7, -2, -4, -7, -7, -5, 0, -7, -6, -6, 0, 1, 3, 2, -1, -3, 1, 1, -3, 1, -2, -3, 0, -1, -4, 0, 0, 2, -3, 0, -2, -8, -1, -5, -4, -6, -3, -4, -1, -5, 0, -6, 0, -5, 0, -1, 2, 3, -2, 0, 3, 3, -3, 2, -3, 4, 2, -3, 3, 2, -6, 1, 0, -4, -4, -2, -4, -4, -8, -6, -5, -4, -1, -3, 1, -5, 0, 4, 0, -3, -1, -1, 1, 2, 0, 5, 1, 1, -2, 0, -4, 0, -5, 1, -7, -6, -1, 0, -5, -3, -6, -4, 0, 0, -5, -1, 0, 2, -3, 0, 2, 4, 4, 0, 3, 0, 3, 3, 0, 3, -2, -1, 2, -3, 0, -5, 0, -1, -4, -7, -3, -4, -6, -7, -4, -3, -3, -1, 0, 0, 1, 0, -2, -2, 2, 1, -2, -3, -2, 0, 2, -3, 0, -1, 0, -2, -4, -6, -3, -5, -2, -6, -4, -3, -4, 0, 0, -6, 0, -3, -5, 0, -4, -3, 0, 0, 3, 0, 4, 4, 0, 1, 3, -3, -3, -3, -3, 1, 0, -5, 0, -6, -2, 2, 0, 2, 0, 0, -3, -5, -3, 0, -1, 2, -4, 0, -2, 3, 0, 4, 0, 1, -4, 0, -3, -1, -4, -2, -1, 1, -5, 2, -3, -4, 0, -1, 2, 0, 1, 0, -4, -3, 2, 1, 0, 1, 0, -1, -1, 0, -1, 2, 3, 3, 3, 2, 0, -3, -2, -2, 0, 2, -5, 2, -1, 2, 0, 1, 3, -2, -4, -4, -3, 1, 3, 0, -5, 2, -1, 0, 0, -4, 0, 3, -3, -3, 3, -1, 3, 3, -4, -1, -4, -1, 0, 2, -3, -4, 3, -4, -4, 2, -3, 1, 1, -4, -2, 0, 3, 1, 0, 3, 3, 4, 3, -4, 0, 1, 1, 0, -4, -4, 1, 1, -4, 0, 0, 0, -4, -1, -2, 4, 2, 4, 1, 0, 3, -4, -1, -5, 0, -1, 0, 2, 2, 3, -3, 3, -5, -1, 0, -5, 1, 0, -4, 2, -2, 1, -4, -3, -5, 4, 4, 0, -3, 5, 2, 0, 3, 1, 0, 4, -3, -3, -2, -1, 1, 2, 2, -4, 0, -1, 0, 3, -3, -3, -3, 1, -3, -1, -1, -3, -3, 3, -3, 5, 4, 0, 5, 5, 4, -2, 2, -1, -2, 5, -3, 0, -2, -4, 0, 3, -5, -2, 0, -1, 1, -1, -1, 1, 4, 1, 0, -3, 0, 2, 3, -2, 1, 3, 5, 5, 2, -3, 4, 4, -2, -1, -2, -3, -3, 4, 2, -4, 0, 0, -3, -1, -2, 2, 0, -4, 0, -1, 2, 3, -1, 3, -2, 4, 1, 4, -1, 2, 5, 0, 0, 4, 0, -1, -4, -2, -2, 2, 1, -3, -1, -5, -4, -2, 1, -4, 4, 3, 3, -3, -3, 0, 2, 5, 5, 5, -2, 0, 6, -1, 5, -1, 1, 4, 1, 3, 0, 4, 1, 0, 2, -4, -1, 2, -1, 0, 2, 2, 4, 2, -2, 0, 1, 5, -3, -1, 0, 5, 0, 6, 1, 0, -1, 3, 0, 3, 0, 0, -4, 0, 3, -2, 2, -1, 2, 1, 2, -3, 1, -2, -1, -2, 0, -2, 3, -3, 0, 0, 0, 1, 4, 0, 1, 3, 4, -2, 4, 4, 0, 0, -2, 3, -2, 0, 0, 0, 2, 2, 0, 0, -4, -2, 3, -1, 3, 1, 1, -3, 0, 4, 6, 5, 0, 5, 0, 0, -1, 2, 3, 1, 1, 4, 4, 1, -2, 3, -1, -1, -4, 0, -1, 2, -4, -4, -4, 4, 3, -3, -2, 0, 4, -1, 5, 0, 3, 0, 0, 3, -1, -1, -3, 2, 2, 0, 0, -1, 4, 0, 0, -5, 2, 1, 2, 0, -5, -4, 1, 0, 4, 2, -2, 3, 1, 6, 0, 5, -1, 3, 6, -1, 1, -2, 1, 0, 5, 2, 4, -1, 1, 0, 3, 1, -1, 2, 2, -3, -4, -4, -3, 2, 2, -3, -1, -3, -1, 5, 4, 6, 3, 5, 0, 1, 5, -2, 3, 0, -1, 0, 4, 1, -4, 0, 3, -4, -1, 0, 1, 1, -1, -4, 1, 3, 0, 4, -2, -2, 4, 4, -2, 4, 0, 6, 2, 1, -1, 5, 0, -1, 1, 0, 0, 4, 4, -2, -4, -2, -3, -2, 0, -1, -5, -2, 3, -2, 4, -1, -1, 5, 4, 5, 4, 3, 0, 0, 1, 4, 1, -3, 0, -1, -1, -1, 2, -1, 3, -4, -4, 2, -1, 1, 0, -4, 1, -3, 0, 1, 3, 3, -1, -1, 1, 4, 0, 0, 3, 3, 0, -1, -2, -2, 0, 3, 4, -3, -3, -4, -4, -3, 0, 2, -4, 2, -5, -4, 0, -3, -1, -2, 1, -4, -4, -6, -5, -1, 0, 1, -4, -4, 1, 0, -5, -6, 1, -2, 1, -5, -3, -1, -1, 1, -3, -4, 0, 3, -1, -3, -4, -2, 0, 2, -5, -5, -2, 0, -3, -5, 0, 1, 0, -6, 0, -6, -6, -1, -6, 0, -6, 0, 0, 1, 0, 3, -3, -2, 0, 0, -3, -1, 0, 1, -4, -5, 1, -1, -4, -1, -5, -1, -1, 0, -6, -6, -4, -3, -4, -1, 0, 0, 0, 2, -1, 3, 2, -2, -2, 0, -1, 0, -4, 2, 0, 0, 1, 3, 0, -3, -3, -6, 1, 0, 0, -1, 0, -2, -4, 0, 0, -7, 0, 1, -3, 0, -3, -2, -1, 1, -3, -2, 3, -1, 0, -4, 0, -2, 4, -2, 0, -3, 0, -3, -3, -2, -4, -1, -6, -7, -3, -1, -7, -6, -5, -1, -4, 0, 0, 0, 2, -1, 0, 0, 0, -3, -1, 2, 1, 3, -3, -3, 0, -1, -3, -1, -3, -4, -5, -3, -3, -3, -8, -8, -8, 0, -7, -1, 2, 0, 1, 0, 3, 1, -1, 4, -3, 2, -3, 2, 0, 3, -3, 1, 0, -5, 0, -5, -4, -6, -4, -7, -8, -8, -9, -9, -2, -3, -6, 0, 1, 3, -2, -3, -3, 4, 1, 0, -3, 5, -2, 3, -3, 0, 2, 3, 3, -3, -6, -1, 0, -6, -8, -1, -5, -1, -6, -6, -3, -2, 1, 1, -5, 0, 2, 4, 0, 0, 5, 0, 5, 0, 1, -3, 2, 0, -3, -1, -1, -2, -3, 0, -7, 0, -6, -3, -8, -4, -1, -8, -6, -5, -3, -5, 1, 3, 4, -1, -3, 3, -1, 2, 4, 0, 3, -1, 0, 0, -2, 4, 2, 0, -1, 0, -7, -2, -3, -7, 0, -5, -9, -6, -3, -2, -5, -2, 1, 1, 1, -3, 0, -1, 2, -2, -1, 0, 1, -1, -2, 2, 2, 2, 3, -1, -6, -6, -7, -1, -2, -2, -7, -5, -6, -5, -5, -4, -6, -5, -6, 1, 2, 0, 1, 0, -2, 4, 1, 5, 0, -2, -3, -3, -2, 0, -5, -5, -5, -2, -4, -2, -4, -7, -4, -4, -5, 0, 1, -1, -6, -2, 0, -2, 0, 0, 4, -3, 3, 2, 4, 1, 4, -1, 4, -1, 1, 0, -4, 1, 1, -4, -4, -3, -1, -6, 0, -4, -5, -3, -5, -6, 0, 1, 2, 3, 4, -3, 3, -1, 0, -1, 2, 2, 5, 1, 3, 2, -2, -3, -3, -4, 2, 0, 0, -3, 0, -3, -1, 1, 0, 0, -3, 1, -2, -1, -1, 1, -3, 1, 4, 0, 2, 4, 5, 2, 0, 0, -2, 3, -3, -2, -4, -2, -3, -1, 0, -4, -2, 3, -5, 2, 0, 0, -4, 1, 1, 3, 0, -3, 0, -2, 0, 0, 0, 0, 0, 0, 0, 3, 3, -1, 2, 1, -4, -3, 0, -3, 0, -2, 1, -2, 2, 0, -1, -4, -2, 0, -2, 1, 2, 2, 2, 0, -1, -1, -2, 0, -2, 0, 3, 4, -2, -1, -2, -3, -4, -5, -1, -2, 3, 1, -4, 0, 1, -3, 0, 4, 1, 0, 2, -3, 0, -4, 1, -1, 4, -1, 2, 0, -1, -2, 5, 2, -1, -4, -3, -1, -3, 3, 1, -4, 2, -2, -2, -1, 1, 4, -1, 3, 0, 2, -3, 2, 3, -2, 0, 2, 0, 0, 2, 5, -3, 2, 0, -2, 3, 0, -1, -2, 0, -3, -4, 0, 2, 1, 1, -1, 4, 0, 3, -3, 0, 3, 0, -4, 0, 5, 1, 2, 3, 1, -1, -3, 4, -2, 0, 0, -1, -3, 2, 3, 2, 2, -3, 1, 0, 5, 0, -2, 0, 3, 0, 4, 0, -2, 2, -1, -2, 1, -1, 5, 4, 0, -2, -2, 2, -2, 1, 3, -3, 3, 3, -1, 2, -2, -3, -3, 0, 0, -1, 0, -2, -2, 3, 1, 0, -1, 0, 3, 0, -1, 4, 3, 3, -1, 0, 1, 1, 4, -3, -1, 0, 0, -3, 4, 4, -2, -1, 4, -3, 1, 0, 6, 0, 4, 0, 6, 4, 0, 1, 5, 4, 2, 3, 2, 2, 3, 0, 4, 4, 0, 4, 0, 4, -1, -3, -2, 1, 0, -2, 1, 0, 1, 4, 2, 0, 3, 6, 3, 4, -1, 0, 2, 3, 0, 0, 5, 3, 3, 5, 1, 0, 0, 4, 0, 5, -1, -1, 0, -2, 1, -1, 0, 4, 4, 5, 0, 2, 2, 7, 7, 2, -1, 1, 3, -1, 5, 1, 2, -2, 5, 3, 1, 0, -2, 0, -1, 2, -3, 2, 5, 2, 1, 0, 4, 2, 4, 0, 7, 0, 4, 1, 8, 7, 5, 0, 0, 4, 6, -2, 1, 5, 5, -1, -2, 1, 0, 0, 2, 0, 0, 0, -2, 4, 6, 6, 0, 6, -1, 6, 8, 8, 8, 5, 0, 0, 5, 2, 6, 1, 4, 3, 0, 3, 5, 5, 1, 3, 4, 1, 1, 0, 1, 1, 0, 4, 3, -2, 6, 7, 0, 6, 8, 1, 7, 3, 7, 1, 3, 2, 1, 4, 0, 0, 2, 4, 3, -2, 1, 2, 3, -2, 2, 3, 3, 6, -2, 0, 0, 5, 0, 0, 6, 2, 5, 4, 3, 8, 5, 5, 6, 1, 0, 0, 3, 6, -1, 0, 4, 4, -1, 0, 3, -3, 4, 4, 2, 0, 6, 6, 6, 5, 2, 1, 1, 7, 0, 1, 1, 2, 2, 5, 6, 5, 2, 1, 5, 6, 0, 6, 1, 2, 1, 2, -1, 2, 1, -1, 4, -1, -1, -1, 0, -1, 6, 6, 1, 8, 6, 5, 8, 6, 5, 8, 4, 0, 0, 7, 7, -1, 0, 5, 4, 3, -1, -2, 5, 4, 0, 3, 0, 0, -1, 5, 3, 4, 6, 0, 0, 0, 1, 8, 8, 2, 8, 3, 3, 0, -1, 0, 6, 0, 3, 2, 1, 1, 5, 3, 1, 0, 1, 2, 4, 4, 6, 4, 4, 2, 2, 1, 2, 4, 3, 3, 8, 5, 6, 1, 1, -1, 1, 1, 4, -1, -2, -1, -2, -2, 3, 2,
    -- filter=0 channel=4
    -9, -9, -11, -5, -9, -2, -7, -2, -5, -6, -2, -1, -8, -9, -7, -8, -2, 0, -4, -4, -7, -3, -6, -9, -6, -9, -3, -4, -7, -5, -9, -8, -9, -2, -1, -4, -8, -7, -7, -9, -1, -8, -5, -4, -7, -3, -7, -5, -4, 0, -6, -6, -7, -9, -6, -5, -7, -9, -9, -2, -9, -11, -10, -14, -4, -10, -2, -6, 0, -7, -6, -7, 0, -5, -3, -2, -7, -3, -7, -5, 0, -1, -2, 0, -5, -6, -4, -6, -5, 1, -1, -6, 0, -5, -3, -10, -5, -2, -8, -1, 0, -3, -5, 0, -4, 2, -2, -5, -5, -3, -4, 0, -1, -5, -2, -3, -4, 1, 1, -4, 1, -1, -6, 0, -4, -2, -3, -2, -10, -3, -6, 0, 0, -2, -2, 1, 4, -2, -6, 1, -2, -4, 0, 0, -4, 0, -1, -2, 0, 0, -1, -3, -1, 2, -1, 0, 0, 0, -7, -3, -4, -4, -7, -4, -6, -2, -4, 1, -1, 1, -2, -6, -8, -3, -8, -5, 0, -3, -6, 0, -5, -5, 0, 1, 3, 5, 0, 2, 1, -4, -3, -5, -9, -7, -9, -4, -2, 0, 1, 0, 2, 0, 0, -3, -3, -1, -5, -3, -9, -4, -6, -4, 0, 1, 1, 0, -3, 4, 3, 0, -6, -4, 0, -2, -7, -7, -3, -7, 0, -2, -4, 2, 2, 1, -2, -2, -3, -5, -5, -7, -4, -1, 1, -2, -4, -4, -4, 2, -4, 1, -3, 2, -5, -8, 0, -3, -2, 0, -3, -5, -1, 0, -1, 0, 6, 0, 1, 0, -2, -7, 0, -3, -5, 0, -4, -8, -7, -1, -4, 0, -2, 0, 1, -1, -3, -6, -7, -7, -4, -1, -4, -1, -3, -3, 5, 5, 4, 0, -1, -3, 0, -7, -7, -2, -5, -7, -5, -6, -1, 0, -2, -7, -2, -1, -6, -1, -4, -1, -7, -5, 0, 1, 0, -5, -3, -2, -1, -1, -3, 2, 0, -4, -3, 0, -1, 0, 0, -2, 0, -5, -3, -5, -2, 0, -6, 0, 0, -4, -2, -4, -3, -2, -3, -1, -6, 0, -6, -2, -4, 4, 0, 5, 4, 2, -5, -2, 0, 0, -5, -3, 0, -2, -3, -6, -5, -5, 0, -6, -1, -5, -2, -4, -6, -4, -3, -6, -2, -3, -1, 0, -5, 0, 3, 3, 3, -4, -4, -3, -7, 0, 3, -1, -4, 0, -4, 2, -5, -6, -1, -6, -2, -7, -6, -1, -3, -3, -4, -4, -7, 1, -1, -4, -1, 1, -4, -3, 1, -3, -6, -8, -4, 0, -5, 2, 2, -1, 0, 4, 2, -2, 1, -3, -5, -1, -3, -1, -5, -3, -1, 0, -6, 2, 0, -5, -3, 3, 1, -5, -6, 1, -1, -3, -3, 2, 3, 0, 0, -2, 2, -3, 0, 1, -3, -2, 1, -2, -5, -2, 0, -8, -9, -3, -6, -4, -1, -1, -1, -1, -1, -1, 0, 1, 0, -4, -1, 1, -1, 5, 2, 0, 0, -1, 0, 0, 4, -3, 0, 0, -2, -1, 0, -9, -4, -7, -3, 0, 2, -3, 0, -3, -2, 1, 0, 3, -2, 0, 1, 0, -2, 3, -2, -3, 0, 1, 5, -1, 0, 4, 1, 0, -3, 3, -4, -5, -3, -5, -3, -3, -4, 2, 3, 1, -1, -1, -1, -1, 0, -4, 2, 0, 5, 3, -2, 6, 5, 3, 3, 0, 4, 2, 5, 2, 2, -3, -1, -5, -5, -5, -4, -1, -2, 1, 0, 0, 5, 0, 5, 0, -1, 2, 2, 0, -1, -1, 2, 3, 5, 3, 4, 9, 6, 7, 4, 1, 5, 0, -3, -9, -3, 4, 2, 4, -1, 1, 6, 4, 1, -1, -1, 1, 4, -2, -2, -8, -4, -3, 0, -2, 6, 0, 0, 2, 8, 1, 8, 2, 5, 4, 0, -9, 1, 4, 0, 6, 4, 3, 0, 2, 0, 2, 4, -1, -2, 2, -3, -12, -6, -2, 1, -1, -2, -3, 0, 4, 6, 2, 8, 1, 6, 5, 2, -7, -3, -2, 2, 4, 5, 1, 5, 2, 5, 1, 0, 4, 2, 0, -6, -7, -6, -6, -3, -3, 1, 1, -4, 2, 7, 1, 1, 6, 0, 0, -1, -1, 0, -1, 6, 5, 2, 6, 5, 0, 6, 1, 3, 6, 4, 0, -3, -5, -6, -6, 1, 2, 0, 3, -2, 5, 8, 7, 8, 4, 0, 5, 0, -8, -1, 6, -2, 1, 2, 3, 1, 4, 3, 4, 3, 0, 5, -1, -3, -4, -3, -3, -1, -1, 1, 0, 4, 3, 3, 2, 1, 5, 6, 0, 0, 0, -3, -2, 0, 5, 6, 6, 2, 2, 1, 6, 2, 8, 6, 4, -2, -2, 0, -3, 3, 6, 5, 3, 4, 0, 3, 0, 5, 0, 6, -1, 1, -5, 1, -3, 5, 2, 3, 0, 2, 0, 0, 3, 5, 6, 8, 4, 4, 6, 1, -4, -2, 2, 0, 1, 2, 2, 9, 2, 1, 7, 3, 3, -6, -2, -3, 0, 3, 5, 2, 3, 1, 0, -2, 0, 7, 4, 2, 6, 4, 6, -1, 2, 0, 0, 6, 1, 8, 0, 6, 6, 3, 0, 1, -5, 0, 0, 2, -3, -2, 1, 6, -1, 0, 1, 0, 5, 6, 6, 9, 9, 2, 2, 5, 5, 1, 3, 4, 4, 4, 5, 3, 1, 2, 2, 1, 2, -2, -5, 0, -1, -2, -2, 0, 6, 5, 3, 3, 4, 7, 2, 2, 9, 7, 8, 1, 9, 4, 4, 1, 4, 4, 5, 3, 7, 6, 1, -2, 0, -4, -5, 0, 2, 0, -1, 5, 3, 4, 4, 8, 7, 3, 4, 3, 2, 9, 2, 5, 8, 1, 2, 2, 3, 9, 6, 1, 0, 2, 3, 0, 0, 3, 0, -2, 0, 3, 3, 6, 5, 4, 1, 5, 5, 6, 7, 5, 6, 8, 1, 4, -1, 3, 7, 3, 3, 0, 4, 0, 3, 0, 2, 2, -1, -4, -1, -1, 5, 0, 3, -1, -1, 3, 0, 0, -1, 5, 2, 5, -1, 4, 5, 4, 0, 3, 0, 2, -2, 3, 0, -2, 1, 0, 4, -2, 0, -1, -6, -9, -4, 1, -3, -2, -2, -3, 3, 2, 1, 0, 1, 1, 2, 0, 5, 3, 5, 5, 5, 5, 3, 0, 0, -1, 3, -4, -5, -1, 0, -2, -7, 0, -2, -4, 0, 0, -2, -1, 0, -2, 5, 4, 2, 0, 5, 3, 1, 3, 7, 4, -1, 3, -2, 3, 0, -1, -3, 0, 0, -3, 1, -6, -3, -6, -1, -4, -3, 4, 4, 3, -1, 5, 0, 0, 3, 5, 0, 5, 1, 6, 7, 0, 6, 5, 4, 7, 0, 5, 3, 0, 5, 4, 1, -4, -2, -4, 1, -2, 3, 2, 0, 1, 4, 1, 6, 7, 9, 4, 2, 4, 0, 8, 6, 6, 0, 8, 7, 3, 6, 6, 7, 3, 5, 4, 5, 1, 1, -5, 2, 1, 4, 6, 2, 5, 1, 4, 7, 1, 8, 8, 7, 1, 1, 3, 0, 1, 0, 4, 6, 8, 4, 6, 3, 6, 3, 5, 4, 6, -1, 2, -1, 4, 2, 2, 2, 5, 3, 6, 4, 5, 7, 1, 5, 7, 7, 1, 2, 3, 1, 6, 6, 4, 4, 7, 13, 2, 6, 3, 0, 1, 5, -3, 3, 4, 0, 5, 10, 7, 9, 4, 3, 9, 0, 3, 1, 5, -1, 9, 7, 9, 2, 3, 8, 7, 4, 11, 6, 6, 2, 8, 5, 3, 0, 4, 1, 5, 1, 8, 6, 6, 7, 5, 10, 6, 4, 6, 0, 2, 2, 3, 8, 11, 6, 8, 6, 7, 8, 4, 12, 8, 8, 6, 5, 2, -1, 3, 6, 0, 8, 11, 10, 8, 11, 8, 12, 11, 8, 3, 8, 7, 9, 9, 10, 6, 5, 4, 11, 9, 5, 11, 5, 8, 4, 5, 6, 6, -1, 4, 8, 4, 5, 5, 9, 9, 14, 10, 9, 5, 5, 7, 8, 3, 6, 3, 3, 2, 2, 4, 4, 7, 8, 6, 6, 4, 9, 3, 2, 5, 2, 6, 10, 4, 9, 3, 1, 8, 7, 12, 14, 12, 9, 8, 10, 7, 3, 6, 0, 1, 6, 7, 8, 8, 6, 10, 5, 3, 2, 10, 9, 2, 3, 6, 4, 8, 4, 6, 1, 5, 11, 12, 10, 10, 2, 0, 7, 2, 3, 7, 1, 1, 4, 10, 10, 6, 8, 10, 4, 10, 6, 10, 2, 3, 4, 1, 5, 10, 9, 6, 3, 4, 5, 8, 4, 7, 6, 3, -3, 0, 4, 3, 7, 6, 1, 1, 8, 12, 11, 7, 8, 3, 8, 3, 6, 7, 3, 2, 5, 4, 5, 11, 5, 7, 9, 4, 7, 0, 3, 3, 0, -5, 0, -4, 0, -3, 1, 1, 10, 10, 11, 3, 10, 10, 6, 10, 6, 11, 5, 3, 4, 9, 6, 9, 4, 6, 4, 8, 4, 0, 1, 2, -2, -4, -2, 0, -1, 3, 0, -1, 4, 7, 6, 10, 10, 6, 7, 6, 8, 4, 8, 7, 7, 13, 8, 9, 7, 3, 4, 0, 4, 0, 0, 0, -2, -8, -6, 0, -1, -3, -1, -3, 0, 8, 7, 3, 5, 7, 9, 12, 9, 10, 6, 2, 12, 7, 7, 7, 5, 11, 7, 8, 0, 1, -3, 1, -4, -2, -3, -6, -3, -6, 1, 0, 0, 0, 4, 6, 6, 10, 9, 12, 7, 4, 0, 2, 9, 11, 8, 13, 14, 13, 4, 5, 9, 3, -1, 2, -6, -7, -2, -1, -6, 0, -2, 2, 4, 1, 11, 7, 11, 11, 16, 8, 8, 6, 3, 2, 12, 8, 9, 12, 15, 9, 5, 7, 9, 7, 0, 4, 0, -5, -10, -9, -6, -8, 0, 2, 4, 8, 11, 11, 9, 13, 15, 12, 15, 9, 3, 10, 10, 12, 7, 16, 9, 7, 5, 9, 9, 7, 6, 1, 1, -5, -11, -12, -4, -9, -5, -1, 3, 5, 12, 14, 16, 17, 13, 9, 9, 9, 6, 8, 6, 15, 14, 15, 13, 11, 13, 11, 8, 8, 3, 4, -1, -9, -6, -11, -12, -6, -5, 2, 0, 1, 8, 6, 9, 13, 11, 12, 11, 10, 1, 6, 11, 12, 14, 16, 12, 12, 6, 12, 9, 6, 4, 0, 2, -6, -6, -5, -9, -7, 0, 6, 6, 1, 7, 5, 7, 14, 10, 8, 10, 12, 1, 9, 11, 12, 12, 12, 10, 17, 15, 15, 9, 5, 11, 4, 0, 0, -2, -9, -2, -2, 6, 9, 8, 8, 8, 10, 7, 16, 10, 8, 13, 11, 0, 6, 12, 8, 12, 15, 13, 15, 15, 15, 7, 14, 9, 9, 4, 2, -1, -1, 1, 0, 1, 10, 11, 11, 11, 11, 13, 13, 15, 15, 8, 6, 6, 2, 9, 12, 14, 13, 12, 12, 11, 12, 13, 11, 11, 5, 8, 1, 0, -2, 5, 8, 11, 8, 8, 10, 14, 11, 7, 15, 13, 9, 7, 6, 5, 7, 6, 13, 7, 10, 11, 11, 13, 13, 15, 15, 12, 8, 7, 5, 8, 4, 1, 7, 5, 12, 11, 9, 13, 12, 13, 15, 9, 8, 9, 5, 0, 3, 6, 7, 12, 10, 14, 10, 7, 13, 8, 15, 8, 11, 13, 14, 13, 3, 8, 11, 8, 14, 7, 11, 13, 10, 10, 14, 9, 6, 9, 2, 4, 5, 9, 7, 5, 8, 13, 6, 10, 13, 14, 15, 11, 16, 15, 7, 14, 14, 11, 15, 16, 14, 15, 12, 8, 13, 13, 9, 10, 6, 11, 6, 7, 4, 5, 6, 14, 5, 13, 10, 9, 15, 14, 17, 12, 12, 11, 14, 16, 15, 10, 12, 14, 12, 9, 13, 12, 11, 14, 9, 10, 6, 5, 8, 10, 3, 5, 10, 12, 7, 8, 14, 11, 15, 14, 16, 15, 9, 15, 14, 12, 10, 17, 11, 12, 16, 13, 9, 10, 14, 9, 12, 10, 6, 8, 9, 8, 4, 8, 11, 12, 6, 7, 14, 12, 13, 14, 15, 9, 12, 11, 9, 9, 10, 9, 13, 8, 7, 9, 12, 12, 6, 13, 5, 10, 6, 10, 12, 7, 6, 12, 5, 12, 7, 9, 13, 7, 8, 10, 14, 7, 6, 9, 13, 10, 4, 10, 11, 10, 8, 10, 12, 7, 12, 7, 6, 6, 5, 6, 10, 2, -13, -9, -11, -10, -9, -6, -12, -11, -6, -10, -6, -12, -9, -8, -10, -5, -10, -9, -12, -13, -7, -12, -6, -9, -10, -14, -8, -7, -9, -14, -16, -16, -14, -11, -8, -5, -12, -5, -9, -10, -5, -5, -10, -7, -12, -7, -10, -12, -2, -7, -8, -4, -8, -9, -10, -12, -4, -10, -12, -8, -12, -11, -10, -11, -10, -9, -11, -7, -2, -6, -7, -3, -9, -5, -4, -9, -5, -3, -9, -9, -4, -8, -9, -9, -4, -7, -3, -5, -7, -1, -6, -8, -5, -10, -6, -8, -17, -13, -10, -10, -2, -6, -6, 0, 0, -3, -4, -2, -2, -6, -7, -4, -6, -3, -7, -5, -4, -3, -8, 0, -6, -1, -1, -8, -8, -8, -9, -9, -8, -9, -4, -8, -5, 0, -5, -5, 0, -3, -5, 0, -2, -6, -2, -3, -3, -1, -7, -3, -5, -2, -1, 0, 0, -1, 1, -3, -2, -8, -4, -8, -7, -8, -11, -10, -6, -7, -4, 0, 2, 0, -4, -7, -8, 0, -7, -9, -9, -1, 0, 0, -7, -5, 0, -2, -2, -3, 0, -2, -9, -6, -6, -7, -11, -12, -11, -1, -5, 1, 1, -2, -1, 0, -7, -2, -7, -6, -6, -7, -3, -5, -1, -6, -3, 0, 0, -3, 0, 2, -5, 0, -7, -4, -9, -11, -10, -2, -8, -1, 0, -2, -5, -2, -4, -4, 2, 2, -7, -6, -8, -6, -3, 0, 2, -6, -3, -6, -4, 0, 0, 0, 1, 1, -2, -6, -9, -12, -3, -8, -7, -2, -1, 3, 0, -2, -1, 1, 0, 3, -3, -5, -6, 0, -2, -1, -7, -5, -6, -3, -4, 1, -1, -5, 0, 0, -1, -4, -3, -8, -6, -5, -5, -2, -4, -3, 2, -1, -2, -2, 1, 4, 2, -4, -7, -3, -7, -8, -2, -2, -1, -2, 1, 1, -1, -1, -5, -1, 0, 0, -6, -5, -8, -4, -1, -6, 0, -7, 2, -2, -2, 2, 0, -1, -3, -4, -9, -8, -6, -6, -2, -1, -6, -3, -3, -1, -3, -2, -4, -2, 0, -5, -2, -8, -5, -2, 0, -5, -4, -1, -6, 0, 4, 0, 1, -4, -4, -7, -8, -5, -2, -6, -3, -1, 0, -3, -6, -5, -6, -2, 0, -4, -5, -4, -3, -5, -8, -3, -3, 0, -7, -3, -4, -5, -1, -3, -1, -6, -3, -5, -5, -9, -5, -4, -7, -5, -2, -4, 0, 0, -5, -5, -9, -3, -3, -8, -2, -8, -5, -8, -7, -1, -7, -7, -6, 0, -1, -2, 0, -2, -4, -4, -2, -3, -4, -2, -8, -3, -7, -5, -1, -1, -2, -7, -9, -5, -9, -7, -1, -5, -4, -9, -4, -6, -2, -4, -5, 1, -8, -9, 0, -6, -5, -11, -9, -9, -4, -5, -9, -6, -4, -1, 0, -3, -6, -5, -9, -4, -8, 0, -7, -8, -3, -5, 0, -6, 0, -6, 0, -7, -4, -3, -7, -2, -3, -8, -9, -8, -4, -2, -4, -5, -3, -5, -1, -7, -6, -4, -1, -2, -1, -2, -3, -2, -4, -3, -2, -5, -6, -3, 0, -2, -4, -2, -7, -9, -2, -6, -13, -9, -11, -5, -3, -8, -3, 0, -3, -4, 1, -4, -6, -7, -3, -4, -3, -12, -11, -7, 0, 0, -4, 1, 0, -1, -7, -8, -6, -5, -6, -3, -7, -6, -3, -6, -5, -7, -8, -7, 0, -7, 0, -6, -2, 0, -6, -3, -2, -12, -5, -1, -7, -7, -3, -2, -5, -5, -8, -5, 0, -4, -2, -9, -13, -8, -13, -5, -11, -6, 0, -8, -6, -5, -4, -3, -4, 3, -3, -5, -1, -3, -6, -7, -2, 0, -1, 0, -2, -8, -7, -8, -6, -6, -8, -10, -14, -12, -12, -12, -8, -4, -8, -6, 0, -5, -1, -6, 0, 0, -4, 2, 0, -6, -9, -4, -3, -2, -3, -5, -4, -8, -8, -2, 0, -5, 0, -4, -6, -17, -14, -16, -6, -7, -8, -8, -8, 0, -4, -1, -3, 1, -4, 0, -2, -4, -4, -2, -7, -1, -1, 0, 0, -2, -5, -3, 0, -6, -7, -10, -12, -18, -11, -16, -6, -5, -5, -3, -2, 0, -3, 1, -5, 0, 0, 0, 0, -5, -4, -6, -8, 0, 1, -2, 0, -1, 0, -3, 0, -5, -4, -4, -9, -12, -10, -7, -8, -1, -2, -1, -4, -6, 0, -3, -1, -4, -7, -1, -3, -12, -6, -2, -5, -8, -1, -3, -3, -1, -1, -2, -3, -2, -7, -9, -5, -7, -9, -5, -8, -4, -7, 0, 0, -1, -4, -3, 0, 0, -7, -2, -3, -8, -9, -8, -8, -5, -6, -8, -2, -9, -6, -7, -3, 0, -3, -4, -5, -7, -10, -7, -9, 0, -4, -3, 1, -1, -1, -1, 0, -4, -3, -8, -10, -8, -5, -3, -8, -7, -8, -1, -3, -8, -5, -6, 0, 0, -8, 0, -4, -5, -7, -4, -1, -6, -3, 1, -1, -2, -8, -1, -1, -5, -9, -4, -7, -10, -10, -4, -12, -12, -7, -8, -11, -4, -12, -6, -1, 0, -6, -6, -5, -2, -3, -3, -4, -8, -3, -6, -7, -3, -9, -7, -7, -5, -4, -4, -7, -11, -11, -5, -7, -8, -4, -7, -3, -12, -12, -3, -5, -2, -7, -4, -1, -9, -8, -11, -4, -6, -8, -11, -10, -6, -5, -10, -10, -6, -6, -3, -7, -9, -10, -9, -12, -10, -9, -8, -8, -7, -7, -7, -3, -6, -5, -2, -8, -10, -9, -3, -9, -5, -3, -8, -7, -5, -3, -10, -3, -12, -10, -8, -12, -9, -11, -13, -4, -5, -2, -2, -5, -4, -7, -8, -5, -4, -9, -9, -1, -5, -8, -3, -2, -3, -2, -7, -7, -11, -8, -7, -11, -11, -7, -6, -11, -5, -11, -10, -12, -4, -10, -8, -2, -3, -12, -7, -4, -10, -9, -6, -10, -5, -5, -4, -12, -6, -5, -4, -6, -10, -9, -11, -11, -5, -6, -6, -6, -10, -8, -12, -4, -10, -11, -10, -8, -10, -11, -8, -10, -12, -11, -12, -10, -7, -9, -7, -9, -6, -7, -11, -13, -9, -5, -12, -7, -12, -9, -13, -9, -9,
    -- filter=0 channel=5
    -1, -8, -3, -3, -1, -2, -4, -6, 0, -5, 3, 0, -2, 1, -3, -2, 0, 1, 0, 0, -1, -3, 3, 0, -4, -7, -4, -1, 0, -4, 1, -5, -1, -5, 2, -3, -3, -4, -4, -3, -1, 1, -1, 6, 8, 9, 8, 8, 6, 7, 2, 9, 10, 6, 0, 0, -4, 0, 1, -6, 0, -2, -6, 0, 2, -1, -2, 1, 0, 3, 3, 0, 6, 4, 8, 4, 13, 6, 12, 13, 12, 14, 16, 16, 6, 8, 9, 5, 0, -1, -5, -1, 1, 1, 1, -5, 3, 2, -4, 3, 5, 2, 4, 6, 5, 4, 11, 12, 8, 15, 11, 13, 15, 12, 15, 17, 8, 10, 8, 5, 5, 0, -1, -2, -3, -2, -5, -1, 2, 1, -3, -3, 4, 1, 1, 6, 9, 6, 14, 13, 18, 22, 20, 15, 17, 14, 20, 11, 17, 14, 11, 10, 7, 5, -3, -4, 1, -2, -3, -3, 1, 3, 2, 4, 5, 3, 9, 3, 7, 11, 10, 18, 17, 22, 20, 21, 17, 14, 19, 13, 11, 14, 14, 8, 8, 4, 0, -2, -3, -4, -4, 1, -1, 3, -1, 6, 3, 1, 4, 5, 11, 11, 15, 18, 17, 19, 20, 19, 16, 22, 17, 15, 15, 16, 10, 11, 7, 2, 6, 4, -1, -2, -2, -2, -1, -2, 2, 0, 5, 5, 1, 7, 5, 6, 9, 13, 17, 12, 20, 16, 18, 16, 18, 15, 18, 12, 15, 11, 7, 3, 8, 4, 2, -3, 1, -4, -2, -3, 0, 5, 6, 4, 9, 5, 3, 6, 7, 6, 14, 14, 17, 12, 16, 17, 12, 16, 10, 15, 11, 8, 9, 8, 2, 4, 1, 0, -1, -4, 0, 2, 2, 0, 6, 5, 7, 8, 10, 8, 10, 4, 4, 8, 8, 12, 9, 6, 9, 14, 9, 13, 12, 5, 3, 6, 2, 0, 0, -3, 0, -1, -3, -3, 1, 0, 0, 5, 5, 4, 1, 6, 3, 1, 6, 2, 6, 11, 5, 5, 10, 8, 4, 9, 7, 8, 3, 7, 2, 5, 4, 4, -4, -3, 0, 1, 2, 5, 2, 7, -1, 1, 6, 6, 0, 5, 2, 4, 5, 5, 6, 7, 4, 10, 7, 6, 0, 4, 1, 0, 5, 5, 0, -2, 5, -1, 1, 2, -2, 3, 4, 0, 2, 4, 0, 0, -1, 1, -2, -1, -3, 1, -2, -4, 0, 3, 2, -2, 0, 1, 3, 7, 6, 0, 3, 2, 0, 3, 1, 4, 5, 4, 2, 0, 0, 5, -1, 0, 2, -2, 1, 0, 0, -5, 1, 0, -3, 1, -2, -1, 3, -1, 6, 6, 0, 0, 0, 3, 2, -1, -1, -2, 3, -3, 1, 0, 1, -1, 2, 0, 2, -3, 1, -2, -6, -2, -3, -5, -4, -7, -4, -5, -3, -1, 0, -2, 1, 2, 1, -2, 1, 0, -4, 2, -3, 0, 3, -3, 0, -2, 0, -4, -3, 0, 2, 0, -4, -7, -3, -8, -1, -3, -4, -5, 1, -2, 4, 2, 2, 6, 1, 0, -1, 3, -1, 3, -2, -1, -3, 0, 3, 1, -1, 4, -3, 3, -3, -5, -3, -1, -5, -2, -2, -7, -5, 1, -3, 1, 0, 0, -1, 4, -2, -2, 3, -1, 2, 4, 0, -3, -1, -3, 1, 0, 4, 4, 2, 0, 3, -2, -2, -3, -1, -3, 1, 0, 0, 2, 4, 7, 6, 7, 6, -2, 0, 0, -4, -1, -2, -4, -4, -3, -2, 5, 3, 0, 0, 4, 9, 0, -1, 2, 5, 4, -1, -4, -5, -1, 0, 1, 8, 2, 6, 1, 5, 0, 0, -2, -4, -2, 0, -2, -5, -4, 4, -1, 5, 1, 2, 6, 4, 2, 8, 5, 1, 3, 0, 3, -3, 2, 5, 2, 8, 1, 9, 6, 0, 2, -3, 3, 0, -2, 0, -4, -2, 2, 0, -3, 1, 0, 4, 2, 9, 8, 3, 7, 2, 1, -1, 3, 3, 4, 4, 7, 9, 8, 10, 1, 7, 6, 0, 0, -6, -9, -7, -6, -3, -5, -3, 4, 5, 0, 5, 4, 5, 13, 8, 3, 1, 6, 3, 2, 1, 7, 3, 4, 8, 1, 2, 7, 4, 4, -4, -5, -4, -7, -10, -4, -3, -5, 0, -1, 0, 6, 6, 6, 6, 11, 6, 7, 11, 5, 2, 2, 10, 2, 2, 9, 4, 9, 6, 5, 0, -1, 1, -2, 0, -11, -12, -3, -4, -2, 1, 0, 3, 3, 5, 6, 9, 11, 7, 11, 9, 2, 7, 3, 5, 10, 9, 3, 6, 11, 9, 2, 7, 2, 0, -2, 1, -5, -4, -3, 0, -3, 2, 0, -1, 1, 8, 4, 6, 9, 7, 11, 5, 3, 8, 11, 6, 12, 10, 8, 2, 10, 11, 3, 7, 8, 1, 0, -1, -9, -5, -3, -1, 0, -2, -1, 4, 7, 3, 3, 11, 11, 11, 9, 3, 11, 13, 8, 7, 10, 6, 2, 7, 8, 9, 6, 7, 7, 3, -5, -1, -6, -11, -11, -3, 0, 2, 2, 4, 6, 10, 6, 10, 14, 9, 13, 4, 5, 6, 13, 13, 8, 9, 4, 8, 5, 6, 4, 0, 6, 4, -2, -1, -12, -4, -5, -1, -6, -3, 5, 6, 0, 10, 12, 13, 11, 11, 8, 12, 8, 9, 12, 9, 13, 12, 4, 3, 1, 3, 1, 4, 2, 1, 0, -2, -11, -11, -3, -9, 2, -3, 5, 4, 5, 6, 6, 9, 5, 7, 10, 12, 4, 4, 8, 7, 11, 5, 7, 2, 2, 3, 5, -1, 3, -1, 0, -9, -8, -5, -11, -2, -3, 2, -3, 4, 6, 9, 1, 7, 7, 6, 5, 9, 9, 2, 7, 4, 5, 6, 5, 1, 0, 4, 5, 5, -3, 1, -3, -8, -5, -4, -10, -3, -3, -1, 0, 3, 5, 7, 7, 6, 4, 3, 5, 5, 2, 4, 6, 2, 8, 0, 2, 1, 6, 2, -2, 0, 1, -3, 0, -2, -5, -7, -6, -5, -1, -1, 0, -1, 4, 3, 2, 0, 4, 6, 0, 1, 5, -1, 2, -2, 0, 1, -1, 0, 0, 0, -1, 0, -1, -3, -7, -7, -5, -6, -10, -11, -14, -12, -12, -13, -8, -16, -9, -14, -12, -12, -4, -8, -7, -5, -8, -8, -7, -12, -5, -7, -8, -11, -14, -9, -11, -11, -7, -11, -9, -13, -14, -6, -12, -11, -11, -13, -5, -5, -5, -4, -6, -1, -7, -7, -3, -6, -3, 0, 1, 0, -5, -10, -10, -4, -11, -8, -11, -13, -7, -7, -8, -4, -12, -10, -9, -4, -8, -4, -7, -7, -2, -1, -6, -4, -1, 0, 0, 5, -1, 0, 0, -2, -4, -7, -5, -11, -6, -13, -9, -6, -6, -13, -5, -3, -6, -11, -8, -2, -1, -7, -1, -4, 0, 2, 0, -2, 4, 1, 6, 7, 2, 2, 4, 0, 2, -5, -2, -9, -6, -11, -6, -7, -6, -7, -6, -2, -6, -11, -3, -3, -1, -1, -1, -4, -3, 0, -1, 1, 9, 4, 8, 4, 5, 9, 7, 5, 5, 2, -4, -2, -9, -5, -11, -3, -10, -13, -7, -6, -6, -9, -9, -9, 0, 1, -3, -3, 0, 0, 7, 2, 10, 5, 10, 5, 5, 8, 3, 4, 0, -1, 0, -6, -3, -1, -7, -4, -7, -7, -8, -7, -1, -2, -3, -3, -6, -4, -7, -2, 3, 3, 7, 6, 6, 4, 4, 8, 2, 5, 1, 5, 4, 2, -3, -4, -1, 0, -5, -7, -3, -4, -3, -4, -10, -2, -3, -5, 0, -4, -2, 0, 1, 0, 6, 2, 2, 5, 5, 2, 8, 3, 4, 6, 1, -1, -3, -2, -3, 1, -2, -5, -1, -3, -8, -10, -2, -6, -9, -8, -5, -2, -7, 0, -3, -1, 2, 3, 3, 8, 1, 4, 3, 6, 0, 0, 0, 1, -3, 2, 0, -6, -5, -1, -6, -3, -6, -8, -10, -7, -6, -3, -3, 0, -1, 1, -2, 2, -5, 0, 3, -1, 2, 0, 1, 3, 0, 0, 1, 2, 0, 0, -2, -6, 0, -1, -1, -5, -10, -6, -6, -10, -9, -4, -7, 0, -1, -2, -1, -3, -3, -8, -5, 4, -4, -2, 0, -1, -3, -4, 0, 1, 0, -3, -8, -10, -6, -8, -9, -4, -5, -7, -7, -4, -9, -2, -2, -1, -3, -5, -2, -8, -2, -6, -4, -3, 1, -2, 0, 0, -1, 1, 0, -1, -1, -7, -8, -4, -4, -5, -7, -7, -10, -3, -3, -8, -7, -1, -8, 0, 1, -4, -3, -7, -6, -1, -7, -6, -3, -3, -6, -8, -4, -2, 0, -7, -5, 0, -2, 0, 0, -8, -9, -3, -7, -2, -4, -2, -5, -9, -4, -1, -4, -2, -8, -1, -2, -9, -8, -7, -2, -5, -8, -5, -7, -7, -3, -2, 0, -7, 0, -1, -7, -2, -4, -3, -1, -4, -5, -9, -5, -8, -5, -8, -7, -2, -2, -2, -8, -3, -6, -3, -1, -3, -8, -3, -9, -2, -7, -5, -6, 0, -4, -1, -6, -1, -7, -5, -3, -10, -7, -11, -10, -7, -6, -3, -2, -2, -8, -3, -1, -3, -7, -5, -4, -2, -3, -8, -2, -11, -3, -5, -3, -4, -3, -2, 1, -8, -4, -2, -6, -9, -5, -5, -4, -2, -9, -6, -4, 0, -2, -2, -3, -5, 0, -3, -4, 0, 0, 0, -8, -5, -7, 1, -3, 2, -6, 1, -5, -6, -3, -3, -8, -10, -3, -10, -5, -7, -3, 0, -4, 2, 4, 4, 0, -2, 4, 0, 0, 0, -3, 0, -6, -3, 0, 4, -1, 3, 3, 0, -1, -6, -2, -6, -4, -10, -4, -5, -7, -4, 0, 0, -4, 3, 1, 4, 5, -1, 1, 3, -2, 3, 0, -4, 1, -5, 1, 0, -4, 2, -3, 2, -2, -3, -3, -4, -11, -9, -8, -1, -6, -7, 0, 0, 0, 3, 4, 1, 5, 1, 0, 3, 0, 2, -6, 0, 0, 3, 0, 2, -1, 0, 0, -2, -4, -6, -7, -6, -10, -13, -2, -7, -7, -3, -5, 1, -2, -1, 6, 1, 7, 1, 3, 2, -2, 0, 1, -3, -2, -1, 5, 3, 0, 1, 5, 0, -3, -2, -7, -3, -9, -13, -8, -6, -10, 0, 0, 0, 3, 4, 4, 5, 4, 7, 6, 5, 1, 2, 4, -2, 0, 0, 2, 3, 0, 4, -2, -1, -4, -4, -5, -10, -11, -14, -8, -6, -9, -1, -5, 0, 3, 0, 2, 4, 8, 7, 7, 7, 2, 1, 6, 4, 0, 5, 0, 3, 7, 0, -1, 0, 0, -7, -5, -5, -9, -11, -14, -12, -8, -7, -7, -1, -5, 1, 4, 0, 3, 1, 5, 5, -1, 4, 0, 2, 8, 3, 7, -2, 1, 0, 3, 3, -1, -6, -7, -10, -7, -15, -10, -6, -10, -7, -4, 0, 2, 2, -1, 0, 5, 2, 3, 4, 5, 5, 1, 1, 1, 2, 0, 5, 0, 0, 6, 3, -3, 0, -2, -5, -13, -15, -13, -5, -2, -6, -6, -6, -3, -3, 0, 5, 2, 0, 1, 5, 7, 2, 3, 8, 7, 3, 2, 3, -1, -2, 5, 4, 1, 0, -4, -8, -15, -10, -11, -10, -11, -5, -8, -3, 0, -1, 4, 3, 0, 8, 9, 0, 0, 6, 2, 0, 2, 1, 2, 4, 1, 0, 0, 0, -5, -1, -3, -11, -15, -15, -14, -9, -4, -7, -2, -5, 1, 0, 0, 6, 0, 2, 4, 3, 4, 0, 0, 0, 3, 1, 4, 4, 0, 2, -5, -3, -7, -5, -10, -6, -10, -10, -10, -8, -8, -10, -7, -5, 1, 1, 1, 1, 2, 2, 0, 5, 0, 1, 0, -3, 4, 0, -2, -4, 1, 2, 1, -5, 0, -6, -13, -11, -11, -15, -10, -10, -7, -8, -1, -2, -3, 4, -4, -3, 3, -3, 2, -1, 3, -1, 0, 3, 1, 0, 1, -2, -3, 0, -1, -5, -1, -4, -6, -12, -17, -12, -14, -9, -12, -11, -6, -1, 0, 1, 1, 0, 0, 4, 2, -5, 0, 0, -5, -1, -1, -2, -4, -5, -1, -3, -6, -7, -8, -8, -9, -14, -9, -13, -14, -10, -13, -13, -3, -6, -5, -4, -1, -2, 0, 0, -8, -3, -8, -1, -2, 0, -1, 1, 0, -7, -3, -9, -5, -10, -9, -9, -12, -8, -14, -11, -16, -14, -10, -13, -17, -9, -13, -19, -13, -11, -8, -12, -11, -11, -8, -8, -8, -13, -10, -12, -13, -8, -11, -8, -16, -14, -17, -17, -18, -18, -12, -10, -13, -16, -12, -8, -14, -9, -13, -7, -10, -6, -10, -8, -9, -9, -5, 0, -7, -8, -7, -4, -10, -10, -10, -12, -9, -17, -12, -13, -12, -11, -15, -7, -8, -12, -11, -10, -13, -11, -11, -3, -8, -2, -8, 0, 1, 2, 0, -4, 3, -3, -2, -5, -3, -1, -11, -11, -7, -14, -8, -7, -7, -8, -8, -13, -8, -5, -6, -7, -6, -8, -10, -9, -2, -5, 0, -3, 4, 3, 4, 1, 2, 0, 6, -1, 1, -2, -2, -11, -3, -11, -13, -9, -10, -11, -7, -8, -7, -13, -14, -12, -10, -2, -3, -1, -5, 0, 1, 7, 9, 4, 9, 3, 5, 9, 7, 6, 1, -5, -1, -8, -6, -10, -12, -5, -13, -15, -7, -9, -11, -5, -11, -8, -3, -3, -5, -1, -2, 5, 7, 7, 10, 12, 7, 12, 8, 4, 9, 2, 3, 0, 0, -3, -2, -8, -10, -9, -10, -7, -6, -7, -8, -7, -3, -7, -4, -5, -1, 0, 1, -1, 8, 11, 4, 4, 6, 6, 9, 2, 7, 2, 4, 6, 1, -1, 1, -3, -7, -10, -11, -5, -5, -11, -12, -11, -8, -6, -2, -1, -1, -2, 3, 4, 6, 2, 10, 4, 2, 11, 6, 4, 6, 7, 4, 4, -1, 0, -2, 1, -9, -1, -10, -9, -12, -8, -3, -3, -10, -2, -6, 0, 0, 0, -3, 1, 2, -2, 6, 8, 5, 4, 10, 9, 3, 2, 7, 3, 0, 0, -6, -2, -8, -8, -7, -8, -3, -9, -8, -7, -7, -2, -1, -1, 1, 0, -2, 3, -1, 0, 8, 3, 2, 3, 4, 7, 7, 1, 4, 5, -1, -5, 0, -7, -1, -8, -10, -3, -7, -3, -9, -2, -1, -10, -3, -5, 2, 0, 2, -2, -1, -2, 0, 2, 9, 7, 2, 8, 6, 0, 2, 0, 0, -4, -1, -4, -8, -4, -5, -10, -6, -9, -9, -1, -3, -6, -4, -1, -3, -1, 2, 0, 0, 1, 0, 0, 3, 2, 3, 0, 4, 1, 1, 0, 2, 0, -2, -4, -2, -5, -9, -8, -9, -1, -7, -4, -5, -8, 0, -6, 0, 1, 1, -3, -1, 4, 4, 3, 1, 5, 4, -2, 0, 3, -1, -1, 2, -1, -4, 1, -1, -3, -7, -3, -5, -1, -6, -4, -8, -1, -4, -5, -3, -3, -3, 0, 3, 1, 0, 3, -1, 3, 1, 3, -2, -3, -3, 2, -1, 0, 2, -2, -2, -3, -5, -1, -2, -1, -1, 0, -1, -3, -2, -2, -3, -3, -4, -3, 1, 0, 1, -1, 2, 2, 3, 5, 2, -3, -4, 1, -3, 3, -3, -3, -2, 0, -7, -5, -1, -1, -2, -2, -1, 0, -2, 3, 0, -2, 1, -2, 0, 3, 0, -1, 2, 0, 4, -1, 0, -3, 0, 0, 0, 2, 3, -3, -1, -7, -8, 0, 0, -1, -2, -5, -5, -4, -1, 0, 3, 3, 0, 0, 5, 2, 6, 2, 7, 0, 9, 0, -1, 2, 4, 3, 6, 0, 1, -3, -3, -5, -9, -8, -6, -4, -8, -8, -7, 0, -1, 4, 1, 8, 8, 6, 6, 7, 2, 11, 9, 9, 6, 1, 0, 0, 3, 0, 3, 2, 2, 1, 1, -1, -7, -6, -6, -7, -1, -9, -6, -5, 0, 0, 0, 6, 9, 13, 4, 5, 10, 9, 9, 11, 8, 6, 8, 9, 9, 8, 4, 8, 1, -2, -3, -2, -3, -9, -10, -3, -7, -6, -2, 1, -1, 0, 5, 3, 4, 12, 8, 7, 9, 7, 11, 5, 5, 1, 4, 9, 4, 6, 2, 8, 2, 3, 1, -2, -7, -1, -11, -9, -2, -4, 0, -1, -1, 0, 7, 2, 9, 7, 14, 9, 6, 9, 12, 7, 5, 9, 5, 9, 5, 9, 10, 6, 3, -1, 0, 0, -6, -7, -9, -3, -9, -3, -5, -4, -3, 2, 8, 7, 10, 6, 11, 17, 7, 12, 12, 6, 5, 6, 6, 11, 7, 9, 5, 5, 9, 4, -1, 2, -3, -10, -9, -8, -5, -9, 0, -5, 1, 0, 2, 9, 11, 13, 14, 9, 12, 10, 9, 9, 8, 8, 13, 5, 8, 7, 7, 7, 3, 4, 0, 2, -6, -5, -7, -10, -10, -4, 0, 0, 0, 2, 6, 8, 7, 10, 8, 14, 12, 10, 11, 14, 13, 12, 15, 16, 10, 11, 4, 5, 9, 5, -1, 1, -5, -1, -4, -10, -3, -2, -2, -2, -2, 0, 6, 3, 9, 6, 6, 6, 12, 10, 9, 5, 11, 11, 8, 13, 13, 9, 3, 6, 6, 4, 0, 0, 1, -7, -6, -9, -7, -5, -2, 0, -2, 1, 7, 2, 3, 5, 9, 13, 12, 5, 10, 7, 11, 7, 8, 8, 12, 2, 4, 9, 8, 11, 0, 2, -4, -10, -7, -13, -7, -2, 1, -2, -1, 6, 5, 7, 8, 15, 12, 7, 14, 5, 13, 10, 15, 12, 12, 7, 6, 8, 10, 8, 4, 3, 2, 0, 0, -9, -14, -11, -2, -6, -2, 3, 0, 5, 9, 9, 8, 13, 7, 11, 12, 7, 9, 12, 9, 8, 6, 6, 5, 10, 7, 11, 0, 6, 2, 0, 1, -2, -5, -11, -9, -1, 0, 4, 4, 1, 5, 4, 11, 6, 14, 6, 6, 7, 7, 10, 9, 9, 9, 4, 3, 8, 9, 5, 3, -1, -1, 0, -2, -9, -9, -3, -8, -7, -3, -1, 2, -1, 5, 6, 2, 7, 4, 10, 7, 11, 6, 3, 7, 5, 2, 8, 3, 6, 3, 6, 7, 5, 4, 0, -3, -4, -9, -7, -7, -6, -2, 0, 3, 1, 8, 4, 8, 10, 7, 5, 5, 10, 4, 1, 1, 7, 7, 8, 9, 2, 6, 5, 0, 3, 0, 0, -5, -8, -4, -8, -8, -3, 1, -5, -5, 3, 5, 3, 6, 5, 7, 2, 0, 4, 6, 6, 4, 6, 1, 1, 6, 1, 6, 0, 2, -2, 2, 1, -5, -9, -9,
    -- filter=0 channel=6
    3, 4, 7, 0, 3, 2, 7, 5, 8, 0, -1, -1, 2, 6, -3, -1, 0, 0, 2, -3, -2, -3, -2, 0, -1, 0, 2, 5, 3, 8, 7, 8, 6, 9, 7, 5, 2, 5, 9, 3, 1, 2, 3, 0, 7, 4, 4, -3, 0, 1, -1, 3, -1, 6, 6, 5, 5, 6, 6, 3, 1, 10, 6, 9, 4, 6, 3, 7, 8, 7, 9, 3, 1, 7, 4, 6, 4, 2, -1, 4, 2, 2, 1, 1, 3, 2, 6, 5, 2, 3, 10, 4, 2, 4, 0, 7, 6, 6, 5, 11, 2, 6, 5, 1, 1, 5, 0, 2, -2, 0, 4, 0, 0, -4, -2, -4, 0, 2, 3, 4, 1, 1, 3, 6, 4, 4, 6, 8, 4, 9, 3, 9, 2, 9, 9, 7, 0, -2, 6, 2, -3, 4, -2, -2, -1, 1, 0, -1, 4, 1, 0, 4, 6, 0, 3, 1, 2, 0, 4, 6, 10, 8, 9, 2, 6, 6, 8, 8, 6, 0, 7, 4, 0, 5, -3, 3, -2, 0, 3, 4, 8, 6, 6, 3, 6, 2, 6, 1, 2, 7, 10, 4, 6, 9, 7, 5, 2, 0, 6, 10, 7, 7, 6, 6, 2, 6, -1, 8, 5, 4, 6, 1, 8, 1, 8, 1, 6, 6, 1, 2, 8, 8, 4, 3, 11, 4, 7, 7, 2, 2, 6, 9, 1, 10, 0, 2, 7, 8, 7, 6, 3, 8, 4, 10, 2, 3, 2, 9, 5, 3, 4, 5, 8, 7, 5, 2, 10, 6, 4, 3, 8, 1, 8, 8, 6, 7, 6, 8, 6, 12, 9, 2, 7, 10, 13, 8, 11, 9, 7, 8, 10, 10, 4, 7, 1, 9, 8, 9, 8, 4, 5, 5, 4, 4, 0, 5, 1, 3, 9, 8, 15, 7, 8, 8, 12, 16, 10, 11, 12, 9, 11, 2, 9, 3, 1, 8, 3, 2, 0, 9, 8, 0, -1, 5, 7, 0, 0, 0, 0, 6, 6, 6, 8, 16, 13, 8, 17, 17, 12, 15, 12, 7, 12, 4, 2, 4, 1, 3, 2, 2, 3, 2, 5, -1, 0, -2, 0, 2, 6, 6, 0, 3, 4, 5, 11, 9, 9, 11, 16, 11, 13, 14, 14, 14, 10, 9, 5, 0, 0, 0, 2, -1, 3, 4, 1, 7, 2, 4, -1, 0, 3, -1, 4, 8, 3, 11, 16, 12, 19, 10, 9, 16, 12, 14, 5, 5, 6, 2, 6, -3, 0, 0, -5, -2, 3, 5, 3, 4, -4, -3, 0, 0, 2, -2, 0, 9, 9, 14, 12, 10, 13, 15, 16, 15, 12, 7, 11, 4, 3, 0, 1, -1, -3, 0, -5, 0, 4, 5, 2, 0, 0, -7, 1, -5, -9, 0, 3, 1, 9, 9, 12, 11, 10, 12, 12, 14, 16, 15, 10, 4, 3, 3, -2, -3, -1, -2, -5, 0, -1, 0, 2, -1, 0, -3, 0, -10, -3, -3, 1, 1, 1, 12, 13, 14, 19, 14, 12, 15, 7, 6, 5, 2, 0, -5, -10, -7, -7, -11, -6, 1, -3, -3, 0, -1, -3, -2, -6, -5, -5, -6, -10, -5, 5, 2, 8, 17, 16, 17, 15, 9, 13, 14, 7, 7, 4, -6, -5, -7, -6, -10, -3, -2, -2, 3, 0, -1, -2, -7, -7, 0, -11, -4, -4, -5, 1, 7, 7, 14, 17, 16, 19, 14, 19, 12, 4, -1, -6, -7, -7, -8, -7, -5, -7, -2, 3, 3, 3, 0, -2, -5, -5, -3, -9, -6, -1, -1, 1, 0, 8, 8, 16, 14, 12, 16, 13, 12, 3, 0, -4, -6, -11, -7, -2, 2, -2, 2, -3, 0, -2, 0, -2, 4, 0, 3, -3, 0, -1, -1, -4, 0, 7, 6, 16, 15, 11, 15, 15, 12, 1, -4, -8, -1, -3, -8, 0, -2, -1, -3, -4, 7, 1, -5, 1, 2, -2, 2, 0, -3, -7, -4, -1, -2, 7, 3, 14, 15, 14, 16, 10, 9, 3, 1, 0, -1, -5, 1, 0, 0, 1, -2, 0, 7, 0, 0, 0, -2, 0, 1, 2, -3, 1, -4, 0, -2, -2, 0, 5, 4, 8, 10, 4, 0, -1, -1, -2, -2, 0, 4, 0, 3, 3, 1, 1, 5, 3, 0, -2, 1, 2, 8, 5, 4, 2, 0, -3, 1, -2, 0, 0, 4, 4, 0, 4, -4, -1, 2, 0, -4, -1, -1, 0, 5, 0, 6, -2, 3, 0, -2, 0, 4, 0, 1, 1, 0, 2, 3, 1, 5, -2, -2, 0, -2, -2, 3, -5, -3, -2, 3, 0, -1, 2, 2, 7, 4, 7, 1, 4, 4, -2, 6, 2, -1, -1, 8, 6, 3, 3, 0, 5, 6, 3, 0, 2, 0, -1, 4, 1, 3, 0, 0, -1, -2, 3, 1, 2, 5, 3, 2, 4, 7, 3, 0, 0, 2, 4, 7, 8, 8, 6, 2, 6, 3, 4, 5, 3, -3, 3, 3, 4, 0, 5, 7, 5, -1, -1, -2, 6, 1, 2, 0, 3, 4, 3, 0, 5, 5, 1, 6, 9, 7, 5, 8, 3, 1, 0, 2, 1, 2, 2, 6, -1, -1, 2, 1, 6, 0, -1, 6, 1, 5, 5, 2, 9, 12, 2, 2, 7, 4, 5, 8, 1, 3, 5, 0, 4, 4, 0, -1, 3, -1, 7, 1, 1, 3, 1, 4, 5, 2, 1, 6, 2, 3, 6, 4, 5, 8, 4, 1, 3, 4, 3, 8, 0, 2, 2, 4, 0, 1, -1, 0, 0, 1, 3, 1, 8, 8, 2, 3, 2, 4, 6, 3, 3, 12, 10, 7, 2, 7, 0, 3, 1, 4, 6, 3, 2, 3, 1, 4, 0, 1, 0, 2, 0, 2, 2, 2, 6, 0, 3, 4, -1, 4, 3, 7, 10, 10, 4, 0, 6, 2, 4, 0, 5, 2, 0, 0, 0, -2, 1, 4, 1, 4, -4, 3, 4, 3, -2, 1, 3, 0, 3, -3, 0, 7, 4, 3, 5, 1, 3, 5, 10, 8, 5, 1, -1, 0, 4, 6, 0, 2, 3, -3, 0, -3, 2, -1, 0, 0, -4, 1, 4, -3, 1, 5, 1, 1, 6, 5, 8, 0, 5, 10, 6, 9, 8, 1, -1, 2, -2, 1, -1, 2, -1, -2, -5, 1, 1, 0, -3, 0, -1, -3, -7, 2, 0, 0, 0, -1, 2, 2, 3, 3, -3, 3, 3, 5, 2, 3, -2, 3, 4, -1, 0, -3, 3, 4, 0, 3, 3, -1, -1, 0, -2, 0, -2, 0, -4, -5, -5, 0, 2, 0, 1, 3, 3, 0, 5, 1, 6, 0, 0, 2, -1, 0, 3, 3, 3, -1, 3, 0, -5, 3, -2, 0, -5, -2, -3, 0, -4, -1, 0, 2, 5, 1, 0, 5, 4, 1, 5, 2, 2, 2, 5, 4, 5, 4, 5, -1, 2, 1, 3, 1, 0, 2, -3, -2, 1, 1, -7, 0, -4, 0, -2, 2, -1, 6, 4, 0, -3, -1, 0, 0, 1, 5, 7, 6, 2, 6, 6, 0, 3, -2, -1, 3, -3, 0, -2, -3, -4, -1, -2, -3, 0, -3, -4, -2, -1, 2, 1, 1, 3, 3, -1, 3, 7, 6, 0, 6, 3, 6, 0, 6, 0, -1, 2, 0, 2, 1, -5, -2, -6, -1, -1, -2, 3, -2, 0, 0, 0, -1, 3, 6, -1, -1, -1, 4, 1, 1, 6, -1, 0, 1, 3, 2, 6, 0, 6, 0, -1, 0, -4, 4, -5, 1, 4, 2, -1, 0, 0, 1, 2, 6, 6, 0, 0, 7, 4, 7, 8, 7, 5, 4, 5, 6, 5, 8, 0, 7, 5, 3, 6, 3, -2, 4, -5, 1, 1, 4, 1, -1, 4, 6, 7, 0, 3, 5, 4, 1, 0, 8, 0, 4, 5, 3, 5, 1, 1, 5, 0, 9, 3, 1, 9, 0, 4, 6, -1, 0, 6, 2, 8, 5, 2, 7, 2, 4, 6, 7, 8, 0, 0, 0, 3, 2, 4, 4, 2, 3, 4, 3, 2, 4, 3, 7, 8, 8, 8, 11, 8, 6, 5, 12, 4, 6, 3, 5, 6, 4, -1, 1, 6, 2, 3, 3, 8, 1, 1, 1, 2, 6, 6, 5, 3, 1, 4, 12, 14, 13, 15, 9, 15, 8, 10, 9, 7, 8, 10, 9, 1, 3, 5, 5, 3, 6, 3, 2, 3, 3, 1, -2, 5, 3, 4, 5, 8, 7, 7, 7, 12, 11, 17, 9, 9, 12, 14, 11, 7, 7, 4, 8, 1, 6, 0, 3, -2, 0, 0, 3, 8, 2, 2, -4, 1, 0, 7, 2, 3, 5, 8, 16, 13, 12, 16, 12, 13, 17, 12, 7, 14, 7, 5, 5, 6, 5, -3, 1, 3, 2, 3, 2, 2, 2, -5, 1, 0, 0, 0, 0, 1, 9, 12, 14, 18, 22, 15, 16, 17, 17, 20, 19, 10, 11, 7, 1, 2, 2, 1, -2, -4, 0, 4, 3, 0, -4, 0, -4, -5, -1, 0, 3, 8, 7, 14, 12, 17, 23, 19, 19, 25, 17, 17, 13, 13, 14, 4, 4, 2, -6, 1, -1, 0, -3, -3, 3, 0, -3, 0, -1, -6, -4, 0, -5, 0, 11, 9, 19, 18, 19, 24, 20, 16, 25, 16, 17, 18, 13, 12, 4, -4, -8, -2, -5, -2, -5, -3, -1, 4, -4, -2, -1, -3, -6, -6, 0, 0, 9, 15, 15, 16, 19, 23, 20, 22, 18, 20, 24, 20, 11, 8, 6, -5, 0, -1, -2, 0, 1, 2, 0, 4, -4, -6, 0, 0, 0, -7, -2, -1, 6, 8, 11, 18, 22, 21, 21, 22, 30, 20, 24, 21, 7, 3, 1, -3, -2, -7, -2, -1, -4, 3, -2, -1, 0, -4, 2, -4, -2, -3, -1, 0, -2, 6, 7, 16, 24, 25, 18, 25, 20, 23, 16, 16, 7, 3, 2, -1, 0, -1, -3, -1, -4, 0, -2, 0, -5, 1, -4, -2, 3, 0, -6, 1, -2, 2, 4, 12, 17, 16, 18, 21, 18, 17, 10, 12, 6, 0, 0, -3, 1, 0, 0, 2, -4, -4, 2, -4, 0, -4, -4, 4, 4, -3, 4, 1, 0, 4, 1, 10, 10, 10, 12, 20, 16, 16, 8, 1, 0, 5, 0, -2, 0, 3, 0, 1, -3, -4, 2, -4, 2, -2, 3, 0, -1, 3, -1, 3, 1, -4, 4, 6, 3, 5, 12, 7, 11, 10, 2, 2, 3, -1, 5, 2, 5, 2, 6, 0, 0, -4, 2, -1, 0, 0, 1, 4, 3, 0, -3, 1, 0, -2, -3, -2, 2, 3, 7, 7, 0, 2, 0, -2, 0, 4, 2, 3, 5, 7, 2, 6, -3, 0, 7, 1, -3, -1, 0, 4, 1, 2, 0, 0, 2, 2, 3, 4, 0, 0, -2, 2, -2, -2, -6, -4, 3, -2, 1, -3, 1, 4, 0, 2, 1, 0, 0, 3, 2, 4, -3, 3, -2, 2, -1, 2, 0, 4, -3, -4, 0, -2, -4, 0, 0, -5, -1, -4, 1, -3, 3, 2, 1, 6, 0, 7, 3, -1, 7, 0, 4, -2, -2, 1, 0, 5, 1, 3, 3, 1, 0, 0, -6, -8, -4, -2, -4, -7, 0, -1, -4, -4, -2, 2, 0, 1, 0, 3, 2, 3, 9, 3, 3, 0, 1, 2, 1, 5, -3, 4, -4, 2, -3, -5, -2, -2, -3, -4, 0, -5, 0, -4, -4, -3, 0, 0, -1, 2, 5, 0, 3, 3, 2, -1, -2, 3, 7, 0, 6, -2, -4, -2, 2, 0, 1, -2, -3, -4, -2, 2, -4, -5, -6, 0, 0, -3, 0, -2, -2, 6, 2, 0, 0, 5, 8, -1, -1, 6, 3, 7, 2, 1, 0, -4, 0, -4, 2, -4, -1, -3, -1, 1, 2, 0, 2, 2, -2, 0, -4, 2, 1, 1, 3, 0, 0, -1, 0, 4, 4, 3, -1, 2, 0, 4, -4, 0, -4, 0, -3, 0, 0, -7, 0, -6, -3, 0, -5, 1, 0, 0, -2, 0, 5, 6, 0, 2, 6, 5, 2, 3, -1, 1, 1, 4, 0, 0, -4, -4, -2, -7, 0, -1, -1, -5, -3, -4, -4, -6, -6, 0, -7, 2, -4, 4, 1, 0, 3, 0, 1, 0, 4, -1, 0, 0, 1, -1, 0, 1, 0, 0, -2, -9, -3, -6, -7, -3, -5, -6, -5, -1, -8, -5, 1, 0, -3, -2, 1, 3, 0, 2, 8, 2, 7, -5, -8, -6, -12, -10, -16, -10, -14, -11, -11, -9, -12, -8, -17, -12, -11, -12, -13, -14, -14, -13, -11, -8, -9, -14, -10, -13, -8, -8, -13, -9, -11, -11, -12, -9, -7, -9, -6, -8, -8, -12, -6, -10, -8, -13, -15, -10, -9, -10, -8, -11, -12, -9, -13, -7, -14, -14, -13, -10, -5, -7, -4, -4, -5, -3, -4, -10, -9, -12, -7, -13, -12, -13, -12, -10, -9, -9, -14, -14, -12, -9, -14, -16, -11, -12, -13, -15, -5, -11, -5, -3, -5, -9, -5, -6, -5, -5, -8, -5, -9, -10, -5, -12, -6, -9, -10, -15, -8, -10, -16, -13, -12, -11, -17, -15, -15, -15, -14, -10, -8, -5, -3, -2, -7, -6, -8, -3, -8, -2, -7, 0, 0, -7, -11, -7, -9, -10, -12, -7, -12, -11, -10, -12, -15, -11, -17, -15, -18, -10, -8, -7, -6, -9, -11, -10, -6, -4, -10, -8, -3, -5, -7, -4, -5, -8, -6, -4, -13, -7, -11, -14, -14, -10, -18, -19, -17, -17, -19, -18, -19, -10, -11, -14, -12, -11, -7, -10, -10, -10, -7, -2, -6, -5, -3, -3, -6, -7, -10, -7, -4, -11, -11, -10, -8, -10, -17, -17, -16, -18, -23, -15, -13, -14, -10, -10, -13, -12, -8, -7, -7, -7, -1, 0, 0, -5, 0, -7, -4, -9, -5, -11, -4, -5, -10, -16, -12, -10, -18, -14, -19, -18, -15, -18, -14, -18, -15, -9, -12, -8, -3, -5, -9, -10, -7, -2, 0, 0, 0, -1, -2, -5, -6, -5, -11, -7, -9, -11, -12, -12, -15, -19, -16, -22, -18, -21, -17, -12, -13, -16, -11, -8, -3, -9, -9, -1, 0, -7, 0, -1, 1, -9, -1, -1, -2, -7, -13, -5, -11, -14, -9, -16, -17, -18, -14, -13, -12, -18, -16, -9, -8, -15, -17, -7, -9, -8, -8, -4, -1, -5, -5, -3, -3, -3, 0, -7, -2, -5, -12, -8, -11, -10, -9, -12, -17, -11, -12, -13, -18, -16, -10, -13, -8, -10, -11, -10, -5, -7, -8, -3, -2, -3, -1, 4, 0, -2, 0, -8, -2, -12, -7, -8, -11, -15, -9, -9, -16, -17, -17, -15, -16, -14, -9, -15, -12, -10, -6, -9, -10, -8, -9, -2, -5, 0, -2, -1, -5, -7, -5, -3, -12, -4, -6, -9, -14, -8, -6, -8, -7, -14, -9, -9, -9, -8, -11, -9, -14, -9, -11, -13, -10, -5, -11, -2, -7, 1, -1, 2, -5, -7, -8, -9, -9, -14, -9, -11, -9, -10, -13, -4, -9, -14, -7, -6, -11, -9, -8, -7, -7, -14, -12, -9, -9, -6, -8, -6, -2, -2, -3, 5, 0, -8, -12, -9, -12, -8, -11, -10, -7, -6, -7, -11, -8, -11, -9, -9, -13, -10, -10, -12, -6, -12, -12, -10, -16, -14, -9, -8, -3, -6, 0, 0, 2, -3, -9, -5, -10, -10, -11, -15, -14, -11, -3, -3, -2, -1, -9, -8, -6, -3, -8, -10, -5, -6, -11, -9, -13, -7, -13, -10, -6, -4, 2, 0, -2, -7, -10, -12, -6, -14, -18, -15, -10, -11, -10, -3, 0, -5, 0, -4, -4, 0, 0, -8, -12, -6, -10, -15, -9, -12, -10, -7, -3, -6, 0, 0, -4, -7, -10, -10, -5, -13, -13, -9, -8, -9, -4, -5, -2, -3, -6, -5, 0, -2, 2, -4, -8, -11, -10, -10, -9, -5, -10, -7, -5, 1, -1, 2, 0, -5, 0, -5, -6, -12, -6, -12, -10, -6, -3, -4, -1, -4, -4, -3, 1, -3, 2, -6, -8, -13, -7, -15, -8, -12, -6, -6, -3, -2, -3, -1, -4, -2, -6, -1, -9, -12, -6, -11, -9, -10, -13, -5, -1, 2, 0, 0, 3, -5, -7, -5, -6, -11, -12, -9, -7, -4, -7, -5, -7, -4, 0, -2, -3, 0, -6, -7, -7, -3, -5, -7, -10, -11, -6, -3, -5, -7, -5, -2, -2, -1, -3, -6, -12, -13, -3, -5, -9, -5, 0, -4, 0, -2, 1, -2, -2, -2, 2, -1, 0, -8, -6, -10, -12, -11, -10, -10, -11, -11, -4, -5, 1, -7, -6, -6, -12, -12, -3, -3, -3, -2, -5, -5, -2, -3, -2, 1, 3, 3, 1, 0, 3, 0, -1, -7, -7, -8, -9, -8, -8, -9, -7, -4, -6, -11, -17, -12, -10, -5, -11, -4, -2, -5, -2, -2, -4, -2, 7, 3, 1, 0, 3, 0, 1, -3, -5, -2, -2, -7, -9, -7, -9, -8, -13, -7, -14, -11, -12, -9, -5, -8, -2, -2, 0, -2, -5, -3, -1, -3, -2, -2, 4, 0, 1, -1, 1, 2, 1, -4, -3, -3, -4, -5, -6, -13, -13, -8, -12, -8, -15, -12, -11, -9, -5, -5, -1, -7, -1, -3, -1, 1, 4, 0, 5, 0, -2, 0, 1, 2, -3, -2, 0, 0, -3, -5, -9, -6, -13, -12, -6, -9, -14, -11, -9, -10, -3, -5, -4, -4, 0, -1, 5, 4, 0, 1, 5, 0, 0, 2, 1, 1, -1, -1, -5, 0, -3, -6, -10, -3, -11, -8, -9, -11, -6, -4, -9, -1, -2, -7, -5, 0, 2, -1, -3, 4, 2, 0, 5, 1, 2, 0, 5, -3, 3, -6, -1, -3, -3, -9, -2, -9, -9, -3, -8, -4, -5, -1, -3, 0, -7, -3, 0, -2, 2, 3, -4, 0, 7, 0, 0, 6, 4, 2, -2, 4, 2, -2, -6, -5, -1, -4, -9, -9, -1, 0, -7, 1, -2, 1, -2, -4, -4, -2, 3, 3, 7, 0, 0, 3, 0, 3, 5, 7, 1, 3, -4, 0, 2, 2, -1, -2, -6, 1, -3, -1, -2, -6, -2, -7, 1, -2, -8, -5, -1, -1, 0, 1, 0, -2, 3, 2, 0, -1, 3, 0, 3, 2, 0, -3, -2, -4, 0, -1, -3, -4, 0, -4, -5, -1, -1, -2, -4, -5, -1, -1, 0, -1, 4, 2, 4, 0, -2, 1, 1, 1, 1, 4, 4, -2, -2, 1, 1, -3, 2, -3, -2, -5, -4, -5, -4, -3, -5, 1, 0, -2, 3, -4, -2, -2, 5, 0, 1, 6, 5, 0, 7,
    -- filter=0 channel=7
    -1, 6, 6, 1, 0, 1, 3, 1, 5, 1, 4, -1, -1, -1, 3, 2, -1, 1, 4, -1, 3, 3, 2, 3, 0, 3, 8, 0, 6, 1, 9, 5, 1, 0, 0, -3, -4, 1, -4, 3, -3, -3, 1, -1, 1, 2, -5, 3, -4, -4, 0, 3, 3, 0, -3, 0, -1, -4, -5, -1, 2, 3, -1, 0, 2, -2, -3, 1, -2, 0, -5, -2, -5, -5, 2, -4, 0, 0, -3, -3, -3, 1, -3, -3, 3, -3, -2, 1, 1, -2, -8, -7, -4, -1, 2, 0, -1, 0, -1, -7, 0, -1, -8, -3, -1, -5, -2, -3, 0, -1, -6, -3, 0, -6, -3, -3, -3, -3, -7, -7, -6, -2, -5, -9, -1, 1, 4, -1, 1, -3, -3, -7, -3, -6, -10, -4, -9, 0, -5, 2, -7, 0, 0, -6, 1, 0, 3, -2, -2, 0, -8, -5, -8, -5, -6, -3, 0, -3, -1, 0, -3, -5, -5, -1, -3, -6, -5, -7, -3, -3, -6, 2, -3, 2, -3, 0, -3, -3, -1, 0, -3, -1, -5, -9, -6, -3, -7, -6, 3, 2, -4, 0, -1, 0, -7, 0, -7, -5, -12, -3, -1, -7, 0, -2, -1, 5, 1, -1, 6, -2, 2, 0, -4, -2, 0, -3, -6, -9, 0, 0, -3, 2, -3, -4, -2, -3, 0, -7, -8, -9, -9, -11, -6, -1, -2, 2, 1, 4, 3, 7, 0, 0, 0, 3, 1, -4, 1, -7, -1, -4, -8, -8, -2, -3, -2, 0, -3, 0, -2, -2, -2, -5, -2, -4, -3, -6, -4, 2, 2, 0, 5, 8, 5, 2, 6, 4, -3, 1, 1, -6, -8, -8, -4, 0, -3, -3, 0, 1, 0, -5, -5, -7, -4, -5, 0, -1, -5, -4, 0, 4, 7, 0, 7, 6, 8, 3, 5, 2, 4, 3, 2, 1, -6, -3, -2, 0, -5, 1, -1, 0, -3, -5, 0, -3, -4, 0, 0, 0, -3, -2, -1, 6, 3, 7, 0, 7, 5, 4, 4, 0, 1, 0, 0, 2, 2, 1, 0, -2, 1, 4, 3, 2, 3, 0, 2, 0, -1, 0, 5, -2, -2, -4, 1, 1, 7, 3, 4, 6, 6, 5, 0, 6, 7, -1, 5, 1, -1, 6, 0, 5, 0, -2, -1, 3, 6, 2, 6, 0, 1, 4, 5, 0, -2, 3, 3, 7, 5, 0, 2, 5, 3, 7, 4, 6, 4, 3, 0, 1, 5, 2, -1, 5, 7, 2, 3, 6, 2, 2, 5, 5, 0, 6, 2, 5, -3, -4, 3, 2, 4, 4, 1, 0, 0, 1, -1, 2, 2, -2, -1, -2, 2, 4, 0, 0, 3, 8, 1, 2, 4, 10, 5, 8, 5, 2, 0, 1, 1, 0, -1, -2, -1, 2, 2, 0, 2, 1, -4, -3, 1, -5, -7, -3, -3, 3, 2, 6, 4, 9, 7, 9, 11, 7, 2, 8, 6, 0, 4, 3, -2, -4, 0, -2, -6, -7, -9, -3, -4, -5, -9, -4, -8, -4, -4, 2, 0, -1, -1, 0, 1, 2, 10, 12, 14, 9, 12, 3, 2, 1, 3, 4, 0, -2, -10, -9, -4, -13, -8, -12, -7, -15, -10, -14, -5, -11, -8, -5, -3, 0, 2, 0, 3, 4, 11, 6, 11, 13, 11, 6, 2, 8, 6, 0, -1, -1, -8, -8, -15, -14, -18, -15, -19, -16, -13, -12, -7, -10, -3, 2, 2, 2, -2, 0, 2, 6, 4, 13, 11, 10, 7, 10, 8, 6, 3, 3, -2, -5, -6, -10, -11, -13, -16, -12, -11, -20, -15, -13, -6, 0, 0, 0, 2, 0, 3, 7, 5, 4, 5, 7, 11, 11, 3, 7, 6, 0, 4, 6, 3, -2, -5, -2, -6, -10, -9, -3, -1, -10, -10, -5, -3, -2, 1, 4, 0, -2, 1, 6, 1, 6, 11, 11, 9, 4, 5, 2, 7, 1, 4, 6, 6, 1, -4, 2, -3, 2, 1, 8, 7, 3, 3, 0, -1, 2, 0, 6, 3, 4, 5, 5, 3, 7, 8, 13, 10, 7, 1, 4, 3, 8, 2, 2, 7, 3, 2, 5, 4, 3, 8, 15, 14, 9, 4, 1, 0, 7, 4, 7, 1, 4, 1, 2, 6, -1, 2, 7, 10, 9, 9, 9, 5, 3, 9, 10, 10, 8, 9, 3, 3, 4, 7, 17, 17, 15, 7, 7, 9, 8, 5, 10, 9, 0, 1, 5, 4, 4, 7, 5, 7, 7, 8, 0, 6, 1, 3, 5, 5, 9, 3, 7, 7, 5, 12, 16, 9, 9, 7, 12, 10, 5, 9, 3, 2, 7, 5, 0, 1, 3, 8, 10, 10, 6, 3, 4, 1, 8, 8, 11, 4, 8, 6, 7, 6, 11, 9, 8, 8, 9, 8, 11, 9, 11, 13, 9, 5, 5, 3, 4, 1, 0, 6, 4, 10, 2, 6, 5, 8, 12, 5, 5, 6, 5, 8, 6, 3, 7, 2, 10, 7, 12, 11, 10, 6, 8, 13, 8, 9, 5, 6, 2, 2, 4, 9, 7, 4, 2, 2, 1, 10, 8, 4, 7, 9, 2, 8, 1, 6, 1, 6, 12, 5, 4, 4, 4, 7, 7, 6, 6, 7, 4, 5, 3, 0, 3, 7, 8, 10, 5, 6, 4, 9, 6, 10, 4, 8, 3, 9, 5, 1, 5, 8, 7, 7, 7, 6, 7, 8, 2, 2, 1, 3, 6, 5, 0, 8, 1, 1, 9, 8, 0, 1, 5, 2, 4, 6, 8, 9, 5, 5, 0, 7, 7, 1, 4, 0, 3, 5, 4, 4, 10, 9, 5, 4, 9, 0, 2, 0, 6, 6, 1, 3, 1, 1, 8, 7, 2, 6, 6, 0, 7, 4, 1, 2, 7, 5, 1, 5, 8, 4, 2, 4, 5, 8, 7, 1, 0, 4, 6, 0, 3, 1, 9, 5, 4, 7, 7, 4, 7, 2, 0, 7, 3, 6, 2, 6, 1, 8, 5, 5, 0, 1, 6, 9, 8, 4, 3, -1, 5, 0, 2, 0, 6, 0, 3, 7, 7, 6, 4, 2, 4, 2, 10, 11, 9, 4, 8, 10, 10, 10, 5, 11, 9, 12, 11, 5, 3, 7, 7, 2, 7, 9, 2, 2, 3, 7, 10, 8, 3, 6, 11, 6, 6, 9, 6, 6, 9, 10, 8, 10, 4, 4, 8, 4, 7, 5, 9, 7, 12, 8, 6, 9, 13, 9, 11, 11, 12, 8, 8, 5, 7, 2, 7, 8, 8, 6, 9, 6, 5, 11, 7, 5, 2, 6, 8, 3, 3, 6, 8, 8, 8, 6, 4, 3, 9, 8, 5, 3, 5, 9, 9, 8, 9, 5, 0, 4, 3, 0, 3, 4, 3, 8, 6, 6, 2, 3, 5, 7, 0, 2, 6, 9, 3, 6, 5, 2, 1, 2, 0, 3, 5, 3, 4, 2, 1, 4, -3, 3, -5, 0, 1, 0, 3, 0, 4, 0, 4, -1, 2, 4, 7, 5, 4, 9, 0, -3, 0, 2, -3, -2, 3, -1, 3, 1, 9, 0, 2, 5, -2, 0, -5, -1, -1, 0, 1, 2, 1, -1, 0, 2, 3, 0, 5, 0, 6, 2, 2, -7, -4, -1, -4, -4, -3, 0, 6, 0, 0, 7, 1, -2, 0, 1, -1, -4, -4, -6, 0, 3, 3, 0, -1, 0, 0, 4, 2, 1, -3, -2, -6, -9, -9, -3, -6, -5, 0, 2, 6, 2, 3, 3, 2, 1, 0, -8, -12, -5, -8, -7, -3, -7, -4, -1, 5, 5, 6, 4, 3, 1, 1, -2, -9, -10, -7, -6, -9, -9, -6, -4, -1, 2, 0, 3, 4, -4, -7, -5, -9, -7, -9, -12, -8, -5, -1, -4, -1, 0, 1, 1, 4, -3, 1, -2, -10, -3, -6, -13, -4, -3, -5, -4, 5, 0, -1, 7, -1, -1, 0, -10, -5, -7, -10, -13, -11, -6, -9, -4, -4, -7, 0, -5, -3, -6, -1, -9, -8, -12, -6, -12, -9, -7, -4, -7, 0, 1, 6, 3, -2, -4, -3, -3, -1, -9, -8, -8, -13, -8, -9, -8, -3, -11, -6, -4, -4, -8, -1, -4, -10, -4, -9, -12, -9, -3, -3, -6, 3, -3, 0, 6, 0, -4, -5, -3, 1, -6, -7, -13, -15, -5, -10, -10, -12, -8, -10, -9, -6, -4, -12, -5, -7, -12, -6, -6, -6, -3, 1, -2, -1, 1, 3, 5, 2, 5, -1, -2, -3, -6, -11, -10, -8, -14, -11, -12, -9, -6, -14, -11, -7, -5, -6, -7, -11, -12, -8, -7, -6, -1, 2, 0, 0, 6, 6, 5, 3, 6, -1, 0, 6, 0, -9, -6, -15, -9, -10, -10, -7, -9, -15, -7, -12, -13, -10, -8, -11, -11, -10, -7, -7, 1, 1, 5, 4, 6, 0, 8, 5, 9, 5, 2, 0, 2, 0, -10, -7, -6, -13, -12, -7, -7, -14, -11, -15, -9, -8, -14, -15, -11, -10, -5, -6, -3, 4, 1, 9, 2, 4, 10, 5, 4, 6, 8, 4, 1, -4, -10, -4, -13, -10, -14, -13, -17, -11, -11, -11, -9, -16, -14, -9, -10, -10, -3, 1, 0, 5, 8, 3, 9, 10, 11, 10, 6, 4, 3, 7, 4, 2, 0, -6, -15, -9, -16, -14, -14, -20, -12, -15, -19, -16, -9, -13, -9, -10, -5, 3, -1, 5, 4, 10, 10, 14, 9, 10, 11, 12, 5, 6, 3, 0, -3, -7, -9, -17, -12, -16, -20, -19, -20, -19, -21, -19, -10, -15, -14, -9, -6, 1, 0, 4, 6, 6, 9, 10, 15, 12, 11, 6, 11, 2, 6, 1, -1, 0, -6, -12, -15, -15, -16, -19, -16, -20, -17, -20, -9, -6, -2, 0, 2, 0, 5, 8, 3, 9, 12, 9, 15, 14, 6, 11, 9, 7, 5, 6, 2, 0, -8, -8, -12, -18, -9, -10, -11, -14, -12, -16, -8, -7, -2, 3, -3, -2, 0, 2, 6, 3, 6, 11, 9, 9, 8, 7, 8, 3, 3, 10, 6, 4, 0, 0, -1, -7, 0, -3, -2, -4, 0, -5, -1, 0, 3, 1, 4, 0, 1, 7, 8, 10, 10, 12, 8, 6, 8, 4, 3, 2, 9, 7, 9, 3, 4, 3, 0, 3, 11, 12, 13, 6, 4, 6, 4, 7, 8, 8, 2, -1, 3, 3, 7, 7, 11, 13, 8, 8, 5, 9, 5, 6, 8, 10, 10, 9, 9, 11, 5, 12, 20, 16, 20, 15, 16, 11, 12, 10, 8, 5, 10, 1, 3, 2, 4, -1, 7, 10, 12, 6, 9, 0, 0, 1, 2, 11, 13, 13, 12, 12, 9, 14, 18, 20, 20, 21, 13, 10, 15, 10, 11, 12, 11, 1, 5, 4, 1, 0, 8, 3, 11, 6, 3, 7, 5, 4, 9, 9, 14, 8, 8, 11, 12, 13, 19, 15, 19, 18, 12, 10, 11, 15, 16, 6, 9, 5, 4, -1, 3, 5, 1, 7, 9, 1, 5, 0, 1, 2, 3, 6, 12, 14, 7, 7, 3, 9, 16, 14, 18, 10, 12, 13, 10, 7, 8, 7, 5, 7, 6, 0, 2, -2, 0, 2, 5, -1, 0, 0, 2, 5, 11, 9, 8, 4, 5, 7, 10, 8, 10, 12, 7, 15, 9, 4, 12, 8, 7, 15, 8, 6, 5, 4, -2, 4, 2, 4, 4, -2, -2, 6, 6, 6, 11, 11, 3, 4, 8, 6, 4, 2, 11, 14, 8, 4, 11, 7, 9, 3, 5, 7, 10, 3, 1, -3, -2, 0, 6, 1, 0, -1, 3, -2, 6, 0, 1, 5, 3, 9, 5, 8, 0, 5, 11, 5, 5, 8, 1, 5, 3, 4, 11, 1, 8, 2, 3, -1, 0, 0, 0, 4, 0, 6, 0, -1, 3, 5, 0, 7, 8, 3, 2, 5, 3, 5, 1, 9, 3, 4, 8, 6, 3, 7, 0, 5, 7, 0, 0, 1, -1, -1, 0, 2, 7, 1, -1, 4, 4, 0, -2, 3, 0, 3, 3, 0, 5, 0, 7, 7, 6, 3, 0, 6, 0, 3, 0, 5, 1, 0, 5, -3, 2, -2, 4, 0, 5, -2, 3, 0, 2, 5, 3, 1, -1, 4, 0, 4, 4, 4, 2, 3, 4, 2, 2, 4, 0, 0, 1, 2, 3, 1, 0, 0, -1, 0, -1, 5, 2, 0, 2, 0, 7, 7, 3, 1, 3, 5, 6, 2, 8, 2, 10, 4, 2, 3, 7, 7, 2, 7, 1, 2, 4, 1, 3, 0, 4, 2, 3, 5, 9, 13, 14, 17, 12, 15, 15, 17, 13, 13, 14, 13, 10, 14, 11, 9, 9, 11, 16, 17, 12, 9, 13, 11, 18, 16, 18, 11, 16, 11, 12, 20, 14, 8, 10, 7, 10, 14, 9, 12, 12, 15, 11, 16, 7, 8, 12, 13, 12, 7, 11, 6, 12, 6, 7, 15, 12, 10, 7, 7, 13, 8, 15, 15, 7, 8, 4, 7, 7, 8, 7, 11, 7, 9, 13, 8, 7, 6, 10, 10, 7, 4, 3, 13, 6, 7, 6, 8, 10, 3, 5, 5, 3, 5, 10, 8, 6, 11, 5, 0, 5, 0, 1, 2, 5, 7, 8, 7, 3, 4, 8, 5, 3, 6, 3, 5, 6, 3, 7, 3, 3, 1, -1, 3, 2, 5, 11, 7, 9, 6, 2, 5, -2, 3, -6, -2, 1, 6, 5, 4, 4, 5, 9, 6, 4, 7, 3, 2, 6, 6, 3, 3, 0, 1, -4, 0, 6, 0, 6, 7, 7, 5, 1, 0, 1, -6, 0, -3, 1, 0, 6, 4, 9, 5, 4, 5, 3, 4, 6, 4, 3, 5, -3, -1, 0, 1, -4, 4, 5, 7, 1, 3, 5, 4, 0, 3, -2, -6, -10, -4, -6, 0, 4, 0, 6, 1, 9, 10, 10, 2, 7, 3, 2, -2, 0, -1, -8, -5, -5, -3, 0, 3, -2, 6, 5, 0, -1, -3, -1, -4, -7, -12, -4, -1, -5, -3, 5, 3, 1, 5, 7, 3, 5, 0, 0, -4, 0, -4, -11, -8, -1, -8, 0, 3, 4, 0, -3, -1, -7, 0, 0, -6, -8, -12, -5, -12, -1, 0, 0, 3, 0, 0, -1, 4, 0, 2, -5, 0, -9, -8, -6, -2, -3, -7, -2, -4, -1, 0, 0, -4, -7, 0, -6, -3, -6, -10, -6, -7, -8, 0, -4, 1, 1, -4, 0, 1, -1, 0, -2, -2, -7, -3, -11, -5, 0, 1, 0, -4, -3, 0, 0, -3, -5, -7, -5, -2, -4, -7, -10, -5, -1, 0, -5, -5, -6, -2, -6, 0, -6, -3, -4, -10, -7, -5, -7, -1, -2, 3, -5, -4, -2, -1, 0, 0, 0, -3, -2, -4, -5, -6, -14, -8, -10, -9, -8, -4, -3, -5, -7, -2, -8, -2, -4, -4, -10, -7, -3, -3, 0, -2, -5, -4, 0, -4, -4, -4, -4, -2, -4, -1, -4, -5, -11, -7, -10, -7, -3, -4, -5, -6, -3, -8, -2, -7, -3, -11, -7, -11, -2, -1, -2, 2, 1, 1, -3, -3, 2, -1, 3, 0, 3, 3, -4, -4, -10, -5, -3, -7, -9, -2, -7, -9, -11, -10, -4, -8, -12, -9, -14, -15, -10, -3, 2, 0, 0, -3, -5, 1, 3, -1, -1, 1, -3, 0, 1, -5, -9, -9, -11, -12, -12, -10, -7, -9, -7, -12, -11, -12, -11, -12, -11, -6, -8, -4, 0, 3, -1, 2, 0, 2, 4, -3, -4, 0, -1, -3, -2, -7, -8, -8, -13, -13, -15, -9, -14, -17, -12, -12, -14, -15, -14, -10, -16, -4, -9, -3, -5, -4, 2, 1, -1, -2, 0, -3, 0, 4, 3, -2, -4, -2, -1, -4, -12, -14, -16, -21, -17, -19, -13, -15, -12, -19, -15, -11, -12, -11, -6, -9, -1, 1, 0, 1, -2, 5, 0, 0, -2, -3, -1, -1, 0, -4, -8, -8, -15, -15, -16, -16, -20, -21, -15, -21, -18, -20, -18, -8, -8, -8, -4, -1, -8, -3, 0, -3, -4, -1, 0, -1, -6, -3, 0, -1, -1, -3, 1, -3, -13, -11, -11, -13, -15, -12, -13, -15, -14, -10, -12, -5, -6, -6, -2, -1, -6, -6, -3, -4, 0, -5, -3, -4, -4, -3, -3, -1, 0, -2, 2, 0, -3, -4, -10, -9, -9, -3, -11, -8, -5, -6, -7, -5, -4, -6, -8, -9, 0, -1, -6, -8, -5, 3, -7, -9, -6, -8, -3, -2, 0, 1, 3, -2, -2, -2, -2, -1, -4, 1, 3, 0, 2, 0, -2, 0, -1, -6, -8, -5, -2, -7, -5, -9, -9, -5, -6, -4, -7, -10, -1, 0, -6, -4, -4, -2, -1, 0, -4, 0, 1, 5, 4, 0, 0, -5, 0, -2, 0, -4, -6, -4, -10, -4, -8, -8, -6, -3, -1, -9, -8, -11, -4, -2, -7, 0, 1, -4, -1, 0, -5, 2, 5, 7, 3, 6, 5, -3, -4, 0, -1, 1, -5, -1, -6, -10, -12, -9, -5, -3, -10, -7, -6, -13, -5, -2, -1, -5, 0, -4, -1, -2, -7, 1, -1, 1, 0, 0, 3, 3, -5, 0, 0, -3, -4, -9, -12, -10, -15, -14, -9, -10, -11, -12, -13, -14, -12, -2, -5, -4, 1, -1, -8, -2, -6, -3, -5, 3, -5, 0, -5, -5, -3, -1, -2, -7, -2, -4, -8, -11, -13, -11, -10, -5, -7, -13, -9, -9, -7, -8, -2, -3, -2, -1, -10, -7, -2, -7, 0, -4, -3, -6, -5, -2, -2, -5, 0, 0, -3, -9, -11, -16, -9, -16, -9, -8, -7, -14, -10, -15, -6, -5, -9, -5, -4, -9, -4, -10, -6, -4, -8, -1, -2, -7, -8, -5, -10, -9, -7, -6, -8, -4, -6, -13, -15, -14, -13, -14, -9, -18, -10, -15, -9, -8, -10, -8, -11, -3, -5, -6, -7, -9, -8, -7, -8, -5, -4, -5, -6, -9, -9, -6, -5, -5, -12, -7, -15, -16, -18, -16, -13, -10, -12, -16, -7, -13, -14, -6, -11, -12, -9, -6, -7, -10, -12, -8, -7, -10, -14, -11, -12, -12, -12, -14, -11, -5, -16, -8, -16, -11, -13, -9, -16, -10, -16, -15, -11, -12, -8, -11, -11, -12, -9, -6, -15, -14, -12, -11, -7, -8, -15, -16, -15, -8, -8, -12, -13, -8, -15, -15, -11, -14, -16, -10, -12, -15, -19, -16, -16, -13, -11, -16, -11, -13, -9, -10, -9, -15, -8, -14, -7, -7, -15, -17, -11, -14, -14, -15, -17, -10, -17, -17, -12, -16, -18, -16, -11, -15, -16, -13, -15, -13, -7, -13, -7, -13, -14, -6, -14, -6, -10, -4, -6, -12, -6, -14, -14, -8, -15, -13, -8, -8, -9, -9, -11, -14, -14, -11,
    -- filter=0 channel=8
    -1, 2, -4, 0, -1, -1, -2, -2, 0, -6, -2, -5, -6, 1, 0, 0, 0, -2, -4, -2, -2, 0, -2, -6, 0, 1, 1, -2, -3, 2, 0, 4, 3, 3, 0, -4, -5, -7, -5, -2, 0, -4, -5, -5, -3, -4, -4, -2, -2, -3, -6, -5, -3, -2, -5, 0, -6, -5, -1, -1, 2, -2, -1, 0, 1, -3, 1, 0, -3, -2, -2, 1, -4, 0, -8, 0, -5, 0, -4, -1, -4, -2, -2, -4, -1, -2, 0, -4, -2, -4, 1, -2, -5, 3, 3, 2, -5, -3, -3, 0, -6, -5, 0, -1, -3, 0, -8, 0, 0, -5, -6, -2, -4, 0, -3, 0, -6, -2, -5, 0, -2, -7, 0, 1, 2, 2, -5, -3, -1, -2, -7, -1, 0, -5, 0, -5, -4, -8, -2, -3, -4, -8, -6, -7, -6, -1, 1, 0, -2, -6, -4, 0, -5, 0, -5, -1, -6, 0, -2, 1, -5, -8, -6, -2, -1, 1, 0, -2, -5, -1, -4, -6, -6, -9, -5, 1, -5, 0, -1, -5, -2, -1, -5, -7, 0, -5, -2, -4, -6, -4, -2, -2, -2, -3, -4, -1, -4, -3, 0, 0, -2, -7, -8, -2, -5, -7, -3, -3, -5, -1, 0, -6, -5, -6, -7, -1, -1, -4, -3, -4, -6, 0, -4, -3, -5, -3, 0, -6, -3, 0, 0, -5, 0, -8, 0, 0, 1, -1, -5, -2, -3, -1, 2, 3, -4, 0, -1, -4, -1, -7, -5, -2, -8, 0, -6, -4, -7, -10, -9, -3, -8, -1, 0, 1, 0, -6, -5, -5, -6, 0, -2, 4, 0, 1, 3, -2, 4, -4, 1, 0, -5, -3, 0, -3, 0, -1, -1, 0, -6, -10, -2, -4, -2, -1, -6, 1, 0, 3, 1, 0, 0, 4, 1, 6, 1, 1, 0, -3, -1, -3, 2, -2, -3, -5, -7, -1, -4, -2, -5, -3, -9, -11, -10, -8, -2, -5, -7, -4, 0, -2, 0, 0, 6, 3, 3, 0, 5, -1, 3, 4, 3, -3, -1, -4, 0, -6, -8, -3, -4, -7, -4, -1, -12, -10, -6, -4, -4, -1, -2, -4, -2, 2, 0, 1, 3, 0, 4, -1, 0, 3, 0, -2, 2, -2, -1, -5, 0, -5, -3, -4, -2, -8, -2, -2, -5, -13, -10, -12, -9, -5, -2, -4, 4, 0, 1, 4, 3, 0, 3, -3, -2, 5, -2, -1, -3, -3, -3, -3, -4, -6, -2, -6, -11, -11, -4, 0, -8, -6, -9, -8, -5, -3, -1, 0, 4, -3, 5, 6, 0, -1, 5, -4, 0, 3, -2, 3, -3, 0, 0, 1, -5, -8, -2, -6, -7, -6, -7, -5, -3, -3, -8, -9, -8, -5, -1, 2, -1, 0, -4, 2, 0, -2, -5, 0, 0, 0, 1, -3, -6, 0, 2, -1, -6, -5, -4, -4, -8, -10, -6, -7, -8, -5, -2, -3, -5, -8, -2, 0, -3, -2, 1, -2, -1, -5, -6, -6, -3, -2, -4, -7, -4, 1, -1, -1, 0, -6, -4, -7, -10, -4, -9, -8, -10, -12, -12, -3, -6, -5, 0, 2, -1, 0, -2, -4, -5, -4, 0, -1, 0, 0, 1, -2, -3, -1, -2, -2, -2, -2, -8, -10, -6, -11, -8, -3, -7, -10, -4, -3, -3, -6, 1, -2, 0, 2, 3, 1, -4, -3, -4, 2, 2, 4, 0, 1, 6, 1, -3, 0, -1, -5, -1, -4, -3, -2, -3, -1, -8, -4, -7, -7, 0, 0, 0, 4, 4, 5, 5, 0, 0, 0, 2, 3, 5, 10, 2, 7, 0, -1, 4, 3, -1, -2, 1, 0, -7, -7, -6, -2, -7, -9, 0, -1, -2, 0, -3, -2, 4, 1, -1, 3, -3, -1, 2, 5, 5, 10, 9, 7, 6, 0, -1, -1, 0, 0, -3, -1, -4, -4, -4, -2, -4, -3, -8, -2, -4, 0, -2, 2, -3, 3, 1, 0, 1, -2, -2, 6, 1, 1, 0, 5, 5, 2, 3, 3, 3, 0, 3, 3, -2, -4, -3, -4, -13, -2, -6, -4, -1, -1, 0, 0, 3, 0, 1, 2, 0, 6, 0, 7, 8, 5, 6, 0, 1, 4, 5, 2, -2, 0, -2, 4, -3, 0, -8, -4, -7, -8, -4, -6, -1, 0, -2, 2, -3, 4, 0, -2, 1, 1, -1, 6, 5, 3, 5, 2, 1, -1, 3, -1, 0, -2, -4, -2, 1, -6, -5, -13, -15, -4, -2, -4, 0, 0, 1, -4, 2, 0, 3, -2, 0, 2, 0, 0, 0, -5, -1, 0, -3, 2, -5, -1, -5, -5, 0, -3, -6, -7, -11, -11, -11, -11, -6, 0, -2, 2, -2, 0, -2, 0, -2, -1, 4, 1, -4, 0, -6, 0, 0, -1, -6, -2, -1, -4, 0, -4, -4, -6, -9, -11, -12, -12, -16, -16, -4, -3, -3, 2, 0, -5, 0, 0, 1, -1, 0, -2, -2, -3, -1, -1, 0, -7, -3, -1, -9, -7, -4, -10, -6, -5, -8, -13, -17, -13, -19, -17, -12, -3, -1, -5, -7, -8, -3, -3, -8, -5, 0, 0, -2, -6, -7, 0, -6, -6, 0, -7, -6, -7, -5, -11, -6, -7, -7, -10, -17, -15, -22, -20, -15, -11, -10, -10, -8, -10, -5, -4, -11, -11, -8, -9, -3, -8, -5, -11, -7, -7, -6, -7, -7, -9, -10, -11, -9, -14, -13, -11, -15, -15, -20, -17, -15, -9, -14, -7, -8, -13, -7, -9, -13, -12, -5, -6, -9, -8, -11, -8, -6, -8, -5, -8, -10, -14, -9, -11, -9, -16, -12, -20, -18, -19, -23, -22, -14, -16, -20, -13, -12, -12, -16, -10, -13, -15, -13, -12, -16, -17, -15, -9, -10, -9, -8, -13, -12, -18, -12, -15, -22, -18, -16, -24, -25, -26, -22, -27, -21, -17, -24, -22, -20, -17, -13, -22, -18, -18, -15, -18, -21, -15, -17, -12, -15, -19, -15, -18, -19, -23, -21, -20, -25, -20, -19, -25, -21, -21, -27, -24, -30, -21, -28, -20, -22, -28, -19, -24, -27, -26, -23, -25, -26, -27, -19, -20, -27, -27, -27, -22, -22, -29, -28, -26, -31, -30, -31, -22, -23, -23, 2, -2, 5, 0, 3, 4, 3, -2, 3, 1, 2, -3, 0, 2, 3, -1, 1, 0, 0, -2, 0, 1, -3, 0, 0, -1, 2, -2, 2, 3, 3, 0, -1, -2, 0, -2, 5, 0, -2, -2, -3, 0, 1, 0, -5, 1, -1, 3, -3, 1, 1, 0, 0, -2, 1, -4, -3, 3, -4, 0, 0, 0, 6, 0, 1, -1, 3, 3, 3, 5, 4, 1, 2, 0, -1, -2, 0, -3, -2, -3, 2, 3, 0, 0, 4, 5, 0, 1, 2, 2, 3, 1, 2, 5, 5, 0, 0, 2, -2, 3, -2, 5, 2, -2, 3, 1, 4, 0, 5, 1, 0, 1, -2, 2, 0, 3, 2, 1, -2, 1, 3, 3, 0, 4, 2, 0, -1, 5, 3, 3, -4, 0, 0, 4, 0, 1, 0, 0, -4, -1, 2, 3, 1, 5, 2, 4, -2, -2, 1, 2, 2, -2, -1, 4, 0, -2, -1, 0, 4, 2, 0, -1, 1, 0, -1, -1, 6, 0, 0, -1, 1, -4, 0, 4, 2, 0, 0, 1, 5, 0, -1, 2, -4, 2, 1, 1, 1, 0, 0, -3, -2, 1, -2, -4, 0, -2, 2, 6, 0, 5, 3, 4, -4, 2, 5, 5, 5, 3, -2, 0, 2, 3, 2, 4, 1, 1, -1, 1, 2, -1, 0, -4, -2, 2, 2, 0, 3, 1, 1, -1, 1, 3, 1, 0, 1, -2, 0, 7, 8, 1, 6, 0, 3, 1, 1, 1, -1, 3, 0, -2, -2, -1, 1, -1, 2, 2, -6, 2, -4, 4, 1, 2, 0, 3, 3, -1, -1, 5, 6, 1, 6, 0, 4, 1, 7, 8, 3, 6, 0, 5, -1, 5, 3, -2, 2, -3, -2, 0, -1, -5, 0, -1, 2, -2, 4, 5, 7, 8, 1, 5, 2, 2, 10, 2, 0, 4, 7, 4, 2, 6, 4, 4, 3, 4, 3, 0, -2, 2, 4, -1, 0, 0, -2, 3, 2, -3, 1, 0, 6, 2, 4, 8, 10, 9, 9, 5, 0, 5, 6, 1, 4, 5, -3, 3, 0, 5, 0, 2, -3, 0, -2, -3, -5, -4, -1, -2, 0, 3, 0, 6, 4, 2, 5, 9, 10, 3, 2, 3, 3, 2, 2, -3, 3, 3, 1, 4, 6, -2, -1, -1, 4, 0, 1, 0, -4, -8, 0, -3, -2, 1, -2, 0, 6, 2, 4, 4, 6, 2, 4, 0, 5, 7, 1, 4, -1, -2, -2, 1, 0, 4, -3, -4, -3, -3, -2, 4, -2, 2, 2, 1, -1, 2, -1, 6, 3, 6, 1, 4, 4, 2, 0, 2, 1, 5, 2, 6, 3, -2, 4, 0, 5, 2, 0, -3, 0, -2, 0, 4, 2, 0, -2, 2, 3, 1, 3, 2, 3, 4, 1, 2, 4, -2, -2, -3, -2, -2, -1, 2, 0, 0, 4, 1, 1, -1, -3, 0, 0, -3, -3, -2, -1, 1, -4, -3, 0, 3, -2, 6, -1, 3, 5, 6, 0, -3, 0, -1, -4, -4, 3, -5, 3, -2, 2, 6, 0, 0, 0, 0, -6, 2, -3, 2, 3, -2, 2, -1, 2, 3, -1, -3, 4, -1, -4, -3, -4, -3, 1, 0, 1, 5, 1, 1, 1, -2, 2, 2, 0, -2, -3, -3, 0, 3, 1, 2, 1, 1, -6, -5, 0, 0, 0, 0, -3, 2, 1, 0, 3, 0, 3, 0, 1, 4, 2, 4, -1, -2, 0, 0, 0, 0, -2, 0, -2, 0, 2, 7, -1, 0, -3, 3, -3, 4, 2, -1, -2, 6, -2, 2, -3, 0, 4, 1, 9, 1, 3, 7, 8, -1, 5, 0, 0, 3, 3, -1, -2, -2, 0, 0, 5, -4, 2, 2, 1, -4, -2, 0, 0, 2, 3, 1, 1, 3, -4, -1, 5, 8, 2, 5, 4, -5, 2, -3, 3, -1, 1, 2, -3, 0, -2, 8, 6, 0, 0, 3, -2, -1, -1, 1, 0, 1, 2, 0, 1, -4, -4, 4, 1, -1, 4, 4, 0, 1, -2, -2, -5, 2, 0, 5, 0, 5, 4, 6, 3, 3, 0, 1, -5, -2, -7, -3, -4, -4, 1, 1, -3, 4, 2, -2, 6, 5, 0, 3, -2, -3, 0, 4, -3, 3, 1, -1, 3, 6, 6, 5, -3, 4, 7, 2, -4, -7, -4, -1, -2, -3, -2, 0, -2, 1, 0, 1, 1, 1, 1, 0, -2, -1, 4, 0, -3, 0, -2, 1, 3, 4, 0, 1, 1, -1, 0, 0, 1, 1, 0, 0, -3, -5, 0, 1, -6, 2, -4, 0, -1, -2, -2, -5, -4, -2, -3, -1, 1, 1, 2, 0, 5, -1, 3, 3, -6, 3, 5, 4, 4, -2, -4, 3, -3, 0, -3, -4, 2, 2, 1, -7, -4, -5, -5, -6, -7, -6, -7, -6, 1, -1, -5, -5, 0, -4, -1, 0, -3, 0, 5, 0, 4, 3, 3, -4, 0, -1, -4, 1, -3, -4, -4, -5, -4, 1, -5, -1, -4, -4, -7, -2, -1, 0, -4, 3, 4, -3, -3, 0, -6, 0, 4, 1, 5, 6, 5, 2, 0, 2, 0, -6, -5, 3, 0, -2, -4, 2, -3, -1, 0, -5, -3, 0, 1, -5, -2, -2, 2, 1, 0, -4, -10, -1, 0, 0, 0, -2, 4, 2, -1, 1, -1, -3, -3, -2, 0, 0, -3, 0, -6, 1, -3, 0, -1, -2, -4, 0, 2, 0, -2, 0, -9, -3, -7, 0, -4, 0, 0, 4, 3, 0, -5, -2, 0, -3, -5, -7, 0, -1, -5, 0, 0, -5, 0, -4, 0, -6, -5, -2, -5, 1, -2, -6, -3, -10, -10, -2, -4, -2, -7, -1, -7, 0, -6, -8, -7, -6, -7, -1, -3, -7, 0, -7, -6, -3, -2, -8, -2, -7, -5, -5, -11, -4, -7, -2, -3, -3, -12, -5, -3, -5, -10, -4, -9, -7, -7, -8, -7, -9, -5, -11, -8, -11, -6, -3, -3, -4, -8, -5, -5, -9, -7, -5, -4, -5, -8, -9, -8, -7, -9, -6, -6, -13, -8, -13, -9, -11, -8, -13, -13, -15, -10, -10, -11, -14, -10, -9, -14, -9, -13, -10, -12, -13, -9, -12, -13, -13, -12, -11, -10, -7, 5, 13, 8, 8, 9, 9, 3, 6, 8, 10, 10, 6, 2, 9, 7, 9, 6, 8, 3, 2, 2, 5, 4, 5, 9, 6, 8, 4, 6, 9, 9, 15, 9, 11, 12, 14, 12, 5, 5, 10, 3, 3, 2, 4, 7, 9, 6, 9, 4, 5, 5, 3, 5, 9, 7, 5, 10, 4, 10, 9, 10, 7, 6, 6, 5, 4, 7, 12, 9, 12, 5, 11, 4, 8, 2, 5, 4, 10, 11, 7, 11, 6, 12, 5, 12, 10, 2, 11, 5, 4, 8, 5, 8, 11, 5, 10, 8, 8, 7, 8, 10, 13, 7, 11, 4, 9, 10, 10, 9, 6, 4, 10, 12, 8, 10, 8, 11, 8, 9, 3, 7, 2, 5, 8, 9, 8, 10, 8, 11, 4, 4, 5, 9, 13, 10, 7, 6, 7, 10, 5, 6, 8, 8, 8, 3, 8, 10, 11, 7, 2, 3, 10, 8, 4, 3, 10, 11, 8, 7, 7, 3, 4, 4, 13, 6, 7, 5, 8, 11, 5, 2, 3, 3, 8, 5, 9, 7, 11, 8, 2, 7, 8, 4, 5, 9, 3, 8, 12, 4, 5, 3, 8, 11, 12, 4, 6, 11, 7, 6, 9, 9, 5, 8, 3, 8, 6, 4, 2, 6, 3, 8, 7, 8, 8, 3, 6, 3, 10, 8, 4, 5, 7, 9, 2, 11, 3, 9, 8, 7, 7, 11, 5, 8, 4, 5, 6, 5, 6, 10, 8, 4, 5, 8, 10, 4, 9, 10, 10, 8, 3, 7, 3, 6, 2, 7, 5, 7, 4, 5, 7, 13, 10, 12, 14, 9, 6, 6, 7, 9, 7, 3, 8, 3, 8, 3, 9, 3, 5, 9, 8, 11, 7, 10, 6, 3, 9, 9, 7, 5, 4, 5, 6, 9, 5, 13, 7, 11, 8, 11, 13, 12, 3, 8, 4, 5, 3, 3, 7, 10, 8, 11, 9, 10, 4, 8, 6, 3, 4, 10, 12, 9, 3, 6, 8, 6, 5, 4, 11, 6, 5, 13, 15, 6, 11, 3, 9, 8, 4, 8, 1, 8, 3, 8, 10, 4, 10, 7, 9, 9, 5, 12, 5, 8, 5, 2, 8, 5, 4, 7, 12, 10, 8, 7, 13, 13, 5, 8, 4, 9, 3, 9, 1, 5, 1, 8, 7, 4, 2, 2, 2, 10, 4, 9, 7, 4, 4, 2, 8, 11, 9, 5, 7, 12, 11, 5, 11, 6, 9, 0, 5, 5, 2, 2, 7, 3, 5, 1, 8, 4, 8, 6, 1, 7, 3, 6, 7, 9, 11, 9, 6, 7, 6, 4, 8, 4, 10, 7, 7, 10, 8, -1, 1, -3, 0, 4, 7, 3, 0, 3, 8, 5, 5, 6, 7, 8, 7, 9, 13, 8, 8, 6, 7, 10, 5, 1, 3, 8, 1, 6, 8, 5, -1, -1, -1, -3, 4, 2, 1, 7, 6, 6, 4, 9, 6, 1, 9, 2, 6, 6, 9, 15, 8, 4, 6, 8, 1, 1, 5, 5, 8, 6, 2, 0, 1, 0, -2, -4, 0, 0, 1, -1, 0, 1, 7, 1, 2, 1, 3, 2, 8, 8, 14, 14, 6, 5, 2, 3, 9, 5, 4, 3, -2, 1, 0, -1, 2, 2, 2, 3, 5, 0, 0, 0, 2, -1, 4, 7, 2, 2, 0, 3, 2, 13, 13, 16, 6, 4, 5, 2, 0, 3, 4, 4, 5, 3, 3, 5, -1, 6, 0, 3, 2, 2, 4, 0, -2, -1, 1, 1, -3, 2, 5, 8, 5, 7, 12, 14, 9, 7, 10, 1, 0, 7, 3, 0, 3, 5, 3, 0, 4, 0, 3, 8, 7, 3, 0, 0, -1, 4, -3, 2, 2, 0, 0, 4, 10, 15, 12, 15, 14, 11, 9, 0, 4, 4, 3, 0, 3, -4, 2, -1, -1, -3, 0, 5, 2, 3, 0, -2, 1, -1, 0, -3, -1, 4, 5, 8, 9, 15, 13, 13, 17, 10, 5, 0, -2, 2, 1, 2, 2, -2, -1, 0, 2, 0, 2, 3, 2, 1, 4, 1, 0, 0, 2, 2, 1, 6, 0, 6, 11, 15, 18, 14, 9, 10, 4, 1, 4, -3, -3, -6, 0, -4, -3, -3, -4, -1, 3, 3, 2, 0, 0, -1, -5, 1, -4, -2, 3, 0, 6, 6, 7, 9, 17, 18, 10, 13, 7, 0, -2, -3, -1, 1, -5, 1, 2, 0, -4, 1, 1, 2, 1, 2, -1, -3, -3, -1, -3, 0, -1, -2, 4, 10, 13, 16, 14, 10, 16, 14, 9, 10, 2, -1, 1, 3, -1, 0, 2, -1, 2, 0, -1, -6, -8, -7, -6, 0, 0, -1, 0, 4, 1, 4, 5, 6, 10, 14, 9, 11, 15, 11, 9, 13, 5, 0, 6, 2, 0, 0, 2, 0, -3, -1, 0, -8, 0, -1, -4, -5, 0, 0, 0, 3, 4, 4, 9, 4, 10, 12, 11, 12, 12, 9, 9, 14, 11, 3, 4, 0, 3, 3, -1, 2, 1, 0, 4, 1, -1, -4, 0, -1, 2, 1, -2, -2, 6, 5, 10, 7, 8, 9, 16, 12, 14, 12, 12, 10, 10, 6, 6, 4, 4, -1, -1, -1, 0, 0, 1, 3, 2, 1, 3, 4, -1, 0, 3, 4, 5, 10, 9, 9, 7, 10, 14, 10, 10, 12, 16, 13, 6, 4, 5, 8, 1, -3, -2, 4, 3, 0, -1, 0, -1, 6, 3, 5, 2, 6, 0, 7, 9, 4, 10, 11, 12, 13, 6, 7, 10, 8, 13, 15, 12, 5, 6, 5, 2, -1, 4, 5, 6, 4, 0, 0, 1, 4, 3, 0, 2, 7, 1, 0, 1, 2, 8, 7, 15, 7, 7, 10, 9, 14, 5, 10, 4, 2, 7, 6, 4, 0, 5, -1, 0, 0, 3, 2, 6, 2, 1, 6, -1, 1, 4, -1, 7, 2, 4, 11, 9, 8, 6, 6, 3, 12, 4, 8, 2, 3, 3, 5, 2, -2, -1, -3, -2, 1, 2, -3, -1, 4, 0, 0, 5, 5, 2, 1, 0, 4, 7, 4, 9, 9, 4, 4, 5, 3, 1, 3, 0, 0, 3, 2, -4, -6, 0, -5, -2, -6, -3, -4, -6, -3, -2, -2, -2, -1, -5, -3, -2, 0, -1, 2, 2, 3, 2,
    -- filter=0 channel=9
    1, 3, 0, 5, 6, 8, 0, 8, 8, 3, 5, 3, 0, 3, 6, 3, 8, 8, 2, 5, 7, 4, 6, 1, 5, 1, 0, 6, 5, 0, 5, 2, 4, 3, 0, 3, 5, 5, 0, 0, -1, 2, 2, 0, 1, -3, 3, 2, 2, 1, -1, 4, 5, 0, 1, 2, 0, 3, 6, 4, 0, 3, 4, -2, 2, -1, 6, 0, 0, 5, 5, 0, -4, -1, -2, -8, -6, 0, -6, 0, -1, 3, -5, 1, -3, -5, 0, -5, 2, 4, 3, 1, 2, -1, 0, 0, 6, 4, 4, 6, -1, 3, -3, -2, -2, -1, -8, -2, 0, -7, -5, 0, -3, -3, -9, -3, 0, -9, -6, -4, 1, -1, 3, 2, 0, 0, 5, 2, 1, 5, 4, 0, 0, -1, 0, 0, 3, -4, -7, 0, -1, -5, -4, -4, 0, -4, -1, -6, -7, -1, -5, -1, -2, 0, 2, -1, -2, 5, -3, 1, 7, 0, -2, -2, 2, 5, 0, 4, 3, 2, 2, -5, -1, -7, 0, 1, 0, 0, -8, -5, -1, -8, -4, -4, 1, -4, -2, 1, -4, -2, 0, 2, 2, 2, 4, 3, 3, 2, 0, -1, 0, -3, 1, 0, -3, -5, -6, -6, -1, -1, -8, -8, 0, -1, -3, -2, 4, 2, 2, 2, 3, -4, 1, 2, 3, -1, 0, -2, -2, 0, 1, 2, -3, 0, -1, -1, 0, -1, -3, 0, -4, -3, -7, -8, 0, 2, -2, 1, 5, 4, 3, -2, 0, -3, -1, -3, 1, 1, 2, -2, 1, 2, 6, 1, 2, -4, -1, 0, 2, 0, 0, 1, -3, -4, -3, -1, -1, -1, -4, 3, 4, 0, 2, 4, 2, 4, -3, 0, 3, 1, 2, 0, 0, -2, 0, 0, 1, 0, 1, 3, -3, -2, -2, 4, 1, -5, -7, 0, -2, -4, 2, -2, 0, -2, 4, -3, 0, 0, -3, -4, 1, 0, 0, -1, 1, 1, 5, 0, 0, 0, -1, -5, 0, 0, 3, 3, 1, 0, -3, 0, -3, 3, -2, 3, 0, 1, -3, -3, 0, -4, 0, -1, 2, 3, 4, 0, 0, 3, 0, -4, 2, -2, 1, -5, -4, 3, 3, 5, 0, 3, 1, 3, 2, -3, -4, -2, 1, -2, -4, -1, -4, -1, -1, -8, 0, 0, -2, 1, -2, -3, -1, -3, -2, -2, -3, -3, 0, 3, 3, 5, 0, -1, 4, -1, 0, 0, 3, -4, -1, 3, 0, -2, -2, 4, -3, -5, -8, 0, -4, 1, 1, 0, 0, -1, -3, -1, -3, 2, -4, 0, 0, -1, 1, 0, -1, -2, -3, -2, 0, 0, -1, 0, 5, 3, -1, 6, -6, -1, -2, -4, -5, -3, -1, 1, 1, 0, 2, 0, 3, -3, 0, 2, 8, 6, 7, 7, 0, 2, 0, 0, -3, -1, 0, 2, 4, 5, 3, 2, -4, -5, -7, -1, -4, -1, -3, -4, 0, 1, 3, 2, 0, 2, 5, 8, 9, 13, 6, 5, 10, 11, 2, 9, 1, 0, 6, 0, 2, 3, 3, 1, 0, -6, -11, -1, 2, 0, 0, -4, 1, 3, 1, 3, 3, 11, 10, 9, 9, 15, 16, 11, 10, 12, 13, 13, 6, 4, 7, 9, 4, 7, 3, 0, 2, -3, -4, -7, -3, -1, 1, -1, 0, 6, 4, 3, 3, 8, 9, 18, 18, 16, 13, 12, 8, 10, 14, 11, 5, 5, 6, 5, 6, 8, 2, -2, -1, -6, -8, -2, -3, -3, 3, -2, -1, 4, 7, 9, 5, 9, 7, 16, 10, 15, 18, 17, 13, 12, 8, 5, 8, 5, 6, 6, 1, 0, 2, -3, 0, -6, -9, 0, -1, -3, -7, 0, 0, 4, 4, 8, 9, 3, 7, 4, 14, 11, 13, 6, 4, 8, 2, 6, 1, 3, 1, 1, 0, 0, -3, 0, -1, -10, -1, -2, -8, -2, -7, -1, -5, 0, 0, 3, 2, 0, 1, 2, 6, 7, 7, 1, 5, -2, -3, 5, 3, -4, -4, -4, -3, -7, -9, 0, -7, -1, -2, -6, -3, -9, -4, -8, -4, -9, -5, -2, -7, -1, -4, -6, 2, 1, -5, -5, -4, -4, -6, 0, 0, -8, -8, -7, -4, -6, -5, -4, 0, 2, 1, -7, -1, -9, -7, -10, -8, -8, -6, -7, -11, -5, -9, -5, -7, -8, -5, -7, -7, -7, -8, -4, -2, -9, -9, -11, -13, -8, -8, -1, 4, -3, 3, 1, 0, -5, -4, -9, -10, -14, -13, -8, -9, -9, -5, -3, -9, -9, -5, -7, -8, -7, -5, -4, -9, -7, -6, -5, -6, -4, -3, 0, 5, 6, 9, 6, 4, -3, -1, -5, -12, -6, -10, -5, -3, -8, -4, -8, -8, -3, -3, -2, -1, -8, -3, -8, -6, -6, -8, -10, -6, 2, 1, 3, 3, 3, 12, 4, 0, 0, -3, -5, -11, -8, -15, -12, -10, -10, -5, -11, -8, -3, -2, -5, -6, -7, -9, -10, -4, -7, -9, -6, -9, 0, -4, 3, 9, 6, 12, 3, 2, 7, 1, -2, -12, -11, -11, -7, -5, -8, -5, -5, -10, -4, -4, -7, -4, -8, -4, -3, -5, -5, -6, -11, -10, -6, 0, 2, 3, 4, 15, 6, 5, 0, -3, -5, -2, -9, -7, -3, -8, -2, -4, -1, -4, -7, 1, 0, -6, -5, -9, -5, -7, -2, -8, -7, -4, -3, -2, 7, 5, 8, 19, 14, 4, 1, 3, 0, -4, -8, -2, -4, -5, -2, -6, 0, -2, -7, -8, -2, -7, -6, -6, -4, -3, -5, -7, -3, -1, -2, 7, 6, 12, 11, 20, 17, 11, 10, 1, 3, 2, 2, -2, -2, 0, -2, -3, 0, 2, -3, 2, -3, 0, -2, 0, -4, -1, 1, -4, -1, 2, 6, 6, 11, 13, 16, 17, 16, 14, 8, 5, 11, 2, 3, -2, 3, 0, 4, 2, 2, -1, 3, 0, 0, 3, -1, 6, 4, -1, 0, 3, 1, 3, 7, 13, 16, 9, 13, 19, 16, 18, 19, 18, 12, 14, 9, 6, 5, 10, 12, 13, 12, 8, 13, 8, 11, 14, 7, 11, 7, 16, 9, 13, 12, 14, 14, 16, 20, 14, 17, 8, 6, 8, 12, 10, 14, 9, 10, 9, 9, 9, 9, 11, 7, 6, 11, 10, 12, 16, 9, 8, 15, 7, 14, 13, 6, 12, 11, 9, 12, 14, 10, 7, 6, 12, 6, 4, 10, 13, 7, 6, 4, 3, 6, 1, 3, 2, 0, 3, 9, 3, 5, 8, 1, 11, 11, 4, 11, 7, 5, 6, 13, 9, 9, 5, 4, 8, 4, 3, 11, 3, 2, 2, 1, -3, -4, -5, -4, -3, 2, -1, 2, 2, -4, -2, 1, 5, 5, 1, 6, 12, 5, 9, 7, 5, 4, 9, 3, 10, 9, 7, 10, 4, 4, 4, -3, -1, -3, 0, -2, -1, -7, -5, -2, -3, -2, -4, -2, 2, 1, 0, 8, 4, 6, 8, 9, 7, 4, 5, 7, 8, 6, 8, 6, 4, 5, 4, -4, -3, -7, -8, -4, -3, -4, -4, -3, -5, -4, 0, -2, 0, 0, 1, 3, 7, 2, 1, 7, 7, 1, 7, 0, 2, 6, 3, 1, 2, 5, 1, -4, 0, -8, -6, -3, -6, -2, -6, -4, -5, -7, -8, -2, -3, 0, -2, 5, 3, 3, 6, 1, 2, 8, 2, 4, 3, 4, 3, 6, 2, 0, 3, 1, -7, -1, -4, -7, -8, -9, -10, -5, -10, -10, -9, -3, 0, 2, 3, 1, 1, 5, 7, 6, 1, 2, 5, 6, 3, 3, 3, 6, 6, 0, -4, -2, -2, -7, -12, -11, -5, -7, -4, -11, -5, -5, -6, -3, -2, 4, 2, 6, 5, 0, 3, -1, 1, 0, 0, -1, 4, 5, -1, 5, 2, 2, -2, -5, -3, -7, -2, -8, -9, -8, -2, -6, -7, -2, -1, 2, 2, 1, 1, 0, 5, -1, 2, 5, 1, -4, 6, 2, -1, -1, 0, 5, 2, 2, 0, -1, -1, -5, -6, -4, 0, 0, -3, -9, -8, -4, 0, -2, 0, 3, 0, 3, -1, 0, 1, 0, 0, 1, 0, 0, -3, 0, 4, 0, -2, 2, 3, -2, -6, -8, -5, -4, -2, -4, 0, -3, -4, 0, -1, -4, 3, 0, -2, 2, 3, -3, -5, -5, 0, -3, -6, -6, -2, 0, 0, -2, 1, -4, -7, -6, -2, -8, -2, -6, -2, -4, -5, -6, -7, -3, -5, -1, -7, -4, -3, 0, -4, -1, -3, -1, 0, -4, -7, -4, 0, -7, -3, -1, -3, -3, -4, -3, -6, -6, -2, 0, -3, 0, -2, -4, 0, 0, -7, -3, -2, -2, -3, 1, -3, -2, -6, -3, -6, -11, -12, -7, -7, -6, 0, -4, -3, -8, -6, -4, -6, -6, -3, -6, -4, 2, -5, -1, -7, -7, -7, -8, -7, -2, -8, -6, -1, -7, -5, -3, -10, -10, -8, -6, -10, -8, -4, -8, -8, -5, -5, -8, -4, -2, -3, -4, -3, 0, -2, 0, -1, -2, -2, -7, -7, -3, -2, -4, -8, -7, -10, -6, -10, -10, -17, -12, -5, -9, -3, -10, -10, -6, 0, -3, -2, 0, -5, -2, -3, -1, 4, 6, 0, 1, 2, 0, -4, -1, -6, -7, -7, -7, -3, -7, -10, -15, -18, -10, -7, -8, -9, -4, -9, -1, -2, -6, 1, -2, -2, 1, 1, 6, 5, 2, -1, 3, -1, 3, 0, -6, -3, 0, -2, -1, -5, -10, -14, -16, -11, -7, -5, -8, -9, -5, -4, -7, 0, -8, -5, 5, 1, 3, 8, 6, 11, 10, 4, 5, 0, 4, 0, -4, -7, -5, -4, -8, -5, -11, -12, -11, -10, -16, -8, -11, -13, -7, -8, -6, -7, -8, 0, -4, 0, 1, 7, 1, 2, 0, -2, 0, -2, -1, -8, -4, -6, -10, -8, -5, -9, -12, -9, -14, -10, -8, -16, -16, -10, -10, -5, -4, -4, -4, -7, -9, -4, -2, 4, 1, -1, -1, -5, -5, -8, -2, -7, -10, -13, -12, -9, -10, -8, -8, -13, -13, -11, -10, -12, -12, -10, -8, -9, -9, -10, -8, -3, -5, -3, -2, -1, -2, -1, -1, -4, -11, -8, -10, -6, -11, -13, -10, -10, -11, -14, -13, -10, -11, -10, -10, -9, -10, -11, -16, -15, -15, -15, -9, -9, -15, -11, -4, -12, -10, -9, -9, -13, -9, -9, -5, -13, -16, -17, -13, -14, -21, -18, -12, -11, -8, -9, -9, -13, -12, -13, -16, -13, -15, -10, -12, -11, -8, -16, -10, -11, -13, -9, -7, -9, -10, -15, -9, -8, -17, -17, -17, -17, -18, -16, -13, -5, -11, -5, -6, -11, -13, -12, -17, -9, -16, -17, -11, -12, -15, -12, -8, -12, -10, -11, -12, -5, -13, -14, -12, -11, -10, -18, -14, -12, -11, -10, -11, -7, -9, 2, -3, -3, -11, -6, -10, -12, -12, -12, -17, -13, -6, -12, -12, -8, -13, -5, -8, -7, -8, -9, -14, -12, -10, -13, -16, -13, -9, -12, -3, -2, -7, 2, -5, -1, -4, -5, -9, -14, -14, -13, -14, -12, -14, -12, -14, -10, -12, -8, -10, -5, -7, -12, -14, -12, -14, -10, -12, -11, -3, -8, -6, 2, 1, 3, 0, 2, 0, -3, -5, -8, -15, -12, -14, -15, -14, -15, -12, -7, -13, -11, -7, -13, -7, -15, -9, -12, -11, -15, -13, -13, -12, -10, 0, 0, 0, 6, 4, 2, -6, -1, -10, -11, -9, -10, -12, -6, -7, -10, -8, -7, -12, -7, -8, -8, -14, -8, -9, -10, -7, -9, -10, -10, -5, -1, 2, 3, 8, 7, 4, 4, -3, -8, -8, -4, -10, -9, -8, -12, -9, -6, -8, -6, -4, -4, -2, -8, -11, -7, -10, -9, -13, -13, -11, -7, -5, 0, 5, 7, 5, 5, 7, 6, -1, 2, -4, -2, -4, -7, -11, -7, -5, -5, -7, -7, -10, -9, -10, -7, -2, -8, -5, -3, -5, -6, -1, -3, -6, -1, 2, 9, 3, 10, 8, 3, 2, 7, 0, 2, -1, -3, -3, 0, -6, -2, -5, 0, -6, 0, -5, 0, -5, 1, -7, -2, 0, 0, -4, -3, 2, 2, 2, 10, 10, 17, 8, 13, 8, 6, 9, 4, 1, 4, 2, 6, 2, 1, 10, 4, 1, 7, 5, 2, 10, 9, 8, 1, 10, 6, 9, 5, 12, 10, 10, 12, 9, 22, 20, 16, 14, 19, 17, 16, 15, 21, 22, 21, 15, 20, 18, 14, 23, 22, 15, 16, 17, 19, 18, 25, 20, 16, 15, 16, 20, 15, 19, 22, 20, 18, 20, 20, 15, 16, 18, 19, 17, 15, 12, 14, 13, 8, 8, 11, 8, 10, 13, 14, 15, 10, 13, 15, 17, 14, 13, 19, 17, 16, 15, 18, 12, 15, 17, 18, 15, 19, 17, 14, 11, 9, 7, 0, 7, 2, 8, 3, 8, 6, 8, 9, 6, 5, 10, 12, 12, 8, 16, 12, 17, 19, 11, 15, 10, 14, 18, 18, 12, 16, 10, 15, 14, 6, 1, 1, 0, 1, 4, 0, -1, 0, 2, 4, -1, 3, 5, 6, 11, 15, 12, 10, 8, 16, 10, 15, 15, 14, 16, 9, 9, 14, 16, 8, 7, 4, 5, -2, 1, -3, 1, -1, 1, -2, 3, 0, 4, 1, 0, 7, 3, 8, 15, 8, 11, 15, 9, 15, 12, 14, 13, 11, 6, 12, 12, 7, 8, 5, 8, 0, -2, -6, -4, -5, 0, -1, -4, -6, -2, -4, 5, 2, 1, 11, 11, 7, 8, 7, 14, 12, 6, 8, 9, 6, 10, 8, 13, 12, 5, 4, 6, -2, 0, -2, -4, -8, -1, -7, -5, -5, 0, 0, -1, 6, 2, 8, 6, 4, 12, 4, 4, 10, 5, 6, 10, 6, 8, 9, 5, 6, 8, 0, 6, -2, 0, -5, -8, -3, -4, 0, -7, -3, -6, 4, -1, 6, 5, 5, 6, 10, 3, 6, 7, 5, 4, 2, 1, 5, 3, 11, 11, 5, 8, 7, 0, 1, 1, 0, 0, 2, 1, 4, -1, -2, -3, -4, 2, 2, 2, 9, 8, 9, 3, 7, 8, 6, 6, 9, 0, 7, 2, 0, 1, 3, 3, 1, 4, -1, -2, 1, 1, 0, 0, -1, -1, -5, 0, -3, 2, 5, 1, 7, 6, 4, 0, 0, 3, 0, 4, 1, 5, 6, 8, 7, 3, 4, 0, 4, -1, 0, 3, 3, 0, -1, 4, -2, 0, -5, 0, -2, 6, 0, 1, 2, 6, 3, 4, 3, 5, 4, 1, 0, 5, 0, 4, 1, 2, 5, -3, 4, 3, -5, 1, -1, -1, 0, 4, 1, 1, -1, 2, 0, -2, 0, 0, -3, 1, -2, -1, 0, 2, -3, -3, -5, -4, 4, 2, 0, 0, -1, -2, 2, -1, -3, -2, -2, 4, -3, 0, 4, 1, -1, -4, -5, 0, -4, 1, 2, 3, -2, 2, 0, -3, -2, -4, -7, -4, 1, 1, -1, -3, 2, 0, -5, -5, -4, -3, -3, -1, 4, 2, 0, 0, 1, -1, 3, -4, 2, 0, 0, 0, 0, 2, -5, -5, -7, -9, -7, -8, -5, -5, 3, -3, 2, 0, 1, 0, 0, -4, 1, -2, 1, 6, 4, 0, 1, -3, 0, 0, 0, -3, -3, 0, 0, 0, -1, -5, -2, -12, -10, -7, -9, -7, -4, -5, -3, -6, 2, 0, -2, -2, 0, 5, 4, 2, 10, 3, 7, 5, 0, 0, 0, -1, -2, 0, 2, -1, -5, -2, -9, -12, -12, -7, -4, -5, -7, 1, 0, -2, -1, -1, 5, 3, 7, 9, 8, 11, 4, 9, 4, 3, 3, 6, 7, 4, -1, -3, -2, -4, -1, -3, -6, -14, -14, -8, -3, -3, 0, 0, 1, -2, -1, 3, 1, 7, 3, 12, 8, 13, 9, 11, 3, 7, 6, 5, 7, 0, -1, -2, -3, 0, -3, -10, -8, -16, -9, -9, -11, -3, -4, 2, -5, 3, 1, -2, 3, 1, 2, 13, 5, 14, 15, 8, 2, 6, 5, 0, 5, 3, 0, 0, 0, -7, -9, -9, -13, -15, -13, -13, -6, -6, -3, 0, 0, -2, -2, 1, 3, 1, -1, 3, 4, 8, 7, 7, 6, 3, 7, 6, 4, -6, 0, -2, -7, -8, -4, -4, -8, -12, -10, -11, -7, -8, -4, -3, 0, -7, -1, -4, 2, -3, -1, 2, 3, 0, 4, 0, 0, -2, -1, -1, 0, -7, -3, -8, -5, -10, -8, -7, -8, -9, -7, -10, -7, -11, -5, -7, -9, -8, -6, -6, -3, -6, -2, -1, 4, -1, -1, -2, 2, -2, 1, -3, -2, -6, -4, -6, -10, -15, -7, -4, -7, -9, -6, -6, -11, -5, -10, -9, -5, -6, -6, -1, -5, -6, -6, 1, -3, 0, -1, -5, 0, 0, -5, 0, -5, -2, -11, -2, -6, -10, -5, -8, -7, -5, -3, -10, -11, -10, -10, -9, -8, -9, -3, -2, -6, -7, -3, -1, 2, 0, 4, 2, -2, -5, -6, -2, 0, -1, -6, -7, -8, -6, -8, -7, -5, -2, -5, 0, -6, -3, -4, -9, -8, -3, -8, -8, -7, -6, 2, -5, -4, 0, 1, 1, 2, -1, -2, -2, -2, -6, -5, -9, -7, -1, -8, -5, -5, -1, 4, 3, 0, -3, -5, -1, -6, -5, -6, -10, 0, -2, -1, -6, -5, 1, -3, -4, -4, -5, -6, -2, -7, -2, -2, -5, -8, -3, -6, -5, -3, -2, 8, 5, -2, -2, -5, -3, -10, -10, -7, -10, -5, -1, -5, 0, -2, 2, 1, 1, 2, -5, 0, -3, -5, -4, -3, -4, -7, -5, -6, -3, 5, 1, 4, 1, 3, 4, 2, 0, -6, -6, -5, 0, -3, -7, 0, -6, 0, 3, -1, 2, -5, -4, -9, -7, -3, -8, -4, -8, -10, -4, -1, 2, 1, 6, 11, 3, 1, -1, 0, 2, -2, -2, -4, -6, -3, -5, -2, -2, -1, 0, 2, 0, -5, -7, -5, -5, -4, -6, -2, -4, -1, -7, -4, 4, 3, 7, 9, 7, 2, 0, -1, -3, -2, 0, 0, 0, 1, -5, -5, 0, -1, 2, 1, -1, 1, -4, -3, -2, 0, -4, -5, 0, -2, -2, 2, 4, 10, 7, 13, 6, 11, 7, 4, 1, 2, 2, 3, 2, 3, -1, 4, -1, 2, 0, 0, 2, 0, 3, 4, -2, 0, 0, 4, 2, 5, 4, 2, 6, 3, 12, 12, 8, 12, 14, 13, 9, 12, 6, 7, 10, 9, 4, 9, 9, 11, 9, 12, 9, 11, 8, 9, 7, 5, 4, 8, 10, 11, 13, 7, 13, 9, 15,

    -- ifmap
    -- channel=0
    158, 159, 165, 166, 160, 156, 162, 159, 158, 159, 161, 160, 161, 166, 169, 170, 167, 162, 160, 160, 156, 149, 150, 148, 149, 143, 140, 141, 143, 137, 126, 116, 
    152, 151, 159, 166, 162, 160, 164, 162, 163, 156, 155, 159, 163, 170, 171, 171, 169, 160, 154, 151, 145, 139, 140, 141, 149, 147, 145, 142, 143, 136, 125, 119, 
    151, 151, 158, 167, 160, 163, 165, 165, 163, 162, 158, 157, 161, 166, 167, 169, 170, 159, 145, 121, 110, 98, 101, 114, 120, 134, 143, 140, 142, 139, 130, 120, 
    155, 155, 160, 174, 167, 167, 169, 169, 165, 165, 167, 191, 177, 157, 162, 164, 158, 149, 104, 103, 98, 92, 80, 74, 86, 83, 113, 132, 140, 140, 136, 127, 
    155, 156, 161, 170, 169, 163, 169, 166, 164, 164, 173, 246, 195, 151, 146, 142, 111, 78, 85, 113, 112, 106, 97, 93, 74, 84, 85, 105, 128, 138, 133, 129, 
    148, 133, 130, 147, 161, 165, 167, 167, 163, 165, 163, 180, 157, 128, 97, 66, 69, 66, 89, 118, 122, 119, 114, 94, 99, 91, 58, 67, 108, 140, 138, 134, 
    127, 109, 47, 88, 153, 170, 168, 170, 169, 166, 164, 147, 129, 127, 100, 68, 78, 72, 83, 132, 146, 124, 105, 107, 115, 85, 63, 46, 79, 132, 141, 134, 
    131, 99, 42, 70, 143, 167, 165, 168, 171, 161, 140, 120, 130, 144, 116, 88, 91, 85, 77, 124, 163, 136, 102, 106, 100, 85, 54, 49, 57, 107, 138, 136, 
    170, 103, 54, 124, 153, 161, 163, 166, 165, 174, 113, 125, 157, 156, 121, 86, 82, 84, 80, 81, 138, 146, 113, 87, 83, 86, 71, 56, 40, 74, 133, 137, 
    180, 134, 94, 154, 174, 158, 156, 153, 207, 237, 207, 156, 174, 148, 125, 93, 86, 74, 59, 76, 137, 143, 133, 106, 86, 87, 84, 75, 50, 40, 95, 132, 
    183, 108, 142, 165, 177, 155, 159, 122, 213, 237, 220, 164, 183, 156, 125, 120, 78, 80, 45, 91, 175, 157, 155, 107, 87, 103, 88, 78, 59, 41, 59, 104, 
    188, 100, 135, 170, 187, 166, 173, 134, 117, 194, 199, 170, 185, 189, 134, 117, 102, 84, 38, 125, 210, 160, 146, 93, 83, 94, 104, 85, 73, 55, 62, 76, 
    189, 90, 127, 175, 174, 166, 178, 159, 97, 168, 168, 137, 186, 216, 160, 123, 120, 115, 50, 150, 194, 155, 123, 91, 84, 84, 95, 86, 84, 73, 79, 73, 
    189, 93, 152, 185, 119, 136, 173, 167, 103, 147, 145, 167, 189, 226, 180, 141, 126, 117, 71, 154, 186, 149, 114, 87, 80, 72, 80, 99, 100, 90, 97, 94, 
    194, 108, 168, 186, 105, 99, 156, 167, 100, 115, 138, 198, 190, 172, 145, 154, 146, 103, 71, 152, 179, 137, 130, 110, 85, 91, 95, 109, 115, 100, 97, 117, 
    197, 132, 172, 184, 130, 78, 140, 155, 115, 130, 143, 230, 242, 145, 135, 131, 121, 108, 95, 144, 168, 152, 112, 87, 71, 87, 105, 112, 120, 103, 121, 136, 
    203, 146, 168, 191, 168, 78, 126, 138, 138, 96, 154, 173, 162, 140, 113, 113, 101, 105, 112, 171, 156, 148, 135, 109, 78, 79, 94, 101, 107, 125, 151, 144, 
    214, 163, 164, 183, 176, 94, 96, 156, 148, 106, 129, 118, 114, 116, 102, 115, 86, 101, 144, 118, 68, 128, 133, 75, 60, 58, 71, 102, 116, 143, 150, 140, 
    212, 178, 167, 173, 176, 124, 86, 141, 153, 135, 104, 77, 134, 124, 129, 147, 85, 92, 150, 132, 117, 107, 75, 64, 44, 65, 86, 133, 155, 160, 154, 151, 
    199, 187, 171, 174, 177, 144, 86, 119, 122, 137, 144, 70, 129, 108, 145, 184, 116, 73, 131, 137, 134, 89, 51, 52, 47, 90, 121, 163, 171, 164, 158, 149, 
    165, 195, 179, 177, 181, 152, 99, 131, 171, 103, 93, 80, 93, 122, 178, 191, 150, 100, 89, 87, 60, 46, 38, 24, 46, 60, 108, 144, 144, 128, 127, 120, 
    117, 195, 177, 178, 181, 138, 83, 150, 245, 219, 133, 134, 149, 176, 190, 194, 168, 125, 110, 61, 35, 34, 49, 58, 61, 58, 69, 72, 78, 69, 59, 55, 
    79, 175, 174, 176, 177, 140, 109, 211, 253, 252, 208, 124, 114, 124, 116, 122, 104, 68, 68, 60, 52, 50, 51, 56, 56, 51, 43, 51, 59, 48, 43, 42, 
    41, 96, 144, 168, 178, 165, 165, 246, 253, 227, 110, 60, 53, 49, 49, 48, 45, 42, 46, 42, 38, 46, 46, 43, 42, 46, 46, 50, 55, 53, 51, 45, 
    29, 29, 59, 131, 166, 132, 194, 254, 241, 141, 61, 50, 50, 51, 49, 50, 47, 42, 39, 34, 35, 39, 38, 42, 45, 56, 62, 59, 56, 50, 46, 51, 
    48, 30, 34, 73, 128, 128, 215, 256, 187, 66, 54, 50, 52, 52, 46, 45, 43, 41, 36, 39, 40, 40, 43, 46, 59, 62, 64, 59, 54, 50, 70, 83, 
    52, 35, 31, 41, 66, 128, 224, 240, 124, 58, 49, 56, 54, 44, 44, 47, 46, 43, 43, 44, 44, 45, 54, 58, 54, 46, 43, 36, 51, 73, 85, 76, 
    50, 35, 29, 35, 44, 78, 202, 211, 97, 65, 54, 48, 58, 48, 40, 45, 47, 48, 47, 46, 51, 39, 39, 48, 47, 39, 28, 40, 67, 67, 46, 51, 
    50, 35, 32, 33, 41, 46, 104, 170, 64, 54, 52, 53, 61, 58, 54, 45, 42, 41, 46, 49, 46, 42, 40, 39, 37, 40, 44, 63, 47, 31, 15, 51, 
    68, 42, 31, 38, 37, 43, 42, 71, 49, 31, 27, 38, 49, 56, 58, 53, 56, 60, 57, 53, 50, 45, 39, 33, 42, 62, 79, 73, 56, 38, 13, 40, 
    61, 49, 35, 43, 39, 42, 44, 40, 42, 27, 23, 30, 27, 29, 36, 47, 56, 62, 66, 75, 69, 49, 43, 43, 60, 85, 109, 93, 60, 26, 29, 20, 
    54, 56, 45, 43, 40, 40, 40, 38, 36, 26, 22, 29, 25, 29, 19, 18, 32, 47, 61, 74, 66, 53, 52, 45, 67, 89, 105, 89, 48, 24, 34, 21, 
    
    -- channel=1
    112, 111, 116, 118, 112, 109, 115, 113, 111, 113, 116, 111, 111, 117, 117, 119, 117, 113, 111, 112, 109, 107, 107, 106, 107, 101, 98, 97, 97, 95, 91, 85, 
    112, 110, 114, 116, 112, 113, 117, 114, 116, 110, 111, 110, 113, 119, 117, 115, 115, 111, 112, 115, 110, 104, 102, 100, 105, 102, 102, 97, 98, 95, 91, 88, 
    110, 109, 111, 111, 106, 115, 117, 117, 115, 115, 114, 109, 111, 115, 114, 113, 116, 114, 111, 96, 90, 78, 77, 85, 86, 96, 103, 99, 99, 98, 95, 89, 
    107, 110, 109, 112, 110, 117, 120, 119, 115, 117, 123, 146, 130, 111, 115, 114, 112, 111, 80, 87, 90, 90, 75, 63, 70, 62, 85, 98, 102, 101, 99, 94, 
    107, 114, 115, 114, 114, 113, 120, 116, 113, 116, 128, 214, 156, 114, 111, 108, 80, 53, 69, 103, 110, 114, 102, 94, 72, 78, 73, 83, 96, 101, 94, 93, 
    109, 104, 100, 112, 115, 113, 116, 115, 111, 116, 118, 138, 122, 102, 75, 50, 58, 56, 83, 113, 121, 122, 116, 96, 100, 91, 58, 58, 84, 105, 98, 95, 
    100, 95, 37, 74, 117, 118, 115, 118, 117, 116, 120, 107, 98, 108, 87, 67, 83, 75, 84, 130, 142, 118, 99, 102, 111, 83, 71, 47, 61, 98, 99, 93, 
    115, 96, 43, 64, 111, 117, 114, 116, 119, 113, 109, 94, 110, 131, 106, 87, 95, 88, 77, 118, 153, 124, 93, 98, 93, 81, 60, 53, 47, 83, 103, 97, 
    161, 105, 58, 121, 124, 113, 117, 122, 121, 135, 89, 105, 141, 143, 111, 80, 81, 85, 78, 71, 125, 135, 103, 79, 77, 82, 73, 57, 35, 59, 106, 103, 
    176, 139, 100, 154, 149, 116, 116, 118, 180, 214, 180, 131, 153, 131, 110, 85, 84, 74, 57, 68, 125, 133, 124, 98, 81, 85, 85, 76, 49, 30, 75, 103, 
    183, 116, 151, 169, 156, 112, 118, 89, 197, 224, 191, 135, 159, 137, 108, 111, 76, 80, 44, 85, 165, 147, 147, 100, 83, 102, 88, 79, 59, 36, 46, 81, 
    191, 108, 144, 175, 167, 120, 123, 93, 95, 182, 171, 142, 161, 171, 119, 107, 98, 84, 38, 121, 201, 152, 139, 89, 80, 93, 104, 87, 75, 53, 55, 56, 
    194, 96, 134, 180, 156, 123, 123, 109, 68, 154, 144, 114, 166, 202, 149, 113, 114, 114, 50, 147, 187, 149, 118, 88, 83, 84, 95, 87, 87, 73, 74, 55, 
    192, 95, 154, 188, 110, 106, 124, 116, 72, 132, 125, 149, 174, 216, 172, 131, 117, 114, 71, 152, 181, 144, 110, 85, 80, 73, 80, 100, 101, 88, 89, 73, 
    196, 107, 167, 186, 109, 89, 119, 122, 74, 106, 123, 185, 180, 165, 140, 143, 136, 100, 71, 152, 175, 133, 128, 109, 86, 93, 96, 110, 116, 96, 85, 95, 
    197, 129, 167, 178, 137, 83, 120, 125, 94, 120, 131, 221, 236, 138, 130, 121, 112, 104, 88, 134, 159, 147, 108, 85, 72, 88, 104, 109, 110, 86, 96, 104, 
    203, 146, 164, 182, 170, 86, 125, 126, 121, 80, 143, 163, 152, 132, 106, 106, 101, 101, 90, 143, 138, 141, 130, 105, 76, 79, 93, 91, 83, 88, 108, 104, 
    215, 166, 167, 184, 182, 102, 96, 149, 137, 93, 116, 105, 102, 105, 91, 110, 91, 103, 128, 96, 56, 120, 126, 69, 56, 56, 70, 93, 94, 112, 116, 110, 
    211, 184, 175, 181, 184, 131, 88, 139, 148, 128, 90, 64, 121, 111, 117, 143, 92, 96, 139, 117, 109, 99, 68, 59, 41, 62, 69, 105, 119, 120, 115, 111, 
    192, 189, 176, 179, 182, 149, 90, 121, 124, 136, 134, 59, 118, 97, 134, 176, 118, 75, 119, 124, 129, 86, 49, 51, 49, 90, 91, 118, 121, 113, 111, 107, 
    156, 193, 178, 173, 181, 157, 103, 135, 175, 105, 90, 77, 90, 118, 173, 182, 148, 100, 78, 77, 61, 52, 46, 33, 57, 71, 100, 125, 123, 109, 113, 105, 
    120, 200, 178, 169, 179, 144, 87, 153, 247, 222, 140, 141, 156, 182, 196, 192, 172, 133, 109, 62, 49, 54, 70, 81, 85, 84, 99, 101, 104, 96, 92, 90, 
    105, 197, 183, 172, 177, 146, 112, 211, 252, 253, 224, 143, 132, 141, 133, 133, 124, 93, 87, 82, 84, 84, 85, 93, 94, 91, 96, 104, 108, 97, 97, 95, 
    89, 137, 168, 174, 182, 170, 166, 245, 251, 231, 136, 88, 80, 76, 75, 72, 79, 81, 81, 82, 86, 90, 89, 87, 89, 93, 94, 96, 96, 94, 95, 90, 
    91, 87, 102, 153, 179, 136, 189, 250, 245, 159, 94, 84, 84, 85, 83, 84, 86, 84, 82, 79, 83, 86, 85, 89, 92, 103, 103, 101, 102, 99, 94, 103, 
    111, 94, 85, 106, 148, 136, 213, 253, 198, 93, 91, 88, 90, 90, 83, 82, 82, 81, 80, 83, 86, 89, 92, 95, 108, 110, 109, 108, 108, 105, 123, 137, 
    114, 99, 86, 83, 95, 145, 229, 245, 143, 92, 87, 94, 92, 82, 82, 83, 84, 83, 86, 88, 90, 97, 106, 110, 105, 97, 95, 91, 108, 130, 138, 125, 
    110, 98, 89, 86, 83, 106, 219, 228, 126, 104, 94, 87, 97, 87, 80, 82, 84, 87, 89, 89, 97, 92, 93, 102, 101, 93, 85, 101, 129, 126, 98, 96, 
    108, 97, 92, 88, 88, 84, 133, 197, 100, 97, 94, 95, 103, 100, 96, 83, 79, 80, 88, 92, 92, 95, 93, 92, 90, 93, 102, 125, 110, 90, 60, 93, 
    124, 100, 88, 91, 87, 89, 79, 107, 89, 77, 71, 82, 93, 100, 102, 92, 94, 99, 99, 97, 95, 94, 88, 83, 91, 112, 132, 131, 116, 97, 64, 85, 
    116, 102, 85, 91, 90, 92, 88, 81, 85, 72, 67, 74, 71, 73, 80, 86, 95, 101, 109, 119, 113, 95, 88, 88, 105, 130, 156, 145, 115, 82, 82, 64, 
    107, 105, 89, 86, 89, 92, 87, 81, 79, 69, 66, 73, 69, 73, 63, 58, 70, 87, 104, 119, 111, 96, 95, 87, 109, 131, 146, 135, 99, 77, 84, 67, 
    
    -- channel=2
    49, 47, 51, 53, 46, 41, 47, 45, 44, 41, 41, 52, 49, 41, 45, 44, 40, 38, 39, 43, 44, 45, 45, 43, 44, 39, 43, 41, 38, 36, 36, 33, 
    51, 40, 45, 56, 49, 43, 47, 45, 46, 38, 41, 54, 52, 41, 40, 33, 30, 33, 41, 50, 53, 55, 52, 48, 50, 46, 45, 38, 34, 31, 32, 34, 
    47, 33, 36, 48, 42, 44, 45, 45, 43, 43, 48, 57, 51, 38, 37, 35, 39, 47, 54, 49, 52, 50, 47, 50, 48, 55, 51, 39, 35, 34, 34, 33, 
    40, 32, 31, 44, 43, 46, 48, 48, 44, 45, 57, 95, 75, 41, 47, 54, 58, 67, 47, 65, 76, 84, 66, 50, 52, 39, 45, 46, 43, 39, 39, 36, 
    41, 48, 49, 47, 43, 40, 47, 44, 41, 42, 59, 164, 107, 56, 60, 71, 50, 31, 56, 98, 111, 118, 105, 93, 67, 70, 47, 45, 48, 46, 36, 36, 
    54, 64, 57, 53, 44, 39, 41, 41, 37, 39, 42, 85, 78, 58, 43, 31, 43, 45, 76, 110, 120, 122, 116, 96, 97, 86, 47, 37, 49, 58, 44, 40, 
    57, 80, 17, 28, 48, 43, 40, 43, 42, 37, 39, 52, 59, 75, 70, 57, 72, 64, 74, 121, 132, 108, 90, 94, 103, 77, 69, 39, 36, 58, 48, 39, 
    90, 92, 38, 41, 56, 42, 36, 39, 49, 51, 51, 49, 77, 107, 93, 79, 88, 82, 69, 107, 140, 112, 81, 88, 84, 74, 58, 49, 32, 50, 51, 39, 
    144, 105, 59, 113, 82, 43, 41, 50, 66, 95, 59, 78, 121, 128, 101, 74, 77, 82, 73, 61, 112, 123, 93, 70, 69, 76, 67, 53, 27, 35, 59, 45, 
    163, 143, 105, 149, 112, 51, 47, 60, 146, 198, 166, 119, 145, 125, 107, 79, 79, 71, 53, 58, 112, 122, 114, 89, 74, 78, 78, 71, 43, 15, 44, 57, 
    175, 122, 158, 168, 122, 50, 51, 47, 179, 226, 188, 131, 155, 132, 104, 104, 69, 77, 40, 77, 154, 137, 138, 92, 77, 96, 79, 73, 59, 33, 31, 46, 
    189, 116, 153, 178, 136, 59, 55, 44, 80, 188, 164, 133, 151, 159, 106, 95, 89, 79, 34, 113, 192, 142, 130, 82, 75, 88, 94, 81, 78, 55, 48, 26, 
    194, 105, 144, 185, 133, 68, 53, 47, 44, 152, 126, 94, 148, 183, 129, 98, 105, 109, 47, 140, 178, 140, 111, 83, 79, 80, 85, 81, 89, 73, 64, 24, 
    193, 103, 163, 192, 98, 66, 58, 50, 39, 120, 103, 127, 155, 200, 157, 117, 107, 109, 68, 147, 174, 136, 104, 80, 76, 70, 72, 94, 99, 81, 69, 34, 
    196, 112, 172, 188, 109, 67, 62, 55, 34, 88, 103, 169, 169, 159, 140, 134, 125, 95, 70, 149, 170, 127, 122, 105, 83, 91, 90, 104, 111, 80, 53, 47, 
    197, 136, 174, 181, 142, 77, 88, 77, 52, 93, 116, 211, 230, 137, 130, 112, 101, 95, 75, 118, 146, 138, 101, 80, 68, 87, 99, 99, 93, 54, 48, 48, 
    204, 160, 178, 188, 172, 90, 126, 113, 82, 37, 133, 155, 141, 117, 88, 90, 92, 87, 58, 104, 109, 126, 118, 97, 72, 77, 94, 82, 55, 45, 55, 46, 
    215, 180, 184, 194, 186, 105, 102, 145, 111, 61, 105, 95, 89, 89, 73, 98, 88, 95, 102, 64, 32, 105, 115, 61, 51, 53, 65, 78, 64, 68, 64, 54, 
    205, 192, 189, 193, 188, 133, 96, 143, 141, 111, 80, 55, 108, 96, 100, 133, 93, 93, 120, 93, 92, 86, 58, 52, 39, 60, 40, 59, 62, 54, 45, 46, 
    180, 187, 181, 185, 184, 152, 99, 132, 130, 135, 126, 51, 108, 86, 123, 168, 118, 73, 103, 105, 118, 78, 44, 50, 52, 93, 60, 68, 64, 52, 50, 46, 
    146, 187, 175, 172, 180, 160, 111, 146, 185, 111, 87, 73, 86, 116, 173, 177, 148, 101, 66, 63, 57, 54, 51, 41, 69, 83, 75, 82, 76, 61, 69, 63, 
    124, 200, 176, 168, 179, 147, 91, 159, 250, 225, 144, 147, 164, 192, 208, 197, 181, 143, 109, 62, 58, 68, 87, 102, 110, 111, 122, 119, 120, 112, 112, 115, 
    133, 213, 192, 177, 182, 150, 113, 209, 247, 252, 232, 157, 149, 162, 156, 152, 148, 119, 104, 101, 111, 110, 115, 125, 131, 130, 135, 141, 142, 132, 137, 132, 
    135, 168, 188, 188, 192, 174, 164, 237, 241, 228, 153, 111, 105, 105, 107, 101, 115, 120, 113, 116, 125, 125, 126, 128, 132, 139, 137, 137, 135, 134, 139, 133, 
    141, 130, 134, 176, 191, 137, 181, 242, 245, 175, 127, 118, 119, 121, 120, 116, 117, 117, 115, 113, 120, 125, 125, 130, 134, 145, 142, 142, 146, 144, 140, 149, 
    162, 140, 124, 136, 167, 143, 209, 249, 205, 118, 128, 125, 127, 127, 121, 115, 113, 112, 113, 117, 123, 131, 134, 138, 150, 152, 147, 149, 154, 152, 167, 182, 
    165, 147, 130, 122, 126, 164, 234, 247, 153, 114, 123, 131, 129, 119, 119, 119, 119, 119, 123, 127, 131, 141, 150, 154, 150, 141, 140, 138, 158, 178, 182, 169, 
    162, 149, 138, 133, 126, 138, 233, 234, 140, 126, 129, 124, 133, 123, 116, 119, 122, 126, 130, 132, 140, 138, 139, 148, 147, 139, 133, 153, 182, 176, 142, 139, 
    161, 147, 143, 141, 138, 125, 159, 211, 119, 121, 128, 130, 139, 135, 131, 120, 118, 120, 130, 135, 136, 139, 138, 136, 135, 138, 151, 178, 164, 140, 103, 136, 
    177, 148, 137, 146, 139, 132, 113, 133, 114, 105, 105, 117, 128, 135, 137, 128, 131, 137, 139, 138, 137, 136, 131, 125, 133, 154, 179, 181, 168, 146, 108, 127, 
    168, 148, 132, 143, 139, 134, 125, 112, 115, 104, 102, 109, 106, 108, 115, 120, 128, 135, 144, 156, 152, 134, 127, 127, 144, 170, 197, 190, 164, 130, 126, 107, 
    160, 149, 132, 134, 134, 132, 123, 115, 114, 105, 101, 108, 104, 108, 98, 89, 100, 118, 137, 152, 145, 131, 130, 123, 145, 167, 182, 175, 145, 124, 129, 110, 
    
    
    others => 0);
end inmem_package;
