library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 18, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 10, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 6, 0, 16, 0, 0, 13, 14, 0, 0, 0, 0, 0, 0, 0, 
    24, 17, 3, 30, 19, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 
    2, 13, 10, 28, 0, 0, 0, 0, 0, 0, 1, 3, 6, 7, 8, 
    5, 0, 19, 22, 0, 0, 0, 0, 0, 0, 3, 7, 3, 11, 13, 
    3, 4, 0, 7, 0, 0, 3, 0, 0, 0, 0, 0, 9, 13, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 5, 0, 0, 0, 9, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 15, 0, 0, 4, 0, 15, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 0, 0, 46, 31, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 14, 2, 0, 0, 0, 1, 6, 0, 
    0, 0, 0, 11, 37, 54, 14, 0, 0, 0, 8, 23, 8, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 4, 0, 0, 2, 26, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 0, 0, 8, 0, 0, 
    23, 25, 0, 0, 2, 0, 19, 3, 0, 0, 0, 0, 0, 0, 0, 
    13, 33, 0, 0, 45, 29, 0, 0, 0, 0, 11, 11, 1, 8, 0, 
    0, 0, 0, 0, 0, 0, 4, 4, 14, 12, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 3, 0, 5, 1, 
    3, 0, 20, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 11, 0, 0, 8, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 23, 1, 0, 0, 0, 8, 2, 0, 
    0, 0, 0, 16, 59, 53, 0, 0, 0, 11, 29, 36, 22, 8, 13, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 10, 0, 0, 10, 
    0, 4, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 0, 0, 15, 11, 0, 
    
    -- channel=6
    49, 50, 49, 49, 50, 45, 54, 61, 52, 40, 34, 36, 37, 43, 43, 
    48, 53, 52, 52, 48, 13, 43, 42, 42, 0, 0, 0, 15, 31, 38, 
    30, 42, 53, 55, 56, 56, 29, 15, 0, 0, 0, 0, 0, 8, 27, 
    0, 0, 48, 51, 38, 17, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 38, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 33, 48, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 41, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 20, 1, 3, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    5, 2, 7, 2, 2, 6, 4, 2, 2, 0, 0, 6, 3, 0, 0, 
    6, 5, 9, 0, 10, 14, 0, 0, 0, 8, 0, 0, 9, 10, 0, 
    0, 24, 6, 1, 10, 6, 0, 0, 9, 37, 0, 0, 0, 15, 12, 
    0, 61, 0, 10, 0, 13, 0, 0, 0, 54, 0, 0, 0, 0, 45, 
    0, 28, 0, 54, 0, 0, 0, 0, 0, 72, 0, 0, 0, 0, 29, 
    0, 7, 0, 18, 43, 0, 0, 0, 0, 130, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 49, 42, 0, 0, 0, 101, 0, 0, 4, 9, 0, 
    0, 0, 0, 0, 37, 50, 0, 0, 0, 65, 0, 0, 17, 2, 0, 
    0, 0, 0, 19, 0, 3, 0, 0, 19, 0, 11, 0, 16, 14, 14, 
    0, 1, 0, 42, 0, 10, 26, 0, 0, 0, 0, 0, 27, 29, 0, 
    37, 0, 0, 112, 0, 0, 39, 0, 0, 0, 0, 9, 12, 6, 0, 
    44, 21, 0, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 46, 63, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 3, 
    0, 0, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    0, 0, 6, 0, 0, 7, 0, 0, 2, 0, 0, 0, 24, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 2, 0, 0, 0, 37, 9, 0, 0, 0, 17, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 8, 8, 6, 0, 0, 
    19, 23, 0, 0, 0, 0, 25, 10, 0, 0, 0, 0, 0, 0, 0, 
    26, 50, 5, 10, 74, 42, 3, 4, 0, 0, 21, 16, 7, 13, 0, 
    0, 3, 4, 0, 0, 0, 19, 15, 15, 29, 0, 0, 0, 7, 21, 
    10, 0, 0, 0, 0, 13, 0, 6, 6, 4, 0, 5, 0, 12, 15, 
    12, 10, 19, 10, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 1, 2, 4, 6, 0, 0, 7, 11, 0, 0, 0, 0, 1, 15, 
    0, 0, 6, 2, 10, 0, 2, 37, 5, 0, 0, 0, 19, 15, 0, 
    0, 0, 0, 44, 82, 69, 12, 0, 0, 0, 21, 33, 12, 0, 0, 
    0, 0, 16, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 13, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 5, 1, 0, 2, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 2, 0, 26, 19, 2, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    9, 8, 11, 6, 6, 12, 9, 8, 5, 2, 4, 15, 12, 3, 0, 
    12, 12, 13, 4, 16, 28, 0, 2, 0, 24, 0, 0, 17, 22, 4, 
    0, 45, 10, 7, 12, 19, 0, 0, 11, 50, 0, 0, 0, 18, 28, 
    0, 71, 7, 16, 0, 28, 0, 0, 0, 62, 0, 0, 0, 0, 62, 
    0, 41, 0, 66, 9, 0, 0, 0, 0, 83, 0, 0, 5, 0, 22, 
    0, 25, 0, 0, 69, 0, 0, 0, 0, 138, 0, 0, 16, 0, 0, 
    0, 0, 8, 0, 65, 48, 0, 0, 0, 115, 0, 0, 9, 18, 0, 
    0, 0, 0, 0, 40, 59, 0, 0, 0, 69, 0, 0, 23, 5, 0, 
    0, 13, 0, 41, 0, 14, 0, 0, 35, 0, 14, 0, 20, 27, 13, 
    0, 8, 0, 59, 0, 0, 42, 0, 0, 0, 0, 4, 42, 38, 0, 
    67, 5, 0, 128, 0, 0, 37, 0, 0, 0, 9, 14, 16, 22, 0, 
    57, 43, 0, 89, 0, 0, 5, 2, 0, 1, 3, 6, 5, 3, 0, 
    0, 50, 78, 0, 0, 0, 0, 0, 0, 3, 8, 6, 0, 4, 14, 
    0, 3, 93, 0, 0, 6, 0, 0, 4, 4, 0, 1, 0, 19, 0, 
    0, 1, 4, 2, 0, 10, 4, 0, 7, 0, 0, 5, 34, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 4, 0, 0, 0, 
    4, 10, 0, 0, 0, 0, 0, 0, 3, 0, 3, 1, 0, 0, 0, 
    4, 8, 0, 0, 0, 0, 11, 2, 0, 0, 0, 3, 0, 0, 0, 
    10, 8, 13, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    8, 7, 17, 0, 1, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 
    5, 2, 14, 0, 2, 0, 5, 20, 18, 8, 10, 13, 18, 9, 7, 
    36, 20, 3, 0, 29, 39, 33, 33, 34, 32, 37, 39, 41, 41, 43, 
    50, 33, 5, 13, 42, 36, 37, 36, 36, 37, 40, 42, 45, 45, 44, 
    56, 45, 22, 43, 34, 36, 37, 37, 38, 41, 46, 49, 49, 49, 58, 
    55, 51, 41, 40, 37, 40, 42, 39, 35, 39, 44, 43, 37, 51, 54, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    33, 37, 36, 37, 37, 33, 39, 43, 38, 27, 22, 23, 30, 34, 35, 
    36, 39, 38, 39, 36, 24, 41, 30, 29, 8, 7, 5, 6, 19, 30, 
    18, 17, 36, 41, 36, 20, 30, 15, 0, 0, 3, 6, 12, 0, 19, 
    30, 0, 36, 35, 33, 17, 13, 7, 0, 0, 18, 2, 10, 4, 0, 
    27, 0, 41, 15, 19, 18, 22, 13, 3, 0, 11, 18, 0, 12, 0, 
    5, 0, 43, 15, 0, 16, 22, 18, 17, 0, 15, 19, 0, 7, 8, 
    9, 2, 19, 45, 0, 0, 8, 15, 22, 0, 22, 10, 0, 0, 8, 
    2, 12, 10, 27, 1, 0, 19, 3, 14, 0, 14, 12, 0, 0, 23, 
    2, 0, 12, 0, 4, 4, 15, 1, 0, 18, 0, 16, 0, 9, 22, 
    0, 0, 22, 0, 10, 0, 0, 11, 0, 4, 14, 0, 0, 10, 30, 
    0, 0, 21, 0, 29, 0, 0, 0, 9, 3, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 11, 0, 0, 0, 34, 0, 0, 0, 19, 0, 0, 0, 20, 0, 
    0, 42, 0, 0, 0, 0, 0, 0, 0, 59, 0, 0, 0, 0, 44, 
    0, 7, 0, 7, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 37, 
    0, 0, 0, 6, 68, 0, 0, 0, 0, 104, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 68, 0, 0, 0, 0, 102, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 50, 0, 0, 0, 71, 0, 0, 13, 1, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 31, 0, 21, 0, 0, 
    0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 18, 7, 0, 
    32, 0, 0, 67, 0, 0, 24, 0, 0, 0, 0, 0, 9, 13, 0, 
    98, 5, 0, 56, 0, 0, 22, 16, 0, 0, 0, 5, 0, 1, 0, 
    0, 83, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 125, 0, 0, 0, 0, 0, 0, 0, 3, 8, 0, 15, 7, 
    0, 1, 14, 21, 0, 25, 9, 0, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 2, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 11, 0, 0, 13, 0, 7, 0, 0, 0, 17, 0, 9, 0, 
    0, 0, 14, 1, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 22, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 4, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 36, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 2, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 34, 15, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    3, 4, 1, 0, 3, 40, 4, 0, 0, 3, 17, 5, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 7, 18, 3, 8, 1, 0, 0, 
    13, 31, 0, 2, 0, 6, 21, 3, 0, 0, 0, 0, 0, 0, 0, 
    15, 38, 0, 15, 51, 27, 0, 2, 0, 15, 22, 7, 10, 8, 0, 
    0, 0, 0, 0, 0, 0, 15, 14, 13, 34, 0, 0, 0, 5, 18, 
    5, 0, 0, 0, 0, 16, 0, 1, 0, 12, 0, 5, 6, 14, 9, 
    3, 9, 10, 8, 6, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    1, 0, 0, 2, 1, 0, 0, 12, 10, 0, 0, 0, 0, 11, 14, 
    0, 0, 0, 16, 0, 0, 11, 29, 1, 0, 0, 0, 11, 7, 0, 
    0, 0, 0, 53, 56, 40, 0, 0, 0, 0, 22, 23, 4, 0, 0, 
    0, 0, 4, 23, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 11, 0, 0, 17, 
    0, 0, 0, 0, 0, 2, 6, 1, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 1, 3, 28, 14, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    20, 0, 0, 0, 31, 11, 7, 0, 0, 0, 6, 0, 0, 0, 0, 
    7, 7, 4, 0, 0, 16, 17, 2, 0, 0, 8, 0, 0, 0, 0, 
    17, 1, 0, 0, 0, 4, 15, 6, 0, 0, 10, 0, 0, 0, 0, 
    17, 21, 0, 0, 0, 9, 6, 0, 0, 0, 4, 0, 0, 0, 0, 
    22, 15, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 12, 14, 0, 9, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    2, 12, 9, 9, 46, 14, 2, 13, 9, 0, 0, 0, 0, 0, 0, 
    0, 7, 25, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 39, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 14, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 9, 21, 12, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 20, 19, 2, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 19, 2, 0, 0, 0, 0, 1, 0, 
    44, 23, 0, 0, 31, 45, 30, 29, 14, 8, 6, 8, 4, 2, 5, 
    3, 35, 7, 0, 34, 3, 5, 6, 3, 0, 0, 0, 7, 12, 0, 
    8, 6, 36, 35, 11, 2, 0, 2, 7, 4, 11, 17, 11, 0, 32, 
    7, 9, 15, 32, 16, 22, 22, 8, 0, 0, 2, 6, 0, 0, 3, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 16, 1, 1, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 23, 4, 0, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 3, 0, 0, 0, 0, 0, 2, 6, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 7, 
    0, 0, 0, 0, 0, 9, 21, 0, 0, 5, 0, 0, 8, 13, 0, 
    0, 0, 0, 12, 0, 0, 17, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 3, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 37, 24, 25, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 
    
    -- channel=20
    61, 65, 65, 66, 64, 63, 68, 72, 66, 48, 38, 43, 51, 58, 56, 
    64, 71, 68, 67, 65, 68, 67, 55, 30, 23, 19, 22, 25, 38, 52, 
    36, 32, 67, 70, 67, 43, 38, 23, 20, 12, 16, 12, 11, 15, 39, 
    25, 25, 63, 68, 59, 38, 34, 16, 6, 6, 23, 15, 9, 10, 22, 
    19, 25, 60, 50, 50, 44, 32, 22, 6, 13, 32, 25, 12, 10, 13, 
    14, 15, 62, 51, 15, 37, 40, 28, 16, 12, 25, 16, 7, 9, 15, 
    25, 13, 39, 58, 17, 36, 22, 25, 17, 3, 22, 19, 9, 12, 20, 
    28, 18, 25, 37, 26, 17, 15, 12, 19, 19, 21, 19, 6, 12, 35, 
    22, 12, 19, 13, 33, 10, 26, 20, 14, 28, 19, 5, 5, 29, 54, 
    16, 14, 17, 5, 22, 16, 19, 26, 20, 10, 0, 0, 7, 42, 51, 
    0, 19, 15, 18, 35, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    30, 29, 30, 31, 32, 28, 33, 34, 34, 29, 20, 20, 22, 26, 28, 
    32, 32, 33, 32, 33, 27, 30, 27, 17, 8, 6, 9, 10, 19, 27, 
    21, 17, 32, 32, 36, 30, 6, 5, 7, 9, 3, 0, 7, 12, 19, 
    6, 20, 32, 33, 28, 15, 16, 6, 4, 13, 0, 6, 0, 4, 19, 
    0, 19, 24, 29, 16, 13, 0, 0, 2, 4, 6, 4, 5, 3, 14, 
    0, 0, 14, 23, 0, 0, 0, 5, 4, 20, 0, 0, 6, 2, 2, 
    0, 1, 5, 23, 19, 5, 7, 0, 2, 20, 0, 0, 2, 5, 5, 
    0, 0, 3, 14, 23, 20, 0, 0, 0, 21, 0, 0, 4, 5, 6, 
    0, 0, 0, 1, 9, 0, 0, 8, 4, 14, 10, 0, 1, 10, 29, 
    0, 0, 0, 2, 1, 0, 0, 8, 5, 3, 0, 0, 9, 28, 25, 
    0, 0, 0, 8, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    24, 29, 29, 29, 26, 27, 30, 30, 25, 16, 11, 14, 22, 26, 24, 
    26, 32, 31, 29, 28, 40, 27, 21, 7, 2, 5, 2, 0, 10, 22, 
    10, 4, 27, 29, 27, 9, 5, 0, 3, 12, 12, 10, 8, 0, 16, 
    11, 8, 23, 27, 23, 8, 21, 11, 5, 2, 14, 5, 2, 1, 4, 
    10, 22, 25, 17, 46, 38, 19, 13, 3, 1, 15, 16, 9, 9, 0, 
    0, 7, 27, 23, 0, 14, 27, 15, 14, 14, 15, 2, 3, 8, 11, 
    5, 10, 1, 29, 9, 18, 14, 15, 11, 10, 5, 6, 1, 6, 13, 
    11, 12, 3, 14, 12, 20, 11, 1, 7, 16, 9, 2, 1, 9, 16, 
    12, 7, 6, 4, 14, 0, 0, 9, 2, 7, 0, 0, 0, 14, 30, 
    6, 7, 10, 1, 7, 9, 5, 23, 8, 3, 0, 0, 7, 24, 17, 
    0, 7, 3, 15, 39, 22, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 10, 0, 
    0, 2, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 14, 22, 0, 32, 0, 2, 0, 30, 0, 5, 0, 0, 27, 
    67, 0, 23, 38, 0, 32, 0, 0, 0, 2, 6, 11, 0, 0, 11, 
    85, 0, 12, 0, 0, 2, 0, 5, 0, 0, 0, 3, 0, 0, 4, 
    65, 0, 48, 0, 5, 0, 10, 0, 0, 0, 0, 0, 0, 0, 7, 
    20, 0, 47, 0, 44, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 57, 13, 0, 36, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 2, 2, 0, 0, 
    0, 0, 4, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 43, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 42, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    
    -- channel=24
    16, 15, 16, 18, 18, 14, 16, 18, 18, 14, 12, 12, 17, 17, 21, 
    19, 16, 15, 17, 17, 19, 17, 9, 13, 20, 22, 12, 7, 17, 20, 
    3, 15, 17, 19, 15, 0, 25, 20, 17, 6, 14, 22, 21, 7, 17, 
    36, 3, 19, 16, 13, 21, 20, 17, 17, 0, 25, 8, 27, 19, 5, 
    47, 4, 22, 8, 23, 0, 16, 19, 14, 3, 21, 23, 18, 30, 0, 
    14, 8, 27, 0, 0, 9, 28, 25, 29, 0, 12, 28, 12, 24, 24, 
    22, 8, 19, 29, 0, 3, 10, 24, 31, 0, 30, 24, 15, 18, 21, 
    11, 28, 12, 33, 5, 0, 13, 7, 31, 0, 25, 24, 9, 6, 26, 
    14, 5, 22, 15, 5, 6, 26, 16, 18, 12, 4, 22, 9, 21, 11, 
    13, 4, 37, 1, 19, 0, 14, 27, 0, 7, 23, 22, 12, 6, 18, 
    3, 5, 34, 0, 50, 14, 0, 4, 26, 25, 23, 17, 5, 8, 17, 
    0, 4, 30, 0, 7, 27, 7, 10, 21, 15, 15, 13, 17, 13, 17, 
    17, 0, 2, 0, 40, 16, 15, 15, 19, 18, 17, 14, 10, 14, 19, 
    24, 12, 0, 27, 28, 14, 21, 14, 14, 13, 12, 13, 20, 9, 4, 
    21, 15, 5, 19, 17, 9, 13, 18, 15, 17, 17, 18, 16, 15, 32, 
    
    -- channel=25
    0, 0, 6, 2, 1, 6, 0, 0, 3, 0, 0, 0, 1, 0, 0, 
    7, 5, 7, 0, 10, 41, 0, 0, 0, 19, 4, 0, 0, 4, 0, 
    0, 2, 3, 1, 5, 0, 0, 0, 20, 39, 0, 0, 0, 1, 9, 
    0, 67, 0, 11, 0, 22, 1, 0, 0, 30, 0, 0, 0, 0, 28, 
    0, 35, 0, 61, 23, 3, 0, 0, 0, 73, 0, 0, 4, 0, 11, 
    0, 1, 0, 0, 13, 0, 0, 0, 0, 130, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 25, 51, 0, 0, 0, 79, 0, 0, 6, 19, 0, 
    0, 0, 0, 0, 31, 28, 0, 0, 0, 40, 0, 0, 13, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 25, 0, 0, 0, 5, 19, 15, 
    0, 0, 0, 37, 0, 0, 33, 0, 0, 0, 0, 0, 30, 22, 0, 
    26, 0, 0, 129, 0, 7, 17, 0, 0, 0, 21, 27, 12, 0, 0, 
    0, 0, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 57, 0, 0, 0, 0, 0, 0, 1, 4, 6, 0, 0, 14, 
    0, 0, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 37, 0, 0, 
    
    -- channel=26
    2, 4, 2, 5, 4, 0, 3, 5, 2, 0, 0, 0, 2, 7, 9, 
    2, 0, 0, 5, 0, 0, 12, 0, 1, 0, 5, 1, 0, 0, 4, 
    2, 0, 1, 6, 0, 0, 30, 8, 0, 0, 13, 17, 20, 0, 0, 
    51, 0, 1, 0, 7, 0, 5, 12, 7, 0, 40, 0, 28, 17, 0, 
    53, 0, 25, 0, 0, 0, 32, 33, 17, 0, 8, 34, 4, 29, 0, 
    31, 0, 41, 0, 0, 15, 40, 25, 43, 0, 36, 46, 0, 17, 19, 
    38, 16, 6, 37, 0, 0, 0, 31, 42, 0, 49, 31, 0, 0, 21, 
    26, 27, 10, 17, 0, 0, 56, 9, 34, 0, 35, 36, 0, 0, 26, 
    31, 0, 62, 0, 9, 0, 22, 6, 0, 11, 0, 45, 0, 1, 0, 
    12, 0, 70, 0, 21, 3, 0, 12, 2, 4, 35, 2, 0, 0, 3, 
    0, 0, 62, 0, 69, 1, 0, 4, 41, 21, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 49, 42, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 83, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 51, 22, 0, 9, 0, 0, 0, 0, 0, 2, 0, 0, 
    21, 0, 0, 0, 3, 0, 0, 2, 0, 0, 4, 0, 0, 5, 32, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 23, 19, 0, 0, 
    22, 0, 0, 0, 0, 7, 20, 22, 33, 42, 50, 52, 55, 55, 56, 
    74, 25, 0, 0, 0, 43, 46, 45, 50, 56, 60, 60, 56, 57, 59, 
    77, 64, 8, 0, 28, 45, 47, 49, 50, 55, 64, 66, 68, 73, 71, 
    74, 72, 55, 29, 49, 53, 49, 46, 47, 52, 61, 61, 56, 67, 74, 
    
    -- channel=28
    8, 13, 13, 10, 10, 14, 10, 10, 11, 7, 1, 8, 8, 4, 5, 
    12, 17, 17, 9, 18, 40, 0, 8, 0, 17, 0, 0, 6, 10, 6, 
    0, 18, 11, 10, 16, 38, 0, 0, 2, 51, 0, 0, 0, 6, 20, 
    0, 58, 6, 19, 7, 18, 10, 0, 0, 56, 0, 0, 0, 0, 44, 
    0, 51, 0, 52, 27, 3, 0, 0, 0, 56, 2, 0, 7, 0, 15, 
    0, 19, 0, 10, 60, 0, 0, 0, 0, 127, 0, 0, 15, 0, 0, 
    0, 0, 0, 0, 74, 40, 6, 0, 0, 119, 0, 0, 6, 17, 0, 
    0, 0, 0, 0, 45, 74, 0, 0, 0, 81, 0, 0, 19, 6, 0, 
    0, 13, 0, 30, 0, 2, 0, 9, 17, 0, 21, 0, 12, 18, 19, 
    0, 9, 0, 56, 0, 0, 21, 11, 0, 0, 0, 0, 31, 39, 0, 
    60, 3, 0, 114, 0, 0, 43, 0, 0, 0, 4, 12, 14, 10, 0, 
    47, 17, 0, 109, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 0, 
    0, 38, 33, 18, 0, 0, 0, 0, 0, 1, 6, 5, 0, 0, 6, 
    0, 0, 70, 0, 0, 2, 0, 0, 1, 2, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 6, 2, 0, 0, 30, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 8, 8, 7, 8, 
    20, 0, 0, 0, 0, 0, 1, 3, 6, 10, 12, 12, 9, 8, 10, 
    21, 15, 0, 0, 0, 2, 2, 5, 5, 8, 13, 15, 15, 21, 16, 
    15, 17, 9, 4, 7, 11, 6, 1, 0, 4, 9, 11, 5, 9, 16, 
    
    -- channel=30
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 6, 0, 0, 16, 9, 0, 
    6, 29, 0, 0, 0, 28, 21, 24, 0, 0, 0, 0, 0, 11, 4, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 4, 0, 0, 6, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 53, 13, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 23, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 18, 4, 0, 5, 2, 1, 0, 7, 
    0, 0, 0, 0, 0, 39, 14, 0, 0, 0, 16, 28, 17, 3, 0, 
    8, 0, 0, 0, 0, 0, 5, 0, 0, 15, 19, 7, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 8, 7, 
    31, 22, 0, 0, 18, 60, 37, 36, 15, 0, 0, 0, 0, 0, 0, 
    0, 25, 20, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 31, 6, 0, 0, 0, 0, 0, 0, 3, 2, 0, 3, 
    0, 0, 2, 40, 9, 12, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 15, 0, 10, 0, 1, 3, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 28, 15, 0, 0, 6, 5, 15, 0, 0, 
    42, 0, 0, 0, 3, 0, 0, 14, 1, 0, 23, 1, 17, 16, 0, 
    46, 0, 23, 0, 0, 1, 20, 22, 10, 0, 0, 29, 0, 17, 0, 
    51, 0, 33, 6, 0, 17, 9, 15, 23, 0, 34, 43, 0, 10, 12, 
    53, 0, 10, 20, 0, 0, 0, 19, 29, 0, 43, 25, 0, 0, 12, 
    36, 0, 29, 3, 0, 0, 49, 5, 20, 0, 22, 29, 0, 0, 9, 
    28, 0, 64, 0, 17, 0, 13, 0, 0, 5, 0, 40, 0, 0, 0, 
    0, 0, 53, 0, 25, 13, 0, 0, 13, 8, 32, 3, 0, 0, 4, 
    0, 0, 47, 0, 34, 9, 0, 4, 42, 19, 0, 0, 0, 0, 9, 
    0, 0, 15, 0, 60, 50, 1, 4, 12, 0, 0, 0, 0, 0, 1, 
    9, 0, 0, 0, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 24, 23, 0, 4, 0, 0, 0, 0, 0, 1, 0, 5, 
    17, 0, 0, 0, 9, 0, 0, 0, 0, 0, 3, 0, 0, 0, 28, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 18, 13, 4, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 2, 7, 6, 12, 6, 12, 0, 0, 
    24, 4, 0, 0, 0, 0, 12, 8, 10, 0, 10, 5, 7, 6, 0, 
    29, 27, 0, 0, 30, 9, 15, 6, 10, 1, 18, 14, 9, 10, 1, 
    26, 33, 0, 0, 0, 3, 22, 11, 15, 13, 24, 13, 9, 12, 3, 
    29, 39, 0, 0, 0, 16, 22, 15, 11, 1, 19, 15, 12, 8, 0, 
    41, 42, 27, 16, 0, 12, 9, 10, 4, 0, 11, 12, 6, 0, 0, 
    40, 39, 37, 26, 20, 0, 7, 21, 6, 6, 12, 9, 1, 0, 0, 
    45, 33, 37, 25, 34, 19, 29, 44, 32, 18, 27, 31, 35, 33, 31, 
    67, 52, 33, 28, 62, 64, 58, 58, 58, 54, 59, 64, 69, 68, 70, 
    75, 59, 38, 49, 65, 59, 59, 56, 58, 61, 67, 69, 71, 73, 77, 
    84, 70, 50, 73, 57, 60, 60, 59, 61, 66, 73, 78, 77, 81, 85, 
    82, 78, 66, 69, 58, 62, 64, 60, 60, 67, 70, 69, 71, 84, 79, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 30, 3, 0, 0, 17, 26, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 15, 16, 0, 2, 2, 0, 0, 
    14, 28, 0, 1, 2, 18, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 22, 0, 18, 39, 15, 0, 0, 0, 20, 17, 4, 7, 6, 0, 
    0, 0, 0, 0, 0, 0, 11, 9, 9, 25, 0, 0, 0, 4, 16, 
    5, 0, 0, 0, 0, 17, 0, 2, 0, 5, 0, 6, 7, 13, 0, 
    3, 7, 11, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 3, 0, 0, 11, 9, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 0, 0, 18, 23, 0, 0, 0, 2, 8, 3, 0, 
    2, 0, 0, 39, 48, 30, 0, 0, 0, 17, 33, 30, 17, 12, 15, 
    0, 0, 2, 9, 0, 0, 0, 0, 0, 3, 2, 3, 7, 2, 2, 
    1, 0, 5, 0, 0, 4, 0, 1, 4, 8, 12, 11, 0, 0, 19, 
    0, 4, 0, 0, 0, 4, 9, 2, 0, 2, 0, 0, 2, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 1, 4, 24, 7, 0, 
    
    -- channel=38
    66, 69, 68, 69, 69, 65, 73, 78, 71, 57, 49, 53, 57, 61, 61, 
    70, 74, 72, 71, 69, 61, 64, 62, 47, 29, 16, 22, 33, 51, 58, 
    44, 55, 73, 74, 72, 61, 46, 30, 17, 10, 6, 6, 10, 24, 51, 
    18, 28, 69, 73, 62, 42, 28, 8, 6, 12, 17, 14, 10, 10, 38, 
    4, 16, 58, 51, 32, 18, 20, 11, 8, 12, 20, 13, 10, 8, 17, 
    0, 12, 56, 43, 28, 24, 26, 19, 11, 7, 11, 11, 9, 6, 7, 
    0, 10, 46, 60, 28, 24, 22, 14, 13, 7, 14, 9, 7, 8, 11, 
    0, 11, 10, 43, 25, 15, 6, 15, 17, 19, 16, 12, 6, 12, 34, 
    0, 1, 0, 18, 17, 20, 26, 16, 14, 32, 24, 11, 9, 31, 50, 
    6, 1, 3, 3, 11, 4, 15, 16, 3, 17, 7, 5, 10, 44, 55, 
    5, 6, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 37, 10, 0, 0, 0, 0, 0, 7, 1, 0, 0, 
    0, 0, 1, 4, 0, 0, 0, 0, 0, 2, 8, 11, 17, 18, 16, 
    23, 0, 0, 0, 0, 11, 9, 8, 10, 14, 20, 22, 15, 15, 30, 
    24, 17, 0, 0, 1, 13, 15, 10, 11, 16, 17, 13, 20, 26, 9, 
    26, 22, 9, 0, 1, 0, 2, 12, 18, 23, 18, 20, 33, 35, 23, 
    
    -- channel=40
    23, 26, 23, 21, 20, 23, 25, 27, 20, 18, 21, 24, 21, 20, 19, 
    19, 27, 24, 22, 22, 0, 6, 19, 28, 2, 0, 0, 14, 20, 16, 
    17, 37, 24, 24, 25, 49, 11, 9, 0, 0, 0, 0, 0, 12, 22, 
    0, 0, 18, 22, 10, 8, 0, 0, 0, 23, 0, 7, 0, 0, 29, 
    0, 0, 2, 13, 0, 0, 0, 0, 2, 11, 0, 0, 0, 0, 13, 
    0, 0, 0, 33, 49, 12, 0, 0, 0, 8, 0, 0, 1, 0, 0, 
    0, 0, 13, 13, 36, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 11, 0, 13, 0, 25, 0, 0, 3, 9, 9, 
    0, 0, 0, 0, 0, 31, 1, 0, 0, 5, 18, 11, 16, 10, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 2, 0, 13, 14, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 21, 0, 0, 0, 4, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 15, 0, 0, 
    51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 4, 0, 
    45, 0, 8, 0, 0, 19, 0, 3, 0, 0, 0, 38, 0, 6, 1, 
    56, 0, 10, 0, 0, 0, 0, 5, 10, 0, 32, 5, 0, 0, 0, 
    14, 0, 15, 0, 0, 0, 34, 0, 16, 0, 8, 11, 0, 0, 11, 
    2, 0, 28, 0, 0, 21, 11, 0, 0, 0, 0, 41, 0, 0, 0, 
    0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 37, 16, 0, 0, 0, 
    0, 0, 32, 0, 0, 0, 0, 0, 33, 25, 0, 0, 0, 0, 11, 
    0, 0, 26, 0, 16, 73, 13, 18, 20, 6, 0, 1, 0, 0, 4, 
    7, 0, 0, 0, 113, 3, 3, 3, 5, 0, 0, 0, 0, 9, 0, 
    23, 1, 0, 7, 32, 0, 7, 0, 1, 0, 1, 3, 18, 0, 0, 
    20, 1, 0, 24, 17, 0, 7, 10, 0, 0, 3, 11, 0, 0, 40, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 50, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 27, 0, 1, 0, 0, 0, 
    0, 49, 0, 0, 0, 0, 16, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 52, 0, 11, 59, 37, 0, 0, 0, 28, 6, 0, 6, 1, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 74, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 31, 0, 0, 0, 39, 0, 0, 2, 13, 5, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 9, 0, 0, 5, 6, 0, 0, 0, 0, 9, 21, 
    0, 0, 0, 17, 0, 0, 9, 21, 0, 0, 0, 0, 20, 19, 0, 
    0, 0, 0, 78, 65, 43, 19, 0, 0, 0, 15, 36, 11, 0, 0, 
    0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 2, 6, 10, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 12, 0, 0, 34, 8, 0, 
    
    -- channel=44
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 0, 4, 0, 4, 4, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 20, 1, 0, 0, 12, 1, 25, 0, 0, 
    63, 0, 0, 0, 7, 0, 6, 10, 2, 0, 29, 1, 16, 18, 0, 
    46, 0, 24, 0, 0, 0, 30, 24, 15, 0, 4, 36, 0, 25, 0, 
    27, 0, 32, 0, 0, 0, 29, 19, 44, 0, 37, 36, 0, 8, 12, 
    20, 29, 0, 32, 0, 0, 9, 18, 44, 0, 44, 26, 0, 0, 18, 
    16, 15, 13, 15, 0, 0, 43, 1, 21, 0, 22, 32, 0, 0, 2, 
    21, 0, 61, 0, 11, 0, 10, 5, 0, 12, 0, 32, 0, 0, 0, 
    0, 0, 68, 0, 34, 0, 0, 15, 8, 2, 29, 0, 0, 0, 1, 
    0, 0, 60, 0, 60, 20, 0, 4, 41, 14, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 78, 28, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 13, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 50, 12, 0, 4, 0, 0, 0, 0, 0, 0, 0, 13, 
    19, 0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 0, 10, 33, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 1, 0, 0, 12, 13, 22, 16, 0, 0, 
    0, 0, 0, 0, 1, 1, 11, 32, 10, 0, 0, 0, 0, 8, 0, 
    4, 24, 5, 0, 1, 10, 0, 0, 0, 0, 0, 0, 1, 4, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 4, 0, 0, 0, 12, 
    0, 0, 0, 17, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 2, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 8, 13, 2, 0, 
    0, 0, 3, 4, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 7, 11, 21, 10, 0, 38, 7, 0, 10, 2, 0, 
    0, 0, 0, 20, 0, 0, 3, 0, 3, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 15, 0, 0, 6, 10, 
    0, 0, 0, 0, 0, 22, 34, 31, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 7, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 1, 40, 0, 16, 0, 0, 0, 9, 0, 0, 0, 0, 9, 
    49, 0, 0, 10, 0, 16, 0, 0, 0, 0, 0, 7, 0, 0, 1, 
    62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 34, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 5, 0, 6, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    28, 26, 29, 28, 29, 24, 30, 35, 30, 22, 19, 21, 22, 22, 23, 
    31, 27, 30, 29, 31, 12, 18, 20, 19, 4, 0, 0, 3, 21, 22, 
    8, 36, 30, 31, 32, 17, 8, 0, 0, 0, 0, 0, 0, 4, 19, 
    0, 8, 25, 31, 16, 18, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 15, 34, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 1, 
    0, 0, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    33, 31, 32, 33, 35, 30, 35, 41, 39, 33, 29, 28, 28, 33, 35, 
    36, 35, 34, 35, 33, 0, 33, 30, 34, 6, 0, 4, 14, 28, 30, 
    21, 34, 34, 37, 35, 18, 22, 22, 6, 0, 0, 0, 0, 17, 20, 
    5, 0, 33, 35, 24, 18, 0, 0, 0, 0, 0, 0, 0, 9, 17, 
    0, 0, 29, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 
    0, 0, 23, 9, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 
    0, 0, 20, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 0, 1, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 10, 0, 5, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    32, 33, 35, 32, 32, 32, 34, 38, 33, 25, 22, 29, 28, 26, 25, 
    35, 36, 36, 32, 35, 37, 10, 28, 13, 14, 0, 0, 18, 31, 27, 
    17, 48, 37, 35, 38, 26, 0, 0, 5, 14, 0, 0, 0, 16, 34, 
    0, 48, 28, 38, 23, 20, 0, 0, 0, 22, 0, 0, 0, 0, 44, 
    0, 10, 0, 37, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 18, 
    0, 0, 0, 19, 30, 0, 0, 0, 0, 67, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 36, 18, 0, 0, 0, 47, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 18, 0, 0, 0, 31, 0, 0, 1, 0, 1, 
    0, 0, 0, 9, 0, 0, 0, 0, 6, 0, 8, 0, 8, 17, 25, 
    0, 0, 0, 2, 0, 0, 2, 0, 0, 0, 0, 0, 20, 33, 18, 
    9, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 5, 46, 0, 0, 0, 32, 11, 2, 3, 4, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 26, 38, 0, 0, 0, 0, 10, 
    0, 71, 0, 6, 0, 30, 0, 0, 0, 10, 0, 0, 0, 0, 24, 
    0, 20, 0, 52, 17, 0, 0, 0, 0, 78, 0, 0, 8, 0, 1, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 115, 0, 0, 2, 0, 6, 
    0, 0, 0, 0, 7, 52, 0, 0, 0, 58, 0, 0, 11, 23, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 21, 0, 0, 10, 0, 0, 
    0, 0, 0, 25, 0, 0, 0, 4, 27, 0, 0, 0, 8, 25, 5, 
    0, 0, 0, 38, 0, 0, 44, 0, 0, 0, 0, 2, 23, 12, 0, 
    29, 0, 0, 126, 0, 0, 0, 0, 0, 0, 34, 29, 10, 3, 0, 
    0, 3, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 65, 0, 0, 2, 0, 0, 0, 7, 11, 10, 0, 0, 26, 
    0, 0, 23, 0, 0, 3, 0, 0, 0, 1, 0, 0, 0, 26, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 0, 6, 44, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 16, 15, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 11, 12, 0, 1, 1, 11, 13, 0, 
    25, 0, 0, 0, 0, 0, 0, 8, 12, 0, 0, 10, 9, 19, 0, 
    21, 0, 0, 0, 0, 0, 0, 6, 16, 0, 2, 11, 9, 17, 18, 
    21, 4, 0, 0, 0, 0, 0, 0, 16, 0, 6, 11, 10, 8, 9, 
    11, 12, 12, 0, 0, 0, 6, 0, 2, 0, 0, 10, 10, 0, 0, 
    14, 9, 20, 0, 0, 0, 0, 1, 4, 0, 0, 10, 3, 0, 0, 
    0, 6, 21, 9, 12, 6, 0, 5, 8, 0, 15, 20, 8, 0, 0, 
    0, 1, 17, 0, 24, 29, 16, 17, 31, 29, 39, 46, 46, 31, 30, 
    39, 13, 18, 0, 12, 34, 36, 38, 50, 55, 60, 61, 63, 63, 64, 
    77, 37, 8, 0, 45, 57, 58, 56, 59, 62, 68, 68, 67, 68, 71, 
    82, 69, 28, 22, 50, 59, 60, 59, 61, 65, 69, 69, 72, 74, 71, 
    79, 74, 58, 47, 56, 56, 59, 60, 60, 63, 67, 68, 66, 76, 82, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=57
    5, 6, 8, 3, 3, 9, 5, 5, 2, 0, 2, 10, 9, 2, 0, 
    6, 10, 9, 2, 10, 17, 0, 0, 0, 16, 0, 0, 11, 15, 2, 
    0, 34, 6, 4, 7, 12, 0, 0, 7, 35, 0, 0, 0, 11, 21, 
    0, 49, 1, 11, 0, 21, 0, 0, 0, 44, 0, 0, 0, 0, 47, 
    0, 20, 0, 49, 0, 0, 0, 0, 0, 62, 0, 0, 0, 0, 15, 
    0, 7, 0, 0, 50, 0, 0, 0, 0, 101, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 49, 29, 0, 0, 0, 81, 0, 0, 3, 8, 0, 
    0, 0, 0, 0, 28, 35, 0, 0, 0, 47, 0, 0, 14, 0, 0, 
    0, 0, 0, 24, 0, 9, 0, 0, 21, 0, 6, 0, 16, 20, 7, 
    0, 0, 0, 39, 0, 0, 28, 0, 0, 0, 0, 3, 30, 22, 0, 
    38, 0, 0, 88, 0, 0, 17, 0, 0, 0, 1, 4, 2, 4, 0, 
    29, 21, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 
    
    -- channel=58
    5, 0, 3, 1, 2, 0, 1, 2, 0, 0, 1, 4, 3, 2, 0, 
    3, 0, 3, 0, 7, 0, 6, 0, 0, 2, 0, 0, 3, 7, 0, 
    0, 17, 3, 0, 2, 0, 0, 7, 17, 0, 0, 2, 0, 15, 0, 
    0, 12, 2, 3, 0, 21, 0, 8, 0, 19, 0, 0, 0, 0, 14, 
    8, 0, 10, 58, 0, 21, 0, 0, 0, 51, 0, 0, 0, 0, 21, 
    46, 0, 16, 3, 0, 36, 0, 0, 0, 27, 0, 5, 0, 0, 7, 
    68, 0, 24, 0, 0, 8, 0, 1, 0, 0, 0, 0, 3, 0, 0, 
    42, 0, 41, 0, 26, 0, 0, 0, 0, 0, 0, 0, 5, 0, 15, 
    7, 0, 8, 0, 12, 16, 0, 0, 21, 0, 0, 0, 4, 1, 0, 
    0, 0, 0, 2, 0, 38, 35, 0, 12, 0, 0, 8, 3, 0, 2, 
    0, 3, 0, 28, 0, 3, 0, 0, 0, 0, 5, 2, 2, 0, 0, 
    0, 7, 21, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 64, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 
    0, 0, 44, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 5, 8, 0, 0, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=62
    0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 3, 0, 0, 4, 50, 3, 0, 0, 11, 22, 4, 0, 0, 1, 
    0, 0, 1, 1, 0, 0, 0, 0, 11, 20, 0, 12, 0, 0, 2, 
    7, 40, 2, 3, 1, 13, 22, 5, 1, 0, 0, 0, 0, 0, 0, 
    24, 39, 3, 17, 67, 29, 0, 6, 0, 24, 21, 8, 11, 11, 0, 
    0, 5, 8, 0, 0, 0, 25, 12, 11, 42, 0, 0, 0, 7, 23, 
    15, 0, 0, 0, 0, 30, 0, 13, 0, 7, 0, 7, 6, 18, 10, 
    14, 14, 12, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    8, 1, 0, 14, 6, 0, 0, 10, 17, 0, 0, 0, 0, 14, 13, 
    0, 0, 3, 15, 0, 0, 22, 33, 0, 0, 0, 0, 16, 11, 0, 
    0, 0, 0, 64, 85, 43, 0, 0, 0, 5, 27, 33, 7, 0, 0, 
    0, 0, 16, 21, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 
    0, 0, 18, 0, 0, 3, 0, 0, 0, 6, 10, 13, 0, 0, 25, 
    0, 0, 0, 0, 0, 2, 8, 0, 0, 2, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 16, 0, 4, 34, 10, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 8, 7, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 6, 8, 8, 10, 11, 13, 3, 0, 
    13, 0, 0, 0, 0, 0, 11, 8, 15, 0, 1, 5, 3, 3, 0, 
    35, 11, 0, 0, 19, 8, 0, 3, 7, 0, 23, 17, 8, 8, 0, 
    23, 26, 0, 0, 0, 0, 19, 7, 14, 2, 23, 11, 7, 3, 1, 
    22, 22, 1, 0, 0, 12, 35, 21, 7, 3, 16, 16, 10, 11, 0, 
    30, 29, 29, 0, 1, 21, 6, 6, 0, 2, 13, 24, 8, 0, 0, 
    30, 31, 29, 11, 17, 7, 0, 4, 14, 17, 23, 9, 0, 0, 0, 
    23, 24, 33, 0, 3, 8, 25, 44, 29, 18, 15, 17, 29, 31, 32, 
    69, 38, 19, 12, 79, 65, 56, 55, 49, 49, 51, 55, 55, 57, 58, 
    66, 59, 19, 49, 71, 48, 50, 49, 50, 51, 53, 55, 61, 63, 56, 
    72, 57, 52, 70, 51, 50, 49, 50, 52, 55, 64, 69, 66, 64, 85, 
    72, 64, 58, 67, 58, 58, 59, 50, 47, 52, 60, 58, 49, 70, 67, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    17, 15, 17, 18, 17, 12, 20, 23, 17, 6, 0, 1, 5, 12, 14, 
    18, 18, 19, 18, 17, 8, 8, 4, 0, 0, 0, 0, 0, 2, 11, 
    0, 5, 20, 20, 22, 12, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 17, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 0, 1, 0, 0, 0, 
    7, 11, 0, 0, 6, 6, 2, 0, 0, 3, 5, 0, 0, 0, 0, 
    20, 16, 0, 0, 10, 1, 1, 0, 0, 19, 12, 0, 3, 1, 0, 
    17, 18, 0, 0, 0, 9, 14, 4, 0, 23, 7, 3, 3, 6, 0, 
    22, 14, 8, 0, 0, 23, 8, 5, 0, 8, 3, 1, 5, 1, 0, 
    27, 28, 15, 7, 7, 0, 0, 5, 3, 0, 5, 0, 0, 0, 0, 
    21, 26, 12, 19, 11, 4, 5, 10, 11, 1, 0, 0, 0, 0, 0, 
    31, 25, 11, 31, 19, 25, 35, 27, 14, 9, 18, 24, 31, 35, 32, 
    52, 34, 16, 40, 36, 27, 32, 30, 30, 33, 37, 39, 39, 41, 41, 
    48, 46, 31, 42, 23, 33, 33, 31, 32, 36, 41, 44, 44, 45, 48, 
    48, 44, 53, 31, 30, 36, 33, 33, 34, 39, 44, 46, 44, 55, 51, 
    46, 44, 41, 32, 33, 36, 36, 33, 36, 39, 40, 39, 46, 53, 40, 
    
    -- channel=67
    31, 29, 31, 32, 34, 28, 36, 42, 40, 33, 24, 23, 22, 25, 28, 
    35, 35, 33, 35, 32, 8, 32, 35, 24, 0, 0, 0, 9, 23, 27, 
    26, 29, 37, 37, 38, 24, 13, 7, 0, 0, 0, 0, 0, 4, 14, 
    0, 0, 37, 38, 34, 11, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 21, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=68
    0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 2, 4, 
    0, 0, 0, 2, 0, 0, 9, 4, 12, 0, 6, 2, 0, 0, 2, 
    17, 0, 0, 1, 0, 6, 24, 4, 0, 0, 13, 6, 27, 0, 0, 
    65, 0, 0, 0, 12, 0, 12, 4, 4, 0, 36, 1, 21, 12, 0, 
    43, 0, 17, 0, 12, 0, 33, 21, 20, 0, 8, 29, 1, 28, 0, 
    4, 0, 22, 0, 0, 0, 41, 21, 51, 0, 35, 32, 0, 13, 6, 
    0, 50, 0, 41, 0, 0, 27, 19, 51, 0, 44, 21, 0, 0, 13, 
    0, 36, 0, 23, 0, 0, 49, 10, 24, 0, 28, 31, 0, 0, 5, 
    15, 0, 40, 0, 0, 0, 14, 12, 0, 23, 0, 38, 0, 0, 0, 
    6, 0, 69, 0, 24, 0, 0, 30, 0, 6, 40, 0, 0, 0, 4, 
    0, 0, 66, 0, 63, 1, 0, 20, 40, 19, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 86, 27, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 33, 62, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 90, 13, 0, 5, 0, 0, 0, 0, 0, 1, 0, 19, 
    20, 0, 0, 19, 5, 0, 0, 0, 0, 0, 5, 0, 0, 15, 34, 
    
    -- channel=69
    0, 0, 0, 2, 3, 0, 0, 0, 1, 0, 0, 0, 0, 5, 7, 
    4, 0, 0, 1, 0, 35, 19, 0, 0, 0, 31, 15, 0, 0, 3, 
    0, 0, 0, 2, 0, 0, 4, 0, 10, 0, 15, 18, 26, 0, 0, 
    56, 4, 2, 0, 10, 0, 30, 22, 11, 0, 26, 0, 14, 15, 0, 
    57, 19, 24, 0, 52, 44, 24, 31, 5, 0, 28, 42, 14, 33, 0, 
    22, 0, 30, 0, 0, 0, 46, 32, 50, 0, 21, 20, 0, 21, 39, 
    42, 10, 0, 22, 0, 4, 0, 33, 28, 0, 26, 34, 11, 12, 28, 
    37, 23, 30, 25, 0, 0, 4, 0, 14, 0, 15, 25, 0, 0, 11, 
    34, 0, 56, 0, 30, 0, 8, 22, 0, 20, 0, 0, 0, 1, 12, 
    0, 0, 53, 0, 10, 3, 0, 43, 14, 0, 0, 0, 0, 0, 0, 
    0, 1, 38, 0, 123, 59, 0, 0, 12, 29, 27, 30, 6, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 1, 2, 1, 11, 8, 10, 
    21, 0, 0, 0, 8, 10, 8, 8, 10, 12, 13, 15, 0, 0, 20, 
    17, 7, 0, 0, 10, 7, 24, 9, 3, 6, 4, 0, 8, 7, 0, 
    25, 6, 1, 0, 0, 0, 0, 5, 15, 24, 17, 9, 18, 31, 30, 
    
    -- channel=70
    5, 2, 3, 2, 3, 3, 7, 9, 7, 9, 10, 9, 4, 4, 3, 
    5, 8, 4, 4, 1, 0, 4, 11, 10, 0, 0, 0, 7, 9, 4, 
    10, 18, 8, 5, 6, 0, 0, 1, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 8, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    3, 0, 0, 0, 0, 3, 0, 0, 0, 1, 4, 5, 3, 1, 1, 
    0, 0, 1, 0, 2, 0, 0, 0, 4, 3, 0, 0, 1, 7, 3, 
    0, 26, 4, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 9, 8, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 2, 2, 12, 
    0, 0, 0, 1, 0, 0, 0, 0, 1, 18, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 5, 4, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 3, 1, 2, 0, 0, 6, 8, 7, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 9, 8, 6, 4, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 3, 4, 6, 2, 
    8, 1, 0, 0, 0, 1, 0, 4, 6, 7, 6, 6, 0, 0, 4, 
    2, 7, 1, 0, 0, 2, 4, 3, 2, 3, 4, 2, 4, 8, 0, 
    0, 4, 10, 0, 4, 5, 0, 0, 3, 4, 3, 6, 8, 0, 0, 
    
    -- channel=72
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 2, 0, 0, 0, 0, 10, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 16, 7, 0, 0, 7, 0, 13, 7, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 33, 18, 18, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 16, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 33, 9, 1, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 24, 0, 21, 0, 0, 8, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 9, 2, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 19, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 4, 20, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 54, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    2, 0, 0, 0, 0, 15, 0, 2, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 2, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 0, 44, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 23, 6, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 0, 0, 0, 16, 31, 37, 33, 2, 0, 0, 0, 0, 0, 0, 
    0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 26, 
    0, 0, 20, 20, 16, 22, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 4, 0, 0, 
    24, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 2, 0, 0, 0, 
    28, 0, 7, 0, 0, 14, 7, 0, 1, 0, 27, 25, 0, 0, 0, 
    18, 17, 0, 1, 0, 0, 17, 5, 19, 0, 38, 2, 0, 0, 0, 
    10, 16, 0, 0, 0, 0, 52, 13, 11, 0, 22, 13, 0, 0, 0, 
    21, 1, 32, 0, 0, 13, 8, 0, 0, 0, 0, 31, 0, 0, 0, 
    18, 6, 44, 0, 15, 0, 0, 0, 0, 10, 25, 0, 0, 0, 0, 
    0, 2, 48, 0, 9, 0, 0, 29, 30, 0, 0, 0, 0, 0, 0, 
    0, 1, 14, 0, 98, 57, 11, 10, 7, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 24, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 79, 16, 0, 0, 0, 0, 0, 0, 4, 4, 0, 26, 
    17, 0, 0, 29, 6, 0, 3, 0, 0, 0, 2, 0, 0, 4, 25, 
    
    -- channel=77
    20, 20, 21, 22, 22, 19, 21, 24, 26, 21, 13, 13, 16, 16, 21, 
    22, 22, 22, 23, 24, 24, 16, 19, 14, 12, 5, 0, 1, 13, 20, 
    12, 15, 22, 24, 24, 18, 10, 5, 3, 4, 0, 0, 0, 0, 15, 
    6, 3, 21, 25, 21, 17, 12, 0, 1, 0, 0, 0, 0, 0, 8, 
    0, 1, 12, 24, 18, 0, 0, 0, 0, 0, 2, 0, 2, 3, 0, 
    0, 0, 6, 6, 0, 0, 2, 1, 2, 5, 0, 0, 1, 2, 0, 
    0, 0, 0, 24, 6, 3, 5, 0, 3, 3, 0, 0, 0, 3, 0, 
    0, 0, 0, 15, 11, 7, 0, 0, 0, 4, 0, 0, 0, 0, 3, 
    0, 0, 0, 2, 0, 0, 0, 6, 1, 2, 4, 0, 0, 5, 14, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 3, 0, 0, 0, 12, 16, 
    0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    0, 0, 4, 4, 4, 2, 1, 2, 1, 0, 0, 0, 0, 4, 3, 
    7, 6, 4, 1, 7, 39, 9, 0, 0, 5, 20, 3, 0, 0, 1, 
    0, 0, 3, 3, 0, 0, 0, 0, 11, 18, 5, 16, 4, 0, 0, 
    15, 31, 4, 5, 0, 14, 20, 9, 1, 0, 0, 0, 0, 0, 0, 
    34, 38, 9, 26, 58, 41, 2, 7, 0, 24, 26, 14, 11, 14, 0, 
    0, 0, 10, 0, 0, 0, 20, 21, 13, 31, 0, 0, 0, 11, 26, 
    29, 0, 0, 0, 0, 19, 0, 13, 2, 1, 0, 10, 8, 17, 15, 
    18, 14, 23, 12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    11, 0, 3, 3, 4, 0, 0, 6, 18, 0, 0, 0, 0, 15, 16, 
    0, 0, 3, 16, 0, 0, 24, 32, 0, 0, 0, 0, 14, 10, 0, 
    0, 0, 0, 56, 81, 49, 0, 0, 0, 7, 26, 28, 5, 0, 0, 
    0, 0, 22, 16, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 
    0, 0, 10, 0, 0, 2, 0, 0, 1, 6, 10, 12, 0, 0, 22, 
    0, 0, 0, 0, 0, 4, 9, 0, 0, 1, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 16, 2, 6, 33, 13, 1, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=81
    16, 15, 18, 19, 20, 16, 16, 20, 20, 13, 8, 9, 15, 15, 19, 
    20, 17, 19, 19, 23, 27, 15, 7, 6, 14, 15, 3, 0, 10, 17, 
    0, 11, 18, 19, 19, 8, 5, 4, 9, 24, 15, 21, 15, 2, 13, 
    14, 17, 16, 20, 12, 23, 20, 17, 17, 15, 15, 8, 12, 5, 11, 
    30, 24, 17, 34, 36, 27, 10, 10, 7, 23, 20, 14, 17, 18, 2, 
    12, 12, 14, 5, 0, 6, 16, 19, 15, 26, 11, 8, 15, 21, 16, 
    19, 6, 0, 15, 13, 17, 12, 20, 14, 23, 12, 11, 15, 20, 16, 
    13, 21, 13, 18, 28, 13, 10, 5, 12, 19, 15, 8, 13, 11, 20, 
    16, 14, 6, 14, 10, 5, 9, 14, 20, 16, 0, 3, 7, 18, 18, 
    17, 17, 13, 21, 2, 10, 23, 27, 5, 2, 8, 10, 16, 20, 17, 
    13, 14, 11, 33, 46, 24, 16, 6, 9, 17, 16, 22, 12, 5, 4, 
    0, 11, 26, 32, 0, 0, 0, 0, 4, 13, 16, 16, 18, 20, 18, 
    18, 0, 20, 3, 1, 15, 14, 15, 19, 21, 23, 21, 17, 19, 26, 
    19, 14, 0, 2, 17, 19, 19, 14, 17, 18, 18, 14, 20, 19, 8, 
    19, 17, 8, 3, 13, 10, 14, 19, 23, 23, 18, 22, 33, 26, 19, 
    
    -- channel=82
    51, 50, 53, 53, 54, 48, 55, 58, 55, 47, 40, 41, 43, 46, 47, 
    54, 52, 55, 55, 54, 45, 50, 47, 39, 22, 15, 15, 22, 39, 46, 
    38, 45, 56, 56, 57, 37, 31, 17, 14, 9, 5, 5, 11, 20, 36, 
    15, 27, 51, 55, 49, 34, 21, 14, 10, 9, 11, 10, 6, 10, 25, 
    7, 15, 46, 43, 27, 23, 10, 9, 6, 9, 10, 12, 8, 8, 17, 
    2, 6, 42, 40, 0, 11, 12, 10, 7, 10, 12, 7, 7, 7, 8, 
    1, 3, 28, 41, 16, 18, 12, 14, 6, 7, 7, 6, 6, 6, 11, 
    2, 0, 15, 30, 26, 13, 10, 6, 10, 12, 10, 4, 4, 10, 23, 
    0, 0, 4, 8, 23, 6, 9, 10, 12, 21, 9, 6, 6, 17, 39, 
    1, 0, 0, 0, 4, 14, 10, 8, 9, 13, 9, 2, 11, 35, 44, 
    0, 1, 0, 0, 9, 6, 5, 0, 2, 2, 0, 0, 0, 0, 4, 
    0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 16, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    45, 0, 0, 0, 6, 0, 14, 3, 0, 0, 10, 0, 0, 0, 0, 
    52, 0, 20, 0, 60, 34, 9, 5, 0, 0, 2, 24, 0, 12, 0, 
    1, 0, 24, 0, 0, 0, 27, 9, 24, 0, 13, 2, 0, 0, 10, 
    12, 0, 0, 21, 0, 0, 0, 18, 15, 0, 13, 4, 0, 0, 2, 
    10, 4, 7, 22, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 31, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 38, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 117, 43, 0, 0, 18, 8, 0, 1, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=84
    2, 2, 0, 0, 0, 0, 0, 1, 0, 2, 11, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 1, 0, 
    13, 19, 0, 0, 0, 28, 15, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 11, 3, 0, 
    0, 0, 3, 0, 0, 0, 2, 0, 12, 0, 0, 0, 0, 0, 0, 
    16, 0, 10, 14, 19, 21, 0, 0, 0, 0, 17, 23, 0, 0, 0, 
    0, 3, 11, 9, 0, 0, 7, 0, 9, 0, 19, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 54, 26, 14, 0, 15, 5, 0, 12, 14, 
    0, 0, 12, 0, 0, 36, 2, 0, 0, 0, 3, 48, 7, 0, 0, 
    5, 0, 13, 0, 1, 5, 0, 0, 0, 35, 45, 2, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 32, 27, 0, 0, 0, 0, 0, 0, 
    15, 6, 0, 0, 73, 46, 12, 9, 1, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 4, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 58, 10, 0, 0, 0, 0, 0, 0, 1, 0, 0, 31, 
    5, 0, 0, 24, 9, 5, 13, 0, 0, 0, 0, 0, 0, 0, 9, 
    
    -- channel=85
    6, 0, 6, 3, 5, 1, 2, 3, 4, 0, 3, 4, 6, 2, 1, 
    6, 0, 3, 1, 8, 0, 7, 0, 3, 11, 0, 0, 1, 7, 0, 
    0, 14, 5, 3, 4, 0, 11, 9, 20, 0, 0, 6, 0, 8, 0, 
    0, 6, 0, 5, 0, 23, 0, 12, 1, 4, 0, 0, 2, 2, 3, 
    20, 0, 12, 52, 0, 19, 0, 0, 0, 48, 0, 2, 0, 0, 13, 
    51, 0, 21, 18, 0, 43, 0, 0, 0, 17, 0, 15, 0, 3, 12, 
    74, 0, 22, 0, 0, 19, 0, 13, 0, 0, 4, 4, 5, 3, 0, 
    54, 0, 39, 0, 17, 0, 1, 0, 0, 0, 4, 0, 3, 0, 15, 
    22, 0, 27, 0, 23, 12, 3, 0, 16, 0, 0, 3, 4, 2, 0, 
    0, 0, 0, 0, 0, 40, 36, 0, 7, 0, 0, 9, 0, 0, 4, 
    0, 5, 0, 17, 3, 2, 0, 0, 8, 8, 7, 9, 5, 0, 11, 
    0, 11, 22, 0, 0, 28, 0, 1, 7, 4, 0, 0, 0, 0, 0, 
    0, 0, 64, 0, 27, 2, 0, 0, 0, 1, 1, 0, 0, 5, 5, 
    0, 2, 22, 0, 16, 2, 1, 0, 2, 0, 0, 0, 4, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 6, 1, 0, 0, 6, 9, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 5, 16, 16, 10, 10, 1, 0, 
    11, 4, 0, 0, 0, 0, 8, 7, 7, 13, 6, 8, 4, 3, 0, 
    16, 23, 0, 0, 18, 22, 16, 8, 7, 10, 18, 11, 9, 5, 4, 
    23, 19, 0, 0, 12, 9, 12, 11, 10, 19, 15, 6, 10, 9, 10, 
    22, 25, 0, 0, 7, 10, 17, 10, 10, 25, 14, 12, 12, 12, 7, 
    26, 27, 17, 0, 4, 20, 10, 8, 2, 12, 7, 11, 11, 8, 0, 
    30, 34, 18, 13, 7, 9, 7, 11, 10, 10, 7, 0, 6, 0, 0, 
    19, 28, 18, 31, 19, 7, 12, 23, 18, 0, 0, 7, 9, 0, 0, 
    29, 28, 20, 33, 27, 32, 30, 24, 15, 17, 25, 28, 33, 32, 28, 
    45, 29, 23, 38, 30, 23, 35, 35, 31, 33, 35, 38, 40, 40, 39, 
    43, 41, 26, 36, 20, 35, 36, 33, 33, 35, 39, 43, 41, 40, 46, 
    43, 44, 44, 22, 23, 37, 36, 36, 35, 39, 41, 41, 41, 48, 45, 
    43, 44, 41, 35, 30, 32, 31, 32, 37, 41, 40, 39, 45, 51, 40, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 3, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 33, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 15, 0, 0, 3, 0, 4, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 0, 0, 2, 8, 
    0, 0, 0, 0, 0, 38, 23, 24, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=88
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=89
    60, 58, 59, 61, 62, 55, 63, 67, 63, 57, 49, 46, 47, 53, 54, 
    60, 59, 61, 64, 59, 43, 63, 57, 50, 18, 17, 22, 28, 41, 52, 
    54, 44, 63, 64, 66, 63, 45, 25, 12, 7, 23, 14, 25, 26, 37, 
    33, 14, 60, 60, 58, 31, 28, 23, 19, 15, 31, 26, 18, 19, 22, 
    20, 19, 62, 32, 25, 34, 32, 22, 22, 0, 22, 28, 13, 17, 23, 
    28, 20, 59, 64, 16, 28, 29, 24, 24, 0, 42, 27, 14, 16, 11, 
    18, 34, 38, 56, 25, 18, 37, 29, 26, 4, 34, 21, 13, 9, 24, 
    22, 15, 27, 36, 29, 25, 46, 29, 23, 23, 31, 25, 10, 26, 33, 
    23, 14, 32, 9, 39, 27, 24, 21, 10, 45, 24, 29, 13, 19, 46, 
    24, 21, 28, 0, 24, 24, 7, 20, 30, 30, 28, 5, 5, 39, 55, 
    4, 22, 30, 0, 22, 16, 16, 22, 20, 10, 0, 0, 0, 4, 7, 
    0, 3, 15, 20, 61, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 46, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 1, 0, 0, 0, 1, 3, 1, 0, 0, 0, 3, 6, 
    0, 0, 0, 3, 0, 9, 14, 4, 3, 0, 13, 4, 0, 0, 4, 
    11, 0, 0, 3, 0, 0, 26, 4, 0, 0, 14, 10, 23, 0, 0, 
    68, 0, 1, 0, 17, 0, 19, 10, 3, 0, 37, 0, 23, 12, 0, 
    57, 0, 20, 0, 29, 0, 34, 29, 14, 0, 15, 35, 4, 31, 0, 
    14, 0, 30, 0, 0, 0, 48, 27, 51, 0, 33, 37, 0, 15, 15, 
    15, 31, 0, 43, 0, 0, 18, 26, 51, 0, 47, 29, 0, 0, 17, 
    12, 37, 2, 31, 0, 0, 37, 0, 28, 0, 29, 33, 0, 0, 7, 
    25, 0, 51, 0, 3, 0, 18, 16, 0, 8, 0, 29, 0, 0, 0, 
    7, 0, 75, 0, 31, 0, 0, 35, 0, 2, 27, 0, 0, 0, 6, 
    0, 0, 64, 0, 88, 21, 0, 8, 42, 21, 0, 0, 0, 0, 1, 
    0, 0, 18, 0, 61, 26, 0, 0, 6, 0, 0, 0, 0, 0, 2, 
    5, 0, 0, 13, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 66, 18, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 14, 32, 
    
    -- channel=91
    73, 76, 76, 75, 75, 74, 77, 83, 78, 67, 61, 63, 64, 65, 65, 
    72, 79, 79, 77, 77, 64, 66, 71, 63, 39, 18, 24, 42, 56, 62, 
    56, 71, 78, 79, 80, 78, 50, 39, 25, 23, 7, 9, 7, 31, 54, 
    8, 34, 68, 80, 68, 58, 27, 14, 9, 31, 16, 20, 10, 7, 48, 
    0, 13, 54, 78, 32, 34, 22, 13, 9, 33, 18, 10, 12, 2, 28, 
    7, 14, 49, 70, 50, 43, 19, 15, 0, 35, 17, 13, 15, 7, 5, 
    7, 3, 45, 58, 50, 40, 25, 19, 4, 33, 11, 7, 12, 11, 7, 
    10, 4, 14, 35, 44, 36, 21, 24, 14, 38, 18, 8, 15, 18, 32, 
    7, 9, 0, 19, 27, 37, 22, 14, 19, 34, 28, 17, 19, 29, 52, 
    18, 11, 0, 16, 5, 28, 31, 6, 13, 29, 15, 9, 13, 48, 60, 
    16, 16, 0, 24, 0, 0, 12, 10, 0, 1, 0, 0, 0, 0, 0, 
    0, 8, 4, 27, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=92
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 6, 8, 0, 
    36, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 24, 0, 27, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 55, 0, 0, 22, 0, 0, 5, 
    0, 0, 0, 20, 0, 0, 0, 0, 44, 0, 11, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 1, 0, 0, 19, 0, 0, 0, 
    0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 
    0, 0, 56, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 
    0, 0, 43, 0, 29, 0, 0, 0, 21, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    
    -- channel=93
    46, 45, 47, 48, 48, 44, 48, 49, 47, 41, 35, 35, 38, 41, 41, 
    47, 46, 48, 49, 48, 53, 48, 40, 29, 27, 29, 25, 25, 36, 42, 
    32, 37, 49, 48, 50, 38, 29, 20, 23, 30, 30, 26, 25, 25, 35, 
    30, 37, 48, 48, 43, 36, 38, 27, 24, 27, 29, 23, 18, 19, 28, 
    35, 48, 48, 46, 57, 44, 31, 23, 17, 24, 36, 29, 24, 22, 20, 
    30, 39, 47, 33, 23, 30, 38, 31, 24, 35, 36, 22, 24, 23, 22, 
    31, 34, 36, 36, 30, 39, 41, 34, 26, 34, 32, 25, 23, 27, 30, 
    34, 33, 35, 39, 38, 43, 29, 23, 27, 33, 31, 23, 21, 27, 32, 
    36, 35, 28, 31, 34, 20, 27, 28, 32, 32, 25, 13, 16, 31, 44, 
    35, 36, 29, 27, 31, 23, 28, 40, 29, 21, 14, 11, 27, 41, 42, 
    33, 36, 28, 41, 54, 43, 35, 26, 24, 16, 16, 19, 19, 22, 22, 
    14, 25, 39, 54, 29, 4, 5, 4, 9, 11, 12, 11, 13, 13, 12, 
    14, 12, 30, 43, 9, 11, 11, 10, 11, 12, 13, 15, 14, 11, 17, 
    10, 10, 17, 22, 15, 13, 13, 11, 10, 11, 11, 9, 9, 13, 11, 
    11, 7, 10, 7, 10, 8, 10, 12, 15, 15, 13, 11, 19, 20, 10, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    3, 25, 0, 0, 51, 12, 1, 0, 0, 27, 6, 0, 0, 0, 0, 
    0, 23, 0, 0, 17, 15, 21, 0, 0, 39, 0, 0, 0, 0, 0, 
    11, 16, 0, 0, 0, 39, 10, 9, 0, 28, 2, 0, 0, 0, 0, 
    22, 34, 0, 9, 0, 11, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    31, 34, 0, 23, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 28, 0, 44, 0, 0, 31, 30, 0, 0, 0, 0, 4, 9, 0, 
    53, 40, 5, 64, 40, 13, 21, 18, 5, 3, 7, 11, 12, 16, 11, 
    11, 43, 36, 57, 3, 7, 6, 5, 3, 5, 10, 14, 18, 17, 19, 
    12, 13, 58, 37, 0, 11, 4, 6, 8, 12, 16, 20, 14, 24, 28, 
    12, 17, 18, 23, 3, 13, 13, 7, 9, 12, 10, 11, 20, 24, 2, 
    
    -- channel=95
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 25, 0, 0, 0, 5, 0, 0, 
    24, 9, 0, 0, 0, 47, 14, 11, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 14, 4, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 10, 
    13, 0, 0, 22, 37, 10, 0, 0, 0, 0, 11, 13, 0, 0, 0, 
    0, 11, 13, 1, 7, 0, 13, 0, 5, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 34, 27, 2, 0, 6, 9, 0, 10, 0, 
    0, 0, 5, 0, 0, 39, 5, 0, 0, 5, 30, 37, 8, 0, 0, 
    1, 0, 2, 0, 11, 0, 0, 0, 7, 34, 31, 2, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 27, 10, 0, 0, 0, 0, 0, 1, 
    50, 3, 0, 0, 86, 51, 33, 30, 11, 0, 0, 0, 0, 0, 0, 
    1, 37, 0, 27, 52, 0, 1, 0, 0, 0, 0, 0, 3, 1, 0, 
    4, 0, 25, 52, 6, 0, 0, 0, 0, 0, 2, 12, 1, 0, 38, 
    4, 0, 8, 47, 17, 17, 17, 0, 0, 0, 1, 0, 0, 0, 6, 
    
    -- channel=96
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=97
    10, 12, 12, 13, 11, 12, 11, 10, 10, 7, 4, 5, 8, 7, 7, 
    10, 11, 12, 13, 14, 35, 12, 9, 0, 10, 14, 5, 0, 3, 9, 
    7, 0, 12, 11, 13, 11, 6, 0, 6, 28, 31, 21, 10, 0, 7, 
    13, 13, 11, 11, 15, 11, 29, 18, 14, 20, 27, 14, 10, 0, 0, 
    31, 40, 15, 17, 60, 42, 31, 20, 8, 13, 33, 20, 17, 8, 0, 
    35, 44, 21, 19, 32, 30, 44, 22, 15, 39, 40, 14, 15, 14, 7, 
    38, 41, 7, 12, 17, 44, 45, 34, 18, 39, 31, 19, 14, 22, 19, 
    48, 46, 15, 18, 18, 55, 35, 20, 19, 35, 32, 17, 14, 22, 12, 
    55, 52, 33, 28, 29, 8, 17, 26, 18, 11, 19, 2, 5, 13, 18, 
    55, 53, 37, 29, 28, 16, 23, 46, 24, 16, 0, 0, 9, 18, 11, 
    49, 51, 33, 63, 72, 47, 50, 41, 23, 6, 11, 21, 18, 14, 13, 
    26, 44, 44, 78, 48, 14, 13, 13, 17, 20, 24, 25, 31, 32, 32, 
    31, 25, 44, 72, 22, 26, 23, 22, 23, 26, 29, 35, 33, 31, 41, 
    32, 24, 34, 47, 27, 27, 27, 24, 25, 29, 30, 30, 28, 43, 34, 
    36, 30, 24, 14, 19, 21, 24, 26, 32, 35, 31, 28, 45, 51, 26, 
    
    -- channel=98
    1, 3, 9, 8, 6, 5, 7, 5, 3, 0, 0, 0, 5, 6, 4, 
    9, 10, 11, 7, 12, 50, 5, 0, 0, 0, 11, 0, 0, 0, 6, 
    0, 0, 6, 6, 3, 0, 0, 0, 1, 26, 3, 14, 1, 0, 7, 
    0, 30, 4, 8, 0, 6, 21, 9, 3, 0, 0, 0, 0, 0, 0, 
    20, 49, 6, 29, 84, 46, 0, 0, 0, 20, 14, 6, 10, 11, 0, 
    0, 5, 7, 0, 0, 0, 20, 8, 4, 56, 0, 0, 0, 9, 19, 
    0, 0, 0, 0, 0, 26, 0, 12, 0, 26, 0, 0, 0, 13, 11, 
    2, 10, 3, 9, 16, 15, 0, 0, 0, 7, 0, 0, 0, 0, 6, 
    2, 0, 0, 13, 0, 0, 0, 0, 16, 0, 0, 0, 0, 14, 23, 
    0, 0, 0, 9, 0, 0, 17, 34, 0, 0, 0, 0, 25, 26, 0, 
    0, 0, 0, 65, 87, 49, 26, 0, 0, 0, 10, 33, 6, 0, 0, 
    0, 0, 19, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 28, 4, 0, 
    
    -- channel=99
    0, 8, 0, 0, 0, 3, 0, 1, 0, 0, 0, 5, 3, 0, 0, 
    0, 7, 1, 0, 1, 41, 0, 3, 0, 13, 0, 0, 0, 8, 2, 
    3, 21, 0, 1, 0, 45, 0, 0, 0, 32, 0, 0, 0, 0, 26, 
    0, 21, 0, 5, 5, 0, 12, 0, 0, 21, 0, 0, 0, 0, 31, 
    0, 36, 0, 0, 36, 0, 0, 0, 2, 2, 1, 0, 9, 0, 0, 
    0, 36, 0, 0, 84, 0, 15, 0, 3, 51, 0, 0, 11, 0, 0, 
    0, 39, 0, 4, 61, 9, 33, 0, 0, 70, 0, 0, 0, 8, 0, 
    0, 30, 0, 9, 0, 55, 0, 2, 0, 47, 0, 0, 8, 2, 0, 
    0, 12, 0, 43, 0, 0, 0, 15, 7, 0, 23, 0, 3, 22, 1, 
    9, 0, 0, 32, 0, 0, 0, 33, 0, 3, 0, 0, 26, 23, 0, 
    74, 0, 0, 47, 0, 0, 10, 15, 0, 0, 0, 0, 0, 11, 0, 
    40, 25, 0, 60, 0, 0, 4, 0, 0, 0, 2, 2, 2, 0, 0, 
    0, 16, 0, 36, 0, 0, 0, 0, 0, 0, 3, 0, 1, 0, 3, 
    0, 0, 0, 62, 0, 0, 0, 0, 0, 0, 0, 5, 0, 5, 0, 
    0, 5, 0, 44, 0, 6, 6, 0, 1, 1, 0, 0, 10, 0, 0, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 10, 14, 11, 6, 5, 21, 23, 23, 
    40, 3, 0, 0, 45, 40, 36, 36, 31, 29, 31, 34, 32, 33, 35, 
    48, 32, 0, 9, 42, 27, 31, 29, 29, 29, 32, 32, 38, 38, 30, 
    50, 40, 18, 35, 24, 28, 30, 30, 29, 32, 40, 42, 43, 36, 59, 
    48, 41, 41, 43, 36, 33, 33, 27, 24, 29, 38, 33, 18, 42, 51, 
    
    -- channel=101
    72, 74, 73, 74, 74, 71, 79, 83, 76, 67, 60, 60, 61, 66, 63, 
    73, 78, 78, 78, 73, 54, 74, 72, 62, 24, 15, 24, 38, 55, 62, 
    60, 64, 78, 79, 79, 71, 46, 30, 16, 5, 8, 2, 15, 32, 51, 
    22, 25, 75, 76, 67, 41, 26, 13, 7, 18, 16, 19, 6, 12, 40, 
    4, 19, 67, 53, 30, 32, 24, 10, 9, 4, 16, 17, 6, 6, 27, 
    5, 12, 62, 59, 25, 30, 19, 16, 7, 0, 22, 12, 9, 4, 6, 
    0, 16, 52, 59, 33, 18, 30, 15, 13, 7, 16, 7, 5, 2, 13, 
    4, 1, 23, 41, 33, 26, 20, 19, 13, 19, 15, 9, 5, 17, 29, 
    0, 1, 4, 12, 26, 26, 19, 10, 12, 36, 25, 14, 8, 22, 54, 
    3, 2, 1, 0, 18, 15, 8, 9, 16, 25, 15, 3, 13, 50, 65, 
    0, 8, 5, 0, 0, 2, 4, 7, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 10, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=102
    12, 15, 12, 12, 10, 13, 15, 16, 11, 8, 7, 7, 6, 3, 0, 
    8, 14, 14, 14, 13, 12, 10, 14, 9, 0, 0, 0, 0, 3, 1, 
    8, 15, 15, 14, 16, 36, 8, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 13, 14, 12, 4, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 9, 15, 13, 5, 7, 0, 0, 0, 1, 0, 0, 0, 0, 
    7, 20, 13, 20, 55, 31, 12, 0, 0, 3, 16, 0, 0, 0, 0, 
    2, 16, 16, 3, 14, 21, 32, 3, 0, 16, 10, 0, 0, 0, 0, 
    14, 14, 0, 1, 0, 37, 19, 10, 0, 15, 9, 0, 0, 0, 0, 
    21, 28, 0, 5, 0, 18, 2, 0, 0, 3, 12, 0, 0, 0, 0, 
    33, 28, 0, 3, 0, 0, 1, 0, 0, 5, 0, 0, 0, 1, 9, 
    33, 29, 3, 18, 0, 0, 12, 26, 0, 0, 0, 0, 0, 0, 0, 
    15, 30, 9, 46, 51, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 24, 57, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    12, 0, 0, 0, 0, 22, 10, 11, 18, 14, 18, 17, 17, 15, 19, 
    27, 10, 0, 0, 14, 14, 15, 15, 15, 17, 17, 15, 20, 23, 14, 
    31, 25, 0, 1, 14, 11, 13, 15, 18, 18, 22, 26, 26, 22, 34, 
    27, 28, 22, 13, 19, 22, 24, 18, 11, 10, 18, 19, 7, 11, 31, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 9, 
    37, 0, 4, 0, 0, 14, 0, 0, 0, 0, 0, 6, 0, 0, 3, 
    53, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 2, 0, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 0, 0, 0, 10, 5, 0, 1, 3, 0, 
    0, 12, 0, 0, 0, 19, 0, 0, 0, 37, 22, 18, 1, 2, 8, 
    0, 18, 0, 0, 0, 9, 14, 5, 11, 45, 13, 13, 4, 0, 18, 
    14, 42, 0, 26, 44, 21, 16, 2, 3, 33, 24, 0, 13, 0, 0, 
    19, 54, 0, 0, 66, 29, 24, 9, 0, 68, 23, 1, 21, 9, 0, 
    18, 39, 9, 0, 38, 42, 50, 20, 4, 73, 18, 3, 12, 23, 6, 
    28, 46, 6, 7, 25, 75, 23, 25, 9, 51, 22, 2, 23, 22, 5, 
    40, 60, 2, 43, 4, 25, 12, 15, 28, 3, 24, 0, 9, 15, 4, 
    56, 58, 14, 49, 20, 8, 32, 35, 10, 22, 2, 2, 21, 18, 0, 
    78, 52, 16, 87, 36, 25, 64, 58, 20, 3, 13, 23, 30, 36, 24, 
    77, 74, 44, 99, 42, 23, 33, 31, 28, 32, 38, 40, 44, 45, 42, 
    40, 63, 72, 72, 14, 36, 34, 33, 33, 37, 43, 47, 49, 50, 56, 
    44, 42, 79, 60, 30, 41, 33, 33, 38, 42, 44, 50, 45, 58, 52, 
    41, 46, 39, 47, 29, 40, 44, 40, 42, 43, 38, 43, 62, 55, 33, 
    
    -- channel=106
    59, 62, 59, 62, 61, 57, 65, 69, 65, 60, 55, 51, 51, 58, 57, 
    59, 64, 61, 66, 57, 33, 72, 65, 59, 16, 16, 26, 31, 42, 54, 
    64, 40, 63, 66, 61, 54, 58, 36, 14, 0, 19, 12, 27, 24, 35, 
    55, 0, 63, 60, 64, 27, 26, 23, 12, 0, 37, 22, 23, 24, 8, 
    35, 0, 72, 17, 21, 27, 43, 31, 23, 0, 19, 39, 8, 24, 15, 
    32, 2, 76, 50, 0, 34, 34, 30, 34, 0, 47, 43, 5, 17, 16, 
    27, 23, 48, 77, 0, 0, 33, 30, 42, 0, 46, 28, 3, 0, 24, 
    23, 16, 29, 46, 4, 0, 58, 26, 32, 0, 31, 34, 0, 16, 34, 
    21, 0, 46, 0, 34, 20, 29, 15, 0, 36, 20, 47, 3, 10, 38, 
    9, 0, 46, 0, 40, 21, 0, 13, 23, 37, 41, 10, 0, 25, 59, 
    0, 8, 45, 0, 23, 13, 0, 22, 37, 14, 0, 0, 0, 0, 2, 
    0, 0, 14, 0, 66, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    3, 1, 1, 5, 5, 0, 4, 5, 5, 4, 4, 0, 2, 8, 8, 
    4, 1, 0, 6, 0, 0, 29, 3, 7, 0, 11, 10, 0, 0, 6, 
    6, 0, 2, 5, 0, 0, 26, 14, 1, 0, 17, 16, 27, 0, 0, 
    62, 0, 10, 0, 7, 0, 8, 21, 7, 0, 34, 4, 22, 21, 0, 
    71, 0, 41, 0, 5, 19, 34, 29, 12, 0, 16, 45, 0, 30, 0, 
    58, 0, 54, 0, 0, 18, 27, 32, 38, 0, 45, 50, 0, 19, 25, 
    65, 9, 22, 30, 0, 0, 7, 32, 46, 0, 57, 35, 0, 0, 26, 
    46, 22, 44, 25, 0, 0, 53, 5, 30, 0, 28, 38, 0, 0, 21, 
    39, 0, 75, 0, 21, 0, 22, 0, 0, 14, 0, 38, 0, 0, 0, 
    2, 0, 72, 0, 44, 10, 0, 13, 19, 4, 32, 6, 0, 0, 13, 
    0, 4, 65, 0, 75, 36, 0, 9, 54, 26, 3, 0, 0, 0, 7, 
    0, 0, 38, 0, 62, 42, 0, 0, 11, 0, 0, 0, 0, 0, 7, 
    17, 0, 0, 0, 88, 3, 5, 2, 3, 0, 0, 0, 0, 0, 0, 
    22, 1, 0, 30, 25, 0, 13, 4, 0, 0, 0, 0, 5, 0, 7, 
    27, 0, 0, 0, 9, 0, 0, 4, 0, 1, 11, 0, 0, 12, 43, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=111
    2, 1, 0, 0, 0, 0, 0, 1, 0, 5, 15, 12, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 4, 12, 0, 
    9, 39, 0, 0, 0, 36, 12, 5, 0, 0, 0, 0, 0, 11, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 6, 3, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 53, 21, 0, 0, 0, 0, 0, 6, 1, 0, 0, 
    0, 0, 22, 0, 17, 0, 8, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 23, 25, 4, 1, 6, 0, 3, 8, 7, 
    0, 0, 0, 0, 0, 45, 3, 0, 0, 0, 15, 31, 11, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 34, 31, 8, 0, 0, 1, 
    6, 0, 0, 0, 0, 0, 0, 33, 11, 0, 0, 0, 0, 2, 0, 
    48, 29, 0, 0, 42, 44, 22, 20, 7, 0, 0, 0, 0, 0, 0, 
    0, 32, 11, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 28, 45, 6, 0, 0, 0, 0, 0, 0, 6, 0, 0, 22, 
    0, 0, 0, 40, 8, 12, 18, 1, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=112
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 17, 0, 0, 0, 0, 0, 0, 
    17, 8, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 
    4, 0, 0, 0, 0, 2, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 24, 26, 8, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 3, 15, 0, 0, 0, 
    0, 0, 0, 0, 10, 7, 0, 0, 0, 34, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 36, 25, 0, 0, 0, 0, 0, 0, 
    31, 6, 0, 0, 38, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 7, 4, 0, 
    0, 0, 23, 27, 2, 0, 0, 0, 0, 0, 0, 4, 0, 0, 28, 
    2, 0, 0, 4, 2, 6, 14, 2, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=113
    8, 6, 11, 7, 9, 7, 11, 14, 9, 0, 0, 3, 7, 10, 11, 
    12, 14, 12, 6, 9, 0, 0, 0, 0, 0, 0, 0, 3, 7, 6, 
    0, 10, 11, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 
    0, 23, 6, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 16, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 12, 0, 0, 6, 8, 0, 0, 0, 0, 0, 3, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 56, 34, 0, 0, 0, 7, 21, 28, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 15, 22, 23, 19, 
    35, 0, 0, 0, 0, 15, 15, 14, 18, 23, 28, 30, 16, 11, 32, 
    29, 25, 0, 0, 0, 17, 27, 19, 14, 19, 21, 11, 21, 29, 3, 
    32, 26, 17, 0, 6, 0, 0, 9, 24, 33, 28, 23, 36, 46, 34, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 9, 6, 4, 9, 6, 0, 
    0, 15, 0, 0, 0, 3, 0, 0, 7, 41, 10, 12, 0, 11, 11, 
    0, 43, 0, 0, 0, 8, 2, 0, 8, 48, 0, 11, 0, 0, 33, 
    0, 48, 0, 28, 20, 24, 2, 0, 0, 59, 16, 0, 10, 0, 18, 
    8, 43, 0, 0, 56, 29, 9, 1, 0, 91, 2, 0, 18, 2, 5, 
    14, 20, 14, 0, 44, 46, 17, 8, 0, 84, 0, 0, 17, 21, 4, 
    24, 21, 15, 0, 29, 53, 0, 16, 0, 55, 7, 0, 24, 18, 7, 
    23, 45, 0, 41, 2, 27, 7, 6, 32, 4, 12, 0, 18, 24, 10, 
    31, 42, 0, 60, 0, 16, 39, 14, 15, 2, 0, 5, 35, 26, 0, 
    62, 39, 0, 98, 9, 13, 52, 24, 0, 0, 14, 24, 31, 24, 7, 
    62, 59, 26, 90, 0, 4, 28, 26, 19, 21, 26, 30, 33, 34, 27, 
    27, 60, 78, 31, 0, 27, 25, 26, 23, 27, 33, 35, 33, 34, 42, 
    23, 36, 89, 0, 8, 32, 23, 26, 30, 31, 32, 32, 30, 43, 28, 
    20, 35, 41, 19, 14, 30, 28, 28, 34, 33, 24, 33, 53, 29, 12, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 7, 0, 
    6, 27, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 5, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 15, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 19, 9, 0, 0, 0, 7, 0, 0, 3, 0, 0, 
    0, 0, 8, 0, 5, 0, 11, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 40, 10, 4, 0, 1, 0, 0, 2, 9, 0, 
    0, 0, 0, 2, 0, 2, 0, 0, 4, 0, 6, 5, 0, 0, 0, 
    0, 0, 0, 0, 6, 4, 0, 0, 0, 35, 11, 1, 8, 0, 0, 
    1, 0, 0, 0, 0, 0, 31, 36, 20, 0, 0, 0, 0, 0, 0, 
    35, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 
    0, 0, 36, 14, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 13, 
    0, 0, 0, 2, 0, 5, 16, 4, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=118
    12, 13, 7, 7, 7, 7, 10, 12, 8, 15, 23, 19, 11, 7, 9, 
    5, 6, 5, 9, 4, 0, 0, 14, 38, 3, 0, 0, 13, 17, 8, 
    27, 35, 9, 10, 9, 41, 38, 22, 0, 0, 0, 0, 0, 11, 12, 
    0, 0, 7, 5, 6, 0, 0, 0, 0, 0, 14, 12, 20, 7, 7, 
    0, 0, 4, 0, 0, 0, 4, 2, 15, 0, 0, 0, 0, 0, 0, 
    7, 0, 11, 21, 55, 24, 0, 0, 0, 0, 11, 25, 0, 0, 0, 
    0, 11, 29, 22, 6, 0, 14, 1, 9, 0, 23, 1, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 37, 31, 21, 0, 24, 14, 0, 10, 12, 
    0, 0, 9, 0, 0, 43, 20, 0, 0, 7, 29, 47, 16, 1, 0, 
    19, 0, 17, 0, 5, 0, 0, 0, 0, 38, 42, 11, 0, 0, 10, 
    6, 0, 24, 0, 0, 0, 0, 31, 20, 0, 0, 0, 0, 2, 9, 
    25, 23, 0, 0, 75, 70, 33, 32, 16, 0, 0, 0, 0, 0, 0, 
    0, 16, 0, 16, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 74, 17, 0, 0, 0, 0, 0, 0, 5, 1, 0, 22, 
    0, 0, 2, 42, 13, 11, 13, 0, 0, 0, 0, 0, 0, 0, 3, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 11, 0, 10, 0, 5, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 30, 15, 0, 0, 5, 11, 15, 0, 0, 
    51, 0, 0, 0, 1, 0, 0, 11, 0, 0, 29, 0, 22, 12, 0, 
    65, 0, 21, 0, 0, 0, 22, 21, 7, 0, 3, 30, 0, 24, 0, 
    42, 0, 34, 0, 0, 15, 22, 21, 29, 0, 30, 47, 0, 15, 13, 
    48, 0, 10, 29, 0, 0, 0, 25, 39, 0, 50, 25, 0, 0, 12, 
    28, 18, 19, 17, 0, 0, 48, 2, 29, 0, 27, 29, 0, 0, 14, 
    28, 0, 58, 0, 2, 0, 18, 0, 0, 0, 0, 42, 0, 0, 0, 
    3, 0, 64, 0, 26, 0, 0, 1, 0, 6, 37, 7, 0, 0, 5, 
    0, 0, 58, 0, 60, 6, 0, 7, 50, 24, 0, 0, 0, 0, 8, 
    0, 0, 28, 0, 52, 53, 0, 0, 13, 0, 0, 0, 0, 0, 1, 
    5, 0, 0, 0, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 42, 28, 0, 6, 0, 0, 0, 0, 0, 3, 0, 0, 
    18, 0, 0, 0, 6, 0, 0, 1, 0, 0, 2, 0, 0, 0, 36, 
    
    -- channel=120
    24, 24, 28, 27, 27, 25, 26, 30, 30, 21, 13, 18, 21, 21, 23, 
    29, 29, 30, 26, 33, 31, 18, 19, 6, 16, 1, 0, 4, 19, 23, 
    1, 22, 29, 28, 30, 4, 0, 0, 14, 14, 0, 0, 0, 6, 19, 
    0, 31, 22, 34, 18, 29, 5, 0, 0, 14, 0, 0, 0, 0, 23, 
    0, 5, 7, 59, 15, 6, 0, 0, 0, 32, 0, 0, 0, 0, 8, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 53, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 11, 17, 0, 0, 0, 26, 0, 0, 0, 5, 0, 
    0, 0, 0, 3, 29, 8, 0, 0, 0, 13, 0, 0, 2, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 9, 21, 
    0, 0, 0, 1, 0, 1, 13, 0, 0, 0, 0, 0, 11, 23, 16, 
    0, 0, 0, 42, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 11, 12, 
    21, 0, 0, 0, 0, 17, 27, 26, 14, 6, 3, 5, 4, 4, 3, 
    4, 18, 0, 0, 0, 0, 0, 3, 5, 5, 3, 1, 0, 0, 0, 
    6, 9, 12, 0, 0, 0, 0, 5, 1, 1, 5, 9, 6, 7, 3, 
    0, 5, 11, 29, 11, 13, 2, 0, 0, 0, 4, 5, 0, 0, 1, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 9, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 8, 0, 2, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 0, 0, 0, 0, 14, 
    6, 0, 0, 0, 4, 0, 0, 0, 0, 6, 0, 0, 4, 0, 1, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 8, 2, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 2, 0, 9, 0, 13, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 9, 0, 0, 13, 6, 0, 0, 
    4, 0, 0, 4, 0, 0, 0, 0, 0, 5, 23, 16, 26, 26, 22, 
    56, 10, 0, 0, 0, 40, 47, 46, 40, 36, 38, 41, 41, 43, 41, 
    50, 54, 16, 0, 20, 34, 35, 36, 38, 40, 42, 42, 41, 42, 42, 
    50, 49, 55, 0, 25, 37, 35, 38, 37, 40, 46, 50, 47, 51, 50, 
    44, 49, 50, 47, 43, 47, 40, 33, 32, 36, 42, 46, 39, 38, 44, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=125
    28, 29, 30, 29, 30, 30, 33, 37, 36, 34, 32, 33, 30, 26, 26, 
    33, 35, 33, 31, 31, 16, 25, 37, 32, 15, 0, 2, 21, 33, 27, 
    27, 48, 34, 33, 33, 24, 11, 13, 4, 0, 0, 0, 0, 14, 27, 
    0, 16, 30, 38, 29, 25, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 9, 36, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 17, 16, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    0, 2, 5, 5, 4, 2, 3, 1, 4, 4, 3, 4, 7, 1, 2, 
    4, 2, 5, 5, 7, 33, 7, 9, 0, 4, 9, 0, 0, 0, 7, 
    2, 0, 3, 2, 0, 0, 0, 0, 0, 10, 3, 11, 4, 0, 4, 
    6, 5, 0, 5, 11, 7, 17, 13, 5, 0, 8, 0, 0, 0, 0, 
    25, 21, 7, 20, 75, 38, 3, 6, 0, 0, 3, 8, 5, 10, 0, 
    0, 4, 9, 0, 0, 0, 17, 3, 5, 20, 9, 0, 0, 10, 10, 
    4, 0, 0, 9, 0, 16, 9, 19, 2, 3, 0, 0, 0, 3, 5, 
    9, 9, 2, 13, 2, 20, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 3, 2, 8, 6, 0, 0, 0, 6, 0, 0, 0, 0, 0, 6, 
    2, 0, 7, 0, 0, 13, 8, 22, 0, 3, 0, 0, 11, 14, 6, 
    0, 0, 0, 23, 76, 41, 41, 18, 27, 8, 5, 29, 13, 0, 1, 
    0, 4, 19, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 9, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 7, 1, 0, 0, 11, 5, 0, 
    
    -- channel=127
    4, 2, 0, 0, 0, 0, 1, 1, 0, 7, 15, 11, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 28, 0, 0, 0, 14, 8, 0, 
    24, 25, 0, 0, 1, 35, 25, 16, 0, 0, 0, 0, 0, 11, 4, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 8, 9, 3, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 8, 
    1, 0, 0, 26, 42, 12, 0, 0, 0, 0, 4, 12, 0, 0, 0, 
    0, 5, 15, 6, 8, 0, 1, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 30, 26, 5, 0, 9, 5, 0, 7, 0, 
    0, 0, 2, 0, 0, 35, 6, 0, 0, 9, 19, 37, 15, 0, 0, 
    6, 0, 0, 0, 0, 4, 0, 0, 0, 28, 32, 4, 0, 0, 2, 
    0, 0, 7, 0, 0, 0, 0, 22, 7, 0, 0, 0, 0, 11, 13, 
    35, 16, 0, 0, 59, 54, 33, 31, 12, 2, 0, 0, 0, 0, 0, 
    0, 26, 0, 16, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 54, 8, 0, 0, 0, 0, 0, 0, 5, 0, 0, 25, 
    0, 0, 8, 35, 13, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
