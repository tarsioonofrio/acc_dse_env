-gN_BRAM_IWGHT=10 -gN_BRAM_IFMAP=2 -gN_BRAM_GOLD=2