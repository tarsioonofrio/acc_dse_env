-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(36-1 downto 0);
        ADDR : in std_logic_vector(9-1 downto 0);
        DO   : out std_logic_vector(36-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(8-1 downto 0);
    signal bram_addr     : std_logic_vector(9-1 downto 0);
    signal bram_di     : std_logic_vector(44-1 downto 0);
    signal bram_do     : std_logic_vector(44-1 downto 0);
    constant bram_par     : std_logic_vector(8-1 downto 0) := "00000000";

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(9-1 downto 0);
    bram_di <= bram_par & DI;
    DO <= bram_do(36-1 downto 0);


    MEM_IWGHT_LAYER0_INSTANCE0 : if BRAM_NAME = "iwght_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffd761ffffffffffffaecbffffffff00001d4000000000ffffca09ffffffff",
            INIT_01 => X"0000271300000000000000cb00000000000001f0000000000000181a00000000",
            INIT_02 => X"fffffafaffffffffffffe634ffffffff000000f300000000fffff3ffffffffff",
            INIT_03 => X"ffffe432ffffffffffffe2e4ffffffff00000bc1000000000000036000000000",
            INIT_04 => X"0000002300000000fffffff0ffffffff00000019000000000000003f00000000",
            INIT_05 => X"ffffffddffffffff0000001200000000fffffff8ffffffff0000001c00000000",
            INIT_06 => X"0000001600000000fffffff7ffffffff0000000d000000000000000900000000",
            INIT_07 => X"ffffffdbfffffffffffffff3fffffffffffffffcffffffff0000000300000000",
            INIT_08 => X"00000048000000000000004700000000ffffffefffffffffffffffcaffffffff",
            INIT_09 => X"0000002c00000000ffffffe4ffffffff0000002b000000000000004400000000",
            INIT_0A => X"0000000900000000ffffffe0ffffffffffffffdbffffffffffffffeaffffffff",
            INIT_0B => X"fffffffbffffffff0000001d000000000000003100000000ffffffe7ffffffff",
            INIT_0C => X"0000000300000000fffffffaffffffff00000033000000000000003d00000000",
            INIT_0D => X"000000110000000000000000000000000000000700000000ffffffeaffffffff",
            INIT_0E => X"fffffffcffffffff000000050000000000000034000000000000000900000000",
            INIT_0F => X"ffffffd4ffffffff0000000e00000000ffffffd6ffffffff0000002100000000",
            INIT_10 => X"ffffffbbfffffffffffffff6ffffffffffffffd0ffffffffffffffbfffffffff",
            INIT_11 => X"0000001f000000000000000d00000000ffffffdfffffffff0000001100000000",
            INIT_12 => X"ffffffdbffffffff0000002100000000ffffffceffffffff0000000200000000",
            INIT_13 => X"0000002100000000ffffffe5ffffffffffffffdcffffffff0000002000000000",
            INIT_14 => X"ffffffeaffffffffffffffd3ffffffffffffffd8ffffffff0000002000000000",
            INIT_15 => X"00000012000000000000000d00000000ffffffdbffffffff0000000000000000",
            INIT_16 => X"00000032000000000000001c00000000fffffff9ffffffff0000001000000000",
            INIT_17 => X"0000001700000000000000350000000000000035000000000000002b00000000",
            INIT_18 => X"ffffffe9ffffffffffffffefffffffffffffffebffffffff0000000a00000000",
            INIT_19 => X"ffffffecffffffffffffffdcffffffff00000009000000000000001e00000000",
            INIT_1A => X"0000001900000000000000230000000000000020000000000000001d00000000",
            INIT_1B => X"0000001f00000000ffffffdefffffffffffffff5fffffffffffffff4ffffffff",
            INIT_1C => X"0000002a00000000fffffffbffffffff0000000600000000fffffff1ffffffff",
            INIT_1D => X"0000002c00000000000000400000000000000030000000000000003100000000",
            INIT_1E => X"0000001b000000000000003300000000ffffffe7ffffffff0000003500000000",
            INIT_1F => X"0000002f00000000ffffffffffffffff00000013000000000000001b00000000",
            INIT_20 => X"ffffffd7ffffffffffffffe9ffffffffffffffe3ffffffff0000000c00000000",
            INIT_21 => X"0000001c0000000000000039000000000000004300000000ffffffcfffffffff",
            INIT_22 => X"0000001400000000fffffffdffffffff00000027000000000000003400000000",
            INIT_23 => X"fffffffbffffffff0000001f000000000000002b000000000000003800000000",
            INIT_24 => X"ffffffd6ffffffffffffffc3ffffffffffffffe3ffffffff0000000c00000000",
            INIT_25 => X"0000001a00000000ffffffbeffffffffffffffc4ffffffffffffffc5ffffffff",
            INIT_26 => X"0000002100000000fffffff2ffffffff00000013000000000000003300000000",
            INIT_27 => X"fffffff0fffffffffffffffeffffffffffffffb8ffffffffffffffecffffffff",
            INIT_28 => X"0000000f00000000ffffffe4ffffffff0000002d000000000000003900000000",
            INIT_29 => X"ffffffb0ffffffffffffffdfffffffff00000028000000000000000400000000",
            INIT_2A => X"fffffff4ffffffff0000003800000000ffffffecffffffffffffffc3ffffffff",
            INIT_2B => X"ffffffebffffffff00000002000000000000003400000000fffffffaffffffff",
            INIT_2C => X"0000000e00000000ffffffdcffffffff0000000100000000ffffffc6ffffffff",
            INIT_2D => X"00000024000000000000001400000000ffffffbcffffffff0000001600000000",
            INIT_2E => X"fffffff4ffffffff00000024000000000000001800000000ffffffc0ffffffff",
            INIT_2F => X"ffffffffffffffffffffffe4ffffffff0000004900000000ffffffd1ffffffff",
            INIT_30 => X"00000016000000000000001700000000ffffffb6ffffffff0000004800000000",
            INIT_31 => X"ffffffcfffffffff0000004c00000000ffffffe8ffffffffffffffcbffffffff",
            INIT_32 => X"ffffffdcffffffffffffffacffffffff0000002c000000000000000a00000000",
            INIT_33 => X"ffffffc8ffffffffffffffebffffffffffffffddffffffff0000005b00000000",
            INIT_34 => X"ffffffe3ffffffffffffffddffffffffffffffe0ffffffffffffffdeffffffff",
            INIT_35 => X"ffffffd0ffffffffffffffe0ffffffffffffffeffffffffffffffff7ffffffff",
            INIT_36 => X"0000000d00000000ffffffd9fffffffffffffffeffffffffffffffe2ffffffff",
            INIT_37 => X"fffffff7ffffffff000000080000000000000020000000000000000600000000",
            INIT_38 => X"fffffffdffffffff0000004800000000ffffffe8ffffffff0000003900000000",
            INIT_39 => X"0000003d0000000000000047000000000000002c000000000000004000000000",
            INIT_3A => X"00000006000000000000000000000000ffffffefffffffffffffffccffffffff",
            INIT_3B => X"ffffffe7ffffffffffffffe4ffffffff00000005000000000000000500000000",
            INIT_3C => X"0000000400000000fffffffdffffffffffffffe7fffffffffffffff3ffffffff",
            INIT_3D => X"fffffffcffffffff00000015000000000000001a00000000ffffffddffffffff",
            INIT_3E => X"ffffffd5ffffffff0000001b00000000ffffffd6ffffffff0000000700000000",
            INIT_3F => X"ffffffe6ffffffff0000001a00000000ffffffd5ffffffffffffffd9ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdcffffffffffffffe4fffffffffffffffbffffffffffffffccffffffff",
            INIT_41 => X"0000001000000000ffffffceffffffffffffffe4ffffffffffffffd4ffffffff",
            INIT_42 => X"0000002700000000fffffffcffffffff0000000400000000ffffffd3ffffffff",
            INIT_43 => X"fffffffaffffffff0000001600000000ffffffddfffffffffffffffbffffffff",
            INIT_44 => X"00000032000000000000002d0000000000000035000000000000000700000000",
            INIT_45 => X"fffffffeffffffffffffffd6ffffffffffffffcdffffffff0000003200000000",
            INIT_46 => X"000000180000000000000000000000000000002800000000fffffff7ffffffff",
            INIT_47 => X"0000002f00000000ffffffe1ffffffff00000049000000000000000c00000000",
            INIT_48 => X"0000001d000000000000002b0000000000000029000000000000000600000000",
            INIT_49 => X"00000010000000000000002c00000000ffffffe8ffffffff0000003a00000000",
            INIT_4A => X"fffffff9ffffffff000000170000000000000017000000000000001700000000",
            INIT_4B => X"0000000a00000000000000270000000000000010000000000000000900000000",
            INIT_4C => X"ffffffe1fffffffffffffff1ffffffffffffffe4ffffffffffffffe9ffffffff",
            INIT_4D => X"fffffffcffffffff0000000900000000ffffffd9ffffffffffffffb8ffffffff",
            INIT_4E => X"00000050000000000000002a000000000000000400000000ffffffc4ffffffff",
            INIT_4F => X"ffffffe4ffffffff0000000300000000ffffffe3ffffffffffffffe8ffffffff",
            INIT_50 => X"0000004e00000000ffffffffffffffff0000001900000000ffffffb8ffffffff",
            INIT_51 => X"ffffffeeffffffff00000023000000000000000a000000000000002100000000",
            INIT_52 => X"0000001300000000ffffffc1ffffffffffffffb6ffffffffffffffd6ffffffff",
            INIT_53 => X"fffffff7fffffffffffffff3ffffffff00000036000000000000003d00000000",
            INIT_54 => X"ffffffe0ffffffffffffffe9ffffffffffffffffffffffffffffffefffffffff",
            INIT_55 => X"00000053000000000000001c00000000ffffffe8fffffffffffffff0ffffffff",
            INIT_56 => X"00000030000000000000001100000000ffffffceffffffff0000001a00000000",
            INIT_57 => X"fffffff5ffffffffffffffccffffffff0000004600000000ffffffbaffffffff",
            INIT_58 => X"0000005500000000ffffffb3ffffffff00000003000000000000000300000000",
            INIT_59 => X"ffffffc6ffffffff0000002900000000ffffffbdffffffffffffffe6ffffffff",
            INIT_5A => X"fffffffcffffffffffffffd1ffffffff0000004f000000000000001900000000",
            INIT_5B => X"fffffffcffffffffffffffbbfffffffffffffff4ffffffff0000004000000000",
            INIT_5C => X"00000038000000000000002e0000000000000002000000000000003500000000",
            INIT_5D => X"0000003a0000000000000037000000000000003f000000000000003500000000",
            INIT_5E => X"ffffffcfffffffffffffffd1ffffffffffffffd7ffffffffffffffd4ffffffff",
            INIT_5F => X"ffffffd1fffffffffffffff4fffffffffffffffdffffffffffffffd9ffffffff",
            INIT_60 => X"0000000a00000000fffffffaffffffff0000001c00000000ffffffe3ffffffff",
            INIT_61 => X"ffffffdeffffffffffffffceffffffffffffffe9ffffffff0000001900000000",
            INIT_62 => X"0000001a00000000ffffffe7ffffffffffffffe5ffffffff0000003100000000",
            INIT_63 => X"0000000c00000000ffffffffffffffffffffffebffffffffffffffd3ffffffff",
            INIT_64 => X"fffffffcfffffffffffffffdffffffffffffffe0fffffffffffffff0ffffffff",
            INIT_65 => X"0000001800000000000000110000000000000018000000000000000d00000000",
            INIT_66 => X"0000001a000000000000002500000000ffffffe5ffffffff0000000300000000",
            INIT_67 => X"000000120000000000000044000000000000000b000000000000003200000000",
            INIT_68 => X"fffffff9ffffffffffffffeaffffffff0000000b000000000000000c00000000",
            INIT_69 => X"0000004600000000fffffff4ffffffff00000030000000000000001a00000000",
            INIT_6A => X"0000000d000000000000004f000000000000003c000000000000000300000000",
            INIT_6B => X"0000000300000000000000040000000000000017000000000000002500000000",
            INIT_6C => X"ffffffd6ffffffffffffffc5ffffffff0000001400000000ffffffccffffffff",
            INIT_6D => X"ffffffd6fffffffffffffff1fffffffffffffff3ffffffffffffffe0ffffffff",
            INIT_6E => X"ffffffd8fffffffffffffff4ffffffff0000000e00000000ffffffffffffffff",
            INIT_6F => X"0000000300000000ffffffc2ffffffff0000000400000000ffffffc6ffffffff",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE0 : if BRAM_NAME = "iwght_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000034400000000000000ced000000000000482b00000000fffff3e3ffffffff",
            INIT_01 => X"fffffc9effffffffffffea15ffffffff0000009b0000000000000f9c00000000",
            INIT_02 => X"fffff35ffffffffffffff7b9ffffffff00001cf800000000000013b300000000",
            INIT_03 => X"000009ee00000000fffffbeefffffffffffffb69ffffffff0000117d00000000",
            INIT_04 => X"000004c70000000000001bfb0000000000001c1d000000000000296600000000",
            INIT_05 => X"00000dbc0000000000000f6400000000ffffe3caffffffff000021c300000000",
            INIT_06 => X"ffffeca2ffffffff0000172600000000fffff3dfffffffff000007e700000000",
            INIT_07 => X"00003b1c0000000000001bb100000000ffffe0d7ffffffff00002d8600000000",
            INIT_08 => X"0000000e000000000000003a000000000000002f000000000000001b00000000",
            INIT_09 => X"0000000100000000fffffffeffffffff0000001600000000fffffff9ffffffff",
            INIT_0A => X"0000000b00000000ffffffc1ffffffffffffffd6fffffffffffffffbffffffff",
            INIT_0B => X"ffffffccfffffffffffffffcffffffffffffffffffffffff0000000800000000",
            INIT_0C => X"000000430000000000000012000000000000000100000000ffffffe8ffffffff",
            INIT_0D => X"00000007000000000000000f0000000000000008000000000000002c00000000",
            INIT_0E => X"00000020000000000000000a0000000000000032000000000000000800000000",
            INIT_0F => X"00000017000000000000001d0000000000000027000000000000002800000000",
            INIT_10 => X"ffffffe9ffffffff00000023000000000000002700000000fffffff8ffffffff",
            INIT_11 => X"ffffffeeffffffff0000002d00000000fffffffffffffffffffffff7ffffffff",
            INIT_12 => X"fffffff2ffffffffffffffd8ffffffff00000003000000000000001e00000000",
            INIT_13 => X"ffffffe5ffffffff0000000800000000ffffffffffffffffffffffe1ffffffff",
            INIT_14 => X"ffffffddffffffffffffffd0ffffffffffffffe7ffffffff0000000400000000",
            INIT_15 => X"ffffffe2ffffffff00000014000000000000001300000000ffffffe8ffffffff",
            INIT_16 => X"ffffffd2fffffffffffffff5ffffffffffffffe0fffffffffffffff6ffffffff",
            INIT_17 => X"fffffff4fffffffffffffffeffffffff0000000200000000fffffff2ffffffff",
            INIT_18 => X"ffffffc6ffffffffffffffe5ffffffffffffffb8ffffffffffffffddffffffff",
            INIT_19 => X"ffffffeeffffffff0000000b00000000fffffff8ffffffffffffffd6ffffffff",
            INIT_1A => X"fffffff4ffffffff0000001b00000000ffffffffffffffff0000000f00000000",
            INIT_1B => X"0000000e00000000ffffffe8ffffffffffffffeffffffffffffffff8ffffffff",
            INIT_1C => X"00000007000000000000000b00000000fffffff7fffffffffffffff5ffffffff",
            INIT_1D => X"0000000a00000000ffffffffffffffffffffffd5ffffffffffffffecffffffff",
            INIT_1E => X"0000000d000000000000001700000000ffffffcaffffffff0000000400000000",
            INIT_1F => X"0000002200000000fffffff8fffffffffffffff7ffffffff0000001700000000",
            INIT_20 => X"0000000500000000ffffffe0fffffffffffffff0ffffffff0000000200000000",
            INIT_21 => X"00000003000000000000001f000000000000000800000000ffffffecffffffff",
            INIT_22 => X"fffffff7ffffffff0000000800000000fffffff2ffffffffffffffdaffffffff",
            INIT_23 => X"0000002d00000000ffffffe0ffffffff0000001e000000000000001400000000",
            INIT_24 => X"0000006f000000000000003100000000ffffffcfffffffff0000001100000000",
            INIT_25 => X"ffffffeaffffffff00000008000000000000000000000000ffffffe2ffffffff",
            INIT_26 => X"fffffffffffffffffffffff6ffffffff0000001f000000000000001400000000",
            INIT_27 => X"0000001d0000000000000024000000000000000600000000ffffffefffffffff",
            INIT_28 => X"ffffffddffffffffffffffe8ffffffff00000007000000000000001700000000",
            INIT_29 => X"0000000100000000fffffff3ffffffff00000014000000000000001600000000",
            INIT_2A => X"fffffff7ffffffff0000000f000000000000000600000000ffffffe5ffffffff",
            INIT_2B => X"0000004800000000000000460000000000000022000000000000001f00000000",
            INIT_2C => X"000000000000000000000016000000000000000b000000000000003900000000",
            INIT_2D => X"ffffffb4ffffffffffffff96ffffffffffffffe9ffffffff0000000a00000000",
            INIT_2E => X"0000001a00000000fffffff8ffffffff0000001200000000ffffffbbffffffff",
            INIT_2F => X"0000001a0000000000000027000000000000001b000000000000001600000000",
            INIT_30 => X"00000031000000000000001c0000000000000029000000000000002a00000000",
            INIT_31 => X"ffffffedffffffffffffffecffffffffffffffecffffffff0000000000000000",
            INIT_32 => X"00000004000000000000000700000000ffffffe5ffffffffffffffeaffffffff",
            INIT_33 => X"ffffffeeffffffffffffffc9fffffffffffffff7fffffffffffffff0ffffffff",
            INIT_34 => X"ffffffd8ffffffffffffffbcffffffffffffffcbffffffffffffffe1ffffffff",
            INIT_35 => X"ffffffedffffffff000000070000000000000031000000000000003900000000",
            INIT_36 => X"ffffffdeffffffffffffffdeffffffff0000000b000000000000000000000000",
            INIT_37 => X"0000002d0000000000000022000000000000004300000000ffffffe9ffffffff",
            INIT_38 => X"ffffffe5fffffffffffffff7ffffffff00000025000000000000004a00000000",
            INIT_39 => X"ffffffb0ffffffffffffffb5ffffffffffffffc0ffffffffffffffcdffffffff",
            INIT_3A => X"ffffffccffffffffffffff9fffffffffffffff83ffffffff0000001e00000000",
            INIT_3B => X"0000002900000000ffffffd1ffffffffffffff85ffffffffffffff61ffffffff",
            INIT_3C => X"0000006a000000000000004b000000000000000e000000000000000d00000000",
            INIT_3D => X"0000003f000000000000002c0000000000000043000000000000007c00000000",
            INIT_3E => X"ffffffecffffffffffffffe9fffffffffffffff4ffffffff0000001b00000000",
            INIT_3F => X"ffffffecfffffffffffffff6ffffffff0000001b000000000000002100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff2ffffffffffffffcaffffffffffffffdefffffffffffffffdffffffff",
            INIT_41 => X"ffffffd4ffffffff0000001a00000000ffffffe6ffffffffffffffdbffffffff",
            INIT_42 => X"ffffffedffffffffffffffe7fffffffffffffff5ffffffffffffffd9ffffffff",
            INIT_43 => X"ffffffefffffffffffffffd1ffffffff0000001400000000fffffff9ffffffff",
            INIT_44 => X"0000003900000000ffffffecffffffff0000000500000000ffffffe6ffffffff",
            INIT_45 => X"000000450000000000000061000000000000005a000000000000001400000000",
            INIT_46 => X"ffffffabffffffffffffffdfffffffffffffffe1ffffffff0000000d00000000",
            INIT_47 => X"000000270000000000000015000000000000000c000000000000002e00000000",
            INIT_48 => X"ffffffadffffffffffffffe1ffffffffffffff86ffffffffffffffefffffffff",
            INIT_49 => X"ffffffcafffffffffffffffdfffffffffffffffdffffffffffffff8cffffffff",
            INIT_4A => X"0000000e0000000000000026000000000000000b000000000000001700000000",
            INIT_4B => X"ffffffe4ffffffff0000001a00000000ffffffe3fffffffffffffff8ffffffff",
            INIT_4C => X"ffffffecffffffffffffffc3ffffffffffffffd4ffffffff0000000300000000",
            INIT_4D => X"fffffff7fffffffffffffff0ffffffffffffffbfffffffffffffffc9ffffffff",
            INIT_4E => X"fffffffdffffffffffffffdaffffffffffffffd0ffffffffffffffb8ffffffff",
            INIT_4F => X"fffffffeffffffff00000023000000000000003200000000ffffffeaffffffff",
            INIT_50 => X"0000001000000000ffffffd8ffffffffffffffc3ffffffffffffffe5ffffffff",
            INIT_51 => X"00000037000000000000000000000000ffffffd1ffffffffffffffc2ffffffff",
            INIT_52 => X"fffffff4ffffffffffffffd4ffffffffffffffe2ffffffff0000002200000000",
            INIT_53 => X"0000002100000000fffffff4ffffffffffffffeeffffffff0000001f00000000",
            INIT_54 => X"fffffff2ffffffffffffffc8ffffffff00000037000000000000004e00000000",
            INIT_55 => X"fffffff2ffffffffffffffe6fffffffffffffff3ffffffffffffffdfffffffff",
            INIT_56 => X"ffffffc5ffffffff000000100000000000000022000000000000001400000000",
            INIT_57 => X"fffffffefffffffffffffff7fffffffffffffff8ffffffffffffffd6ffffffff",
            INIT_58 => X"00000025000000000000001f00000000fffffffdffffffff0000000600000000",
            INIT_59 => X"ffffffe7ffffffff00000011000000000000001500000000ffffffeaffffffff",
            INIT_5A => X"0000001f000000000000003400000000ffffffb9ffffffffffffffd1ffffffff",
            INIT_5B => X"0000001a00000000000000330000000000000006000000000000000f00000000",
            INIT_5C => X"0000000b00000000000000160000000000000014000000000000006d00000000",
            INIT_5D => X"0000003100000000fffffff4ffffffff0000000f000000000000003500000000",
            INIT_5E => X"ffffffc6ffffffffffffff9affffffffffffffd4ffffffff0000003100000000",
            INIT_5F => X"fffffffaffffffffffffff95ffffffffffffffa0ffffffffffffffdfffffffff",
            INIT_60 => X"0000001000000000fffffff1fffffffffffffff2fffffffffffffffcffffffff",
            INIT_61 => X"ffffffdfffffffffffffffecffffffffffffffebffffffff0000001700000000",
            INIT_62 => X"ffffffffffffffffffffffe4ffffffff0000000000000000fffffffcffffffff",
            INIT_63 => X"0000000b00000000fffffff6ffffffff0000000d00000000ffffffebffffffff",
            INIT_64 => X"ffffffebffffffffffffffe0fffffffffffffffeffffffffffffffe7ffffffff",
            INIT_65 => X"0000001d00000000000000370000000000000039000000000000001600000000",
            INIT_66 => X"0000000300000000ffffffdcffffffff0000002b000000000000002f00000000",
            INIT_67 => X"00000007000000000000000a000000000000001700000000ffffffdbffffffff",
            INIT_68 => X"0000003d0000000000000048000000000000001a000000000000001300000000",
            INIT_69 => X"0000003e000000000000008a0000000000000052000000000000005d00000000",
            INIT_6A => X"0000000a00000000000000400000000000000047000000000000003700000000",
            INIT_6B => X"ffffffe2ffffffffffffffddffffffff0000001500000000fffffff5ffffffff",
            INIT_6C => X"ffffffd5ffffffffffffffbffffffffffffffff9ffffffffffffffa8ffffffff",
            INIT_6D => X"ffffffaeffffffffffffffa0ffffffffffffffbcffffffffffffffeaffffffff",
            INIT_6E => X"0000001c000000000000000900000000fffffffaffffffff0000000800000000",
            INIT_6F => X"fffffff0ffffffffffffffd8ffffffff0000003f000000000000004500000000",
            INIT_70 => X"ffffffeaffffffff00000008000000000000001500000000ffffffe5ffffffff",
            INIT_71 => X"ffffffc5ffffffff00000012000000000000000c000000000000002500000000",
            INIT_72 => X"ffffffd6ffffffffffffffc6ffffffffffffffc1ffffffffffffffccffffffff",
            INIT_73 => X"0000000a000000000000000a000000000000002a00000000ffffffd2ffffffff",
            INIT_74 => X"ffffffc7ffffffff0000000b000000000000000000000000ffffffc4ffffffff",
            INIT_75 => X"fffffff4ffffffffffffffe3ffffffff0000000200000000fffffff0ffffffff",
            INIT_76 => X"ffffffffffffffff000000000000000000000038000000000000000e00000000",
            INIT_77 => X"0000002e000000000000001e000000000000001c000000000000002c00000000",
            INIT_78 => X"ffffffdcffffffffffffffcdffffffff0000002e00000000fffffffdffffffff",
            INIT_79 => X"fffffff4ffffffff0000000700000000ffffffeffffffffffffffff5ffffffff",
            INIT_7A => X"ffffffd5ffffffff00000001000000000000000100000000ffffffc3ffffffff",
            INIT_7B => X"0000000800000000ffffffe4ffffffff0000000f00000000fffffffaffffffff",
            INIT_7C => X"00000033000000000000001800000000ffffffeeffffffff0000003e00000000",
            INIT_7D => X"ffffffe7ffffffff000000050000000000000005000000000000000600000000",
            INIT_7E => X"ffffffeaffffffffffffffeefffffffffffffffdffffffff0000001800000000",
            INIT_7F => X"ffffffc5ffffffffffffffd6ffffffffffffffd5fffffffffffffffeffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE1 : if BRAM_NAME = "iwght_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff89ffffffffffffff98ffffffffffffff87ffffffffffffffbaffffffff",
            INIT_01 => X"fffffff3ffffffff0000001e00000000ffffffa2ffffffffffffff9cffffffff",
            INIT_02 => X"ffffffeeffffffff000000030000000000000013000000000000000100000000",
            INIT_03 => X"fffffff4ffffffffffffffe7ffffffffffffffecffffffff0000003e00000000",
            INIT_04 => X"0000001100000000ffffffd6ffffffff00000010000000000000001700000000",
            INIT_05 => X"0000004f000000000000003000000000fffffff5ffffffff0000003a00000000",
            INIT_06 => X"0000001300000000fffffff9fffffffffffffff2ffffffffffffffffffffffff",
            INIT_07 => X"fffffffeffffffffffffffdffffffffffffffff2fffffffffffffffcffffffff",
            INIT_08 => X"0000003d000000000000001e00000000ffffffd7ffffffff0000000b00000000",
            INIT_09 => X"0000001b000000000000002e000000000000002f00000000fffffff2ffffffff",
            INIT_0A => X"0000000700000000fffffff0ffffffff00000049000000000000003500000000",
            INIT_0B => X"0000000b00000000fffffffffffffffffffffff3ffffffff0000000800000000",
            INIT_0C => X"ffffffd0ffffffff0000001d00000000ffffffe8fffffffffffffff3ffffffff",
            INIT_0D => X"ffffff76ffffffffffffff9bffffffffffffffa1ffffffffffffffd7ffffffff",
            INIT_0E => X"ffffffaaffffffffffffffc3ffffffffffffff96ffffffffffffff8bffffffff",
            INIT_0F => X"ffffffd5ffffffffffffff9cffffffffffffff77fffffffffffffff1ffffffff",
            INIT_10 => X"ffffff86ffffffffffffffdeffffffffffffff40ffffffffffffff32ffffffff",
            INIT_11 => X"ffffffddfffffffffffffffaffffffffffffffecffffffffffffff87ffffffff",
            INIT_12 => X"fffffff7ffffffffffffffd3fffffffffffffff8ffffffffffffffffffffffff",
            INIT_13 => X"ffffffddffffffffffffffe4ffffffff0000000800000000fffffffeffffffff",
            INIT_14 => X"0000002f000000000000001a00000000fffffff5fffffffffffffff8ffffffff",
            INIT_15 => X"0000000e0000000000000022000000000000001a00000000ffffffd9ffffffff",
            INIT_16 => X"00000000000000000000001d00000000ffffffefffffffff0000000d00000000",
            INIT_17 => X"fffffffbffffffffffffffffffffffffffffffeafffffffffffffff2ffffffff",
            INIT_18 => X"ffffffccffffffff0000000500000000ffffffe4fffffffffffffff1ffffffff",
            INIT_19 => X"0000001500000000ffffffcaffffffff00000014000000000000000000000000",
            INIT_1A => X"fffffff3ffffffff00000031000000000000000c000000000000000000000000",
            INIT_1B => X"0000003500000000fffffffffffffffffffffffbffffffff0000001500000000",
            INIT_1C => X"ffffffdeffffffffffffffdcfffffffffffffff2ffffffff0000000c00000000",
            INIT_1D => X"0000000a00000000fffffff1fffffffffffffffaffffffff0000001300000000",
            INIT_1E => X"ffffffe4fffffffffffffffcffffffff00000026000000000000000800000000",
            INIT_1F => X"0000000100000000ffffffe2ffffffff00000019000000000000001300000000",
            INIT_20 => X"00000028000000000000001400000000ffffffe6fffffffffffffffaffffffff",
            INIT_21 => X"ffffffdeffffffffffffffe7ffffffff0000000a000000000000000200000000",
            INIT_22 => X"0000001100000000ffffffdcffffffffffffffeffffffffffffffff7ffffffff",
            INIT_23 => X"000000000000000000000019000000000000000800000000fffffff1ffffffff",
            INIT_24 => X"ffffffcdffffffffffffffdfffffffffffffffc9fffffffffffffffdffffffff",
            INIT_25 => X"0000004f000000000000003e00000000ffffffa7ffffffffffffff93ffffffff",
            INIT_26 => X"00000020000000000000000d0000000000000044000000000000001500000000",
            INIT_27 => X"ffffffffffffffff0000002e0000000000000028000000000000002c00000000",
            INIT_28 => X"ffffffc5ffffffffffffffe4ffffffffffffffeaffffffffffffffd1ffffffff",
            INIT_29 => X"fffffff5ffffffffffffffedffffffffffffffd0fffffffffffffff8ffffffff",
            INIT_2A => X"ffffffeeffffffff0000000b00000000fffffff9ffffffff0000000000000000",
            INIT_2B => X"ffffffe2ffffffff000000160000000000000007000000000000001300000000",
            INIT_2C => X"ffffffddffffffff000000120000000000000018000000000000002000000000",
            INIT_2D => X"0000001d00000000000000030000000000000009000000000000001300000000",
            INIT_2E => X"0000000000000000000000120000000000000028000000000000002c00000000",
            INIT_2F => X"ffffffe8ffffffff000000140000000000000004000000000000001000000000",
            INIT_30 => X"0000000a0000000000000017000000000000001800000000fffffff1ffffffff",
            INIT_31 => X"ffffffc3fffffffffffffffbffffffffffffffcaffffffffffffffe6ffffffff",
            INIT_32 => X"ffffffa4ffffffffffffffafffffffffffffffcdffffffffffffffcfffffffff",
            INIT_33 => X"00000013000000000000003e000000000000002400000000fffffff3ffffffff",
            INIT_34 => X"ffffffebffffffff00000006000000000000002a00000000fffffff8ffffffff",
            INIT_35 => X"0000002400000000fffffff5ffffffffffffffdeffffffff0000002a00000000",
            INIT_36 => X"00000008000000000000000b000000000000001800000000ffffffefffffffff",
            INIT_37 => X"0000000800000000ffffffdbffffffff00000006000000000000002200000000",
            INIT_38 => X"0000000c00000000fffffff2ffffffff0000001300000000ffffffd7ffffffff",
            INIT_39 => X"ffffffd7ffffffff00000011000000000000000100000000fffffffeffffffff",
            INIT_3A => X"ffffffc9ffffffffffffffcaffffffffffffffc9ffffffffffffffdaffffffff",
            INIT_3B => X"ffffffd7ffffffffffffffd9ffffffff0000000000000000fffffffbffffffff",
            INIT_3C => X"ffffffdfffffffff0000001d000000000000000600000000ffffffd0ffffffff",
            INIT_3D => X"ffffffedffffffff00000006000000000000000a00000000fffffff8ffffffff",
            INIT_3E => X"00000026000000000000000e000000000000001600000000fffffffeffffffff",
            INIT_3F => X"0000000000000000000000280000000000000004000000000000000e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffdfffffffffffffff4ffffffffffffffecffffffff0000000500000000",
            INIT_41 => X"0000001e000000000000001300000000ffffffddffffffff0000002500000000",
            INIT_42 => X"ffffffd6ffffffff0000001e000000000000000600000000ffffffe5ffffffff",
            INIT_43 => X"ffffffefffffffffffffffd2ffffffff0000000e000000000000000c00000000",
            INIT_44 => X"00000005000000000000001700000000ffffffe6ffffffff0000001b00000000",
            INIT_45 => X"ffffffeaffffffff0000001600000000ffffffe4fffffffffffffff2ffffffff",
            INIT_46 => X"ffffffcaffffffff0000000100000000fffffffcffffffffffffffe2ffffffff",
            INIT_47 => X"0000002700000000ffffffe8fffffffffffffffafffffffffffffff0ffffffff",
            INIT_48 => X"ffffffc2ffffffffffffffc2ffffffffffffffb5ffffffffffffffbeffffffff",
            INIT_49 => X"00000050000000000000005000000000ffffffd4ffffffffffffffebffffffff",
            INIT_4A => X"00000040000000000000009b0000000000000071000000000000004d00000000",
            INIT_4B => X"ffffffe5ffffffff00000073000000000000009300000000000000b300000000",
            INIT_4C => X"ffffffebffffffff00000008000000000000000a00000000fffffff1ffffffff",
            INIT_4D => X"fffffff8fffffffffffffffdfffffffffffffffdfffffffffffffff5ffffffff",
            INIT_4E => X"0000001e0000000000000014000000000000000500000000ffffffeaffffffff",
            INIT_4F => X"0000000500000000fffffff5fffffffffffffffdffffffffffffffffffffffff",
            INIT_50 => X"00000010000000000000001200000000ffffffd2ffffffff0000001300000000",
            INIT_51 => X"ffffffe3ffffffff0000003b00000000fffffff1ffffffffffffffcfffffffff",
            INIT_52 => X"fffffff1ffffffffffffffe6ffffffff00000019000000000000001800000000",
            INIT_53 => X"0000003300000000fffffff4ffffffff0000000d000000000000000a00000000",
            INIT_54 => X"fffffffaffffffff0000001200000000ffffffe1fffffffffffffffeffffffff",
            INIT_55 => X"ffffffecffffffffffffffe9ffffffff00000038000000000000003700000000",
            INIT_56 => X"0000002b000000000000002200000000ffffffdaffffffff0000001f00000000",
            INIT_57 => X"00000075000000000000005200000000fffffff3ffffffff0000002100000000",
            INIT_58 => X"00000066000000000000008b0000000000000037000000000000002800000000",
            INIT_59 => X"000000230000000000000010000000000000001f000000000000006b00000000",
            INIT_5A => X"fffffffeffffffff00000016000000000000001200000000fffffff5ffffffff",
            INIT_5B => X"0000002000000000ffffffd8ffffffffffffffe1ffffffffffffffdbffffffff",
            INIT_5C => X"00000034000000000000001600000000ffffffe4ffffffff0000001d00000000",
            INIT_5D => X"00000031000000000000000e000000000000000900000000ffffffdbffffffff",
            INIT_5E => X"ffffffe4ffffffff0000002500000000ffffffe4ffffffffffffffecffffffff",
            INIT_5F => X"ffffffeaffffffff00000004000000000000000900000000ffffffc4ffffffff",
            INIT_60 => X"0000000a00000000ffffffddffffffffffffffccfffffffffffffff0ffffffff",
            INIT_61 => X"ffffffe0fffffffffffffffaffffffff0000001f000000000000001b00000000",
            INIT_62 => X"0000001f00000000000000380000000000000040000000000000000000000000",
            INIT_63 => X"ffffffd5ffffffff0000002800000000ffffffefffffffff0000000b00000000",
            INIT_64 => X"fffffff5ffffffffffffffeeffffffffffffffefffffffffffffffdeffffffff",
            INIT_65 => X"00000018000000000000000600000000fffffff0fffffffffffffff3ffffffff",
            INIT_66 => X"ffffffd9fffffffffffffffcffffffff00000006000000000000001000000000",
            INIT_67 => X"fffffff8ffffffffffffffceffffffff0000000800000000ffffffefffffffff",
            INIT_68 => X"0000000a00000000fffffff5fffffffffffffff4fffffffffffffffcffffffff",
            INIT_69 => X"000000220000000000000020000000000000001900000000ffffffe6ffffffff",
            INIT_6A => X"ffffffe3fffffffffffffff9ffffffff0000003b000000000000002e00000000",
            INIT_6B => X"0000003b0000000000000008000000000000000900000000ffffffdbffffffff",
            INIT_6C => X"fffffff0ffffffff0000004f000000000000005e000000000000002c00000000",
            INIT_6D => X"0000003b00000000000000470000000000000055000000000000001600000000",
            INIT_6E => X"0000003800000000000000340000000000000051000000000000001700000000",
            INIT_6F => X"ffffffedffffffff0000002700000000ffffffd9fffffffffffffffcffffffff",
            INIT_70 => X"ffffffc5ffffffffffffffdbffffffff00000028000000000000000b00000000",
            INIT_71 => X"00000034000000000000003b000000000000002500000000ffffffe6ffffffff",
            INIT_72 => X"0000001400000000fffffffcffffffffffffffe4ffffffff0000001700000000",
            INIT_73 => X"fffffff8fffffffffffffff8ffffffff00000017000000000000000c00000000",
            INIT_74 => X"00000035000000000000000000000000ffffffecffffffffffffffecffffffff",
            INIT_75 => X"0000001b00000000fffffff2ffffffffffffffdeffffffff0000000200000000",
            INIT_76 => X"0000000200000000fffffff9ffffffff00000038000000000000003500000000",
            INIT_77 => X"ffffffecfffffffffffffff6ffffffff00000025000000000000002300000000",
            INIT_78 => X"00000028000000000000000a00000000ffffffeeffffffff0000000000000000",
            INIT_79 => X"0000005d00000000000000630000000000000038000000000000002200000000",
            INIT_7A => X"0000007b000000000000003f0000000000000006000000000000006000000000",
            INIT_7B => X"0000001200000000000000300000000000000001000000000000000a00000000",
            INIT_7C => X"ffffffd9fffffffffffffff3ffffffff00000004000000000000005c00000000",
            INIT_7D => X"0000002c000000000000000100000000fffffff7ffffffffffffffe7ffffffff",
            INIT_7E => X"ffffffd5ffffffffffffffc5ffffffffffffffc6ffffffffffffffe1ffffffff",
            INIT_7F => X"ffffffe4fffffffffffffff4fffffffffffffffbffffffffffffffddffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE1;


    MEM_IWGHT_LAYER1_INSTANCE2 : if BRAM_NAME = "iwght_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001900000000ffffffe8ffffffffffffffd2ffffffff0000001b00000000",
            INIT_01 => X"00000023000000000000000200000000fffffff8ffffffffffffffe3ffffffff",
            INIT_02 => X"0000001d000000000000002e0000000000000030000000000000002000000000",
            INIT_03 => X"0000000700000000fffffff8ffffffff00000002000000000000000700000000",
            INIT_04 => X"0000000500000000ffffffefffffffff00000019000000000000002800000000",
            INIT_05 => X"ffffffebffffffff00000003000000000000001d000000000000000100000000",
            INIT_06 => X"ffffffc5ffffffffffffffc8ffffffffffffffd6ffffffff0000001f00000000",
            INIT_07 => X"ffffffc1ffffffffffffffa0ffffffffffffffa9ffffffffffffffb7ffffffff",
            INIT_08 => X"00000027000000000000001200000000ffffffc8ffffffffffffffdaffffffff",
            INIT_09 => X"0000001600000000fffffffcffffffff00000003000000000000002300000000",
            INIT_0A => X"0000001000000000fffffffaffffffff0000001f00000000ffffffe1ffffffff",
            INIT_0B => X"fffffffdffffffff000000030000000000000026000000000000002d00000000",
            INIT_0C => X"fffffff7ffffffff0000001800000000ffffffe5fffffffffffffff9ffffffff",
            INIT_0D => X"0000000000000000ffffffe4fffffffffffffff3ffffffff0000000100000000",
            INIT_0E => X"ffffffdbffffffffffffffe7ffffffffffffffcdfffffffffffffffdffffffff",
            INIT_0F => X"ffffffc8ffffffffffffffd5fffffffffffffff5ffffffffffffffcdffffffff",
            INIT_10 => X"0000000d00000000ffffffd5ffffffffffffffd2ffffffffffffffe3ffffffff",
            INIT_11 => X"0000001300000000ffffffebfffffffffffffffcffffffff0000000b00000000",
            INIT_12 => X"0000000a0000000000000040000000000000002d000000000000002e00000000",
            INIT_13 => X"fffffff7ffffffff0000001e000000000000001a000000000000003500000000",
            INIT_14 => X"0000003800000000000000080000000000000033000000000000003100000000",
            INIT_15 => X"00000029000000000000003500000000fffffff1ffffffff0000000b00000000",
            INIT_16 => X"ffffffe6ffffffffffffffe5fffffffffffffff4ffffffffffffffe7ffffffff",
            INIT_17 => X"fffffffcffffffff0000000a00000000fffffff2ffffffff0000000000000000",
            INIT_18 => X"0000000500000000000000190000000000000015000000000000000000000000",
            INIT_19 => X"0000000a000000000000000a000000000000000900000000fffffff8ffffffff",
            INIT_1A => X"ffffffd8ffffffffffffffd8ffffffff0000000b000000000000000100000000",
            INIT_1B => X"ffffffdeffffffffffffffddffffffff0000000900000000ffffffdbffffffff",
            INIT_1C => X"0000000e00000000ffffffd2fffffffffffffff1ffffffffffffffd0ffffffff",
            INIT_1D => X"0000003e00000000000000160000000000000030000000000000000a00000000",
            INIT_1E => X"0000003600000000000000370000000000000035000000000000001d00000000",
            INIT_1F => X"00000025000000000000000800000000ffffffefffffffff0000001900000000",
            INIT_20 => X"00000016000000000000002400000000fffffffeffffffff0000001d00000000",
            INIT_21 => X"ffffffe2ffffffffffffffd9ffffffffffffffaafffffffffffffff2ffffffff",
            INIT_22 => X"ffffffd0ffffffffffffffbfffffffffffffff97ffffffffffffffd9ffffffff",
            INIT_23 => X"0000001b000000000000001400000000ffffffd9ffffffffffffffdeffffffff",
            INIT_24 => X"0000001100000000000000260000000000000014000000000000003200000000",
            INIT_25 => X"00000028000000000000000600000000fffffff7ffffffffffffffefffffffff",
            INIT_26 => X"0000000c00000000000000490000000000000051000000000000003000000000",
            INIT_27 => X"000000510000000000000040000000000000004c000000000000003e00000000",
            INIT_28 => X"ffffffecffffffff00000011000000000000002300000000fffffffaffffffff",
            INIT_29 => X"fffffff8ffffffffffffffd1ffffffff00000034000000000000000600000000",
            INIT_2A => X"00000036000000000000001f000000000000002b000000000000000c00000000",
            INIT_2B => X"0000002600000000000000310000000000000026000000000000002d00000000",
            INIT_2C => X"fffffff5ffffffffffffffdfffffffff0000001e000000000000001400000000",
            INIT_2D => X"fffffffdfffffffffffffff8ffffffffffffffe4ffffffff0000002600000000",
            INIT_2E => X"ffffffe5ffffffffffffffd5fffffffffffffff9ffffffffffffffc5ffffffff",
            INIT_2F => X"0000000000000000ffffffe1ffffffff00000041000000000000001400000000",
            INIT_30 => X"0000001b000000000000000f00000000ffffffcbffffffff0000002500000000",
            INIT_31 => X"000000210000000000000036000000000000000a000000000000002200000000",
            INIT_32 => X"0000000c00000000fffffff8ffffffff00000024000000000000002a00000000",
            INIT_33 => X"ffffffe2fffffffffffffff8ffffffff00000009000000000000001b00000000",
            INIT_34 => X"00000017000000000000001a000000000000001b00000000fffffff7ffffffff",
            INIT_35 => X"ffffffacfffffffffffffff1ffffffffffffffd8ffffffff0000000800000000",
            INIT_36 => X"ffffff8bffffffffffffffc4ffffffffffffffb7ffffffffffffffd6ffffffff",
            INIT_37 => X"fffffff3ffffffffffffff89ffffffffffffffafffffffffffffffd7ffffffff",
            INIT_38 => X"0000000800000000fffffff9fffffffffffffff9ffffffff0000000600000000",
            INIT_39 => X"00000005000000000000000100000000ffffffe2ffffffff0000000000000000",
            INIT_3A => X"0000000600000000fffffff6ffffffff00000019000000000000000b00000000",
            INIT_3B => X"ffffffedffffffff0000000d000000000000000b00000000fffffff0ffffffff",
            INIT_3C => X"00000039000000000000002f00000000ffffffe7fffffffffffffff7ffffffff",
            INIT_3D => X"ffffffc5ffffffff0000001400000000ffffffedffffffffffffffecffffffff",
            INIT_3E => X"0000001000000000fffffff3ffffffff0000001200000000fffffff6ffffffff",
            INIT_3F => X"0000001e000000000000001a00000000ffffffdaffffffff0000002d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000005000000000000000500000000fffffffbffffffffffffffdfffffffff",
            INIT_41 => X"fffffffdffffffff0000001d000000000000002d000000000000000a00000000",
            INIT_42 => X"ffffffdfffffffffffffffd0ffffffff00000022000000000000002a00000000",
            INIT_43 => X"ffffff60ffffffffffffff1dffffffffffffff7affffffffffffffb5ffffffff",
            INIT_44 => X"ffffff13ffffffffffffff67ffffffffffffff0fffffffffffffff31ffffffff",
            INIT_45 => X"00000012000000000000000b000000000000001700000000ffffff0fffffffff",
            INIT_46 => X"0000000100000000000000020000000000000002000000000000000300000000",
            INIT_47 => X"00000021000000000000000300000000ffffffe3ffffffff0000000500000000",
            INIT_48 => X"0000001600000000fffffff6fffffffffffffffaffffffff0000003000000000",
            INIT_49 => X"fffffff4ffffffff00000010000000000000001200000000ffffffc7ffffffff",
            INIT_4A => X"ffffffc3ffffffffffffffdfffffffffffffffc4ffffffffffffffb8ffffffff",
            INIT_4B => X"ffffffc0ffffffffffffffdaffffffff0000001800000000ffffffd2ffffffff",
            INIT_4C => X"0000002900000000ffffffeeffffffffffffffcbffffffff0000000600000000",
            INIT_4D => X"fffffff9ffffffff0000002600000000ffffffd2ffffffff0000000800000000",
            INIT_4E => X"ffffffebfffffffffffffff1ffffffff0000000900000000fffffff1ffffffff",
            INIT_4F => X"fffffffcffffffffffffffe6fffffffffffffff4ffffffff0000000200000000",
            INIT_50 => X"fffffffaffffffff0000000000000000fffffff5fffffffffffffff0ffffffff",
            INIT_51 => X"ffffffd9ffffffffffffffebffffffff0000000900000000ffffffbaffffffff",
            INIT_52 => X"0000000500000000fffffffcfffffffffffffffeffffffff0000000d00000000",
            INIT_53 => X"fffffffeffffffff0000001400000000ffffffd8ffffffffffffffe3ffffffff",
            INIT_54 => X"000000310000000000000031000000000000001a00000000ffffffdeffffffff",
            INIT_55 => X"0000002a00000000ffffffc8ffffffffffffffd4fffffffffffffffcffffffff",
            INIT_56 => X"ffffffffffffffff0000002100000000ffffffddffffffff0000001100000000",
            INIT_57 => X"0000000a0000000000000014000000000000002d00000000ffffffe1ffffffff",
            INIT_58 => X"0000004100000000000000100000000000000000000000000000003e00000000",
            INIT_59 => X"0000009e000000000000002100000000ffffffeeffffffff0000001600000000",
            INIT_5A => X"00000023000000000000004c00000000ffffffdeffffffff0000001500000000",
            INIT_5B => X"000000120000000000000050000000000000003e000000000000000900000000",
            INIT_5C => X"ffffffe9ffffffffffffffd6ffffffffffffffebfffffffffffffffaffffffff",
            INIT_5D => X"000000010000000000000023000000000000000e000000000000000b00000000",
            INIT_5E => X"fffffffbffffffffffffffeefffffffffffffff3ffffffff0000001400000000",
            INIT_5F => X"ffffffe0ffffffff0000001500000000fffffffefffffffffffffffdffffffff",
            INIT_60 => X"ffffffeefffffffffffffffeffffffff00000002000000000000000200000000",
            INIT_61 => X"0000002800000000ffffffe9ffffffffffffffe7fffffffffffffff6ffffffff",
            INIT_62 => X"0000000e0000000000000025000000000000003300000000fffffff8ffffffff",
            INIT_63 => X"ffffffe0fffffffffffffff3ffffffff0000000b00000000ffffffd5ffffffff",
            INIT_64 => X"00000010000000000000002000000000fffffff3ffffffff0000001600000000",
            INIT_65 => X"0000005700000000000000340000000000000014000000000000001900000000",
            INIT_66 => X"00000001000000000000001b000000000000003f000000000000003800000000",
            INIT_67 => X"00000046000000000000007500000000000000a5000000000000005a00000000",
            INIT_68 => X"000000270000000000000011000000000000007b000000000000008c00000000",
            INIT_69 => X"00000018000000000000000000000000fffffffcffffffff0000005500000000",
            INIT_6A => X"fffffff5ffffffff00000018000000000000003100000000fffffffaffffffff",
            INIT_6B => X"ffffffe6fffffffffffffff4ffffffff00000029000000000000001c00000000",
            INIT_6C => X"ffffffd5ffffffffffffffe7ffffffff0000000c00000000ffffffc8ffffffff",
            INIT_6D => X"ffffffcfffffffff00000009000000000000000e000000000000000e00000000",
            INIT_6E => X"ffffffeaffffffffffffffbfffffffff00000018000000000000000000000000",
            INIT_6F => X"ffffffa6ffffffffffffffd3ffffffffffffffe9ffffffffffffffedffffffff",
            INIT_70 => X"0000000400000000000000420000000000000032000000000000001500000000",
            INIT_71 => X"ffffffecffffffffffffffe2fffffffffffffffbffffffff0000000400000000",
            INIT_72 => X"ffffffbeffffffffffffffc4ffffffffffffffd0ffffffff0000001800000000",
            INIT_73 => X"0000000100000000fffffff0ffffffff00000011000000000000000700000000",
            INIT_74 => X"00000007000000000000000000000000ffffffd3ffffffff0000000300000000",
            INIT_75 => X"fffffff9fffffffffffffff6ffffffff00000013000000000000003500000000",
            INIT_76 => X"ffffffffffffffff0000002500000000fffffff3ffffffff0000001f00000000",
            INIT_77 => X"fffffff0ffffffff000000050000000000000036000000000000001a00000000",
            INIT_78 => X"fffffff7ffffffff000000200000000000000021000000000000001000000000",
            INIT_79 => X"ffffffe7ffffffff00000000000000000000001f00000000fffffff6ffffffff",
            INIT_7A => X"0000000d00000000fffffff4fffffffffffffffffffffffffffffff3ffffffff",
            INIT_7B => X"ffffffdaffffffffffffffc9ffffffffffffffe6fffffffffffffff9ffffffff",
            INIT_7C => X"fffffff2ffffffffffffffd9ffffffffffffffe7ffffffffffffffb8ffffffff",
            INIT_7D => X"0000003400000000fffffffaffffffffffffff93ffffffffffffffbdffffffff",
            INIT_7E => X"00000017000000000000003e000000000000000300000000ffffffefffffffff",
            INIT_7F => X"fffffff2fffffffffffffff4ffffffff0000001b00000000fffffff3ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE2;


    MEM_IWGHT_LAYER1_INSTANCE3 : if BRAM_NAME = "iwght_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffdbfffffffffffffff3fffffffffffffff6ffffffffffffffe9ffffffff",
            INIT_01 => X"fffffff1fffffffffffffff6ffffffffffffffe1ffffffffffffffe8ffffffff",
            INIT_02 => X"fffffff6fffffffffffffff1ffffffffffffffeeffffffff0000000200000000",
            INIT_03 => X"fffffff4ffffffff0000000d000000000000000800000000ffffffe7ffffffff",
            INIT_04 => X"0000000400000000ffffffe7ffffffff00000000000000000000000f00000000",
            INIT_05 => X"0000002400000000000000000000000000000015000000000000002800000000",
            INIT_06 => X"0000000f000000000000000000000000fffffffcffffffff0000000b00000000",
            INIT_07 => X"ffffffe5fffffffffffffff5ffffffff0000000b00000000fffffff7ffffffff",
            INIT_08 => X"fffffff6fffffffffffffff6ffffffff0000001c000000000000001600000000",
            INIT_09 => X"ffffffe8ffffffffffffffadffffffffffffffcefffffffffffffffcffffffff",
            INIT_0A => X"ffffff9effffffffffffff98ffffffffffffffb0ffffffffffffffa3ffffffff",
            INIT_0B => X"0000002e000000000000000f0000000000000026000000000000000700000000",
            INIT_0C => X"0000002d0000000000000017000000000000001d000000000000002800000000",
            INIT_0D => X"ffffffcaffffffffffffffd7ffffffffffffffdbffffffff0000001200000000",
            INIT_0E => X"0000001c00000000ffffffd8fffffffffffffffcffffffff0000000f00000000",
            INIT_0F => X"00000034000000000000001000000000ffffffd8ffffffff0000000d00000000",
            INIT_10 => X"0000000f00000000ffffffffffffffff00000005000000000000001500000000",
            INIT_11 => X"0000004800000000ffffffe9ffffffff0000000000000000ffffffe2ffffffff",
            INIT_12 => X"0000002000000000000000410000000000000034000000000000002c00000000",
            INIT_13 => X"0000007400000000000000460000000000000032000000000000003800000000",
            INIT_14 => X"ffffffedffffffffffffffecfffffffffffffffcffffffff0000001d00000000",
            INIT_15 => X"fffffff1fffffffffffffff1ffffffff0000000100000000ffffffe8ffffffff",
            INIT_16 => X"00000012000000000000002f000000000000004000000000ffffffebffffffff",
            INIT_17 => X"fffffffeffffffffffffffecffffffffffffffe2ffffffff0000002400000000",
            INIT_18 => X"0000001d00000000fffffff7ffffffffffffffe2ffffffffffffffeeffffffff",
            INIT_19 => X"0000001c0000000000000012000000000000000f000000000000001e00000000",
            INIT_1A => X"fffffffffffffffffffffffcffffffff0000001a00000000fffffff7ffffffff",
            INIT_1B => X"ffffffe5fffffffffffffffeffffffffffffffe3ffffffffffffffdeffffffff",
            INIT_1C => X"0000001d00000000000000060000000000000011000000000000000a00000000",
            INIT_1D => X"0000000e00000000000000400000000000000022000000000000004d00000000",
            INIT_1E => X"0000000b000000000000001900000000ffffffd5ffffffffffffffe5ffffffff",
            INIT_1F => X"0000000b000000000000001c00000000fffffffcffffffffffffffe1ffffffff",
            INIT_20 => X"0000001200000000000000160000000000000015000000000000000300000000",
            INIT_21 => X"ffffffdafffffffffffffff5ffffffff00000003000000000000001500000000",
            INIT_22 => X"0000000f000000000000000e00000000ffffffbcffffffff0000000b00000000",
            INIT_23 => X"ffffffadfffffffffffffff1ffffffff0000003900000000ffffffffffffffff",
            INIT_24 => X"00000035000000000000002400000000ffffffb5ffffffffffffff8fffffffff",
            INIT_25 => X"0000002b0000000000000034000000000000003b000000000000005100000000",
            INIT_26 => X"fffffff6ffffffff0000000e00000000fffffffbffffffff0000000f00000000",
            INIT_27 => X"ffffffecffffffffffffffe7ffffffffffffffe7ffffffffffffffefffffffff",
            INIT_28 => X"ffffffc5ffffffffffffffbfffffffffffffffe8ffffffff0000000e00000000",
            INIT_29 => X"0000001e000000000000000e000000000000002a000000000000000600000000",
            INIT_2A => X"0000002e0000000000000045000000000000000b000000000000003700000000",
            INIT_2B => X"ffffffe3ffffffffffffffe0ffffffff0000000b000000000000002e00000000",
            INIT_2C => X"0000003c00000000fffffffeffffffff0000000000000000ffffffd5ffffffff",
            INIT_2D => X"0000001a000000000000000b0000000000000017000000000000002800000000",
            INIT_2E => X"ffffffffffffffff00000045000000000000003f000000000000000b00000000",
            INIT_2F => X"ffffffd8ffffffff0000000d0000000000000016000000000000001400000000",
            INIT_30 => X"0000003600000000ffffffe2ffffffff00000017000000000000000700000000",
            INIT_31 => X"fffffff7ffffffff0000000a000000000000001800000000fffffffcffffffff",
            INIT_32 => X"ffffffb2ffffffffffffffedffffffffffffffc7ffffffffffffffd6ffffffff",
            INIT_33 => X"fffffffdffffffffffffffe5ffffffffffffffc0ffffffffffffffb2ffffffff",
            INIT_34 => X"ffffffe2ffffffff00000002000000000000000900000000fffffffdffffffff",
            INIT_35 => X"0000004b0000000000000012000000000000000f00000000fffffff9ffffffff",
            INIT_36 => X"fffffff5ffffffff0000001a000000000000006d000000000000005b00000000",
            INIT_37 => X"ffffffeaffffffffffffffc1ffffffffffffff9effffffff0000001700000000",
            INIT_38 => X"fffffff0ffffffffffffffd1ffffffffffffffd9ffffffffffffffd8ffffffff",
            INIT_39 => X"0000000000000000ffffffe3ffffffff00000016000000000000000200000000",
            INIT_3A => X"fffffffdffffffff0000001100000000fffffff2ffffffffffffffe5ffffffff",
            INIT_3B => X"00000035000000000000001800000000fffffff6ffffffff0000001200000000",
            INIT_3C => X"0000000200000000ffffffedffffffff00000020000000000000001d00000000",
            INIT_3D => X"ffffffe9ffffffffffffffdcffffffffffffffe3fffffffffffffffbffffffff",
            INIT_3E => X"00000000000000000000001400000000fffffffaffffffff0000000400000000",
            INIT_3F => X"fffffff4ffffffff0000000f00000000ffffffebffffffffffffffd3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002b000000000000001e000000000000002500000000ffffffefffffffff",
            INIT_41 => X"fffffff8ffffffff0000000a0000000000000025000000000000001100000000",
            INIT_42 => X"ffffffd3ffffffffffffffe5ffffffff00000003000000000000001f00000000",
            INIT_43 => X"000000300000000000000015000000000000001700000000ffffffc7ffffffff",
            INIT_44 => X"ffffffc5ffffffff000000600000000000000057000000000000003300000000",
            INIT_45 => X"00000007000000000000002600000000ffffffb4ffffffffffffff9cffffffff",
            INIT_46 => X"0000000800000000ffffffd9ffffffffffffffbaffffffff0000001300000000",
            INIT_47 => X"0000000400000000ffffff58ffffffffffffff21ffffffffffffff10ffffffff",
            INIT_48 => X"0000000b00000000ffffffd5fffffffffffffffcfffffffffffffffeffffffff",
            INIT_49 => X"0000003d00000000000000190000000000000012000000000000000200000000",
            INIT_4A => X"fffffffffffffffffffffff4fffffffffffffff9ffffffff0000000400000000",
            INIT_4B => X"ffffffe2ffffffffffffffe8ffffffff0000001d000000000000000a00000000",
            INIT_4C => X"0000000d00000000ffffffe9ffffffffffffffebfffffffffffffff5ffffffff",
            INIT_4D => X"00000023000000000000002d0000000000000003000000000000000a00000000",
            INIT_4E => X"ffffffe2fffffffffffffff5ffffffff0000004e000000000000003100000000",
            INIT_4F => X"ffffffd8ffffffff0000001400000000ffffffe8fffffffffffffffdffffffff",
            INIT_50 => X"00000027000000000000001c0000000000000034000000000000002000000000",
            INIT_51 => X"0000007d000000000000006c00000000fffffffdffffffff0000002500000000",
            INIT_52 => X"ffffff7effffffffffffff4affffffffffffff89ffffffff0000004500000000",
            INIT_53 => X"fffffff5ffffffff0000002e0000000000000019000000000000002e00000000",
            INIT_54 => X"ffffff09fffffffffffffef4fffffffffffffffeffffffffffffffd0ffffffff",
            INIT_55 => X"fffffffcffffffffffffffcdffffffffffffffcfffffffffffffff28ffffffff",
            INIT_56 => X"0000004900000000ffffffd8ffffffffffffffd1ffffffffffffffebffffffff",
            INIT_57 => X"ffffffe9ffffffffffffffd6ffffffff00000055000000000000004600000000",
            INIT_58 => X"fffffff5ffffffff00000007000000000000000b00000000ffffffddffffffff",
            INIT_59 => X"00000027000000000000000d0000000000000013000000000000000000000000",
            INIT_5A => X"fffffff3ffffffffffffffebffffffff0000003d000000000000002e00000000",
            INIT_5B => X"ffffffaaffffffffffffff8cffffffffffffffadffffffffffffffa2ffffffff",
            INIT_5C => X"ffffffecfffffffffffffff5ffffffff0000000f00000000fffffffeffffffff",
            INIT_5D => X"0000000f00000000fffffff9ffffffffffffffefffffffff0000001d00000000",
            INIT_5E => X"ffffffd0ffffffffffffffd5fffffffffffffffaffffffffffffffecffffffff",
            INIT_5F => X"0000002000000000ffffffd4ffffffffffffffeaffffffff0000000000000000",
            INIT_60 => X"00000005000000000000002000000000ffffffedffffffffffffffffffffffff",
            INIT_61 => X"fffffff5fffffffffffffff6ffffffff0000002d00000000ffffffd4ffffffff",
            INIT_62 => X"0000002a00000000ffffffdeffffffffffffffefffffffff0000001c00000000",
            INIT_63 => X"ffffffeaffffffff0000002f00000000ffffffdfffffffffffffffe8ffffffff",
            INIT_64 => X"ffffffe1ffffffff00000000000000000000002700000000ffffffc9ffffffff",
            INIT_65 => X"0000001800000000fffffffaffffffff0000002000000000ffffffffffffffff",
            INIT_66 => X"0000003200000000000000150000000000000012000000000000002f00000000",
            INIT_67 => X"ffffffe2ffffffffffffffe9fffffffffffffffbffffffff0000001300000000",
            INIT_68 => X"ffffffe7ffffffffffffffceffffffffffffffc7ffffffffffffffe6ffffffff",
            INIT_69 => X"0000001c000000000000006f00000000ffffffa2ffffffffffffffd4ffffffff",
            INIT_6A => X"0000007900000000000000090000000000000062000000000000004b00000000",
            INIT_6B => X"00000015000000000000009b000000000000001d000000000000005300000000",
            INIT_6C => X"00000011000000000000002c00000000ffffffebffffffffffffffe7ffffffff",
            INIT_6D => X"ffffffeaffffffffffffffedffffffff0000001500000000fffffffdffffffff",
            INIT_6E => X"0000000700000000ffffffeaffffffffffffffecfffffffffffffff0ffffffff",
            INIT_6F => X"000000050000000000000018000000000000000000000000ffffffedffffffff",
            INIT_70 => X"ffffffc9ffffffff000000030000000000000027000000000000001c00000000",
            INIT_71 => X"0000003a00000000ffffffccffffffffffffffd2ffffffff0000000500000000",
            INIT_72 => X"ffffffe3fffffffffffffff8fffffffffffffffcffffffffffffffe6ffffffff",
            INIT_73 => X"ffffffe1ffffffffffffffe5ffffffff0000001700000000fffffff6ffffffff",
            INIT_74 => X"0000000d00000000fffffff2ffffffff00000013000000000000002900000000",
            INIT_75 => X"ffffffb0ffffffffffffffeeffffffffffffffe4ffffffffffffffddffffffff",
            INIT_76 => X"ffffffc3ffffffffffffff94ffffffffffffffc7ffffffffffffffceffffffff",
            INIT_77 => X"0000001a0000000000000067000000000000005700000000ffffffefffffffff",
            INIT_78 => X"0000004800000000000000150000000000000076000000000000006c00000000",
            INIT_79 => X"0000001500000000fffffffbffffffff00000018000000000000008200000000",
            INIT_7A => X"0000000f0000000000000015000000000000001600000000fffffffeffffffff",
            INIT_7B => X"0000000d000000000000000600000000ffffffeaffffffffffffffdfffffffff",
            INIT_7C => X"ffffffebffffffff00000017000000000000002900000000ffffffd6ffffffff",
            INIT_7D => X"0000000100000000ffffffdaffffffff0000001d000000000000002900000000",
            INIT_7E => X"fffffff0ffffffff0000000b000000000000000b00000000ffffffecffffffff",
            INIT_7F => X"fffffff4ffffffff0000000f00000000fffffff1ffffffff0000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE3;


    MEM_IWGHT_LAYER1_INSTANCE4 : if BRAM_NAME = "iwght_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000018000000000000001600000000ffffffe8ffffffff0000001100000000",
            INIT_01 => X"fffffffcffffffff0000000c0000000000000017000000000000001700000000",
            INIT_02 => X"0000000000000000ffffffe7ffffffff00000005000000000000000c00000000",
            INIT_03 => X"ffffffefffffffffffffffe6fffffffffffffffffffffffffffffffdffffffff",
            INIT_04 => X"ffffffefffffffff0000001300000000ffffffebffffffff0000000e00000000",
            INIT_05 => X"fffffffdffffffff000000080000000000000013000000000000000600000000",
            INIT_06 => X"0000000600000000000000070000000000000009000000000000000c00000000",
            INIT_07 => X"fffffff8ffffffffffffffecffffffffffffffe5ffffffff0000000d00000000",
            INIT_08 => X"ffffffe3ffffffffffffffe5ffffffffffffffeaffffffff0000000a00000000",
            INIT_09 => X"fffffff9ffffffff0000001300000000fffffff3ffffffffffffffeeffffffff",
            INIT_0A => X"fffffff2fffffffffffffff2ffffffff0000000600000000fffffff1ffffffff",
            INIT_0B => X"ffffffebffffffffffffffe2ffffffff0000001300000000ffffffedffffffff",
            INIT_0C => X"ffffffecffffffff0000000d00000000ffffffedfffffffffffffff1ffffffff",
            INIT_0D => X"fffffff2ffffffff0000000600000000ffffffe6ffffffffffffffe2ffffffff",
            INIT_0E => X"ffffffecffffffffffffffeffffffffffffffff5ffffffffffffffe2ffffffff",
            INIT_0F => X"0000000e000000000000000500000000fffffffdffffffffffffffe4ffffffff",
            INIT_10 => X"fffffff1ffffffff0000000500000000fffffff8ffffffff0000000800000000",
            INIT_11 => X"ffffffeeffffffffffffffdeffffffff0000000f00000000fffffffcffffffff",
            INIT_12 => X"fffffff2ffffffff00000014000000000000001b000000000000001400000000",
            INIT_13 => X"fffffff9ffffffff0000000900000000fffffff7fffffffffffffffcffffffff",
            INIT_14 => X"0000000f00000000ffffffeffffffffffffffff4fffffffffffffff7ffffffff",
            INIT_15 => X"ffffffe4fffffffffffffff4ffffffff00000000000000000000000500000000",
            INIT_16 => X"00000006000000000000000300000000ffffffeaffffffffffffffffffffffff",
            INIT_17 => X"fffffffeffffffff00000006000000000000001300000000fffffff5ffffffff",
            INIT_18 => X"00000007000000000000000d00000000fffffffaffffffffffffffedffffffff",
            INIT_19 => X"ffffffeaffffffffffffffefffffffff00000012000000000000000c00000000",
            INIT_1A => X"00000016000000000000000700000000ffffffeeffffffff0000001300000000",
            INIT_1B => X"0000000e00000000ffffffe1ffffffffffffffe8ffffffffffffffebffffffff",
            INIT_1C => X"ffffffebfffffffffffffff8ffffffffffffffebffffffff0000000b00000000",
            INIT_1D => X"ffffffe7ffffffffffffffe4ffffffff0000001600000000ffffffecffffffff",
            INIT_1E => X"fffffffeffffffff0000000600000000fffffff3fffffffffffffff0ffffffff",
            INIT_1F => X"ffffffe4ffffffffffffffe8fffffffffffffff3fffffffffffffffdffffffff",
            INIT_20 => X"ffffffe6ffffffff0000000200000000fffffff9ffffffff0000000500000000",
            INIT_21 => X"0000000c00000000000000190000000000000017000000000000000800000000",
            INIT_22 => X"fffffff8ffffffffffffffe6ffffffff00000016000000000000001100000000",
            INIT_23 => X"0000000b00000000ffffffeeffffffffffffffeeffffffff0000001a00000000",
            INIT_24 => X"00000013000000000000001200000000ffffffe1ffffffffffffffe8ffffffff",
            INIT_25 => X"fffffff9ffffffff0000001100000000fffffff1fffffffffffffff6ffffffff",
            INIT_26 => X"000000180000000000000015000000000000002500000000fffffff1ffffffff",
            INIT_27 => X"ffffffbdfffffffffffffff7fffffffffffffff6ffffffff0000000b00000000",
            INIT_28 => X"fffffff8ffffffffffffffe5ffffffffffffffb6ffffffffffffffbbffffffff",
            INIT_29 => X"fffffff6fffffffffffffff5ffffffff00000007000000000000000200000000",
            INIT_2A => X"0000002500000000ffffffd7fffffffffffffffbffffffff0000002700000000",
            INIT_2B => X"ffffffecffffffffffffffecffffffff00000007000000000000001500000000",
            INIT_2C => X"000000030000000000000000000000000000000700000000fffffffdffffffff",
            INIT_2D => X"000000090000000000000007000000000000000b00000000fffffffbffffffff",
            INIT_2E => X"ffffffceffffffffffffffe3fffffffffffffff5ffffffff0000002300000000",
            INIT_2F => X"ffffffd8fffffffffffffffeffffffff0000000900000000fffffff2ffffffff",
            INIT_30 => X"0000003a000000000000001d000000000000000b000000000000003400000000",
            INIT_31 => X"fffffffcfffffffffffffff4ffffffff00000011000000000000001100000000",
            INIT_32 => X"0000000d000000000000005d000000000000000c00000000ffffffcaffffffff",
            INIT_33 => X"00000002000000000000001b0000000000000007000000000000001300000000",
            INIT_34 => X"ffffffe6ffffffffffffffe0ffffffff0000001a000000000000002700000000",
            INIT_35 => X"000000110000000000000006000000000000002700000000fffffff2ffffffff",
            INIT_36 => X"0000000c00000000ffffffe4ffffffff0000000b00000000ffffffeeffffffff",
            INIT_37 => X"0000001800000000fffffffafffffffffffffff6ffffffff0000001300000000",
            INIT_38 => X"fffffffcffffffffffffffecfffffffffffffffafffffffffffffff9ffffffff",
            INIT_39 => X"0000000c00000000ffffffd9ffffffff0000000400000000ffffffe0ffffffff",
            INIT_3A => X"fffffff7ffffffff0000001a000000000000000f00000000fffffffaffffffff",
            INIT_3B => X"ffffffe2fffffffffffffffbffffffff0000000500000000fffffff2ffffffff",
            INIT_3C => X"ffffffebffffffffffffffc0ffffffffffffffb9ffffffffffffffceffffffff",
            INIT_3D => X"00000043000000000000005b000000000000000d000000000000002700000000",
            INIT_3E => X"000000770000000000000067000000000000004e000000000000005a00000000",
            INIT_3F => X"0000007000000000000000380000000000000034000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000040000000000000002c000000000000004d000000000000005000000000",
            INIT_41 => X"0000001c000000000000002f000000000000002a000000000000001500000000",
            INIT_42 => X"ffffffbeffffffff000000140000000000000003000000000000001d00000000",
            INIT_43 => X"00000007000000000000002a00000000ffffffcfffffffffffffffb5ffffffff",
            INIT_44 => X"fffffff1ffffffffffffffe4fffffffffffffff8ffffffffffffffe7ffffffff",
            INIT_45 => X"0000004500000000fffffff1ffffffffffffffd7ffffffff0000000200000000",
            INIT_46 => X"00000045000000000000005a0000000000000058000000000000007100000000",
            INIT_47 => X"0000000800000000ffffffe8fffffffffffffff6ffffffff0000003f00000000",
            INIT_48 => X"ffffffe7ffffffffffffffd4fffffffffffffff2ffffffff0000001400000000",
            INIT_49 => X"ffffffeefffffffffffffff8fffffffffffffff4fffffffffffffff9ffffffff",
            INIT_4A => X"0000000d000000000000001500000000fffffff4ffffffff0000000500000000",
            INIT_4B => X"fffffffeffffffff000000280000000000000014000000000000000000000000",
            INIT_4C => X"ffffffc2ffffffffffffffd9ffffffff0000003e000000000000003e00000000",
            INIT_4D => X"ffffffd8ffffffffffffffcefffffffffffffffcffffffffffffffdbffffffff",
            INIT_4E => X"0000001400000000fffffffaffffffffffffffdefffffffffffffff9ffffffff",
            INIT_4F => X"0000000100000000fffffff6ffffffffffffffddffffffffffffffe2ffffffff",
            INIT_50 => X"fffffff9ffffffffffffffebffffffff00000024000000000000001100000000",
            INIT_51 => X"00000017000000000000001c0000000000000009000000000000001400000000",
            INIT_52 => X"0000003700000000000000070000000000000025000000000000002600000000",
            INIT_53 => X"000000360000000000000024000000000000003c000000000000001300000000",
            INIT_54 => X"ffffffeeffffffffffffffefffffffffffffffe4ffffffffffffffefffffffff",
            INIT_55 => X"0000000d00000000ffffffd2fffffffffffffff0ffffffffffffffe2ffffffff",
            INIT_56 => X"ffffffeaffffffffffffffe3ffffffffffffffacffffffff0000001600000000",
            INIT_57 => X"0000001800000000ffffffefffffffff0000000600000000ffffffcbffffffff",
            INIT_58 => X"ffffffb6ffffffffffffffe4fffffffffffffff4fffffffffffffff7ffffffff",
            INIT_59 => X"ffffffd0ffffffffffffffc0ffffffffffffffb3ffffffffffffffe2ffffffff",
            INIT_5A => X"0000001000000000fffffff7ffffffffffffffeaffffffff0000001000000000",
            INIT_5B => X"0000000100000000fffffffdfffffffffffffff4fffffffffffffff9ffffffff",
            INIT_5C => X"00000007000000000000000800000000fffffff3ffffffff0000001d00000000",
            INIT_5D => X"0000000b00000000ffffffefffffffffffffffe8ffffffff0000002300000000",
            INIT_5E => X"00000004000000000000001400000000fffffffbffffffff0000000e00000000",
            INIT_5F => X"00000007000000000000001f000000000000001a00000000ffffffe6ffffffff",
            INIT_60 => X"00000016000000000000000500000000fffffffbffffffff0000002f00000000",
            INIT_61 => X"ffffffdaffffffff000000010000000000000025000000000000000f00000000",
            INIT_62 => X"ffffffccffffffffffffffc6ffffffffffffffe8ffffffffffffffddffffffff",
            INIT_63 => X"0000000500000000ffffffffffffffff00000009000000000000001900000000",
            INIT_64 => X"fffffff5ffffffff0000001000000000fffffff9ffffffff0000000b00000000",
            INIT_65 => X"fffffff6fffffffffffffffbfffffffffffffff1fffffffffffffff4ffffffff",
            INIT_66 => X"0000001600000000000000040000000000000021000000000000000b00000000",
            INIT_67 => X"ffffffe3ffffffff000000030000000000000035000000000000001300000000",
            INIT_68 => X"ffffffe1ffffffff0000001100000000ffffffedffffffff0000000e00000000",
            INIT_69 => X"ffffffa2ffffffff0000000e0000000000000002000000000000001000000000",
            INIT_6A => X"ffffff9fffffffffffffffabffffffffffffffe3ffffffffffffffa2ffffffff",
            INIT_6B => X"ffffffc7ffffffffffffffb5ffffffffffffffb5ffffffffffffffcaffffffff",
            INIT_6C => X"0000001100000000ffffffdcffffffffffffffd5ffffffff0000000600000000",
            INIT_6D => X"fffffff6ffffffff00000008000000000000000c00000000fffffffaffffffff",
            INIT_6E => X"0000000300000000ffffffe7ffffffffffffffbfffffffff0000000a00000000",
            INIT_6F => X"0000002f000000000000000a000000000000001d00000000fffffffbffffffff",
            INIT_70 => X"fffffff9ffffffff00000010000000000000001f000000000000004200000000",
            INIT_71 => X"fffffff9ffffffffffffffd6ffffffff0000002f00000000ffffffd8ffffffff",
            INIT_72 => X"0000000b00000000ffffffc6ffffffffffffffd1fffffffffffffffaffffffff",
            INIT_73 => X"fffffff4ffffffff0000000d000000000000001000000000fffffff5ffffffff",
            INIT_74 => X"fffffff6ffffffff0000000000000000ffffffdaffffffff0000002000000000",
            INIT_75 => X"ffffffe1fffffffffffffffeffffffffffffffb3ffffffffffffffc9ffffffff",
            INIT_76 => X"fffffff5fffffffffffffff9ffffffffffffffe4ffffffffffffffa2ffffffff",
            INIT_77 => X"0000000c00000000fffffff7fffffffffffffff7ffffffff0000002700000000",
            INIT_78 => X"0000000200000000fffffff0ffffffffffffffd9ffffffff0000001200000000",
            INIT_79 => X"0000001800000000ffffffd6ffffffffffffffbfffffffffffffffcdffffffff",
            INIT_7A => X"fffffffcffffffff00000053000000000000001d000000000000000b00000000",
            INIT_7B => X"0000002900000000fffffffeffffffff00000026000000000000004100000000",
            INIT_7C => X"00000000000000000000001b0000000000000022000000000000003a00000000",
            INIT_7D => X"ffffffd0ffffffffffffffd6fffffffffffffff3ffffffffffffffd9ffffffff",
            INIT_7E => X"0000000200000000ffffffe4ffffffffffffffefffffffffffffffe4ffffffff",
            INIT_7F => X"0000001000000000fffffffbffffffff0000000c000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE4;


    MEM_IWGHT_LAYER1_INSTANCE5 : if BRAM_NAME = "iwght_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000400000000ffffffdaffffffffffffffbbffffffff0000000400000000",
            INIT_01 => X"fffffffbfffffffffffffff0ffffffff0000000b00000000ffffffd1ffffffff",
            INIT_02 => X"ffffffc0ffffffffffffffd1fffffffffffffff9fffffffffffffff0ffffffff",
            INIT_03 => X"0000001f00000000ffffffd3ffffffffffffffe7ffffffffffffffdcffffffff",
            INIT_04 => X"ffffffd1ffffffff0000001c00000000fffffff1ffffffff0000000600000000",
            INIT_05 => X"ffffffe8ffffffffffffffe9fffffffffffffffeffffffffffffffd8ffffffff",
            INIT_06 => X"ffffffaaffffffffffffffb5ffffffffffffffc2ffffffffffffffe4ffffffff",
            INIT_07 => X"0000004900000000ffffffe8ffffffff00000011000000000000003000000000",
            INIT_08 => X"0000003b000000000000006800000000ffffffdeffffffff0000005700000000",
            INIT_09 => X"0000002000000000fffffff9ffffffff0000001e000000000000001600000000",
            INIT_0A => X"000000540000000000000041000000000000000b000000000000002300000000",
            INIT_0B => X"ffffffdeffffffffffffffdbffffffff0000004a000000000000004600000000",
            INIT_0C => X"0000000500000000ffffffd2ffffffffffffffd7ffffffff0000000400000000",
            INIT_0D => X"ffffffebffffffff0000001a00000000ffffffdcffffffffffffffdfffffffff",
            INIT_0E => X"fffffff0ffffffff0000001100000000ffffffd6ffffffffffffffc5ffffffff",
            INIT_0F => X"000000340000000000000043000000000000005b000000000000000c00000000",
            INIT_10 => X"ffffffe9ffffffffffffffe8ffffffffffffffdfffffffffffffffb5ffffffff",
            INIT_11 => X"00000023000000000000000200000000ffffffbfffffffffffffffb6ffffffff",
            INIT_12 => X"fffffffcffffffffffffffd5ffffffffffffffe9ffffffff0000000800000000",
            INIT_13 => X"0000001b000000000000000300000000ffffffe9fffffffffffffffaffffffff",
            INIT_14 => X"ffffffe0ffffffff0000001200000000fffffff8fffffffffffffff2ffffffff",
            INIT_15 => X"fffffffdffffffff00000008000000000000000d00000000ffffffe1ffffffff",
            INIT_16 => X"ffffffdbffffffff0000000c0000000000000024000000000000001200000000",
            INIT_17 => X"ffffffd8ffffffffffffffffffffffffffffffccffffffffffffffb6ffffffff",
            INIT_18 => X"000000000000000000000037000000000000001400000000ffffffc3ffffffff",
            INIT_19 => X"ffffffe5ffffffffffffffefffffffffffffffd1ffffffff0000000200000000",
            INIT_1A => X"0000000d000000000000001c00000000fffffff7fffffffffffffff3ffffffff",
            INIT_1B => X"0000001e000000000000001b0000000000000015000000000000001400000000",
            INIT_1C => X"ffffffccffffffff0000001500000000ffffffeeffffffffffffffedffffffff",
            INIT_1D => X"00000000000000000000000b00000000ffffffdaffffffffffffffc1ffffffff",
            INIT_1E => X"00000011000000000000003600000000fffffff3ffffffff0000004400000000",
            INIT_1F => X"0000001a00000000000000410000000000000066000000000000001500000000",
            INIT_20 => X"00000053000000000000001a0000000000000029000000000000001500000000",
            INIT_21 => X"0000003a000000000000001e0000000000000024000000000000004100000000",
            INIT_22 => X"0000000500000000fffffff1ffffffff00000017000000000000000f00000000",
            INIT_23 => X"0000001400000000fffffff3fffffffffffffff7ffffffff0000000800000000",
            INIT_24 => X"ffffffb7ffffffffffffffc5ffffffffffffffeeffffffff0000001900000000",
            INIT_25 => X"0000001400000000ffffffe8fffffffffffffffeffffffff0000000d00000000",
            INIT_26 => X"ffffffd6ffffffffffffffd1ffffffff00000034000000000000003c00000000",
            INIT_27 => X"ffffffdffffffffffffffff1fffffffffffffffbffffffffffffffb9ffffffff",
            INIT_28 => X"ffffffceffffffff00000017000000000000002b000000000000002300000000",
            INIT_29 => X"fffffff4ffffffffffffffd8ffffffff00000033000000000000000800000000",
            INIT_2A => X"0000000e00000000ffffffd7ffffffffffffffc6ffffffff0000004400000000",
            INIT_2B => X"0000003d00000000000000080000000000000034000000000000004500000000",
            INIT_2C => X"0000004400000000000000370000000000000087000000000000009c00000000",
            INIT_2D => X"ffffffcaffffffff0000000f000000000000000f000000000000008100000000",
            INIT_2E => X"fffffff7fffffffffffffff9ffffffff0000001b000000000000001500000000",
            INIT_2F => X"ffffffadffffffffffffffbaffffffff00000026000000000000003000000000",
            INIT_30 => X"ffffffe8ffffffffffffffd7ffffffff0000000e00000000ffffffceffffffff",
            INIT_31 => X"ffffffe2ffffffffffffffe4ffffffff00000007000000000000002c00000000",
            INIT_32 => X"ffffffcfffffffffffffffbcfffffffffffffffdffffffff0000000600000000",
            INIT_33 => X"ffffff8cffffffffffffffc1ffffffffffffffbdffffffffffffffaeffffffff",
            INIT_34 => X"ffffffd1fffffffffffffff0ffffffffffffffedffffffffffffffeaffffffff",
            INIT_35 => X"ffffffe4fffffffffffffff0fffffffffffffffbffffffffffffffe8ffffffff",
            INIT_36 => X"0000002900000000ffffffebffffffff0000000b000000000000002200000000",
            INIT_37 => X"fffffffaffffffff00000017000000000000000000000000fffffffdffffffff",
            INIT_38 => X"fffffff8fffffffffffffff6ffffffff0000001a000000000000000900000000",
            INIT_39 => X"00000000000000000000000000000000fffffffffffffffffffffff5ffffffff",
            INIT_3A => X"ffffffc0fffffffffffffffeffffffffffffffd8ffffffffffffffd3ffffffff",
            INIT_3B => X"ffffffe7ffffffffffffffcafffffffffffffff1ffffffffffffffa8ffffffff",
            INIT_3C => X"ffffffe8ffffffffffffffeeffffffffffffffdaffffffffffffffe0ffffffff",
            INIT_3D => X"ffffffe8ffffffffffffffc4ffffffffffffffedffffffffffffffe3ffffffff",
            INIT_3E => X"0000001000000000fffffff0ffffffffffffffd8ffffffffffffffeeffffffff",
            INIT_3F => X"ffffffdeffffffffffffffdbfffffffffffffff1ffffffff0000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001500000000ffffffddffffffffffffffc6ffffffffffffffe2ffffffff",
            INIT_41 => X"ffffffeaffffffffffffffd6fffffffffffffffcffffffff0000001f00000000",
            INIT_42 => X"00000030000000000000002500000000fffffff9ffffffff0000000200000000",
            INIT_43 => X"0000000c000000000000002f0000000000000006000000000000003a00000000",
            INIT_44 => X"000000250000000000000026000000000000002d000000000000004200000000",
            INIT_45 => X"ffffffe7ffffffff0000000c000000000000001400000000ffffffe9ffffffff",
            INIT_46 => X"0000001b00000000fffffffcffffffff0000000700000000fffffff4ffffffff",
            INIT_47 => X"0000000d00000000ffffffebfffffffffffffffcffffffffffffffefffffffff",
            INIT_48 => X"0000003700000000ffffffebffffffffffffffc6fffffffffffffffdffffffff",
            INIT_49 => X"fffffffeffffffff000000240000000000000002000000000000001700000000",
            INIT_4A => X"ffffffe4ffffffffffffffefffffffff0000002c000000000000001900000000",
            INIT_4B => X"0000001a00000000fffffff5ffffffffffffffc1ffffffffffffffe9ffffffff",
            INIT_4C => X"ffffffe2ffffffff0000001f000000000000001d00000000ffffffd0ffffffff",
            INIT_4D => X"fffffffefffffffffffffff0ffffffffffffffc9ffffffffffffffefffffffff",
            INIT_4E => X"fffffffeffffffff0000001700000000ffffffe9ffffffffffffffe8ffffffff",
            INIT_4F => X"ffffffaaffffffff0000000400000000fffffff0fffffffffffffff4ffffffff",
            INIT_50 => X"ffffffc4ffffffffffffff90fffffffffffffff5ffffffffffffffc1ffffffff",
            INIT_51 => X"ffffffe2ffffffffffffffe0ffffffffffffffb5ffffffff0000000100000000",
            INIT_52 => X"ffffffe2ffffffff00000039000000000000001e00000000ffffffdfffffffff",
            INIT_53 => X"ffffffdcffffffffffffffbfffffffff0000001f00000000ffffffffffffffff",
            INIT_54 => X"fffffffffffffffffffffffbffffffffffffffc8ffffffffffffffc4ffffffff",
            INIT_55 => X"ffffffcbfffffffffffffffcffffffffffffffedffffffffffffffe6ffffffff",
            INIT_56 => X"fffffff5ffffffffffffffcfffffffff0000000200000000fffffff4ffffffff",
            INIT_57 => X"0000002e000000000000003300000000ffffffd8ffffffff0000002300000000",
            INIT_58 => X"ffffffe5ffffffff0000001700000000ffffffe4ffffffff0000000400000000",
            INIT_59 => X"0000000900000000ffffffe5ffffffffffffffe9ffffffff0000000b00000000",
            INIT_5A => X"0000000000000000000000220000000000000020000000000000001200000000",
            INIT_5B => X"0000001800000000fffffff5ffffffff0000001a000000000000002700000000",
            INIT_5C => X"fffffffbfffffffffffffff3ffffffff00000019000000000000002500000000",
            INIT_5D => X"fffffffdffffffff0000000800000000ffffffeefffffffffffffff9ffffffff",
            INIT_5E => X"ffffffd9ffffffff0000000000000000ffffffdcffffffffffffffeeffffffff",
            INIT_5F => X"fffffff1fffffffffffffff7fffffffffffffff9ffffffff0000001100000000",
            INIT_60 => X"0000000800000000ffffffe4ffffffffffffffe1ffffffffffffffefffffffff",
            INIT_61 => X"ffffffdeffffffffffffffdeffffffff00000008000000000000000600000000",
            INIT_62 => X"fffffff7ffffffffffffffefffffffffffffffecffffffff0000000600000000",
            INIT_63 => X"0000001900000000000000410000000000000056000000000000001300000000",
            INIT_64 => X"fffffff4ffffffff0000001b0000000000000032000000000000000d00000000",
            INIT_65 => X"fffffff6ffffffff0000001600000000fffffff8ffffffffffffffefffffffff",
            INIT_66 => X"ffffffe5ffffffff0000001c000000000000000e00000000fffffff4ffffffff",
            INIT_67 => X"ffffff8affffffff00000028000000000000005c000000000000004400000000",
            INIT_68 => X"ffffff81ffffffffffffffc0ffffffffffffffacffffffffffffff8effffffff",
            INIT_69 => X"ffffffbcffffffffffffffbfffffffffffffffcdffffffffffffffabffffffff",
            INIT_6A => X"fffffffaffffffff0000001a0000000000000015000000000000001000000000",
            INIT_6B => X"0000001b00000000ffffffffffffffff0000000800000000fffffffaffffffff",
            INIT_6C => X"0000000000000000ffffffccffffffffffffffeaffffffffffffffe7ffffffff",
            INIT_6D => X"ffffffd3fffffffffffffff7ffffffffffffffe5ffffffffffffffc6ffffffff",
            INIT_6E => X"00000013000000000000000f00000000fffffffaffffffffffffffe2ffffffff",
            INIT_6F => X"fffffff5ffffffff000000140000000000000006000000000000001700000000",
            INIT_70 => X"0000001e00000000ffffffedffffffffffffffeeffffffffffffffedffffffff",
            INIT_71 => X"0000002a000000000000002a00000000fffffff4ffffffff0000000d00000000",
            INIT_72 => X"0000002400000000000000120000000000000028000000000000001f00000000",
            INIT_73 => X"0000000300000000000000050000000000000017000000000000000200000000",
            INIT_74 => X"000000460000000000000025000000000000001c000000000000001200000000",
            INIT_75 => X"00000024000000000000003d000000000000003a000000000000003500000000",
            INIT_76 => X"0000002d00000000000000180000000000000031000000000000001d00000000",
            INIT_77 => X"ffffffeaffffffffffffffdaffffffff00000018000000000000002900000000",
            INIT_78 => X"ffffffe3ffffffffffffffecffffffff0000000300000000ffffffe9ffffffff",
            INIT_79 => X"fffffffafffffffffffffff3ffffffffffffffebffffffffffffffd8ffffffff",
            INIT_7A => X"ffffffaeffffffffffffffc9ffffffffffffffe8ffffffffffffffbaffffffff",
            INIT_7B => X"ffffffd6ffffffffffffffcbffffffffffffffd7ffffffffffffffb7ffffffff",
            INIT_7C => X"fffffffaffffffff000000340000000000000008000000000000000500000000",
            INIT_7D => X"ffffffdbffffffff000000020000000000000027000000000000002800000000",
            INIT_7E => X"fffffff3ffffffff00000011000000000000001100000000ffffffddffffffff",
            INIT_7F => X"ffffffeefffffffffffffff1ffffffffffffffe3ffffffff0000001500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE5;


    MEM_IWGHT_LAYER1_INSTANCE6 : if BRAM_NAME = "iwght_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000028000000000000001400000000fffffffefffffffffffffffcffffffff",
            INIT_01 => X"fffffff2ffffffffffffffecfffffffffffffff0ffffffff0000002000000000",
            INIT_02 => X"fffffff4fffffffffffffffcfffffffffffffff4ffffffffffffffefffffffff",
            INIT_03 => X"ffffffe1fffffffffffffffcffffffff00000014000000000000001d00000000",
            INIT_04 => X"ffffffeeffffffffffffffdafffffffffffffff6ffffffff0000001800000000",
            INIT_05 => X"00000023000000000000001b000000000000001d000000000000002100000000",
            INIT_06 => X"ffffffddffffffff000000040000000000000024000000000000000b00000000",
            INIT_07 => X"000000280000000000000019000000000000000800000000fffffff2ffffffff",
            INIT_08 => X"0000003100000000000000470000000000000039000000000000002600000000",
            INIT_09 => X"0000002f000000000000002b000000000000001e000000000000001c00000000",
            INIT_0A => X"0000002b0000000000000032000000000000004100000000fffffffdffffffff",
            INIT_0B => X"000000130000000000000004000000000000001c00000000ffffffe1ffffffff",
            INIT_0C => X"fffffffdffffffffffffffd0ffffffff0000001500000000fffffffcffffffff",
            INIT_0D => X"0000002200000000ffffffeffffffffffffffff3ffffffffffffffe7ffffffff",
            INIT_0E => X"00000016000000000000000e0000000000000018000000000000001700000000",
            INIT_0F => X"ffffffffffffffffffffffefffffffff0000000400000000ffffffe1ffffffff",
            INIT_10 => X"0000000c0000000000000000000000000000001800000000fffffff2ffffffff",
            INIT_11 => X"fffffff7fffffffffffffff8ffffffffffffffd4fffffffffffffffaffffffff",
            INIT_12 => X"0000001100000000fffffffdffffffffffffffebffffffff0000001000000000",
            INIT_13 => X"fffffff6fffffffffffffff7fffffffffffffff6ffffffff0000001d00000000",
            INIT_14 => X"000000460000000000000003000000000000000e00000000fffffffaffffffff",
            INIT_15 => X"00000068000000000000003f000000000000002f000000000000004000000000",
            INIT_16 => X"0000007600000000000000520000000000000049000000000000004600000000",
            INIT_17 => X"000000180000000000000025000000000000001c000000000000001000000000",
            INIT_18 => X"0000001f0000000000000007000000000000004e000000000000003100000000",
            INIT_19 => X"ffffffd9ffffffffffffffe1ffffffffffffffdaffffffff0000002400000000",
            INIT_1A => X"0000001400000000ffffffe6ffffffffffffffdeffffffff0000000000000000",
            INIT_1B => X"0000003b000000000000002e000000000000000900000000fffffff0ffffffff",
            INIT_1C => X"fffffffeffffffff0000000000000000ffffffe9ffffffff0000002f00000000",
            INIT_1D => X"0000000600000000ffffffd7ffffffffffffffd0fffffffffffffff1ffffffff",
            INIT_1E => X"0000001f000000000000001c0000000000000012000000000000002800000000",
            INIT_1F => X"0000003f000000000000001e0000000000000011000000000000002300000000",
            INIT_20 => X"ffffffc7ffffffff000000260000000000000032000000000000002600000000",
            INIT_21 => X"00000015000000000000001100000000ffffffbeffffffffffffffb3ffffffff",
            INIT_22 => X"ffffffd1fffffffffffffff1ffffffff00000000000000000000001900000000",
            INIT_23 => X"ffffffecffffffff0000000300000000ffffffdcfffffffffffffff5ffffffff",
            INIT_24 => X"0000000c00000000ffffffe6ffffffff0000000b00000000ffffffe3ffffffff",
            INIT_25 => X"ffffffd9fffffffffffffffaffffffffffffffd7ffffffff0000000600000000",
            INIT_26 => X"0000001b00000000ffffffe3ffffffff0000000700000000ffffffe7ffffffff",
            INIT_27 => X"fffffff0ffffffff00000005000000000000000b000000000000001c00000000",
            INIT_28 => X"ffffffe7ffffffff00000018000000000000000300000000fffffff1ffffffff",
            INIT_29 => X"ffffff9effffffff0000001100000000fffffff7ffffffff0000001300000000",
            INIT_2A => X"0000001e000000000000001400000000ffffff99ffffffffffffff91ffffffff",
            INIT_2B => X"0000000e00000000ffffffecfffffffffffffff9ffffffff0000000b00000000",
            INIT_2C => X"0000000e00000000ffffffd7ffffffffffffffb5ffffffffffffffdeffffffff",
            INIT_2D => X"0000000f000000000000000f00000000fffffff3ffffffff0000001d00000000",
            INIT_2E => X"ffffffc7ffffffffffffffb7ffffffffffffffc3ffffffff0000002b00000000",
            INIT_2F => X"ffffffb0ffffffff00000004000000000000000e00000000ffffffebffffffff",
            INIT_30 => X"00000042000000000000004c00000000ffffffecffffffffffffffc9ffffffff",
            INIT_31 => X"fffffff9ffffffffffffffcdffffffffffffffd0ffffffff0000000f00000000",
            INIT_32 => X"fffffff1ffffffff000000090000000000000016000000000000001f00000000",
            INIT_33 => X"fffffff6ffffffff0000001c000000000000000d000000000000001600000000",
            INIT_34 => X"ffffffcdffffffffffffffcfffffffffffffffccffffffff0000000e00000000",
            INIT_35 => X"00000002000000000000001b000000000000003d000000000000000700000000",
            INIT_36 => X"ffffffd8ffffffffffffffdffffffffffffffff1ffffffffffffffefffffffff",
            INIT_37 => X"fffffff2fffffffffffffff8ffffffff0000000000000000fffffffcffffffff",
            INIT_38 => X"0000004100000000ffffffe4ffffffffffffffeaffffffffffffffd7ffffffff",
            INIT_39 => X"ffffff80ffffffffffffff94ffffffff00000013000000000000003500000000",
            INIT_3A => X"000000150000000000000065000000000000003200000000ffffffdcffffffff",
            INIT_3B => X"ffffffe7ffffffff0000003d0000000000000002000000000000002500000000",
            INIT_3C => X"fffffffdffffffff00000026000000000000001900000000ffffffd4ffffffff",
            INIT_3D => X"00000024000000000000001c000000000000001f000000000000002600000000",
            INIT_3E => X"fffffff9ffffffff00000018000000000000002f000000000000003000000000",
            INIT_3F => X"0000001f000000000000001c00000000ffffffd9fffffffffffffff9ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000600000000ffffffedffffffffffffffebffffffff0000000600000000",
            INIT_41 => X"00000042000000000000001e000000000000000200000000fffffff5ffffffff",
            INIT_42 => X"000000390000000000000050000000000000002d000000000000001800000000",
            INIT_43 => X"0000001c00000000000000120000000000000013000000000000001f00000000",
            INIT_44 => X"0000001900000000ffffffeaffffffffffffffe9ffffffff0000001800000000",
            INIT_45 => X"00000010000000000000000b00000000ffffffeefffffffffffffff4ffffffff",
            INIT_46 => X"ffffffcfffffffffffffffd6ffffffffffffffc9ffffffffffffffe9ffffffff",
            INIT_47 => X"0000001000000000ffffffdafffffffffffffff5ffffffff0000000600000000",
            INIT_48 => X"00000015000000000000000b00000000ffffffebffffffff0000000000000000",
            INIT_49 => X"fffffff3fffffffffffffff4ffffffff0000000c00000000ffffffe9ffffffff",
            INIT_4A => X"fffffffefffffffffffffffdffffffff00000009000000000000001d00000000",
            INIT_4B => X"ffffffefffffffff0000002e00000000fffffffaffffffffffffffecffffffff",
            INIT_4C => X"00000011000000000000002f000000000000003a00000000ffffffecffffffff",
            INIT_4D => X"0000000000000000ffffffeefffffffffffffff1ffffffff0000000400000000",
            INIT_4E => X"ffffffe3ffffffff0000000600000000fffffff8ffffffffffffffd7ffffffff",
            INIT_4F => X"fffffff2ffffffffffffffefffffffff00000001000000000000000800000000",
            INIT_50 => X"ffffffc3ffffffffffffffd0ffffffffffffff98ffffffffffffffa1ffffffff",
            INIT_51 => X"ffffff5affffffffffffff54ffffffff0000000400000000ffffffffffffffff",
            INIT_52 => X"ffffff58ffffffffffffff3fffffffffffffff30ffffffffffffff9affffffff",
            INIT_53 => X"0000001f00000000ffffff60ffffffffffffff0affffffffffffff90ffffffff",
            INIT_54 => X"00000027000000000000001a0000000000000004000000000000000000000000",
            INIT_55 => X"000000310000000000000042000000000000005200000000ffffffe5ffffffff",
            INIT_56 => X"0000000e00000000fffffffdffffffff0000001f00000000ffffffeaffffffff",
            INIT_57 => X"ffffffecffffffff0000000b000000000000001500000000ffffffffffffffff",
            INIT_58 => X"fffffff0ffffffffffffffe2ffffffff00000018000000000000000200000000",
            INIT_59 => X"0000000b00000000ffffffeefffffffffffffff2ffffffff0000000d00000000",
            INIT_5A => X"ffffffdeffffffff000000140000000000000000000000000000002300000000",
            INIT_5B => X"ffffffeaffffffff0000000300000000fffffffdffffffffffffffebffffffff",
            INIT_5C => X"ffffffe0ffffffff000000200000000000000036000000000000001c00000000",
            INIT_5D => X"ffffff52ffffffffffffff66ffffffffffffffceffffffffffffffbdffffffff",
            INIT_5E => X"ffffffc0ffffffffffffffacffffffffffffff91ffffffffffffff88ffffffff",
            INIT_5F => X"0000000700000000ffffffc2ffffffffffffffbeffffffffffffffecffffffff",
            INIT_60 => X"0000003f00000000ffffffe6ffffffff00000000000000000000000400000000",
            INIT_61 => X"fffffff7fffffffffffffff6ffffffffffffffe2ffffffff0000003f00000000",
            INIT_62 => X"00000016000000000000000a000000000000002c000000000000003700000000",
            INIT_63 => X"ffffffeffffffffffffffff3ffffffff0000003e000000000000004a00000000",
            INIT_64 => X"0000000100000000000000080000000000000013000000000000000a00000000",
            INIT_65 => X"0000002b00000000000000030000000000000012000000000000002d00000000",
            INIT_66 => X"00000040000000000000002f0000000000000058000000000000004d00000000",
            INIT_67 => X"0000007000000000000000500000000000000054000000000000003200000000",
            INIT_68 => X"0000000d0000000000000012000000000000002300000000ffffffefffffffff",
            INIT_69 => X"0000001000000000fffffff5ffffffffffffffffffffffff0000001d00000000",
            INIT_6A => X"ffffffffffffffff0000001f00000000fffffff4ffffffff0000000e00000000",
            INIT_6B => X"ffffffeeffffffff0000000b000000000000002c000000000000000b00000000",
            INIT_6C => X"0000000000000000fffffff2ffffffff00000014000000000000001300000000",
            INIT_6D => X"00000002000000000000001e0000000000000017000000000000001c00000000",
            INIT_6E => X"0000001400000000fffffff4ffffffffffffffe1ffffffffffffffeaffffffff",
            INIT_6F => X"ffffffe6ffffffff000000070000000000000000000000000000001500000000",
            INIT_70 => X"ffffffe7ffffffffffffffb4ffffffffffffffcbfffffffffffffffaffffffff",
            INIT_71 => X"fffffff3ffffffffffffffe3ffffffffffffffebffffffff0000000600000000",
            INIT_72 => X"fffffff6ffffffff0000000d00000000ffffffeaffffffff0000000b00000000",
            INIT_73 => X"0000001000000000fffffff3ffffffff00000002000000000000000000000000",
            INIT_74 => X"0000002300000000000000370000000000000065000000000000001e00000000",
            INIT_75 => X"ffffffd3ffffffffffffffc5ffffffff00000014000000000000004400000000",
            INIT_76 => X"ffffffc9ffffffffffffffc9ffffffffffffffc9ffffffffffffffb8ffffffff",
            INIT_77 => X"00000035000000000000000100000000fffffffdffffffff0000001200000000",
            INIT_78 => X"0000003300000000ffffffe2ffffffff00000015000000000000004500000000",
            INIT_79 => X"0000002c00000000000000250000000000000041000000000000002a00000000",
            INIT_7A => X"ffffffefffffffffffffffd9ffffffffffffffeefffffffffffffffcffffffff",
            INIT_7B => X"fffffff4ffffffff0000001e000000000000001e00000000fffffff9ffffffff",
            INIT_7C => X"fffffff5ffffffffffffffe2ffffffff00000015000000000000000a00000000",
            INIT_7D => X"ffffffc3fffffffffffffff1fffffffffffffff5ffffffffffffffe8ffffffff",
            INIT_7E => X"ffffffefffffffff0000001b00000000ffffffe8ffffffffffffffd7ffffffff",
            INIT_7F => X"0000000b00000000ffffffecffffffff0000000000000000ffffffffffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE6;


    MEM_IWGHT_LAYER1_INSTANCE7 : if BRAM_NAME = "iwght_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe1ffffffffffffffd5fffffffffffffff9ffffffff0000000500000000",
            INIT_01 => X"00000022000000000000001700000000ffffffe4ffffffff0000000200000000",
            INIT_02 => X"0000002400000000000000410000000000000025000000000000002a00000000",
            INIT_03 => X"00000037000000000000000900000000fffffff8ffffffff0000002600000000",
            INIT_04 => X"00000047000000000000003500000000ffffffd3ffffffff0000001700000000",
            INIT_05 => X"0000003f0000000000000039000000000000005500000000ffffffddffffffff",
            INIT_06 => X"0000002a000000000000003d000000000000004a000000000000004600000000",
            INIT_07 => X"0000002200000000fffffff7ffffffff0000001a00000000fffffffbffffffff",
            INIT_08 => X"0000000600000000ffffffe9fffffffffffffff5ffffffff0000000000000000",
            INIT_09 => X"0000004b00000000ffffffe1ffffffffffffffdcffffffffffffffd7ffffffff",
            INIT_0A => X"0000005a00000000000000380000000000000038000000000000004d00000000",
            INIT_0B => X"0000003b000000000000003b0000000000000026000000000000003b00000000",
            INIT_0C => X"ffffffe1fffffffffffffffdffffffffffffffe6ffffffffffffffd8ffffffff",
            INIT_0D => X"0000002700000000ffffffecffffffff00000021000000000000000000000000",
            INIT_0E => X"0000002400000000fffffffeffffffff00000003000000000000002500000000",
            INIT_0F => X"fffffffdffffffff0000001d000000000000000a00000000ffffffedffffffff",
            INIT_10 => X"ffffffeeffffffffffffffc1fffffffffffffff1fffffffffffffffcffffffff",
            INIT_11 => X"ffffffdbffffffff0000001b00000000ffffffe8ffffffffffffffddffffffff",
            INIT_12 => X"0000000300000000000000230000000000000014000000000000000400000000",
            INIT_13 => X"0000000700000000ffffffe6ffffffff0000000500000000ffffffe1ffffffff",
            INIT_14 => X"000000290000000000000006000000000000001900000000fffffffcffffffff",
            INIT_15 => X"ffffffd3fffffffffffffff3fffffffffffffff4ffffffffffffffd2ffffffff",
            INIT_16 => X"ffffffdbffffffffffffffbfffffffffffffffefffffffffffffffeeffffffff",
            INIT_17 => X"00000034000000000000002e000000000000002900000000fffffffcffffffff",
            INIT_18 => X"fffffff8ffffffff00000011000000000000001a000000000000003000000000",
            INIT_19 => X"0000003a00000000000000480000000000000011000000000000002d00000000",
            INIT_1A => X"fffffffeffffffff000000140000000000000048000000000000003d00000000",
            INIT_1B => X"fffffffafffffffffffffffffffffffffffffff6ffffffff0000004d00000000",
            INIT_1C => X"fffffff5fffffffffffffff5ffffffffffffffe8ffffffff0000001400000000",
            INIT_1D => X"0000001800000000fffffff5fffffffffffffffdfffffffffffffff6ffffffff",
            INIT_1E => X"0000000c000000000000000400000000ffffffefffffffff0000001200000000",
            INIT_1F => X"ffffffe3fffffffffffffff5ffffffffffffffe8ffffffff0000001400000000",
            INIT_20 => X"0000001e000000000000001500000000ffffffdcffffffff0000001b00000000",
            INIT_21 => X"0000000000000000fffffff2ffffffffffffffe8ffffffff0000000300000000",
            INIT_22 => X"0000001400000000ffffffe7fffffffffffffff1ffffffff0000001300000000",
            INIT_23 => X"0000002a00000000ffffffffffffffffffffffdcffffffff0000000200000000",
            INIT_24 => X"0000003200000000ffffffebfffffffffffffffaffffffff0000000700000000",
            INIT_25 => X"0000005f0000000000000048000000000000002b000000000000005b00000000",
            INIT_26 => X"00000014000000000000002e0000000000000023000000000000002800000000",
            INIT_27 => X"00000028000000000000002f000000000000000b000000000000001300000000",
            INIT_28 => X"00000091000000000000006c000000000000000b000000000000004c00000000",
            INIT_29 => X"00000048000000000000002d000000000000000f000000000000003d00000000",
            INIT_2A => X"000000080000000000000038000000000000003e000000000000001800000000",
            INIT_2B => X"ffffffd9ffffffffffffffeaffffffff0000000d000000000000002b00000000",
            INIT_2C => X"00000007000000000000000f0000000000000010000000000000000600000000",
            INIT_2D => X"fffffff7ffffffff0000001000000000fffffff6ffffffff0000002700000000",
            INIT_2E => X"fffffff8ffffffff00000002000000000000002100000000ffffffe0ffffffff",
            INIT_2F => X"0000002d000000000000000c0000000000000025000000000000003000000000",
            INIT_30 => X"fffffff5ffffffff0000002100000000ffffffddfffffffffffffff5ffffffff",
            INIT_31 => X"0000000800000000fffffffeffffffffffffffdbffffffffffffffe8ffffffff",
            INIT_32 => X"fffffff0ffffffff0000000200000000ffffffeaffffffffffffffd5ffffffff",
            INIT_33 => X"ffffffb0fffffffffffffff3ffffffffffffffe9ffffffffffffffdeffffffff",
            INIT_34 => X"ffffffecfffffffffffffffbffffffffffffffc2ffffffffffffffe2ffffffff",
            INIT_35 => X"ffffffeaffffffffffffffe8ffffffff0000000600000000fffffff2ffffffff",
            INIT_36 => X"00000000000000000000000d00000000fffffffafffffffffffffff7ffffffff",
            INIT_37 => X"0000001900000000fffffff5ffffffff00000015000000000000001700000000",
            INIT_38 => X"000000090000000000000019000000000000001a00000000ffffffe5ffffffff",
            INIT_39 => X"000000070000000000000025000000000000000e00000000ffffffebffffffff",
            INIT_3A => X"00000015000000000000001e000000000000000600000000fffffff0ffffffff",
            INIT_3B => X"fffffff6ffffffffffffffdeffffffffffffffd6fffffffffffffff5ffffffff",
            INIT_3C => X"0000000d00000000ffffffdaffffffffffffffdeffffffffffffffd9ffffffff",
            INIT_3D => X"ffffffe4ffffffffffffffceffffffffffffffe7ffffffff0000002100000000",
            INIT_3E => X"0000000600000000ffffffb2ffffffffffffffc6ffffffffffffffe8ffffffff",
            INIT_3F => X"0000000a00000000ffffffcaffffffffffffffb7ffffffffffffffc7ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000047000000000000004e0000000000000018000000000000003100000000",
            INIT_41 => X"0000006700000000000000630000000000000063000000000000003800000000",
            INIT_42 => X"fffffffafffffffffffffff8ffffffffffffffffffffffffffffffe4ffffffff",
            INIT_43 => X"0000000d000000000000001a00000000ffffffedffffffff0000000e00000000",
            INIT_44 => X"fffffff9ffffffff00000022000000000000001500000000ffffffefffffffff",
            INIT_45 => X"0000001b0000000000000008000000000000001c000000000000003000000000",
            INIT_46 => X"ffffffccfffffffffffffff7ffffffff00000037000000000000003100000000",
            INIT_47 => X"fffffff3fffffffffffffffaffffffffffffffe6ffffffff0000000400000000",
            INIT_48 => X"ffffffe4ffffffffffffffe7ffffffffffffffc9ffffffffffffffbfffffffff",
            INIT_49 => X"ffffffc4ffffffffffffffecffffffff0000001500000000ffffffdfffffffff",
            INIT_4A => X"ffffffebffffffff0000002000000000fffffff5ffffffffffffffe9ffffffff",
            INIT_4B => X"ffffffd4ffffffffffffffeeffffffffffffffc2ffffffffffffffe7ffffffff",
            INIT_4C => X"ffffffdaffffffff0000000200000000fffffffeffffffffffffffb0ffffffff",
            INIT_4D => X"ffffffc4ffffffffffffffaeffffffffffffffb8fffffffffffffffbffffffff",
            INIT_4E => X"ffffffa5ffffffffffffffc8ffffffffffffff98ffffffffffffffbbffffffff",
            INIT_4F => X"ffffffebffffffff0000000f00000000ffffffa0ffffffffffffff95ffffffff",
            INIT_50 => X"0000000f00000000000000050000000000000009000000000000002600000000",
            INIT_51 => X"00000053000000000000001a000000000000000d000000000000000500000000",
            INIT_52 => X"00000000000000000000002a000000000000005d000000000000002300000000",
            INIT_53 => X"0000001700000000000000310000000000000052000000000000004000000000",
            INIT_54 => X"0000001500000000ffffffe7ffffffffffffffe2ffffffff0000000d00000000",
            INIT_55 => X"00000030000000000000000a00000000fffffffeffffffff0000002400000000",
            INIT_56 => X"0000000100000000ffffffe5fffffffffffffff3ffffffff0000000100000000",
            INIT_57 => X"0000000e00000000ffffffd7fffffffffffffff8fffffffffffffff2ffffffff",
            INIT_58 => X"fffffffaffffffff0000001700000000ffffffdbffffffffffffffe4ffffffff",
            INIT_59 => X"000000050000000000000028000000000000001d00000000ffffffe7ffffffff",
            INIT_5A => X"0000001e0000000000000007000000000000000e000000000000003700000000",
            INIT_5B => X"0000003000000000fffffffcfffffffffffffff0fffffffffffffffcffffffff",
            INIT_5C => X"00000025000000000000002600000000ffffffffffffffffffffffecffffffff",
            INIT_5D => X"ffffffd5ffffffffffffffe5fffffffffffffffbffffffffffffffe6ffffffff",
            INIT_5E => X"ffffffe9ffffffffffffffddffffffffffffffe5ffffffff0000000700000000",
            INIT_5F => X"ffffffd3ffffffffffffffafffffffffffffffb0ffffffffffffffedffffffff",
            INIT_60 => X"0000003700000000ffffff9fffffffffffffffdffffffffffffffff1ffffffff",
            INIT_61 => X"ffffff90ffffffffffffffe4fffffffffffffff9ffffffff0000004700000000",
            INIT_62 => X"ffffff47ffffffffffffffbbffffffff0000002d00000000ffffff57ffffffff",
            INIT_63 => X"0000001400000000ffffffa2ffffffff00000027000000000000003d00000000",
            INIT_64 => X"00000026000000000000001700000000fffffff5ffffffff0000000000000000",
            INIT_65 => X"fffffff1ffffffff00000039000000000000002600000000fffffff2ffffffff",
            INIT_66 => X"ffffffebffffffff0000000500000000fffffffbfffffffffffffff5ffffffff",
            INIT_67 => X"0000000f00000000ffffffebffffffff0000000d00000000fffffff1ffffffff",
            INIT_68 => X"ffffffd4fffffffffffffff9fffffffffffffff7ffffffff0000000500000000",
            INIT_69 => X"000000220000000000000011000000000000001d000000000000002e00000000",
            INIT_6A => X"0000000100000000ffffffe3ffffffff00000001000000000000002100000000",
            INIT_6B => X"0000000b00000000ffffffecfffffffffffffff3fffffffffffffff4ffffffff",
            INIT_6C => X"ffffffa5ffffffff0000003000000000fffffff7ffffffff0000000700000000",
            INIT_6D => X"ffffff8bfffffffffffffffeffffffffffffffb3ffffffffffffff96ffffffff",
            INIT_6E => X"fffffff9ffffffff00000008000000000000003b00000000ffffffa1ffffffff",
            INIT_6F => X"ffffffb3ffffffff0000002b000000000000001000000000ffffffefffffffff",
            INIT_70 => X"fffffff6fffffffffffffff1ffffffff0000002a00000000ffffffe7ffffffff",
            INIT_71 => X"00000008000000000000001100000000ffffffe3ffffffff0000003200000000",
            INIT_72 => X"ffffffddffffffff000000310000000000000008000000000000000200000000",
            INIT_73 => X"ffffffefffffffff000000140000000000000031000000000000002e00000000",
            INIT_74 => X"ffffffd2fffffffffffffffbffffffff0000001c00000000ffffffd5ffffffff",
            INIT_75 => X"000000440000000000000012000000000000001c000000000000001b00000000",
            INIT_76 => X"00000010000000000000000b0000000000000055000000000000003000000000",
            INIT_77 => X"0000000e000000000000000c000000000000000f000000000000000400000000",
            INIT_78 => X"fffffffeffffffffffffffdcffffffffffffffecffffffffffffffc5ffffffff",
            INIT_79 => X"ffffffd8fffffffffffffffaffffffffffffffeffffffffffffffff1ffffffff",
            INIT_7A => X"0000000a0000000000000014000000000000002c000000000000001700000000",
            INIT_7B => X"0000002700000000000000180000000000000034000000000000002f00000000",
            INIT_7C => X"ffffffb6ffffffffffffffe3ffffffff00000006000000000000002a00000000",
            INIT_7D => X"ffffffc7ffffffffffffffd5ffffffffffffffc6ffffffffffffffebffffffff",
            INIT_7E => X"ffffffd6ffffffff0000000900000000ffffffdeffffffffffffffe3ffffffff",
            INIT_7F => X"0000000900000000ffffffe0fffffffffffffff7ffffffff0000000a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE7;


    MEM_IWGHT_LAYER1_INSTANCE8 : if BRAM_NAME = "iwght_layer1_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff5ffffffff0000000100000000fffffffeffffffffffffffe2ffffffff",
            INIT_01 => X"0000002f00000000000000100000000000000024000000000000001000000000",
            INIT_02 => X"000000290000000000000018000000000000002d000000000000002400000000",
            INIT_03 => X"0000003900000000fffffffdffffffff00000019000000000000002500000000",
            INIT_04 => X"0000001f000000000000002a00000000fffffff6fffffffffffffffdffffffff",
            INIT_05 => X"0000000800000000ffffffe7ffffffff00000024000000000000002500000000",
            INIT_06 => X"0000001b00000000fffffff8fffffffffffffff2ffffffff0000000c00000000",
            INIT_07 => X"ffffffdefffffffffffffff1ffffffff0000000600000000ffffffecffffffff",
            INIT_08 => X"ffffffddffffffffffffffe5ffffffff0000000a00000000ffffffe0ffffffff",
            INIT_09 => X"0000000f00000000ffffffe5fffffffffffffff7ffffffff0000001900000000",
            INIT_0A => X"00000008000000000000001100000000ffffffe9fffffffffffffff6ffffffff",
            INIT_0B => X"0000000b00000000ffffffeaffffffffffffffecffffffffffffffffffffffff",
            INIT_0C => X"fffffff7ffffffff00000014000000000000000d000000000000000c00000000",
            INIT_0D => X"00000020000000000000001900000000fffffffeffffffff0000001300000000",
            INIT_0E => X"0000000800000000ffffffe2ffffffff0000001e000000000000003100000000",
            INIT_0F => X"0000000a00000000fffffffbffffffff0000001b00000000fffffff3ffffffff",
            INIT_10 => X"ffffffedfffffffffffffffefffffffffffffff8ffffffff0000002d00000000",
            INIT_11 => X"ffffffe9fffffffffffffffdffffffffffffffddffffffffffffffd4ffffffff",
            INIT_12 => X"fffffffefffffffffffffffdffffffff0000001b000000000000000300000000",
            INIT_13 => X"ffffffe4ffffffff0000000100000000fffffff3ffffffff0000000d00000000",
            INIT_14 => X"fffffff2ffffffff0000000c00000000fffffffbffffffff0000002400000000",
            INIT_15 => X"ffffffd4ffffffffffffffdbfffffffffffffffdffffffff0000001200000000",
            INIT_16 => X"ffffffecffffffffffffffdeffffffffffffffdcffffffffffffffdeffffffff",
            INIT_17 => X"ffffffdcffffffffffffffe7ffffffff0000001300000000ffffffe6ffffffff",
            INIT_18 => X"0000000600000000000000100000000000000000000000000000000e00000000",
            INIT_19 => X"ffffff76ffffffff0000001700000000ffffffedffffffff0000002300000000",
            INIT_1A => X"ffffff86ffffffffffffff9effffffffffffff8affffffffffffff60ffffffff",
            INIT_1B => X"ffffff96ffffffffffffffaaffffffffffffffa3ffffffffffffffbfffffffff",
            INIT_1C => X"0000001200000000ffffff74ffffffffffffff7bffffffffffffff87ffffffff",
            INIT_1D => X"00000045000000000000001b0000000000000034000000000000001100000000",
            INIT_1E => X"ffffffc0fffffffffffffff5fffffffffffffffcffffffff0000004600000000",
            INIT_1F => X"0000002c0000000000000010000000000000001f000000000000001a00000000",
            INIT_20 => X"ffffffc9fffffffffffffffeffffffff0000002f000000000000000e00000000",
            INIT_21 => X"fffffff8ffffffff00000010000000000000000900000000ffffffdcffffffff",
            INIT_22 => X"ffffffc1ffffffff000000390000000000000027000000000000001500000000",
            INIT_23 => X"00000020000000000000002200000000ffffffc5ffffffffffffffc2ffffffff",
            INIT_24 => X"00000030000000000000000100000000fffffffbffffffff0000002300000000",
            INIT_25 => X"0000000000000000ffffff94ffffffffffffff81ffffffffffffffb5ffffffff",
            INIT_26 => X"0000004600000000000000360000000000000013000000000000000000000000",
            INIT_27 => X"000000630000000000000058000000000000005e000000000000003500000000",
            INIT_28 => X"ffffffdcffffffff00000016000000000000001500000000ffffffccffffffff",
            INIT_29 => X"ffffffe7ffffffffffffffe1ffffffffffffffd8ffffffffffffffdcffffffff",
            INIT_2A => X"ffffffcefffffffffffffffefffffffffffffff7ffffffff0000000800000000",
            INIT_2B => X"0000002a00000000ffffffc6ffffffffffffffd3ffffffff0000000900000000",
            INIT_2C => X"0000000b00000000ffffffecffffffff0000003d000000000000003300000000",
            INIT_2D => X"ffffffdeffffffffffffffdeffffffffffffffdfffffffff0000002100000000",
            INIT_2E => X"ffffffe7ffffffffffffffe3fffffffffffffff9fffffffffffffff9ffffffff",
            INIT_2F => X"ffffffe7ffffffff0000000300000000fffffffafffffffffffffffcffffffff",
            INIT_30 => X"0000001a000000000000004a0000000000000028000000000000000b00000000",
            INIT_31 => X"00000012000000000000000e000000000000000b00000000fffffff7ffffffff",
            INIT_32 => X"ffffffdaffffffffffffffdfffffffff0000000400000000fffffff5ffffffff",
            INIT_33 => X"00000007000000000000001f000000000000000300000000ffffffccffffffff",
            INIT_34 => X"000000510000000000000020000000000000003c000000000000003b00000000",
            INIT_35 => X"000000280000000000000024000000000000002a000000000000005000000000",
            INIT_36 => X"0000002600000000ffffffeffffffffffffffff9ffffffff0000005c00000000",
            INIT_37 => X"ffffffdaffffffffffffffdeffffffffffffffdffffffffffffffff4ffffffff",
            INIT_38 => X"ffffffe2ffffffff00000000000000000000002800000000ffffffafffffffff",
            INIT_39 => X"ffffffeeffffffffffffffe7ffffffffffffffecffffffffffffffd9ffffffff",
            INIT_3A => X"fffffff0ffffffff0000001e000000000000001c00000000ffffffeeffffffff",
            INIT_3B => X"ffffffcdffffffffffffffe2ffffffff0000001200000000fffffffaffffffff",
            INIT_3C => X"0000002e0000000000000032000000000000000000000000ffffffe0ffffffff",
            INIT_3D => X"ffffffd3ffffffff00000001000000000000001b000000000000001d00000000",
            INIT_3E => X"fffffffbffffffff0000001e00000000ffffffdaffffffffffffffa9ffffffff",
            INIT_3F => X"0000000800000000000000040000000000000013000000000000002900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000a00000000fffffffbffffffff00000007000000000000000000000000",
            INIT_41 => X"fffffff5ffffffff0000001f000000000000001400000000fffffffdffffffff",
            INIT_42 => X"fffffff7ffffffff0000002d000000000000004500000000fffffff1ffffffff",
            INIT_43 => X"0000000300000000fffffffcffffffff0000001600000000fffffff3ffffffff",
            INIT_44 => X"0000000500000000ffffffeeffffffffffffffe7ffffffffffffffecffffffff",
            INIT_45 => X"0000002000000000ffffffeeffffffff0000000500000000ffffffe4ffffffff",
            INIT_46 => X"fffffff2fffffffffffffff9ffffffff0000001d000000000000003000000000",
            INIT_47 => X"0000000300000000fffffff7ffffffffffffffedffffffffffffffeaffffffff",
            INIT_48 => X"fffffffafffffffffffffff0ffffffff00000019000000000000001000000000",
            INIT_49 => X"0000001a0000000000000010000000000000001c000000000000002f00000000",
            INIT_4A => X"000000150000000000000027000000000000000d000000000000002100000000",
            INIT_4B => X"ffffffebffffffff0000001b000000000000002d00000000fffffff2ffffffff",
            INIT_4C => X"ffffffe5ffffffff000000260000000000000021000000000000001d00000000",
            INIT_4D => X"ffffffafffffffffffffffb3ffffffff0000002000000000fffffffeffffffff",
            INIT_4E => X"ffffffb6ffffffffffffffc1ffffffffffffffa2ffffffffffffffbdffffffff",
            INIT_4F => X"ffffffb8ffffffff0000000400000000ffffffebffffffffffffffa3ffffffff",
            INIT_50 => X"ffffffceffffffffffffffd6ffffffffffffffbaffffffffffffffd0ffffffff",
            INIT_51 => X"ffffffc7ffffffff0000000200000000ffffffddfffffffffffffffaffffffff",
            INIT_52 => X"00000000000000000000000300000000ffffffeeffffffff0000000a00000000",
            INIT_53 => X"fffffff9ffffffffffffffe7ffffffff00000004000000000000000b00000000",
            INIT_54 => X"ffffffceffffffffffffffdcffffffff0000000900000000ffffffecffffffff",
            INIT_55 => X"0000002b00000000ffffffe7ffffffffffffffe1ffffffff0000001500000000",
            INIT_56 => X"0000001e000000000000003d00000000ffffffdbfffffffffffffff2ffffffff",
            INIT_57 => X"00000001000000000000000a00000000fffffffbffffffffffffffefffffffff",
            INIT_58 => X"ffffffe4ffffffffffffffe0ffffffff00000000000000000000002900000000",
            INIT_59 => X"0000002b000000000000000e00000000ffffffd1ffffffffffffffd3ffffffff",
            INIT_5A => X"ffffffdeffffffff0000000700000000ffffffd6ffffffff0000000600000000",
            INIT_5B => X"00000048000000000000000a000000000000000400000000fffffff3ffffffff",
            INIT_5C => X"0000002f0000000000000040000000000000002d000000000000000100000000",
            INIT_5D => X"0000004100000000000000150000000000000044000000000000006100000000",
            INIT_5E => X"0000000c000000000000003a0000000000000008000000000000002000000000",
            INIT_5F => X"ffffffdfffffffffffffffe3ffffffff0000000b000000000000000700000000",
            INIT_60 => X"fffffff8ffffffff0000001100000000fffffff1ffffffffffffffd8ffffffff",
            INIT_61 => X"ffffffd6fffffffffffffff7ffffffff00000012000000000000002000000000",
            INIT_62 => X"ffffffbcffffffffffffff95ffffffffffffffdcffffffffffffffc5ffffffff",
            INIT_63 => X"ffffffbdffffffffffffffb3ffffffffffffff9dffffffffffffffccffffffff",
            INIT_64 => X"fffffffaffffffff000000010000000000000011000000000000002100000000",
            INIT_65 => X"ffffffbafffffffffffffff7ffffffffffffffe4ffffffff0000001200000000",
            INIT_66 => X"fffffff2ffffffff0000000000000000ffffffffffffffffffffffafffffffff",
            INIT_67 => X"ffffffdafffffffffffffffcffffffffffffffdefffffffffffffffbffffffff",
            INIT_68 => X"00000003000000000000001e00000000fffffff0ffffffffffffffe1ffffffff",
            INIT_69 => X"ffffffb0ffffffffffffffc5ffffffffffffffd7fffffffffffffff8ffffffff",
            INIT_6A => X"0000002300000000ffffffb6ffffffffffffffb1ffffffffffffffedffffffff",
            INIT_6B => X"fffffff5ffffffff00000022000000000000000c000000000000002500000000",
            INIT_6C => X"ffffffeaffffffff00000009000000000000000f00000000fffffff4ffffffff",
            INIT_6D => X"0000004a00000000000000330000000000000042000000000000003100000000",
            INIT_6E => X"0000003e000000000000002a000000000000002c000000000000004600000000",
            INIT_6F => X"0000000600000000ffffffd2ffffffffffffffe5ffffffff0000001400000000",
            INIT_70 => X"fffffffdffffffffffffffc1fffffffffffffffbfffffffffffffff0ffffffff",
            INIT_71 => X"ffffffc4ffffffffffffffe8ffffffffffffffc3ffffffffffffffc4ffffffff",
            INIT_72 => X"fffffff4ffffffffffffffc2ffffffffffffffc8ffffffffffffffe3ffffffff",
            INIT_73 => X"00000044000000000000003f000000000000000700000000ffffffb9ffffffff",
            INIT_74 => X"ffffffebffffffff000000130000000000000007000000000000001a00000000",
            INIT_75 => X"ffffffebffffffffffffffe9ffffffff0000001000000000ffffffe5ffffffff",
            INIT_76 => X"ffffffeaffffffff0000001000000000ffffffe4ffffffff0000000b00000000",
            INIT_77 => X"0000001400000000fffffff8ffffffffffffffefffffffff0000001d00000000",
            INIT_78 => X"ffffffe1ffffffff000000350000000000000031000000000000001900000000",
            INIT_79 => X"fffffff5ffffffffffffffd7ffffffffffffffefffffffff0000002a00000000",
            INIT_7A => X"ffffffecffffffffffffffe7ffffffffffffffebfffffffffffffff1ffffffff",
            INIT_7B => X"fffffff6ffffffff000000170000000000000013000000000000000d00000000",
            INIT_7C => X"fffffffcffffffffffffffeeffffffffffffffd0ffffffffffffffe1ffffffff",
            INIT_7D => X"0000001300000000fffffff9ffffffff0000002b000000000000001b00000000",
            INIT_7E => X"ffffffd1ffffffffffffffbaffffffffffffffc7ffffffffffffffeaffffffff",
            INIT_7F => X"00000025000000000000000000000000ffffffccffffffffffffffe1ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE8;


    MEM_IWGHT_LAYER1_INSTANCE9 : if BRAM_NAME = "iwght_layer1_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffceffffffff0000003800000000fffffff8ffffffffffffffb7ffffffff",
            INIT_01 => X"ffffffe1ffffffffffffffcfffffffffffffffa6ffffffff0000000100000000",
            INIT_02 => X"ffffff9bffffffffffffffccffffffffffffffb8ffffffffffffffc1ffffffff",
            INIT_03 => X"00000000000000000000003100000000ffffffa0ffffffffffffff8effffffff",
            INIT_04 => X"ffffffd8ffffffff0000000e0000000000000005000000000000001900000000",
            INIT_05 => X"ffffffcdfffffffffffffffcffffffff0000000f00000000fffffffbffffffff",
            INIT_06 => X"00000002000000000000001400000000ffffffdcffffffffffffffa2ffffffff",
            INIT_07 => X"ffffffdeffffffffffffffb8ffffffffffffffd2ffffffffffffffdfffffffff",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE9;


    MEM_IWGHT_LAYER2_INSTANCE0 : if BRAM_NAME = "iwght_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffd64fffffffffffff0f4ffffffff00001d59000000000000122900000000",
            INIT_01 => X"fffffbe7ffffffff00001dd400000000fffffa11ffffffff000027ec00000000",
            INIT_02 => X"0000157600000000ffffea4bffffffff00000b130000000000001a0d00000000",
            INIT_03 => X"0000445400000000ffffe85dffffffff000028d800000000ffffeaddffffffff",
            INIT_04 => X"0000025400000000fffff10efffffffffffff086ffffffff0000105900000000",
            INIT_05 => X"fffff3cbffffffff00002d9400000000000026b8000000000000042d00000000",
            INIT_06 => X"00000396000000000000050600000000fffff815ffffffff00002c6400000000",
            INIT_07 => X"0000085100000000fffffd34ffffffffffffe25effffffff00002b5400000000",
            INIT_08 => X"00000dcd00000000ffffee74ffffffff0000212f0000000000003ee100000000",
            INIT_09 => X"fffffbfffffffffffffff3d5ffffffff00003ae8000000000000215c00000000",
            INIT_0A => X"000010f100000000ffffd6a7fffffffffffff49cffffffffffffdb76ffffffff",
            INIT_0B => X"00004dae00000000000043e200000000fffff867fffffffffffffed3ffffffff",
            INIT_0C => X"00000f2e0000000000002f4b00000000fffffc31ffffffff0000158100000000",
            INIT_0D => X"00002ede00000000fffffc82ffffffff000027540000000000001ca800000000",
            INIT_0E => X"000042c300000000000006aa00000000fffffb18fffffffffffff033ffffffff",
            INIT_0F => X"000003ed000000000000335600000000fffffe8dffffffff000023ac00000000",
            INIT_10 => X"00000016000000000000001c0000000000000017000000000000000f00000000",
            INIT_11 => X"ffffffc0ffffffffffffffceffffffff0000000f00000000fffffffbffffffff",
            INIT_12 => X"ffffffe5ffffffffffffffdfffffffffffffffdbffffffffffffffb2ffffffff",
            INIT_13 => X"fffffff3fffffffffffffffbffffffffffffffe2ffffffff0000002300000000",
            INIT_14 => X"0000001c0000000000000031000000000000001600000000ffffffc9ffffffff",
            INIT_15 => X"0000002800000000000000220000000000000038000000000000000c00000000",
            INIT_16 => X"fffffff2ffffffff0000001f000000000000002a000000000000003700000000",
            INIT_17 => X"ffffffb3ffffffffffffffadffffffffffffffe9fffffffffffffff9ffffffff",
            INIT_18 => X"ffffffe6fffffffffffffffeffffffffffffffd9ffffffffffffffb3ffffffff",
            INIT_19 => X"ffffffc9fffffffffffffffcfffffffffffffff8fffffffffffffff0ffffffff",
            INIT_1A => X"ffffffd2ffffffffffffffedffffffffffffffb8ffffffffffffffc2ffffffff",
            INIT_1B => X"0000000900000000ffffffedffffffff0000000600000000ffffffe5ffffffff",
            INIT_1C => X"ffffffe6ffffffffffffffc6ffffffffffffffaafffffffffffffff2ffffffff",
            INIT_1D => X"fffffff6ffffffff0000002c00000000ffffffccffffffffffffff8cffffffff",
            INIT_1E => X"0000000c0000000000000039000000000000001e000000000000002300000000",
            INIT_1F => X"fffffffffffffffffffffff2ffffffff00000016000000000000000c00000000",
            INIT_20 => X"00000038000000000000001100000000ffffffefffffffff0000001300000000",
            INIT_21 => X"fffffff8ffffffff0000000500000000fffffff3ffffffff0000002200000000",
            INIT_22 => X"0000000a00000000fffffff8ffffffff00000000000000000000001d00000000",
            INIT_23 => X"fffffff4ffffffff0000000300000000fffffffeffffffff0000002100000000",
            INIT_24 => X"0000001d0000000000000056000000000000003f00000000ffffffedffffffff",
            INIT_25 => X"0000000d0000000000000007000000000000000400000000fffffffaffffffff",
            INIT_26 => X"0000000600000000fffffffdffffffff0000003b00000000ffffffdcffffffff",
            INIT_27 => X"fffffff9fffffffffffffff8ffffffff00000000000000000000000d00000000",
            INIT_28 => X"fffffff7ffffffffffffffb5ffffffffffffffdaffffffffffffffe5ffffffff",
            INIT_29 => X"ffffffefffffffff0000003500000000ffffffd4ffffffffffffffefffffffff",
            INIT_2A => X"0000000c00000000000000210000000000000028000000000000000700000000",
            INIT_2B => X"0000004600000000000000060000000000000046000000000000004300000000",
            INIT_2C => X"0000005400000000000000320000000000000022000000000000006a00000000",
            INIT_2D => X"00000010000000000000001d0000000000000009000000000000006000000000",
            INIT_2E => X"ffffffddfffffffffffffff7ffffffffffffffdfffffffffffffffcfffffffff",
            INIT_2F => X"00000007000000000000000c00000000ffffffffffffffffffffffddffffffff",
            INIT_30 => X"0000000800000000ffffffffffffffff00000011000000000000001700000000",
            INIT_31 => X"fffffff8fffffffffffffff5ffffffffffffffeffffffffffffffff0ffffffff",
            INIT_32 => X"0000001600000000000000340000000000000000000000000000000c00000000",
            INIT_33 => X"00000056000000000000003e0000000000000037000000000000002700000000",
            INIT_34 => X"fffffff8ffffffffffffffdfffffffff0000000000000000ffffffffffffffff",
            INIT_35 => X"00000007000000000000002200000000ffffffb5ffffffffffffffe7ffffffff",
            INIT_36 => X"0000001a000000000000001000000000ffffffebffffffffffffffebffffffff",
            INIT_37 => X"ffffffefffffffff00000043000000000000001d000000000000000800000000",
            INIT_38 => X"ffffffb8ffffffffffffffe1ffffffffffffffe2ffffffff0000000400000000",
            INIT_39 => X"ffffffd6ffffffffffffff92ffffffffffffffc0ffffffffffffffc2ffffffff",
            INIT_3A => X"ffffffffffffffffffffffe8ffffffffffffffceffffffffffffffe8ffffffff",
            INIT_3B => X"000000430000000000000006000000000000000600000000ffffffbfffffffff",
            INIT_3C => X"fffffff0ffffffff0000000800000000ffffffbaffffffff0000001f00000000",
            INIT_3D => X"0000001500000000fffffff7fffffffffffffff4ffffffff0000002700000000",
            INIT_3E => X"0000000d00000000fffffff9ffffffff0000000e000000000000001d00000000",
            INIT_3F => X"00000013000000000000000c0000000000000016000000000000000100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002a00000000000000140000000000000015000000000000001f00000000",
            INIT_41 => X"00000030000000000000000000000000ffffffffffffffff0000001a00000000",
            INIT_42 => X"0000001100000000000000300000000000000023000000000000001700000000",
            INIT_43 => X"fffffffdffffffff0000001a000000000000004b000000000000004100000000",
            INIT_44 => X"ffffffe8ffffffffffffffdeffffffffffffffe7ffffffffffffffebffffffff",
            INIT_45 => X"ffffffd6fffffffffffffff9ffffffffffffffe8ffffffffffffffacffffffff",
            INIT_46 => X"0000003d00000000fffffff7ffffffffffffffdbffffffff0000000800000000",
            INIT_47 => X"0000002500000000000000080000000000000010000000000000003400000000",
            INIT_48 => X"00000026000000000000000f0000000000000017000000000000001e00000000",
            INIT_49 => X"0000000800000000ffffffecffffffff00000000000000000000001000000000",
            INIT_4A => X"00000012000000000000001c00000000ffffffe0ffffffffffffffdbffffffff",
            INIT_4B => X"0000002f000000000000002e00000000fffffffcfffffffffffffffcffffffff",
            INIT_4C => X"ffffffefffffffff0000000700000000ffffffe8fffffffffffffff9ffffffff",
            INIT_4D => X"ffffffc1ffffffffffffffc6ffffffffffffffd5ffffffffffffffdbffffffff",
            INIT_4E => X"ffffffbcffffffffffffffdaffffffffffffffd7ffffffffffffffb4ffffffff",
            INIT_4F => X"fffffff8ffffffffffffffe5ffffffffffffffdeffffffffffffffc2ffffffff",
            INIT_50 => X"0000000700000000fffffff6ffffffffffffffe4ffffffff0000001e00000000",
            INIT_51 => X"0000002200000000fffffff3fffffffffffffff8ffffffff0000001000000000",
            INIT_52 => X"0000003f00000000ffffffdcfffffffffffffff1ffffffff0000001500000000",
            INIT_53 => X"ffffffe5ffffffff000000070000000000000015000000000000005300000000",
            INIT_54 => X"ffffffe7fffffffffffffff2ffffffff00000000000000000000000400000000",
            INIT_55 => X"000000030000000000000018000000000000001700000000fffffffdffffffff",
            INIT_56 => X"0000001e000000000000001b00000000ffffffefffffffff0000002900000000",
            INIT_57 => X"0000000900000000ffffffffffffffffffffffe9ffffffff0000000f00000000",
            INIT_58 => X"ffffffe9ffffffff0000000c0000000000000007000000000000000300000000",
            INIT_59 => X"0000000100000000ffffffeffffffffffffffffbffffffffffffffe4ffffffff",
            INIT_5A => X"fffffff1ffffffff0000000c0000000000000008000000000000000700000000",
            INIT_5B => X"ffffffcaffffffff0000001700000000fffffffcffffffff0000000800000000",
            INIT_5C => X"ffffffd0ffffffff00000000000000000000001e000000000000001600000000",
            INIT_5D => X"0000000800000000ffffffecffffffffffffffdcffffffffffffffedffffffff",
            INIT_5E => X"0000000e000000000000001e0000000000000019000000000000000c00000000",
            INIT_5F => X"fffffff3ffffffffffffffdeffffffffffffffadffffffffffffffe9ffffffff",
            INIT_60 => X"0000002800000000fffffffcfffffffffffffff2ffffffffffffffeeffffffff",
            INIT_61 => X"fffffff9ffffffff000000010000000000000017000000000000004200000000",
            INIT_62 => X"ffffffb8ffffffffffffffc6ffffffff0000001600000000ffffffdfffffffff",
            INIT_63 => X"00000017000000000000001f000000000000002f00000000ffffffedffffffff",
            INIT_64 => X"ffffffe3ffffffff00000007000000000000000000000000fffffff4ffffffff",
            INIT_65 => X"0000001b000000000000000800000000fffffffeffffffffffffffd3ffffffff",
            INIT_66 => X"fffffffaffffffff0000000b0000000000000032000000000000003c00000000",
            INIT_67 => X"ffffffdaffffffff00000030000000000000002400000000fffffff8ffffffff",
            INIT_68 => X"0000000000000000fffffff6ffffffffffffffd6ffffffffffffffe6ffffffff",
            INIT_69 => X"000000300000000000000020000000000000000c00000000fffffffaffffffff",
            INIT_6A => X"0000001400000000000000280000000000000030000000000000002200000000",
            INIT_6B => X"0000000000000000ffffffeefffffffffffffffcffffffff0000001e00000000",
            INIT_6C => X"0000000f00000000ffffffffffffffff0000000700000000ffffffebffffffff",
            INIT_6D => X"fffffff9ffffffff00000001000000000000000b000000000000000a00000000",
            INIT_6E => X"ffffffffffffffff00000004000000000000002300000000ffffffe3ffffffff",
            INIT_6F => X"0000000300000000000000090000000000000003000000000000000100000000",
            INIT_70 => X"fffffff6ffffffffffffffeeffffffffffffffc2ffffffff0000001000000000",
            INIT_71 => X"fffffff2ffffffff0000000000000000ffffffeeffffffff0000001a00000000",
            INIT_72 => X"000000300000000000000007000000000000000d00000000fffffffaffffffff",
            INIT_73 => X"00000019000000000000000e00000000ffffffe1ffffffffffffffdcffffffff",
            INIT_74 => X"0000001000000000fffffffefffffffffffffffaffffffff0000004300000000",
            INIT_75 => X"0000002c00000000ffffffe5ffffffff00000004000000000000003a00000000",
            INIT_76 => X"ffffffe2ffffffff0000000900000000ffffffd7ffffffffffffffafffffffff",
            INIT_77 => X"ffffffffffffffff0000000300000000ffffffb0ffffffffffffff90ffffffff",
            INIT_78 => X"00000001000000000000001400000000fffffff2ffffffffffffffffffffffff",
            INIT_79 => X"0000000700000000fffffffcffffffff0000000b000000000000000200000000",
            INIT_7A => X"00000030000000000000002b00000000ffffffe6ffffffff0000000600000000",
            INIT_7B => X"00000041000000000000002c000000000000002900000000fffffff0ffffffff",
            INIT_7C => X"ffffffd3ffffffff0000001d00000000fffffffdffffffff0000000d00000000",
            INIT_7D => X"ffffffc5ffffffffffffffd3ffffffff0000000a00000000ffffffddffffffff",
            INIT_7E => X"00000006000000000000002e000000000000001400000000ffffffabffffffff",
            INIT_7F => X"ffffffadffffffff0000000c0000000000000018000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE0;


    MEM_IWGHT_LAYER2_INSTANCE1 : if BRAM_NAME = "iwght_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff8cffffffffffffffa3ffffffffffffffd8ffffffffffffffccffffffff",
            INIT_01 => X"ffffffdfffffffffffffffb5ffffffffffffffe5ffffffffffffff73ffffffff",
            INIT_02 => X"ffffffcfffffffffffffffcdfffffffffffffff4ffffffff0000002e00000000",
            INIT_03 => X"ffffffe9ffffffffffffff9effffffffffffffeeffffffffffffffd8ffffffff",
            INIT_04 => X"00000000000000000000001900000000ffffffedffffffffffffffcaffffffff",
            INIT_05 => X"00000025000000000000002b000000000000000b000000000000004600000000",
            INIT_06 => X"fffffff3ffffffffffffffc7ffffffff0000001c000000000000001400000000",
            INIT_07 => X"00000010000000000000000f000000000000001400000000ffffffc4ffffffff",
            INIT_08 => X"ffffffecffffffff000000100000000000000008000000000000000b00000000",
            INIT_09 => X"000000620000000000000017000000000000000c000000000000003300000000",
            INIT_0A => X"0000002a00000000000000490000000000000038000000000000000500000000",
            INIT_0B => X"ffffffbcffffffff00000006000000000000001f00000000ffffffddffffffff",
            INIT_0C => X"fffffff8ffffffffffffffeaffffffffffffffa6ffffffffffffffb3ffffffff",
            INIT_0D => X"ffffffdbffffffffffffffe6ffffffff0000002100000000fffffff4ffffffff",
            INIT_0E => X"00000021000000000000000800000000fffffffdffffffff0000002c00000000",
            INIT_0F => X"fffffffdffffffffffffffd4ffffffff00000024000000000000003500000000",
            INIT_10 => X"0000002b0000000000000019000000000000002700000000ffffffc8ffffffff",
            INIT_11 => X"ffffffccffffffff0000000000000000fffffffdffffffff0000000800000000",
            INIT_12 => X"00000024000000000000002600000000ffffffc4ffffffffffffffcbffffffff",
            INIT_13 => X"000000190000000000000022000000000000002d00000000fffffff5ffffffff",
            INIT_14 => X"ffffffcaffffffff0000000d000000000000001c000000000000004500000000",
            INIT_15 => X"fffffff5ffffffffffffffe0ffffffffffffffceffffffffffffffa5ffffffff",
            INIT_16 => X"ffffffcfffffffffffffffe3ffffffffffffffddfffffffffffffff9ffffffff",
            INIT_17 => X"00000005000000000000001f0000000000000028000000000000003900000000",
            INIT_18 => X"ffffffe5ffffffffffffffeeffffffff0000000800000000fffffff8ffffffff",
            INIT_19 => X"00000014000000000000000c000000000000000700000000ffffffedffffffff",
            INIT_1A => X"fffffff6ffffffff0000000500000000ffffffc6ffffffffffffffccffffffff",
            INIT_1B => X"0000001f000000000000003500000000ffffffe6fffffffffffffff3ffffffff",
            INIT_1C => X"0000001000000000000000100000000000000020000000000000002600000000",
            INIT_1D => X"0000001000000000ffffffc4ffffffffffffffdaffffffffffffffb7ffffffff",
            INIT_1E => X"0000000d000000000000000700000000fffffff8ffffffffffffffdbffffffff",
            INIT_1F => X"0000003600000000000000010000000000000021000000000000000d00000000",
            INIT_20 => X"fffffff1ffffffff0000000c00000000ffffffc9ffffffffffffffccffffffff",
            INIT_21 => X"ffffffe6ffffffffffffffebffffffff0000000f00000000ffffffebffffffff",
            INIT_22 => X"fffffffcffffffff00000000000000000000001800000000fffffff4ffffffff",
            INIT_23 => X"0000004c00000000ffffffd5ffffffff00000008000000000000002400000000",
            INIT_24 => X"fffffffaffffffff0000002d00000000ffffffe4fffffffffffffff5ffffffff",
            INIT_25 => X"ffffffdbffffffffffffffe5ffffffff0000003900000000ffffffc7ffffffff",
            INIT_26 => X"0000003600000000ffffffe2ffffffff00000014000000000000003400000000",
            INIT_27 => X"ffffffd8ffffffff000000390000000000000004000000000000000200000000",
            INIT_28 => X"0000000300000000ffffffccffffffff00000004000000000000002500000000",
            INIT_29 => X"fffffffcffffffff000000000000000000000020000000000000001d00000000",
            INIT_2A => X"ffffffe1fffffffffffffffcffffffff00000023000000000000001900000000",
            INIT_2B => X"00000031000000000000000e000000000000000b000000000000000300000000",
            INIT_2C => X"ffffffa1ffffffff0000004800000000fffffff4ffffffffffffffe4ffffffff",
            INIT_2D => X"ffffffddffffffff00000005000000000000001500000000ffffff88ffffffff",
            INIT_2E => X"fffffff4ffffffffffffffc2ffffffff00000005000000000000000300000000",
            INIT_2F => X"ffffffb7ffffffff0000002200000000fffffffcffffffff0000000400000000",
            INIT_30 => X"0000000900000000ffffffdbffffffffffffffe8ffffffffffffff9fffffffff",
            INIT_31 => X"ffffffdefffffffffffffffafffffffffffffffeffffffff0000000d00000000",
            INIT_32 => X"00000028000000000000000f00000000ffffffdeffffffff0000001f00000000",
            INIT_33 => X"00000000000000000000003e00000000fffffffbffffffffffffffdaffffffff",
            INIT_34 => X"fffffff8ffffffff0000003000000000ffffffddffffffff0000002000000000",
            INIT_35 => X"ffffffa9ffffffffffffffecffffffff0000001700000000fffffff8ffffffff",
            INIT_36 => X"ffffffe9ffffffffffffffb8ffffffff0000000300000000fffffff8ffffffff",
            INIT_37 => X"00000009000000000000001100000000ffffffe7ffffffff0000001500000000",
            INIT_38 => X"00000027000000000000000100000000fffffff9fffffffffffffff8ffffffff",
            INIT_39 => X"ffffffcbffffffff0000000600000000fffffff5ffffffff0000001600000000",
            INIT_3A => X"ffffffe5ffffffffffffffffffffffff0000002b00000000ffffffc4ffffffff",
            INIT_3B => X"0000003100000000ffffffabffffffffffffffeaffffffff0000003600000000",
            INIT_3C => X"00000047000000000000008600000000ffffffc2ffffffffffffffe4ffffffff",
            INIT_3D => X"0000000100000000000000190000000000000000000000000000000b00000000",
            INIT_3E => X"ffffffb7ffffffff0000000d000000000000001f00000000ffffffedffffffff",
            INIT_3F => X"fffffff9ffffffff0000001300000000ffffffe2ffffffff0000000a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000000700000000ffffffedffffffff0000000000000000",
            INIT_41 => X"ffffffe6fffffffffffffff6fffffffffffffffcffffffff0000000f00000000",
            INIT_42 => X"ffffffdaffffffff0000000f00000000ffffffc1ffffffffffffffd3ffffffff",
            INIT_43 => X"ffffffdfffffffffffffffccffffffffffffffe3ffffffffffffffc8ffffffff",
            INIT_44 => X"0000000b00000000fffffff2ffffffff00000006000000000000000c00000000",
            INIT_45 => X"fffffff8ffffffff0000000500000000ffffffedffffffff0000001000000000",
            INIT_46 => X"0000000c00000000ffffffe4ffffffff00000014000000000000000b00000000",
            INIT_47 => X"00000001000000000000002a00000000ffffffe2ffffffff0000003100000000",
            INIT_48 => X"00000022000000000000002200000000fffffffdffffffffffffffafffffffff",
            INIT_49 => X"ffffffefffffffff000000260000000000000034000000000000003800000000",
            INIT_4A => X"0000000c00000000ffffffd9fffffffffffffffaffffffffffffffe9ffffffff",
            INIT_4B => X"0000000e000000000000004200000000fffffff1fffffffffffffff5ffffffff",
            INIT_4C => X"0000000d0000000000000002000000000000000d000000000000002200000000",
            INIT_4D => X"ffffffd7ffffffff000000320000000000000011000000000000000500000000",
            INIT_4E => X"ffffffe9ffffffff00000002000000000000000200000000fffffff2ffffffff",
            INIT_4F => X"ffffffd6ffffffffffffffbeffffffffffffffecfffffffffffffff3ffffffff",
            INIT_50 => X"fffffff7ffffffffffffffe1ffffffffffffffcbffffffffffffffe8ffffffff",
            INIT_51 => X"00000029000000000000003800000000ffffffe2fffffffffffffff7ffffffff",
            INIT_52 => X"ffffffa6fffffffffffffffaffffffff0000000f000000000000000200000000",
            INIT_53 => X"ffffffbfffffffff000000090000000000000027000000000000004800000000",
            INIT_54 => X"0000000800000000ffffffe9ffffffffffffffdfffffffff0000001300000000",
            INIT_55 => X"ffffffc1ffffffff0000001200000000ffffffecffffffffffffffc2ffffffff",
            INIT_56 => X"00000006000000000000000200000000fffffffbffffffff0000001400000000",
            INIT_57 => X"0000000a000000000000000400000000ffffffdffffffffffffffff0ffffffff",
            INIT_58 => X"0000001e0000000000000001000000000000002000000000ffffffd0ffffffff",
            INIT_59 => X"ffffffd5ffffffff0000002b00000000ffffffe9ffffffff0000000800000000",
            INIT_5A => X"ffffffc8ffffffffffffffd3ffffffff0000000800000000ffffffd8ffffffff",
            INIT_5B => X"ffffffcbffffffffffffffe5ffffffffffffffe6ffffffffffffffeaffffffff",
            INIT_5C => X"ffffffd6ffffffff0000000500000000fffffffeffffffff0000001d00000000",
            INIT_5D => X"0000000c00000000fffffff6fffffffffffffffcffffffff0000000300000000",
            INIT_5E => X"ffffffdcffffffffffffffc5ffffffffffffffe4ffffffffffffffe8ffffffff",
            INIT_5F => X"0000002a00000000fffffffffffffffffffffff0fffffffffffffff3ffffffff",
            INIT_60 => X"00000002000000000000001300000000ffffffeeffffffff0000000d00000000",
            INIT_61 => X"ffffffc6ffffffff0000004a000000000000003300000000fffffffaffffffff",
            INIT_62 => X"0000003200000000ffffffe3ffffffff00000016000000000000003300000000",
            INIT_63 => X"0000001900000000fffffff3ffffffffffffffc3ffffffffffffffe0ffffffff",
            INIT_64 => X"ffffffdffffffffffffffffffffffffffffffff1ffffffffffffffeeffffffff",
            INIT_65 => X"ffffffdcffffffffffffffd2ffffffff00000013000000000000000a00000000",
            INIT_66 => X"0000001800000000fffffffeffffffffffffffc1ffffffffffffffc1ffffffff",
            INIT_67 => X"ffffffe4ffffffff00000022000000000000000c00000000ffffffd2ffffffff",
            INIT_68 => X"ffffffebffffffff0000000500000000fffffff7fffffffffffffff3ffffffff",
            INIT_69 => X"0000000100000000ffffffe8ffffffff0000001300000000fffffff6ffffffff",
            INIT_6A => X"ffffffdfffffffffffffffd1ffffffffffffffe6ffffffffffffffe1ffffffff",
            INIT_6B => X"0000000b00000000ffffffe8fffffffffffffff4ffffffffffffffdfffffffff",
            INIT_6C => X"ffffffd9ffffffffffffffb9ffffffffffffffd2fffffffffffffff6ffffffff",
            INIT_6D => X"000000270000000000000036000000000000000900000000fffffff1ffffffff",
            INIT_6E => X"0000001c000000000000003e000000000000002c000000000000002400000000",
            INIT_6F => X"000000180000000000000025000000000000001a000000000000002900000000",
            INIT_70 => X"ffffffe4ffffffff0000000000000000ffffffebfffffffffffffff1ffffffff",
            INIT_71 => X"0000000800000000000000030000000000000006000000000000001a00000000",
            INIT_72 => X"ffffffe4ffffffff0000000600000000ffffffe9ffffffffffffffebffffffff",
            INIT_73 => X"ffffffd9ffffffffffffffc9fffffffffffffff5ffffffff0000001b00000000",
            INIT_74 => X"fffffffdffffffff00000001000000000000002e000000000000001a00000000",
            INIT_75 => X"fffffff4fffffffffffffffaffffffff0000001a000000000000001500000000",
            INIT_76 => X"000000340000000000000012000000000000001a00000000ffffffe3ffffffff",
            INIT_77 => X"00000018000000000000000f0000000000000012000000000000001800000000",
            INIT_78 => X"00000008000000000000000e0000000000000003000000000000000700000000",
            INIT_79 => X"000000170000000000000030000000000000001b000000000000000100000000",
            INIT_7A => X"0000000100000000000000300000000000000027000000000000003100000000",
            INIT_7B => X"ffffffdbffffffff0000000000000000fffffff6ffffffffffffffd2ffffffff",
            INIT_7C => X"ffffffc6ffffffffffffffc7ffffffffffffffc8ffffffffffffffecffffffff",
            INIT_7D => X"ffffffefffffffff0000000a00000000fffffffffffffffffffffff4ffffffff",
            INIT_7E => X"fffffff8ffffffffffffffefffffffff00000015000000000000000000000000",
            INIT_7F => X"0000000200000000fffffff7fffffffffffffff5ffffffffffffffeaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE1;


    MEM_IWGHT_LAYER2_INSTANCE2 : if BRAM_NAME = "iwght_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000ffffffebffffffffffffffefffffffff0000000200000000",
            INIT_01 => X"00000040000000000000001a000000000000001c000000000000003700000000",
            INIT_02 => X"00000019000000000000002f0000000000000029000000000000002f00000000",
            INIT_03 => X"fffffff7ffffffff0000000c0000000000000026000000000000002300000000",
            INIT_04 => X"0000000400000000fffffff9fffffffffffffff1ffffffff0000000000000000",
            INIT_05 => X"ffffffb3ffffffffffffffa6fffffffffffffff9ffffffff0000003400000000",
            INIT_06 => X"ffffffe8ffffffff0000000000000000ffffffe7ffffffffffffffebffffffff",
            INIT_07 => X"00000001000000000000000a0000000000000028000000000000000900000000",
            INIT_08 => X"fffffffefffffffffffffff4fffffffffffffffefffffffffffffff8ffffffff",
            INIT_09 => X"0000000c00000000fffffff2fffffffffffffff6ffffffff0000000000000000",
            INIT_0A => X"0000001600000000000000270000000000000005000000000000001700000000",
            INIT_0B => X"00000035000000000000002c0000000000000029000000000000002800000000",
            INIT_0C => X"ffffffefffffffff0000001a00000000fffffffbffffffff0000002c00000000",
            INIT_0D => X"ffffffb6ffffffffffffffd6ffffffffffffffd9ffffffffffffffb9ffffffff",
            INIT_0E => X"fffffff1ffffffffffffff97ffffffffffffffe1ffffffffffffffe1ffffffff",
            INIT_0F => X"00000042000000000000001400000000fffffff8ffffffff0000001700000000",
            INIT_10 => X"0000001b00000000ffffffe8ffffffff00000070000000000000007c00000000",
            INIT_11 => X"fffffffbfffffffffffffff0ffffffffffffffe3ffffffff0000000300000000",
            INIT_12 => X"0000001e0000000000000004000000000000000e00000000ffffffdaffffffff",
            INIT_13 => X"ffffffc6ffffffffffffffd4fffffffffffffff7ffffffff0000001600000000",
            INIT_14 => X"00000024000000000000000100000000ffffffefffffffffffffffbcffffffff",
            INIT_15 => X"ffffffdfffffffff0000002a0000000000000008000000000000004000000000",
            INIT_16 => X"ffffffb4ffffffffffffffe5ffffffffffffffe3ffffffffffffffb3ffffffff",
            INIT_17 => X"ffffffe8ffffffffffffffdcfffffffffffffff9fffffffffffffff9ffffffff",
            INIT_18 => X"0000002500000000fffffffeffffffff0000000100000000ffffffeeffffffff",
            INIT_19 => X"fffffff3ffffffffffffff8affffffff00000019000000000000001b00000000",
            INIT_1A => X"00000025000000000000002600000000ffffffedfffffffffffffff5ffffffff",
            INIT_1B => X"0000000f000000000000006b000000000000002c000000000000002500000000",
            INIT_1C => X"0000001300000000ffffffecffffffff0000001c000000000000000400000000",
            INIT_1D => X"ffffffdbfffffffffffffff8fffffffffffffff7ffffffffffffffe8ffffffff",
            INIT_1E => X"ffffffd8ffffffffffffffedffffffffffffffe4ffffffff0000002200000000",
            INIT_1F => X"fffffffbffffffff00000017000000000000000600000000ffffffb2ffffffff",
            INIT_20 => X"ffffffecffffffffffffffbcffffffffffffffe4ffffffff0000003f00000000",
            INIT_21 => X"0000001a000000000000000b000000000000000100000000ffffffffffffffff",
            INIT_22 => X"0000001b00000000ffffffefffffffff00000025000000000000001d00000000",
            INIT_23 => X"ffffffeeffffffff0000000900000000ffffffd9ffffffff0000000800000000",
            INIT_24 => X"ffffffe9ffffffff00000015000000000000002d00000000fffffff5ffffffff",
            INIT_25 => X"0000002700000000000000010000000000000008000000000000001500000000",
            INIT_26 => X"ffffffe3ffffffffffffffc4ffffffffffffffecfffffffffffffffaffffffff",
            INIT_27 => X"fffffff3fffffffffffffff9ffffffffffffffe0ffffffff0000000e00000000",
            INIT_28 => X"ffffffe7fffffffffffffff4ffffffffffffffc9ffffffffffffffb2ffffffff",
            INIT_29 => X"00000038000000000000000300000000ffffffd2ffffffffffffffeeffffffff",
            INIT_2A => X"ffffffffffffffff0000001b0000000000000072000000000000003600000000",
            INIT_2B => X"0000003a000000000000007000000000fffffff9ffffffff0000002b00000000",
            INIT_2C => X"0000001b00000000fffffff4ffffffff00000014000000000000003b00000000",
            INIT_2D => X"0000000500000000ffffffe3ffffffffffffffadffffffffffffffc8ffffffff",
            INIT_2E => X"00000014000000000000001800000000ffffffd5ffffffff0000001300000000",
            INIT_2F => X"ffffffdeffffffff00000009000000000000001500000000fffffffcffffffff",
            INIT_30 => X"fffffff4ffffffff0000000700000000fffffffaffffffff0000000800000000",
            INIT_31 => X"fffffffbffffffff000000010000000000000010000000000000000f00000000",
            INIT_32 => X"ffffffe9ffffffffffffffecffffffff00000015000000000000000400000000",
            INIT_33 => X"0000000400000000ffffffd8ffffffff00000002000000000000000100000000",
            INIT_34 => X"00000021000000000000001f000000000000000300000000ffffffe7ffffffff",
            INIT_35 => X"ffffffd2fffffffffffffff7ffffffff00000008000000000000001100000000",
            INIT_36 => X"0000001100000000000000110000000000000026000000000000001e00000000",
            INIT_37 => X"0000000d000000000000001900000000ffffffdafffffffffffffffeffffffff",
            INIT_38 => X"ffffffd2ffffffffffffffeeffffffff0000001900000000ffffffeaffffffff",
            INIT_39 => X"fffffffffffffffffffffffaffffffff0000000b000000000000001c00000000",
            INIT_3A => X"0000000a0000000000000012000000000000001300000000fffffff5ffffffff",
            INIT_3B => X"fffffffbffffffffffffffefffffffffffffffd3ffffffff0000000800000000",
            INIT_3C => X"ffffffcafffffffffffffff5ffffffffffffffd5ffffffffffffffd7ffffffff",
            INIT_3D => X"fffffffcffffffff0000001a00000000ffffffe2ffffffffffffffbfffffffff",
            INIT_3E => X"0000001500000000fffffff1ffffffff0000000200000000fffffff7ffffffff",
            INIT_3F => X"0000000500000000000000130000000000000013000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c00000000fffffff5fffffffffffffffdffffffff0000002400000000",
            INIT_41 => X"ffffffcdffffffff0000000200000000fffffff4ffffffffffffffd2ffffffff",
            INIT_42 => X"0000000400000000ffffffc1ffffffffffffffffffffffff0000003000000000",
            INIT_43 => X"00000016000000000000000400000000ffffffc8ffffffff0000001400000000",
            INIT_44 => X"0000004b000000000000001b00000000ffffffecffffffff0000000600000000",
            INIT_45 => X"fffffffbffffffff0000001e00000000fffffff1ffffffffffffffe0ffffffff",
            INIT_46 => X"00000018000000000000001a0000000000000013000000000000001100000000",
            INIT_47 => X"ffffffe7fffffffffffffffbffffffff00000009000000000000000100000000",
            INIT_48 => X"0000000800000000ffffffeaffffffff0000002700000000fffffffcffffffff",
            INIT_49 => X"0000000900000000ffffffd7fffffffffffffff3ffffffff0000001700000000",
            INIT_4A => X"ffffffe3fffffffffffffff3ffffffffffffffffffffffffffffffe1ffffffff",
            INIT_4B => X"0000002100000000fffffff7ffffffff00000028000000000000000c00000000",
            INIT_4C => X"0000004600000000000000510000000000000011000000000000002c00000000",
            INIT_4D => X"00000008000000000000001900000000ffffffcaffffffff0000006900000000",
            INIT_4E => X"ffffffb7ffffffff0000000400000000fffffff3ffffffffffffffbbffffffff",
            INIT_4F => X"fffffffaffffffffffffffedfffffffffffffffeffffffff0000000700000000",
            INIT_50 => X"0000000300000000fffffffbfffffffffffffffcffffffff0000001200000000",
            INIT_51 => X"ffffffdbfffffffffffffffffffffffffffffff6ffffffff0000000100000000",
            INIT_52 => X"ffffffedffffffffffffffd3ffffffff0000000800000000ffffffe6ffffffff",
            INIT_53 => X"ffffffc8ffffffffffffffddffffffffffffffa8ffffffffffffffdeffffffff",
            INIT_54 => X"0000001400000000fffffffaffffffff0000000d000000000000001500000000",
            INIT_55 => X"000000100000000000000002000000000000000c000000000000000800000000",
            INIT_56 => X"0000003800000000ffffffc6ffffffffffffffeeffffffff0000001f00000000",
            INIT_57 => X"00000000000000000000001400000000ffffffb8ffffffffffffffd3ffffffff",
            INIT_58 => X"fffffff7ffffffff00000009000000000000000000000000ffffffe6ffffffff",
            INIT_59 => X"ffffffe4ffffffffffffff91fffffffffffffffbffffffff0000003900000000",
            INIT_5A => X"0000000000000000ffffffcaffffffffffffffeeffffffffffffffe3ffffffff",
            INIT_5B => X"000000160000000000000001000000000000001800000000fffffff3ffffffff",
            INIT_5C => X"fffffff5fffffffffffffffaffffffff00000000000000000000000500000000",
            INIT_5D => X"fffffff5ffffffff0000001d000000000000000200000000fffffff9ffffffff",
            INIT_5E => X"ffffffe9ffffffff00000002000000000000000000000000fffffff5ffffffff",
            INIT_5F => X"fffffff7ffffffff0000000800000000ffffffefffffffff0000001c00000000",
            INIT_60 => X"ffffffdbffffffff0000000000000000ffffffedffffffffffffffcfffffffff",
            INIT_61 => X"ffffffefffffffff0000000b0000000000000012000000000000000d00000000",
            INIT_62 => X"ffffffddffffffff00000019000000000000001000000000fffffff3ffffffff",
            INIT_63 => X"000000030000000000000023000000000000002e000000000000002500000000",
            INIT_64 => X"ffffffeaffffffff0000000000000000fffffff9fffffffffffffff3ffffffff",
            INIT_65 => X"ffffffb0ffffffff0000000a000000000000000100000000ffffffc1ffffffff",
            INIT_66 => X"fffffff7fffffffffffffff8ffffffffffffffbcffffffffffffffd7ffffffff",
            INIT_67 => X"ffffffedffffffffffffffdbffffffffffffffd3ffffffffffffffd6ffffffff",
            INIT_68 => X"0000000f00000000ffffffd6ffffffffffffffc7ffffffffffffffe6ffffffff",
            INIT_69 => X"ffffffdcffffffff0000000300000000ffffffd7ffffffffffffffddffffffff",
            INIT_6A => X"fffffff2ffffffff0000002500000000fffffff9ffffffffffffffe3ffffffff",
            INIT_6B => X"ffffffe8ffffffff00000035000000000000000e000000000000000200000000",
            INIT_6C => X"fffffff5ffffffff0000000a0000000000000017000000000000002400000000",
            INIT_6D => X"ffffffeeffffffffffffffeafffffffffffffff8ffffffff0000000600000000",
            INIT_6E => X"ffffffd4fffffffffffffff6ffffffffffffffe3ffffffffffffffb3ffffffff",
            INIT_6F => X"0000001d0000000000000000000000000000003b000000000000002f00000000",
            INIT_70 => X"000000240000000000000024000000000000001a000000000000001c00000000",
            INIT_71 => X"00000015000000000000001200000000fffffffaffffffff0000000900000000",
            INIT_72 => X"0000004400000000ffffffe0fffffffffffffff2ffffffffffffffecffffffff",
            INIT_73 => X"0000001d000000000000000100000000fffffffaffffffff0000001300000000",
            INIT_74 => X"ffffffe8ffffffff0000000600000000fffffff4fffffffffffffff8ffffffff",
            INIT_75 => X"0000000900000000ffffffd7ffffffff0000000a00000000fffffffdffffffff",
            INIT_76 => X"0000002b000000000000000f0000000000000010000000000000002500000000",
            INIT_77 => X"0000000b000000000000002f000000000000000d000000000000001c00000000",
            INIT_78 => X"0000000800000000ffffffeafffffffffffffffbfffffffffffffff5ffffffff",
            INIT_79 => X"ffffffd1ffffffffffffffcbffffffffffffffeaffffffffffffffeaffffffff",
            INIT_7A => X"0000002a000000000000000500000000ffffffeafffffffffffffff9ffffffff",
            INIT_7B => X"0000000a00000000ffffffd6ffffffffffffffeaffffffffffffffdbffffffff",
            INIT_7C => X"0000000700000000ffffffe6ffffffffffffffdbffffffff0000001b00000000",
            INIT_7D => X"ffffffd5ffffffffffffff9fffffffffffffff9cffffffff0000000e00000000",
            INIT_7E => X"ffffffedffffffff0000002e000000000000001f000000000000002c00000000",
            INIT_7F => X"ffffffcbffffffffffffffb9ffffffffffffffafffffffff0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE2;


    MEM_IWGHT_LAYER2_INSTANCE3 : if BRAM_NAME = "iwght_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002b000000000000002f00000000fffffff7ffffffff0000000700000000",
            INIT_01 => X"ffffffa7ffffffffffffffe9ffffffffffffffc8ffffffffffffffc7ffffffff",
            INIT_02 => X"0000001e00000000fffffff7fffffffffffffff8ffffffffffffffc5ffffffff",
            INIT_03 => X"fffffffbffffffffffffffe4ffffffff00000000000000000000002100000000",
            INIT_04 => X"ffffffd8ffffffff000000470000000000000017000000000000002900000000",
            INIT_05 => X"fffffffbffffffff0000000600000000ffffffe2ffffffffffffffdcffffffff",
            INIT_06 => X"0000000b00000000000000130000000000000014000000000000003400000000",
            INIT_07 => X"0000000900000000ffffffd9ffffffff00000012000000000000002c00000000",
            INIT_08 => X"0000002400000000fffffffbffffffffffffffc9ffffffff0000001b00000000",
            INIT_09 => X"ffffffcaffffffff0000000800000000ffffffd8ffffffffffffffd8ffffffff",
            INIT_0A => X"0000000600000000ffffffffffffffff00000011000000000000003400000000",
            INIT_0B => X"ffffffb2ffffffffffffffb7ffffffffffffffcfffffffffffffffd6ffffffff",
            INIT_0C => X"00000020000000000000000700000000ffffffd9ffffffff0000000000000000",
            INIT_0D => X"0000003200000000000000170000000000000017000000000000000800000000",
            INIT_0E => X"ffffffedffffffffffffffe5ffffffffffffffdfffffffff0000001100000000",
            INIT_0F => X"ffffffd5ffffffffffffffe5fffffffffffffff3ffffffffffffffccffffffff",
            INIT_10 => X"00000000000000000000000a00000000fffffff0fffffffffffffff5ffffffff",
            INIT_11 => X"0000002100000000fffffffbffffffff00000032000000000000000700000000",
            INIT_12 => X"ffffffe9ffffffffffffffddffffffffffffffddfffffffffffffff3ffffffff",
            INIT_13 => X"ffffffddffffffff000000040000000000000013000000000000001b00000000",
            INIT_14 => X"0000005d000000000000008300000000fffffff2ffffffffffffffe2ffffffff",
            INIT_15 => X"0000003300000000fffffff6ffffffffffffffbcffffffff0000002600000000",
            INIT_16 => X"ffffffecffffffff00000022000000000000001900000000fffffffbffffffff",
            INIT_17 => X"00000000000000000000000c00000000ffffffabffffffffffffffd1ffffffff",
            INIT_18 => X"00000000000000000000000a00000000ffffffeefffffffffffffff8ffffffff",
            INIT_19 => X"0000001600000000000000110000000000000001000000000000001500000000",
            INIT_1A => X"00000012000000000000000e000000000000000f000000000000000300000000",
            INIT_1B => X"0000001c000000000000005a0000000000000013000000000000000000000000",
            INIT_1C => X"ffffffcfffffffff0000000b00000000ffffffecffffffffffffffe3ffffffff",
            INIT_1D => X"ffffffd6ffffffff0000000100000000fffffff8ffffffffffffffc5ffffffff",
            INIT_1E => X"fffffffbffffffff0000002700000000fffffff8fffffffffffffffcffffffff",
            INIT_1F => X"ffffffe0ffffffff0000000f00000000ffffffffffffffffffffffecffffffff",
            INIT_20 => X"ffffffefffffffff000000040000000000000025000000000000002300000000",
            INIT_21 => X"ffffffffffffffff0000000800000000ffffffe2ffffffff0000000100000000",
            INIT_22 => X"ffffffdbffffffffffffffbefffffffffffffffcffffffff0000004600000000",
            INIT_23 => X"fffffff6fffffffffffffff6ffffffff0000001a000000000000001400000000",
            INIT_24 => X"ffffffe7fffffffffffffff8ffffffff00000006000000000000000600000000",
            INIT_25 => X"0000001000000000000000090000000000000026000000000000003000000000",
            INIT_26 => X"ffffffdaffffffffffffffc6ffffffff0000000e000000000000001100000000",
            INIT_27 => X"0000000a00000000fffffffaffffffffffffffeeffffffff0000001200000000",
            INIT_28 => X"0000002b00000000ffffffe4ffffffff0000001700000000fffffffcffffffff",
            INIT_29 => X"0000000c000000000000001a00000000fffffff7ffffffff0000001700000000",
            INIT_2A => X"0000001100000000000000390000000000000048000000000000001d00000000",
            INIT_2B => X"fffffff2fffffffffffffff6ffffffff0000001a000000000000001600000000",
            INIT_2C => X"fffffff9ffffffffffffff88ffffffffffffffcbffffffff0000002300000000",
            INIT_2D => X"ffffffd9ffffffffffffffecffffffff0000000a00000000ffffffdfffffffff",
            INIT_2E => X"00000012000000000000001d0000000000000027000000000000003a00000000",
            INIT_2F => X"0000000a00000000ffffffd6ffffffffffffffe1ffffffff0000002100000000",
            INIT_30 => X"0000001f00000000fffffffdffffffff0000002600000000ffffffdbffffffff",
            INIT_31 => X"fffffff4ffffffff0000000000000000fffffff4ffffffff0000002500000000",
            INIT_32 => X"00000061000000000000002900000000fffffff9ffffffff0000001500000000",
            INIT_33 => X"ffffffeeffffffff0000004c000000000000000a00000000ffffffddffffffff",
            INIT_34 => X"0000001200000000ffffffd8ffffffff0000000500000000ffffffd2ffffffff",
            INIT_35 => X"0000000000000000ffffffceffffffff0000000e000000000000002200000000",
            INIT_36 => X"ffffffd8ffffffffffffffe7ffffffffffffffeffffffffffffffff8ffffffff",
            INIT_37 => X"fffffffcffffffff00000021000000000000002d000000000000001200000000",
            INIT_38 => X"ffffffe8fffffffffffffffefffffffffffffffdffffffff0000001000000000",
            INIT_39 => X"ffffffecffffffff000000050000000000000025000000000000000400000000",
            INIT_3A => X"ffffffd1ffffffffffffffb1ffffffffffffffeeffffffffffffffe5ffffffff",
            INIT_3B => X"ffffffdcfffffffffffffff5fffffffffffffffafffffffffffffffeffffffff",
            INIT_3C => X"ffffffefffffffffffffffe8fffffffffffffffeffffffff0000003400000000",
            INIT_3D => X"fffffffcffffffffffffffd4ffffffffffffffb6ffffffffffffffb0ffffffff",
            INIT_3E => X"0000001f000000000000000e00000000fffffff1ffffffff0000002200000000",
            INIT_3F => X"ffffffecfffffffffffffff6ffffffffffffffaeffffffff0000002500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000170000000000000000000000000000000f00000000ffffffffffffffff",
            INIT_41 => X"0000000b00000000000000240000000000000011000000000000000500000000",
            INIT_42 => X"00000030000000000000001f000000000000000e00000000fffffffeffffffff",
            INIT_43 => X"ffffffeeffffffff000000160000000000000007000000000000004b00000000",
            INIT_44 => X"0000000200000000000000450000000000000002000000000000001500000000",
            INIT_45 => X"fffffff1ffffffff0000000b00000000ffffffeeffffffff0000004000000000",
            INIT_46 => X"ffffffffffffffff0000001d000000000000000a00000000fffffffbffffffff",
            INIT_47 => X"0000000400000000ffffffffffffffff00000011000000000000000000000000",
            INIT_48 => X"0000000000000000ffffffc6ffffffff0000000e00000000fffffffcffffffff",
            INIT_49 => X"ffffffefffffffffffffffd4ffffffffffffffe5fffffffffffffff9ffffffff",
            INIT_4A => X"fffffffaffffffffffffffffffffffffffffffffffffffffffffffe9ffffffff",
            INIT_4B => X"fffffff2ffffffff00000027000000000000001e00000000fffffffaffffffff",
            INIT_4C => X"ffffffe5ffffffff00000025000000000000001b00000000ffffffe6ffffffff",
            INIT_4D => X"0000001c0000000000000024000000000000002300000000ffffffe4ffffffff",
            INIT_4E => X"0000002b000000000000000c0000000000000006000000000000001a00000000",
            INIT_4F => X"0000000500000000ffffffd0ffffffffffffffe8ffffffffffffffdbffffffff",
            INIT_50 => X"ffffffccffffffff0000000c00000000ffffffeafffffffffffffff5ffffffff",
            INIT_51 => X"0000001c00000000000000090000000000000002000000000000000d00000000",
            INIT_52 => X"0000000900000000fffffffbffffffffffffffeaffffffffffffffd7ffffffff",
            INIT_53 => X"fffffff4ffffffff0000001a00000000ffffffeaffffffff0000000300000000",
            INIT_54 => X"00000043000000000000003a0000000000000041000000000000000000000000",
            INIT_55 => X"ffffffe3ffffffff00000015000000000000003f000000000000002d00000000",
            INIT_56 => X"ffffffdffffffffffffffff9ffffffff00000002000000000000003100000000",
            INIT_57 => X"ffffffe4ffffffffffffffdcffffffff0000000400000000ffffffe3ffffffff",
            INIT_58 => X"0000002700000000000000080000000000000017000000000000003a00000000",
            INIT_59 => X"0000002e0000000000000033000000000000002e000000000000000000000000",
            INIT_5A => X"0000000e00000000ffffffe0ffffffffffffffceffffffff0000002400000000",
            INIT_5B => X"fffffff1ffffffff000000550000000000000029000000000000002f00000000",
            INIT_5C => X"ffffffdcffffffffffffffd9ffffffffffffffb9ffffffffffffffd4ffffffff",
            INIT_5D => X"ffffffe4ffffffffffffffffffffffff0000000800000000ffffffeeffffffff",
            INIT_5E => X"000000110000000000000004000000000000002700000000ffffffefffffffff",
            INIT_5F => X"ffffffffffffffff0000001100000000fffffff0ffffffff0000001700000000",
            INIT_60 => X"00000000000000000000000200000000fffffffbffffffff0000001100000000",
            INIT_61 => X"0000002500000000fffffff2fffffffffffffff0fffffffffffffffdffffffff",
            INIT_62 => X"ffffffdcffffffff0000000c0000000000000025000000000000002400000000",
            INIT_63 => X"ffffffc6ffffffffffffffccffffffffffffffc2ffffffff0000002000000000",
            INIT_64 => X"fffffff9ffffffff00000006000000000000000a000000000000000000000000",
            INIT_65 => X"0000002b0000000000000011000000000000000e000000000000002300000000",
            INIT_66 => X"fffffff6ffffffffffffffe3ffffffffffffffd4ffffffff0000001500000000",
            INIT_67 => X"0000001e0000000000000007000000000000000300000000ffffffdcffffffff",
            INIT_68 => X"fffffffeffffffff00000058000000000000001b00000000fffffff6ffffffff",
            INIT_69 => X"ffffffebffffffff0000003b00000000ffffffeeffffffff0000002000000000",
            INIT_6A => X"0000002e00000000ffffffe4ffffffffffffffefffffffffffffffc7ffffffff",
            INIT_6B => X"fffffff5fffffffffffffff0ffffffff0000000200000000fffffff6ffffffff",
            INIT_6C => X"fffffffaffffffffffffffcaffffffffffffffffffffffff0000001c00000000",
            INIT_6D => X"00000003000000000000001f000000000000002000000000ffffffeaffffffff",
            INIT_6E => X"fffffffeffffffff000000010000000000000014000000000000002400000000",
            INIT_6F => X"0000002c000000000000003d000000000000003d000000000000002400000000",
            INIT_70 => X"ffffffc6ffffffff000000270000000000000016000000000000003f00000000",
            INIT_71 => X"ffffffd1ffffffff0000003500000000ffffffc5ffffffffffffffc4ffffffff",
            INIT_72 => X"ffffffebffffffff0000000e00000000ffffffefffffffff0000001800000000",
            INIT_73 => X"00000041000000000000001600000000fffffff8ffffffffffffffe3ffffffff",
            INIT_74 => X"00000024000000000000000f000000000000000200000000ffffffc7ffffffff",
            INIT_75 => X"ffffffe4ffffffffffffffe3ffffffff0000000000000000ffffffdbffffffff",
            INIT_76 => X"fffffff0ffffffff000000220000000000000024000000000000002f00000000",
            INIT_77 => X"ffffffe7fffffffffffffffdffffffff0000002a000000000000000c00000000",
            INIT_78 => X"000000200000000000000022000000000000001300000000fffffff6ffffffff",
            INIT_79 => X"ffffffe8ffffffff000000140000000000000038000000000000001800000000",
            INIT_7A => X"ffffffc7ffffffff0000001d000000000000000f00000000ffffffdbffffffff",
            INIT_7B => X"0000001500000000fffffff1ffffffff0000000e00000000fffffffdffffffff",
            INIT_7C => X"00000009000000000000003000000000ffffffeafffffffffffffff6ffffffff",
            INIT_7D => X"000000150000000000000012000000000000001300000000ffffffbdffffffff",
            INIT_7E => X"0000001100000000fffffffbffffffffffffffffffffffffffffffeaffffffff",
            INIT_7F => X"ffffffe3ffffffffffffffdafffffffffffffffaffffffffffffffd9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE3;


    MEM_IWGHT_LAYER2_INSTANCE4 : if BRAM_NAME = "iwght_layer2_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000045000000000000003900000000ffffffe7ffffffff0000001200000000",
            INIT_01 => X"0000005d00000000ffffffcfffffffff00000016000000000000002300000000",
            INIT_02 => X"fffffffefffffffffffffffbffffffff0000000f000000000000001400000000",
            INIT_03 => X"000000070000000000000017000000000000002200000000ffffffd3ffffffff",
            INIT_04 => X"0000001a00000000000000380000000000000003000000000000000000000000",
            INIT_05 => X"0000000b0000000000000013000000000000001d000000000000001e00000000",
            INIT_06 => X"fffffff3ffffffff0000001f00000000ffffffebffffffffffffffeaffffffff",
            INIT_07 => X"00000028000000000000002d0000000000000023000000000000000100000000",
            INIT_08 => X"fffffff3ffffffff0000000d00000000ffffffecffffffff0000000000000000",
            INIT_09 => X"00000000000000000000001a000000000000000c00000000fffffffaffffffff",
            INIT_0A => X"ffffffccfffffffffffffff0ffffffff00000004000000000000000200000000",
            INIT_0B => X"fffffff8ffffffffffffffd4ffffffffffffffe4ffffffffffffffcbffffffff",
            INIT_0C => X"0000001c0000000000000026000000000000000d00000000fffffffaffffffff",
            INIT_0D => X"0000004000000000000000340000000000000044000000000000002700000000",
            INIT_0E => X"0000000b00000000ffffffffffffffffffffffe5ffffffffffffffeeffffffff",
            INIT_0F => X"00000005000000000000000b0000000000000025000000000000001900000000",
            INIT_10 => X"fffffff1ffffffffffffffe4ffffffffffffffebfffffffffffffff8ffffffff",
            INIT_11 => X"ffffffeaffffffffffffffeefffffffffffffff0ffffffff0000000100000000",
            INIT_12 => X"ffffffecffffffffffffffe9ffffffff00000009000000000000001100000000",
            INIT_13 => X"ffffffecffffffffffffffe4ffffffffffffffd0ffffffffffffffe8ffffffff",
            INIT_14 => X"fffffffafffffffffffffffeffffffff0000003600000000ffffffedffffffff",
            INIT_15 => X"ffffffdeffffffffffffffdfffffffffffffffb2fffffffffffffff4ffffffff",
            INIT_16 => X"fffffff5ffffffff0000002e00000000fffffff7ffffffff0000000200000000",
            INIT_17 => X"fffffff7ffffffffffffffedfffffffffffffffaffffffff0000000a00000000",
            INIT_18 => X"0000000000000000fffffff9ffffffff0000002b00000000fffffff7ffffffff",
            INIT_19 => X"fffffff8ffffffffffffffe9ffffffff0000001800000000fffffffbffffffff",
            INIT_1A => X"0000000900000000fffffffdffffffff0000001c00000000ffffffe6ffffffff",
            INIT_1B => X"0000001d00000000000000190000000000000012000000000000000000000000",
            INIT_1C => X"ffffffe9ffffffffffffffe0ffffffff00000011000000000000002700000000",
            INIT_1D => X"00000017000000000000000c000000000000000e000000000000004b00000000",
            INIT_1E => X"ffffffe3fffffffffffffffcffffffffffffffccffffffffffffffd3ffffffff",
            INIT_1F => X"0000000000000000fffffff8ffffffff0000001c000000000000000600000000",
            INIT_20 => X"00000006000000000000000800000000fffffffbfffffffffffffff4ffffffff",
            INIT_21 => X"000000150000000000000034000000000000000700000000fffffffaffffffff",
            INIT_22 => X"000000390000000000000006000000000000004b000000000000003000000000",
            INIT_23 => X"00000008000000000000002d000000000000001b000000000000000700000000",
            INIT_24 => X"0000001000000000ffffffd2ffffffff00000033000000000000000700000000",
            INIT_25 => X"ffffffbeffffffffffffffe8ffffffff00000015000000000000001d00000000",
            INIT_26 => X"0000001e00000000fffffff2ffffffff00000008000000000000001e00000000",
            INIT_27 => X"fffffffcfffffffffffffff9ffffffffffffffe0ffffffff0000000800000000",
            INIT_28 => X"fffffff7ffffffff0000000000000000fffffff3ffffffff0000000300000000",
            INIT_29 => X"fffffff8fffffffffffffffeffffffff0000000f000000000000000500000000",
            INIT_2A => X"0000002f000000000000003900000000fffffff2ffffffffffffffefffffffff",
            INIT_2B => X"ffffffefffffffffffffffedffffffff00000027000000000000003600000000",
            INIT_2C => X"0000000a00000000fffffffefffffffffffffffdffffffffffffffedffffffff",
            INIT_2D => X"00000003000000000000001900000000fffffffffffffffffffffff3ffffffff",
            INIT_2E => X"fffffff4ffffffffffffffddffffffffffffffeeffffffff0000001000000000",
            INIT_2F => X"0000000000000000000000100000000000000006000000000000000f00000000",
            INIT_30 => X"fffffff7fffffffffffffff2fffffffffffffffeffffffff0000001000000000",
            INIT_31 => X"00000019000000000000000e000000000000003000000000ffffffd6ffffffff",
            INIT_32 => X"ffffffb5ffffffffffffffc9ffffffffffffffe8ffffffff0000001900000000",
            INIT_33 => X"0000001700000000ffffffe4ffffffffffffffceffffffffffffffb9ffffffff",
            INIT_34 => X"00000002000000000000001300000000fffffff9ffffffff0000001600000000",
            INIT_35 => X"fffffffaffffffffffffffe8ffffffffffffffeffffffffffffffffcffffffff",
            INIT_36 => X"000000060000000000000025000000000000000600000000fffffffeffffffff",
            INIT_37 => X"ffffffecffffffffffffffebffffffffffffffecffffffff0000001b00000000",
            INIT_38 => X"0000000e0000000000000008000000000000000500000000fffffffaffffffff",
            INIT_39 => X"00000013000000000000001d000000000000001e00000000fffffffcffffffff",
            INIT_3A => X"000000170000000000000028000000000000003f000000000000002100000000",
            INIT_3B => X"ffffffebfffffffffffffff4ffffffffffffffcbffffffff0000001200000000",
            INIT_3C => X"0000000f00000000000000210000000000000002000000000000001600000000",
            INIT_3D => X"ffffffe3ffffffffffffffe2ffffffffffffffc6fffffffffffffffeffffffff",
            INIT_3E => X"00000012000000000000000100000000ffffffdcffffffffffffffe3ffffffff",
            INIT_3F => X"00000022000000000000002e000000000000003000000000ffffffebffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000100000000fffffff4ffffffff00000012000000000000001200000000",
            INIT_41 => X"00000000000000000000002e0000000000000043000000000000002600000000",
            INIT_42 => X"00000002000000000000000100000000ffffffdfffffffff0000001700000000",
            INIT_43 => X"0000000500000000ffffffeafffffffffffffffdfffffffffffffffaffffffff",
            INIT_44 => X"fffffff4fffffffffffffffdffffffff00000000000000000000000000000000",
            INIT_45 => X"00000018000000000000000f00000000fffffff6fffffffffffffff5ffffffff",
            INIT_46 => X"00000000000000000000000c00000000ffffffc3ffffffff0000001300000000",
            INIT_47 => X"ffffffebfffffffffffffff5ffffffff0000000400000000ffffffeeffffffff",
            INIT_48 => X"ffffffd8ffffffffffffffebffffffffffffffeefffffffffffffff5ffffffff",
            INIT_49 => X"00000019000000000000001b000000000000003300000000ffffffe7ffffffff",
            INIT_4A => X"00000014000000000000003c000000000000002e000000000000002700000000",
            INIT_4B => X"0000001100000000ffffffedffffffff00000061000000000000003100000000",
            INIT_4C => X"0000001300000000ffffffe4ffffffff0000002400000000fffffffaffffffff",
            INIT_4D => X"fffffffbffffffff000000190000000000000017000000000000002c00000000",
            INIT_4E => X"ffffffe7fffffffffffffff1fffffffffffffffbffffffff0000000500000000",
            INIT_4F => X"fffffffbfffffffffffffff4ffffffff0000000000000000ffffffe4ffffffff",
            INIT_50 => X"fffffffaffffffff0000000200000000fffffffbffffffffffffffe4ffffffff",
            INIT_51 => X"ffffffe8fffffffffffffffaffffffff00000006000000000000000000000000",
            INIT_52 => X"ffffffd7ffffffffffffffedfffffffffffffffeffffffff0000000300000000",
            INIT_53 => X"0000003300000000fffffff8ffffffffffffffffffffffffffffffe8ffffffff",
            INIT_54 => X"0000000800000000000000080000000000000036000000000000003e00000000",
            INIT_55 => X"ffffffadfffffffffffffffeffffffff0000001900000000ffffffebffffffff",
            INIT_56 => X"fffffffbffffffff000000150000000000000007000000000000000900000000",
            INIT_57 => X"ffffffd2ffffffffffffffe4fffffffffffffff1ffffffff0000002600000000",
            INIT_58 => X"ffffffe0ffffffffffffffd9ffffffffffffffb7ffffffffffffffe5ffffffff",
            INIT_59 => X"fffffffeffffffffffffffefffffffff0000000d000000000000002700000000",
            INIT_5A => X"0000000300000000ffffffe2fffffffffffffff0fffffffffffffff3ffffffff",
            INIT_5B => X"00000021000000000000001f00000000fffffffcffffffffffffffeaffffffff",
            INIT_5C => X"ffffffcbffffffff0000002c00000000ffffffefffffffffffffffedffffffff",
            INIT_5D => X"00000047000000000000000b000000000000000a00000000ffffffdcffffffff",
            INIT_5E => X"ffffffe3fffffffffffffff7ffffffffffffffedffffffff0000001400000000",
            INIT_5F => X"fffffff3fffffffffffffff1fffffffffffffffbfffffffffffffff9ffffffff",
            INIT_60 => X"0000003300000000000000020000000000000005000000000000003b00000000",
            INIT_61 => X"00000006000000000000000d00000000ffffffd8ffffffff0000001d00000000",
            INIT_62 => X"ffffffdfffffffff0000001b000000000000000e000000000000000100000000",
            INIT_63 => X"ffffffd2ffffffffffffffeafffffffffffffff8ffffffff0000000200000000",
            INIT_64 => X"0000001e000000000000001b00000000fffffffbffffffffffffffdfffffffff",
            INIT_65 => X"00000022000000000000001400000000fffffffaffffffff0000000400000000",
            INIT_66 => X"ffffffecffffffff00000002000000000000002c000000000000000d00000000",
            INIT_67 => X"0000001400000000ffffffdfffffffffffffffddffffffff0000000300000000",
            INIT_68 => X"fffffff9ffffffffffffffffffffffffffffffd9ffffffffffffffdcffffffff",
            INIT_69 => X"fffffffdffffffffffffffeaffffffff00000012000000000000003000000000",
            INIT_6A => X"ffffffbaffffffffffffffd7fffffffffffffff0ffffffffffffffd8ffffffff",
            INIT_6B => X"ffffffe6ffffffffffffffe1ffffffff00000017000000000000002500000000",
            INIT_6C => X"0000001a000000000000000f00000000ffffffb9fffffffffffffff9ffffffff",
            INIT_6D => X"0000000f00000000ffffffe2ffffffffffffffdcffffffff0000002800000000",
            INIT_6E => X"0000000700000000fffffffdfffffffffffffff6ffffffffffffffe4ffffffff",
            INIT_6F => X"0000000d00000000000000080000000000000016000000000000002100000000",
            INIT_70 => X"ffffffecffffffff0000001300000000fffffff8fffffffffffffffdffffffff",
            INIT_71 => X"ffffffdaffffffff00000002000000000000000e00000000fffffffaffffffff",
            INIT_72 => X"0000001d00000000000000000000000000000000000000000000002f00000000",
            INIT_73 => X"0000002b00000000000000430000000000000009000000000000001200000000",
            INIT_74 => X"ffffffedfffffffffffffff4ffffffffffffffadffffffff0000000600000000",
            INIT_75 => X"ffffffeaffffffff0000000000000000ffffffefffffffffffffffd3ffffffff",
            INIT_76 => X"ffffffeaffffffffffffffb8ffffffffffffffdeffffffffffffffddffffffff",
            INIT_77 => X"0000005600000000ffffffebffffffff0000000e00000000fffffff4ffffffff",
            INIT_78 => X"0000001a00000000fffffffdffffffff0000004c000000000000005c00000000",
            INIT_79 => X"ffffffcbffffffff0000000f00000000ffffffccffffffff0000001f00000000",
            INIT_7A => X"0000001200000000000000220000000000000013000000000000004100000000",
            INIT_7B => X"ffffffcafffffffffffffff0ffffffff00000014000000000000001300000000",
            INIT_7C => X"00000012000000000000002c00000000ffffffdfffffffffffffffc8ffffffff",
            INIT_7D => X"ffffffd3ffffffffffffffdfffffffffffffffc4ffffffff0000001700000000",
            INIT_7E => X"fffffffffffffffffffffffcfffffffffffffff0ffffffffffffffe4ffffffff",
            INIT_7F => X"00000007000000000000002800000000fffffff9fffffffffffffff6ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE4;


    MEM_IWGHT_LAYER2_INSTANCE5 : if BRAM_NAME = "iwght_layer2_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff1ffffffff000000010000000000000008000000000000000500000000",
            INIT_01 => X"0000002200000000ffffffd6ffffffff0000001f000000000000001f00000000",
            INIT_02 => X"ffffffecffffffff0000002d00000000fffffffefffffffffffffff2ffffffff",
            INIT_03 => X"ffffffd0fffffffffffffff7ffffffff0000000d00000000fffffffdffffffff",
            INIT_04 => X"0000000200000000ffffffcdffffffffffffffebffffffffffffffdaffffffff",
            INIT_05 => X"fffffff2ffffffff00000012000000000000002b00000000fffffffdffffffff",
            INIT_06 => X"ffffffe3ffffffffffffffadfffffffffffffff3ffffffffffffffd0ffffffff",
            INIT_07 => X"00000026000000000000004000000000ffffffc0fffffffffffffff1ffffffff",
            INIT_08 => X"fffffffdffffffff0000000900000000fffffffbffffffff0000002e00000000",
            INIT_09 => X"fffffffdffffffff0000000000000000fffffffdffffffffffffffedffffffff",
            INIT_0A => X"0000001b00000000ffffffe2fffffffffffffffcffffffff0000000000000000",
            INIT_0B => X"0000001300000000ffffffecffffffffffffffd7ffffffff0000001000000000",
            INIT_0C => X"ffffffd5ffffffffffffffdfffffffffffffffe9ffffffffffffffbdffffffff",
            INIT_0D => X"ffffffe2ffffffffffffffc8ffffffff0000002800000000ffffffd8ffffffff",
            INIT_0E => X"ffffffceffffffff0000000900000000ffffffe0ffffffff0000001a00000000",
            INIT_0F => X"fffffffbffffffffffffffe6ffffffffffffffebffffffff0000003200000000",
            INIT_10 => X"fffffff3ffffffffffffffe2ffffffffffffffd2ffffffffffffffe2ffffffff",
            INIT_11 => X"000000070000000000000047000000000000002f00000000fffffffeffffffff",
            INIT_12 => X"fffffffcfffffffffffffffeffffffff0000001d000000000000002800000000",
            INIT_13 => X"ffffffe0ffffffff0000001800000000ffffffd4ffffffff0000000f00000000",
            INIT_14 => X"fffffff5ffffffffffffffe4ffffffff0000000600000000fffffff1ffffffff",
            INIT_15 => X"fffffffaffffffffffffffd2ffffffffffffffe3ffffffff0000000300000000",
            INIT_16 => X"0000000000000000fffffff7ffffffff00000008000000000000002f00000000",
            INIT_17 => X"fffffff2ffffffffffffffe4ffffffffffffffd9ffffffff0000002d00000000",
            INIT_18 => X"ffffffcefffffffffffffff1ffffffff00000018000000000000002200000000",
            INIT_19 => X"ffffffd4ffffffffffffffdaffffffffffffffeeffffffffffffffd4ffffffff",
            INIT_1A => X"ffffffb8ffffffffffffffc4ffffffffffffffc2ffffffffffffffdfffffffff",
            INIT_1B => X"0000002000000000ffffffceffffffffffffffc5ffffffffffffffebffffffff",
            INIT_1C => X"00000017000000000000000a000000000000000a000000000000002400000000",
            INIT_1D => X"0000002a00000000fffffff8ffffffff00000027000000000000001100000000",
            INIT_1E => X"ffffffc5fffffffffffffffeffffffff0000000c000000000000002800000000",
            INIT_1F => X"fffffff7ffffffffffffffc4ffffffffffffffcdffffffffffffffe3ffffffff",
            INIT_20 => X"0000000000000000fffffff7ffffffffffffffffffffffffffffffd8ffffffff",
            INIT_21 => X"0000000400000000ffffffe7ffffffffffffffefffffffffffffffeaffffffff",
            INIT_22 => X"fffffff8ffffffff0000001e00000000fffffffdffffffff0000001000000000",
            INIT_23 => X"0000001e00000000fffffff4ffffffff00000008000000000000001200000000",
            INIT_24 => X"ffffffc6ffffffff0000000300000000fffffffaffffffffffffffecffffffff",
            INIT_25 => X"fffffffeffffffff0000002200000000fffffff5ffffffffffffffccffffffff",
            INIT_26 => X"0000000000000000ffffffe6ffffffffffffffe8ffffffff0000000200000000",
            INIT_27 => X"000000270000000000000006000000000000000700000000fffffff9ffffffff",
            INIT_28 => X"0000002b000000000000001d0000000000000037000000000000005d00000000",
            INIT_29 => X"ffffffb6ffffffffffffffd7ffffffffffffffc2ffffffff0000001300000000",
            INIT_2A => X"0000000000000000ffffffd5ffffffffffffffe8fffffffffffffff0ffffffff",
            INIT_2B => X"00000008000000000000001400000000fffffff6ffffffffffffffddffffffff",
            INIT_2C => X"00000024000000000000000b000000000000000d000000000000000200000000",
            INIT_2D => X"000000020000000000000018000000000000000100000000ffffffffffffffff",
            INIT_2E => X"0000001e0000000000000023000000000000000800000000fffffffcffffffff",
            INIT_2F => X"ffffffbaffffffffffffffd2ffffffffffffffe0ffffffff0000000000000000",
            INIT_30 => X"fffffffbffffffffffffffb9ffffffffffffffe7ffffffffffffffdbffffffff",
            INIT_31 => X"ffffffc3ffffffff000000110000000000000025000000000000000400000000",
            INIT_32 => X"0000001e00000000ffffffedffffffff0000001d00000000fffffff8ffffffff",
            INIT_33 => X"00000017000000000000001000000000fffffff7fffffffffffffffeffffffff",
            INIT_34 => X"00000025000000000000001f0000000000000043000000000000002300000000",
            INIT_35 => X"00000000000000000000000d0000000000000000000000000000001c00000000",
            INIT_36 => X"fffffff9fffffffffffffffefffffffffffffff4fffffffffffffff3ffffffff",
            INIT_37 => X"00000004000000000000001300000000fffffff6fffffffffffffff6ffffffff",
            INIT_38 => X"ffffffeeffffffff000000000000000000000007000000000000000000000000",
            INIT_39 => X"00000017000000000000000b000000000000000900000000fffffff8ffffffff",
            INIT_3A => X"00000019000000000000000700000000fffffff6ffffffff0000000b00000000",
            INIT_3B => X"0000001800000000000000150000000000000016000000000000000200000000",
            INIT_3C => X"0000000000000000ffffffdaffffffff0000000100000000ffffffe8ffffffff",
            INIT_3D => X"00000004000000000000002d000000000000000a00000000fffffffbffffffff",
            INIT_3E => X"ffffffd1ffffffffffffffcfffffffffffffffe0ffffffff0000001900000000",
            INIT_3F => X"0000000f00000000000000160000000000000024000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff9fffffffffffffff7ffffffff0000000f000000000000002a00000000",
            INIT_41 => X"ffffffd1ffffffffffffffd4ffffffffffffffe2ffffffffffffffcfffffffff",
            INIT_42 => X"0000000b00000000fffffff3fffffffffffffffaffffffff0000000600000000",
            INIT_43 => X"fffffff3ffffffffffffffd7ffffffff0000000900000000fffffff4ffffffff",
            INIT_44 => X"ffffffd5ffffffff0000000e00000000ffffffc8ffffffffffffffb6ffffffff",
            INIT_45 => X"0000001200000000ffffffa1ffffffffffffffeaffffffffffffffe3ffffffff",
            INIT_46 => X"0000002900000000000000550000000000000018000000000000001e00000000",
            INIT_47 => X"0000002f0000000000000013000000000000001a000000000000002a00000000",
            INIT_48 => X"0000001500000000fffffff7ffffffffffffffeafffffffffffffffdffffffff",
            INIT_49 => X"0000001f000000000000000c000000000000000700000000fffffffaffffffff",
            INIT_4A => X"0000000900000000000000230000000000000055000000000000004f00000000",
            INIT_4B => X"ffffffd5ffffffffffffffffffffffff00000003000000000000002500000000",
            INIT_4C => X"0000000b00000000fffffff2ffffffffffffffcaffffffffffffffa2ffffffff",
            INIT_4D => X"fffffff1ffffffffffffffe3ffffffff0000000300000000ffffffc7ffffffff",
            INIT_4E => X"fffffffbffffffffffffffa2ffffffffffffffa0ffffffffffffffbcffffffff",
            INIT_4F => X"000000470000000000000047000000000000000900000000ffffffeeffffffff",
            INIT_50 => X"ffffffddffffffffffffffdbfffffffffffffff0ffffffff0000003100000000",
            INIT_51 => X"fffffffdffffffff000000110000000000000018000000000000002700000000",
            INIT_52 => X"0000002300000000000000120000000000000025000000000000000f00000000",
            INIT_53 => X"fffffffbffffffff0000003d00000000ffffffecffffffff0000001600000000",
            INIT_54 => X"ffffffd7ffffffff0000000f000000000000001e00000000ffffffdcffffffff",
            INIT_55 => X"ffffffe8fffffffffffffff6ffffffffffffffdfffffffffffffff8bffffffff",
            INIT_56 => X"fffffffcffffffffffffffedffffffffffffffcdffffffffffffffdaffffffff",
            INIT_57 => X"0000001b00000000ffffffe3ffffffff0000000400000000fffffff9ffffffff",
            INIT_58 => X"00000001000000000000002800000000fffffff3ffffffff0000000500000000",
            INIT_59 => X"0000001500000000000000170000000000000028000000000000000f00000000",
            INIT_5A => X"00000020000000000000001800000000fffffffdffffffffffffffe9ffffffff",
            INIT_5B => X"ffffffbeffffffffffffffbbffffffff0000000e000000000000000f00000000",
            INIT_5C => X"fffffffeffffffff0000000d000000000000000400000000ffffffe9ffffffff",
            INIT_5D => X"00000046000000000000002a0000000000000010000000000000002700000000",
            INIT_5E => X"ffffffebfffffffffffffff7ffffffff00000033000000000000004a00000000",
            INIT_5F => X"ffffffceffffffffffffffd3ffffffffffffffc9ffffffff0000002100000000",
            INIT_60 => X"fffffff9ffffffff00000001000000000000001b000000000000000700000000",
            INIT_61 => X"ffffffe4ffffffffffffffedffffffffffffffedffffffff0000000a00000000",
            INIT_62 => X"0000000600000000fffffff4ffffffffffffffebffffffff0000001000000000",
            INIT_63 => X"ffffffe3ffffffff0000001a000000000000000600000000fffffffeffffffff",
            INIT_64 => X"ffffffdafffffffffffffff3ffffffffffffffe6ffffffffffffffbdffffffff",
            INIT_65 => X"0000002700000000fffffffcffffffff0000000500000000ffffffdfffffffff",
            INIT_66 => X"0000000500000000000000180000000000000022000000000000000600000000",
            INIT_67 => X"ffffffcfffffffffffffffd5ffffffff0000001e000000000000000d00000000",
            INIT_68 => X"ffffffeaffffffffffffffdbfffffffffffffff0ffffffff0000000400000000",
            INIT_69 => X"ffffffe0ffffffffffffffeaffffffffffffffd9ffffffffffffffe0ffffffff",
            INIT_6A => X"00000008000000000000000000000000ffffffeaffffffffffffffe6ffffffff",
            INIT_6B => X"0000000000000000ffffffc6ffffffffffffffd8ffffffff0000000900000000",
            INIT_6C => X"0000002200000000ffffffeaffffffff0000003000000000fffffffeffffffff",
            INIT_6D => X"ffffffb2ffffffffffffffc3fffffffffffffff0ffffffff0000001500000000",
            INIT_6E => X"00000023000000000000003a000000000000003b00000000fffffff8ffffffff",
            INIT_6F => X"00000010000000000000001d0000000000000025000000000000004200000000",
            INIT_70 => X"fffffff5ffffffffffffffeaffffffff0000001c00000000fffffff8ffffffff",
            INIT_71 => X"0000000a00000000fffffff7fffffffffffffff9ffffffffffffffe1ffffffff",
            INIT_72 => X"fffffff2ffffffffffffffe6ffffffffffffffeefffffffffffffffaffffffff",
            INIT_73 => X"00000008000000000000001900000000ffffffe5ffffffffffffffecffffffff",
            INIT_74 => X"ffffffe3ffffffffffffffe7ffffffffffffffd1ffffffff0000001000000000",
            INIT_75 => X"0000000b00000000000000000000000000000026000000000000002000000000",
            INIT_76 => X"0000000a000000000000001200000000fffffffbffffffff0000000e00000000",
            INIT_77 => X"fffffff3ffffffff0000000e00000000fffffff6ffffffff0000001200000000",
            INIT_78 => X"ffffffdcffffffffffffffefffffffff0000000300000000ffffffe0ffffffff",
            INIT_79 => X"00000028000000000000001a00000000ffffffd7ffffffffffffffa2ffffffff",
            INIT_7A => X"0000000800000000000000000000000000000009000000000000001b00000000",
            INIT_7B => X"0000000100000000ffffffeffffffffffffffffaffffffff0000004500000000",
            INIT_7C => X"00000001000000000000000700000000ffffffe0ffffffffffffffeeffffffff",
            INIT_7D => X"0000001a00000000fffffff2ffffffffffffffc3fffffffffffffff9ffffffff",
            INIT_7E => X"00000021000000000000000e0000000000000020000000000000000b00000000",
            INIT_7F => X"ffffffeeffffffff000000030000000000000028000000000000000a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE5;


    MEM_IWGHT_LAYER2_INSTANCE6 : if BRAM_NAME = "iwght_layer2_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000100000000ffffffeeffffffff0000000d00000000fffffff5ffffffff",
            INIT_01 => X"0000000000000000ffffffefffffffff00000010000000000000001300000000",
            INIT_02 => X"0000002c000000000000002b000000000000000100000000ffffffd1ffffffff",
            INIT_03 => X"fffffff6ffffffff000000070000000000000012000000000000002100000000",
            INIT_04 => X"fffffffcffffffffffffffe6ffffffffffffffe4ffffffffffffffdaffffffff",
            INIT_05 => X"000000140000000000000027000000000000001300000000fffffff4ffffffff",
            INIT_06 => X"0000002000000000ffffffe5ffffffff0000001c000000000000003c00000000",
            INIT_07 => X"ffffffc0ffffffffffffffeaffffffffffffffebffffffff0000001900000000",
            INIT_08 => X"ffffffebffffffff0000002100000000fffffff5ffffffffffffffbfffffffff",
            INIT_09 => X"ffffffc5ffffffffffffff8dffffffff0000001d000000000000000c00000000",
            INIT_0A => X"ffffffc9ffffffff000000060000000000000000000000000000000300000000",
            INIT_0B => X"ffffffddffffffffffffffe4fffffffffffffffaffffffff0000000e00000000",
            INIT_0C => X"fffffff8ffffffffffffffdbffffffff0000000400000000ffffffc8ffffffff",
            INIT_0D => X"0000000800000000fffffff4ffffffffffffffdefffffffffffffff6ffffffff",
            INIT_0E => X"fffffff4ffffffff000000220000000000000012000000000000003400000000",
            INIT_0F => X"0000001700000000ffffffe6ffffffffffffffbfffffffffffffffe7ffffffff",
            INIT_10 => X"0000002300000000000000030000000000000016000000000000003500000000",
            INIT_11 => X"ffffffdeffffffffffffffffffffffff00000013000000000000003000000000",
            INIT_12 => X"0000000c0000000000000003000000000000003a00000000ffffffc3ffffffff",
            INIT_13 => X"0000001c00000000ffffffffffffffffffffffd0ffffffffffffffecffffffff",
            INIT_14 => X"0000001300000000000000000000000000000018000000000000000900000000",
            INIT_15 => X"ffffffdbfffffffffffffff9fffffffffffffffcffffffff0000001200000000",
            INIT_16 => X"00000020000000000000001f00000000fffffff9ffffffff0000000f00000000",
            INIT_17 => X"ffffffa3ffffffffffffffeaffffffff0000000000000000fffffffbffffffff",
            INIT_18 => X"ffffffd4ffffffffffffffdfffffffff0000000200000000fffffff4ffffffff",
            INIT_19 => X"ffffffecffffffff00000013000000000000001c000000000000002400000000",
            INIT_1A => X"0000001e000000000000001700000000ffffffdfffffffffffffffe5ffffffff",
            INIT_1B => X"fffffffcfffffffffffffff8ffffffff0000000d000000000000003900000000",
            INIT_1C => X"fffffffcfffffffffffffff5ffffffff0000001a000000000000001800000000",
            INIT_1D => X"fffffffdffffffff00000006000000000000001700000000ffffffffffffffff",
            INIT_1E => X"ffffffd6fffffffffffffff9ffffffff0000002100000000fffffffaffffffff",
            INIT_1F => X"fffffffdffffffffffffffdfffffffffffffffc7ffffffffffffffddffffffff",
            INIT_20 => X"0000004c000000000000001c0000000000000011000000000000002700000000",
            INIT_21 => X"ffffffeefffffffffffffff1ffffffffffffffcfffffffff0000002100000000",
            INIT_22 => X"0000001b0000000000000041000000000000002b000000000000005400000000",
            INIT_23 => X"fffffffaffffffffffffffe4fffffffffffffff8fffffffffffffffeffffffff",
            INIT_24 => X"0000002c000000000000000200000000fffffffaffffffff0000001700000000",
            INIT_25 => X"ffffffe4ffffffff0000001400000000fffffff8fffffffffffffff9ffffffff",
            INIT_26 => X"00000010000000000000001f000000000000000300000000fffffffeffffffff",
            INIT_27 => X"0000003000000000000000200000000000000032000000000000001100000000",
            INIT_28 => X"0000000200000000fffffffbfffffffffffffff2ffffffffffffffedffffffff",
            INIT_29 => X"00000042000000000000001f0000000000000018000000000000000500000000",
            INIT_2A => X"00000011000000000000001b00000000ffffffdcffffffff0000001c00000000",
            INIT_2B => X"ffffffe5ffffffff0000002f00000000fffffff7ffffffffffffffdcffffffff",
            INIT_2C => X"0000002b000000000000002300000000fffffff8ffffffffffffffe4ffffffff",
            INIT_2D => X"fffffffdffffffff000000000000000000000000000000000000000d00000000",
            INIT_2E => X"fffffff5ffffffff0000000200000000fffffff0ffffffff0000002300000000",
            INIT_2F => X"0000000300000000ffffffecffffffff0000003100000000ffffffebffffffff",
            INIT_30 => X"00000005000000000000000c000000000000000f000000000000001e00000000",
            INIT_31 => X"fffffff9ffffffff0000001e0000000000000021000000000000002500000000",
            INIT_32 => X"00000000000000000000000f00000000ffffffdeffffffff0000000700000000",
            INIT_33 => X"0000002600000000ffffffe4ffffffffffffffdeffffffffffffffebffffffff",
            INIT_34 => X"00000029000000000000000c000000000000001b000000000000000c00000000",
            INIT_35 => X"0000001100000000fffffff2ffffffffffffffddffffffff0000000900000000",
            INIT_36 => X"0000000f000000000000001f0000000000000033000000000000003700000000",
            INIT_37 => X"ffffffcbffffffffffffffc6ffffffff0000001b000000000000003500000000",
            INIT_38 => X"0000000a000000000000000300000000ffffffe7ffffffffffffffc6ffffffff",
            INIT_39 => X"0000001c000000000000001e0000000000000023000000000000002600000000",
            INIT_3A => X"00000002000000000000000f000000000000000a000000000000000200000000",
            INIT_3B => X"ffffffedffffffffffffffeafffffffffffffff3ffffffff0000000b00000000",
            INIT_3C => X"00000014000000000000001300000000ffffffeefffffffffffffff7ffffffff",
            INIT_3D => X"fffffffdfffffffffffffffdffffffff00000003000000000000000800000000",
            INIT_3E => X"ffffffe4ffffffff00000002000000000000000c000000000000000100000000",
            INIT_3F => X"0000001d00000000000000000000000000000014000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffc9ffffffff00000034000000000000001c000000000000002b00000000",
            INIT_41 => X"0000002c00000000000000130000000000000036000000000000000400000000",
            INIT_42 => X"ffffffd8fffffffffffffff9ffffffff0000001700000000fffffff6ffffffff",
            INIT_43 => X"ffffffddffffffff0000000400000000ffffffefffffffffffffffb0ffffffff",
            INIT_44 => X"00000008000000000000003100000000fffffff2ffffffffffffffd8ffffffff",
            INIT_45 => X"000000040000000000000006000000000000000f00000000ffffffe9ffffffff",
            INIT_46 => X"ffffffbfffffffffffffffe5ffffffffffffffceffffffffffffffeaffffffff",
            INIT_47 => X"0000000e00000000ffffffedffffffffffffffe6ffffffffffffffc7ffffffff",
            INIT_48 => X"0000000d0000000000000011000000000000000500000000fffffff0ffffffff",
            INIT_49 => X"fffffff3fffffffffffffffcffffffff00000015000000000000000500000000",
            INIT_4A => X"fffffff0ffffffff0000000d00000000ffffffe7ffffffff0000002300000000",
            INIT_4B => X"fffffffcffffffff0000001c0000000000000011000000000000000800000000",
            INIT_4C => X"fffffffaffffffff0000000d0000000000000023000000000000000d00000000",
            INIT_4D => X"ffffffcbfffffffffffffff8fffffffffffffffcfffffffffffffff3ffffffff",
            INIT_4E => X"0000002a000000000000000a00000000ffffffefffffffffffffffecffffffff",
            INIT_4F => X"fffffff4fffffffffffffff7fffffffffffffff0ffffffff0000000000000000",
            INIT_50 => X"ffffffe8ffffffffffffffe5ffffffff0000001000000000ffffffd0ffffffff",
            INIT_51 => X"ffffffdaffffffff0000000a00000000ffffffe4ffffffffffffffe8ffffffff",
            INIT_52 => X"00000032000000000000000000000000fffffff7ffffffff0000000600000000",
            INIT_53 => X"000000210000000000000000000000000000003c000000000000001f00000000",
            INIT_54 => X"ffffffecffffffffffffffe9ffffffffffffffe4fffffffffffffffeffffffff",
            INIT_55 => X"0000002700000000000000200000000000000038000000000000003a00000000",
            INIT_56 => X"0000001900000000fffffff1ffffffff0000000400000000fffffffcffffffff",
            INIT_57 => X"fffffffdffffffff0000001000000000ffffffe7ffffffff0000000000000000",
            INIT_58 => X"0000002a00000000fffffff9ffffffffffffffc6ffffffff0000001800000000",
            INIT_59 => X"ffffffa5ffffffffffffffc8ffffffffffffffd1ffffffff0000000000000000",
            INIT_5A => X"0000001300000000fffffff1ffffffff0000000f00000000ffffffeeffffffff",
            INIT_5B => X"000000160000000000000029000000000000000000000000fffffffbffffffff",
            INIT_5C => X"0000000700000000fffffff8ffffffffffffffeffffffffffffffffbffffffff",
            INIT_5D => X"00000024000000000000002b000000000000000b000000000000000b00000000",
            INIT_5E => X"00000006000000000000001d0000000000000003000000000000001b00000000",
            INIT_5F => X"0000001e000000000000001c000000000000002d000000000000000100000000",
            INIT_60 => X"0000002100000000fffffff9fffffffffffffffbffffffff0000000c00000000",
            INIT_61 => X"00000037000000000000001d000000000000002300000000fffffffdffffffff",
            INIT_62 => X"ffffffdbffffffff000000110000000000000022000000000000002b00000000",
            INIT_63 => X"0000000f000000000000002d000000000000000a00000000ffffffffffffffff",
            INIT_64 => X"ffffffe9ffffffff0000001e0000000000000029000000000000000600000000",
            INIT_65 => X"fffffff2ffffffff0000000c00000000ffffffdcffffffffffffffdaffffffff",
            INIT_66 => X"0000003f000000000000004500000000ffffffeffffffffffffffffcffffffff",
            INIT_67 => X"0000001f000000000000003b000000000000004c000000000000004900000000",
            INIT_68 => X"ffffffe7ffffffff0000001b0000000000000001000000000000002000000000",
            INIT_69 => X"fffffffdffffffffffffffdbffffffff0000000c00000000ffffffe7ffffffff",
            INIT_6A => X"ffffffe5ffffffffffffffdffffffffffffffff1ffffffffffffffdbffffffff",
            INIT_6B => X"00000034000000000000001700000000ffffffe3ffffffff0000000000000000",
            INIT_6C => X"fffffffcffffffffffffffeaffffffffffffffe0ffffffff0000001d00000000",
            INIT_6D => X"fffffffefffffffffffffffaffffffffffffffd8ffffffffffffffdeffffffff",
            INIT_6E => X"ffffffe2ffffffff0000002300000000fffffffeffffffff0000001b00000000",
            INIT_6F => X"0000001000000000fffffff1fffffffffffffff9ffffffff0000000b00000000",
            INIT_70 => X"fffffff5ffffffff0000000f000000000000000e000000000000001000000000",
            INIT_71 => X"0000000900000000ffffffe0ffffffff00000009000000000000000200000000",
            INIT_72 => X"ffffffc0ffffffffffffff96ffffffffffffffa1ffffffffffffffe7ffffffff",
            INIT_73 => X"0000001f00000000000000130000000000000030000000000000001500000000",
            INIT_74 => X"ffffffefffffffff00000000000000000000002d000000000000000a00000000",
            INIT_75 => X"00000007000000000000001600000000fffffffbfffffffffffffff1ffffffff",
            INIT_76 => X"0000001e00000000000000240000000000000019000000000000001400000000",
            INIT_77 => X"000000000000000000000006000000000000002f00000000fffffff3ffffffff",
            INIT_78 => X"ffffffe9ffffffff00000019000000000000002200000000ffffffecffffffff",
            INIT_79 => X"00000025000000000000000400000000fffffffaffffffff0000000600000000",
            INIT_7A => X"0000001f0000000000000032000000000000000300000000ffffffeeffffffff",
            INIT_7B => X"fffffff3ffffffff0000002600000000ffffffefffffffff0000000900000000",
            INIT_7C => X"0000004200000000fffffff2ffffffff00000018000000000000001a00000000",
            INIT_7D => X"00000024000000000000000800000000ffffffe5ffffffff0000003000000000",
            INIT_7E => X"00000015000000000000002b0000000000000027000000000000001700000000",
            INIT_7F => X"0000000500000000ffffffccfffffffffffffff8ffffffff0000000800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE6;


    MEM_IWGHT_LAYER2_INSTANCE7 : if BRAM_NAME = "iwght_layer2_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff9ffffffff0000001800000000ffffffe2ffffffff0000000100000000",
            INIT_01 => X"ffffffe2ffffffffffffffe3fffffffffffffff8ffffffffffffffdfffffffff",
            INIT_02 => X"000000080000000000000032000000000000001f000000000000002200000000",
            INIT_03 => X"0000000000000000fffffffaffffffff0000002e000000000000000300000000",
            INIT_04 => X"ffffffc4fffffffffffffff5ffffffffffffffe3ffffffff0000000e00000000",
            INIT_05 => X"fffffff7ffffffffffffffe1ffffffff0000003600000000fffffff7ffffffff",
            INIT_06 => X"0000001c000000000000001200000000fffffff6ffffffff0000002e00000000",
            INIT_07 => X"ffffffe8ffffffff000000030000000000000005000000000000000000000000",
            INIT_08 => X"fffffffbfffffffffffffff3ffffffff0000000e00000000fffffff0ffffffff",
            INIT_09 => X"0000003100000000000000340000000000000007000000000000002c00000000",
            INIT_0A => X"ffffffd7ffffffff0000000200000000ffffffeeffffffff0000004000000000",
            INIT_0B => X"0000002200000000000000270000000000000031000000000000001a00000000",
            INIT_0C => X"00000027000000000000000b00000000fffffffeffffffff0000002600000000",
            INIT_0D => X"0000000000000000fffffffdffffffffffffffecffffffff0000002c00000000",
            INIT_0E => X"fffffff2ffffffff00000007000000000000000d00000000ffffffe7ffffffff",
            INIT_0F => X"fffffffeffffffffffffffecffffffff00000018000000000000004600000000",
            INIT_10 => X"00000001000000000000000900000000fffffff8ffffffff0000000000000000",
            INIT_11 => X"00000014000000000000000a0000000000000011000000000000000500000000",
            INIT_12 => X"00000019000000000000000a0000000000000002000000000000002900000000",
            INIT_13 => X"ffffffedffffffffffffffefffffffffffffffafffffffff0000003000000000",
            INIT_14 => X"fffffff4ffffffff0000001400000000ffffffceffffffffffffffe0ffffffff",
            INIT_15 => X"ffffffedffffffffffffffedffffffff0000000500000000ffffffd8ffffffff",
            INIT_16 => X"fffffff7ffffffff0000001600000000fffffff2ffffffff0000001a00000000",
            INIT_17 => X"0000000e000000000000000800000000fffffffbffffffffffffffddffffffff",
            INIT_18 => X"0000002400000000fffffff1ffffffff00000007000000000000001700000000",
            INIT_19 => X"ffffffddffffffff0000001f00000000ffffffe1ffffffffffffffe8ffffffff",
            INIT_1A => X"ffffffccffffffffffffffffffffffff00000042000000000000001700000000",
            INIT_1B => X"ffffffc8ffffffffffffffb0ffffffff00000003000000000000002400000000",
            INIT_1C => X"ffffffe1ffffffff0000000a00000000ffffffe7ffffffffffffffe4ffffffff",
            INIT_1D => X"ffffffe7ffffffff0000000a00000000ffffffdbfffffffffffffff8ffffffff",
            INIT_1E => X"ffffffcaffffffff00000002000000000000002000000000ffffffc6ffffffff",
            INIT_1F => X"00000004000000000000002000000000fffffff2ffffffff0000000600000000",
            INIT_20 => X"fffffffdfffffffffffffff2ffffffff0000000d000000000000000700000000",
            INIT_21 => X"ffffffbcffffffffffffffb6ffffffffffffffedffffffffffffffefffffffff",
            INIT_22 => X"0000003500000000000000500000000000000018000000000000001000000000",
            INIT_23 => X"0000002000000000fffffff7ffffffff0000000500000000fffffff3ffffffff",
            INIT_24 => X"00000020000000000000000c000000000000001b000000000000003c00000000",
            INIT_25 => X"00000016000000000000001000000000ffffffe2fffffffffffffff6ffffffff",
            INIT_26 => X"fffffff7fffffffffffffff9ffffffffffffffe0ffffffffffffffe3ffffffff",
            INIT_27 => X"ffffffc2ffffffffffffffcdffffffff0000001c00000000ffffffe2ffffffff",
            INIT_28 => X"fffffffaffffffff0000000a00000000fffffff1ffffffffffffffe2ffffffff",
            INIT_29 => X"000000000000000000000015000000000000001100000000ffffffdeffffffff",
            INIT_2A => X"ffffffe0fffffffffffffff6ffffffffffffffe5ffffffff0000001300000000",
            INIT_2B => X"fffffff6ffffffffffffffedfffffffffffffffbfffffffffffffff0ffffffff",
            INIT_2C => X"0000001400000000fffffffcffffffffffffffdcffffffff0000000100000000",
            INIT_2D => X"0000002100000000fffffff4fffffffffffffff7ffffffff0000003b00000000",
            INIT_2E => X"ffffffeeffffffff0000001f00000000fffffffaffffffff0000000900000000",
            INIT_2F => X"ffffffe5fffffffffffffff0ffffffffffffffc2ffffffff0000000300000000",
            INIT_30 => X"ffffffe9ffffffff0000000000000000ffffffeaffffffffffffffb1ffffffff",
            INIT_31 => X"ffffffd2ffffffff0000000f000000000000002000000000fffffff7ffffffff",
            INIT_32 => X"0000002a00000000fffffff1ffffffff00000019000000000000004700000000",
            INIT_33 => X"ffffffeaffffffff0000000000000000fffffff9ffffffff0000002700000000",
            INIT_34 => X"0000000d00000000ffffffd8fffffffffffffffaffffffff0000002300000000",
            INIT_35 => X"fffffff8ffffffff0000002c00000000ffffffd3ffffffffffffffd1ffffffff",
            INIT_36 => X"fffffffeffffffffffffffe4ffffffff0000001400000000fffffff7ffffffff",
            INIT_37 => X"00000020000000000000000800000000ffffffc0fffffffffffffffbffffffff",
            INIT_38 => X"ffffffe0ffffffffffffffbcffffffffffffffe5ffffffffffffffcaffffffff",
            INIT_39 => X"00000024000000000000000200000000fffffffdffffffff0000001500000000",
            INIT_3A => X"0000002c00000000000000130000000000000024000000000000001000000000",
            INIT_3B => X"ffffffebffffffff0000000300000000ffffffbeffffffff0000002200000000",
            INIT_3C => X"00000033000000000000000c00000000ffffffa1ffffffffffffffd3ffffffff",
            INIT_3D => X"00000051000000000000000a0000000000000004000000000000002c00000000",
            INIT_3E => X"00000024000000000000000000000000ffffffdaffffffffffffffdcffffffff",
            INIT_3F => X"00000029000000000000001000000000fffffff5ffffffff0000000600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffddffffffff0000000b00000000fffffff9ffffffffffffffdbffffffff",
            INIT_41 => X"0000000500000000ffffffdaffffffff0000000900000000fffffff2ffffffff",
            INIT_42 => X"00000029000000000000000100000000fffffffaffffffff0000001400000000",
            INIT_43 => X"ffffffe8ffffffffffffffb9ffffffffffffffdcffffffff0000000600000000",
            INIT_44 => X"0000001a00000000fffffffcfffffffffffffff8ffffffff0000003400000000",
            INIT_45 => X"ffffffe9ffffffffffffffd3ffffffff0000001f000000000000001e00000000",
            INIT_46 => X"0000000200000000ffffffd6fffffffffffffff6fffffffffffffffaffffffff",
            INIT_47 => X"ffffffccfffffffffffffff6ffffffff00000009000000000000000200000000",
            INIT_48 => X"ffffffc7ffffffffffffffbdffffffffffffffdfffffffffffffffc2ffffffff",
            INIT_49 => X"ffffffe7fffffffffffffff4ffffffffffffffcdffffffffffffffcfffffffff",
            INIT_4A => X"ffffffdfffffffffffffffd1ffffffff0000000000000000fffffffeffffffff",
            INIT_4B => X"0000000d00000000ffffffdfffffffffffffffe9ffffffff0000000000000000",
            INIT_4C => X"0000002b00000000000000240000000000000002000000000000001000000000",
            INIT_4D => X"0000003e000000000000003a00000000fffffff4ffffffff0000003900000000",
            INIT_4E => X"fffffffaffffffffffffffd8ffffffff00000012000000000000002300000000",
            INIT_4F => X"ffffffd9ffffffffffffffe5ffffffff0000000500000000ffffffe9ffffffff",
            INIT_50 => X"00000013000000000000000a00000000fffffff9ffffffff0000000d00000000",
            INIT_51 => X"ffffffeeffffffff0000002300000000fffffff7ffffffffffffffe1ffffffff",
            INIT_52 => X"ffffffc4ffffffffffffffbdffffffffffffffa6ffffffffffffffd5ffffffff",
            INIT_53 => X"ffffffb3ffffffff00000008000000000000002600000000fffffff7ffffffff",
            INIT_54 => X"fffffffbffffffffffffffc2ffffffff0000000e00000000ffffffdcffffffff",
            INIT_55 => X"0000002300000000ffffffd9fffffffffffffffbffffffffffffffecffffffff",
            INIT_56 => X"0000002e000000000000000900000000ffffffcdfffffffffffffff4ffffffff",
            INIT_57 => X"0000000b00000000000000140000000000000021000000000000002800000000",
            INIT_58 => X"fffffff3ffffffffffffffedffffffffffffffedffffffff0000001000000000",
            INIT_59 => X"fffffff8fffffffffffffffbffffffffffffffecffffffffffffffffffffffff",
            INIT_5A => X"ffffffbcffffffffffffffe7ffffffff00000005000000000000000b00000000",
            INIT_5B => X"ffffffc7ffffffffffffff93ffffffffffffffbeffffffffffffffabffffffff",
            INIT_5C => X"ffffffebffffffff0000001c0000000000000019000000000000000d00000000",
            INIT_5D => X"fffffffdffffffff00000011000000000000000b00000000fffffff3ffffffff",
            INIT_5E => X"0000000c000000000000002e0000000000000008000000000000000000000000",
            INIT_5F => X"0000000600000000000000220000000000000025000000000000003b00000000",
            INIT_60 => X"00000019000000000000002100000000fffffffcffffffff0000000900000000",
            INIT_61 => X"000000460000000000000000000000000000001e000000000000003d00000000",
            INIT_62 => X"0000001900000000ffffffe7ffffffffffffffd5ffffffffffffffe6ffffffff",
            INIT_63 => X"0000002c000000000000002500000000ffffffd7ffffffffffffffefffffffff",
            INIT_64 => X"fffffff9fffffffffffffff9ffffffff0000000b00000000ffffffbfffffffff",
            INIT_65 => X"ffffffffffffffff000000250000000000000026000000000000000600000000",
            INIT_66 => X"fffffffcffffffff0000001a000000000000000d000000000000001a00000000",
            INIT_67 => X"ffffffe7ffffffff0000000200000000fffffff1ffffffff0000000c00000000",
            INIT_68 => X"ffffffe6ffffffffffffffc8ffffffffffffffcafffffffffffffffeffffffff",
            INIT_69 => X"ffffffebffffffffffffffe0ffffffffffffffedffffffffffffffe1ffffffff",
            INIT_6A => X"ffffffd8ffffffffffffff79ffffffffffffffd8ffffffffffffffdeffffffff",
            INIT_6B => X"ffffffcfffffffffffffffe7ffffffffffffffdaffffffffffffffdbffffffff",
            INIT_6C => X"ffffffe6fffffffffffffff2ffffffff0000002d00000000ffffffe6ffffffff",
            INIT_6D => X"ffffffc0ffffffffffffffb2ffffffffffffffcaffffffff0000002d00000000",
            INIT_6E => X"000000000000000000000018000000000000001e000000000000000600000000",
            INIT_6F => X"ffffffe1fffffffffffffffcffffffff0000001600000000fffffff6ffffffff",
            INIT_70 => X"fffffff6ffffffffffffffecfffffffffffffff0fffffffffffffff2ffffffff",
            INIT_71 => X"0000000b00000000000000080000000000000012000000000000000000000000",
            INIT_72 => X"0000001e000000000000001b0000000000000019000000000000001e00000000",
            INIT_73 => X"fffffff7ffffffff000000150000000000000010000000000000001000000000",
            INIT_74 => X"ffffff9afffffffffffffffdffffffffffffffebffffffff0000002200000000",
            INIT_75 => X"fffffff1ffffffffffffffdeffffffff00000009000000000000001a00000000",
            INIT_76 => X"0000000700000000ffffffcdffffffffffffffd2ffffffff0000000a00000000",
            INIT_77 => X"ffffffdaffffffff00000024000000000000000900000000fffffff8ffffffff",
            INIT_78 => X"0000000800000000fffffff7ffffffff0000000700000000ffffffe6ffffffff",
            INIT_79 => X"00000016000000000000002d00000000ffffffdffffffffffffffffeffffffff",
            INIT_7A => X"fffffffbffffffff00000032000000000000004a00000000ffffffffffffffff",
            INIT_7B => X"fffffff3fffffffffffffffeffffffff0000001900000000ffffffefffffffff",
            INIT_7C => X"0000002600000000ffffffe5ffffffffffffffe6ffffffff0000000600000000",
            INIT_7D => X"fffffffcfffffffffffffffbffffffff0000001700000000fffffff5ffffffff",
            INIT_7E => X"fffffffbffffffff0000000c0000000000000006000000000000000d00000000",
            INIT_7F => X"0000000800000000fffffffeffffffff0000001e00000000fffffff8ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE7;


    MEM_IWGHT_LAYER2_INSTANCE8 : if BRAM_NAME = "iwght_layer2_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000027000000000000003b0000000000000045000000000000005700000000",
            INIT_01 => X"0000001900000000fffffff7ffffffff00000019000000000000003200000000",
            INIT_02 => X"ffffffe7ffffffffffffffdaffffffffffffffe0ffffffff0000000900000000",
            INIT_03 => X"ffffffe7ffffffffffffffb8ffffffffffffffd1ffffffffffffffcfffffffff",
            INIT_04 => X"0000000800000000fffffff4ffffffffffffffcbffffffff0000000600000000",
            INIT_05 => X"ffffffecffffffffffffffd8ffffffffffffffb5ffffffffffffffc9ffffffff",
            INIT_06 => X"fffffff6fffffffffffffff0ffffffffffffffe7ffffffff0000001800000000",
            INIT_07 => X"ffffffd6ffffffffffffffbfffffffffffffffceffffffffffffffdaffffffff",
            INIT_08 => X"ffffffefffffffffffffffe4fffffffffffffffcffffffffffffffc5ffffffff",
            INIT_09 => X"fffffffbfffffffffffffff3ffffffffffffffffffffffff0000000600000000",
            INIT_0A => X"00000007000000000000000400000000ffffffecffffffff0000001600000000",
            INIT_0B => X"000000050000000000000009000000000000000000000000fffffffbffffffff",
            INIT_0C => X"ffffffedffffffff0000001d000000000000000400000000fffffff8ffffffff",
            INIT_0D => X"00000000000000000000001300000000ffffffe9ffffffffffffffdfffffffff",
            INIT_0E => X"fffffff8fffffffffffffff7fffffffffffffffbffffffff0000001300000000",
            INIT_0F => X"0000002200000000ffffffe3fffffffffffffff6fffffffffffffff2ffffffff",
            INIT_10 => X"fffffffefffffffffffffff6ffffffff00000025000000000000002e00000000",
            INIT_11 => X"fffffff2ffffffff00000024000000000000000d000000000000000b00000000",
            INIT_12 => X"00000009000000000000001f0000000000000022000000000000001300000000",
            INIT_13 => X"00000011000000000000000200000000fffffff3ffffffff0000001100000000",
            INIT_14 => X"0000000c0000000000000021000000000000001400000000ffffffe3ffffffff",
            INIT_15 => X"fffffff8ffffffff000000050000000000000023000000000000000600000000",
            INIT_16 => X"0000002d0000000000000056000000000000000200000000ffffffffffffffff",
            INIT_17 => X"fffffffcffffffff0000001b000000000000002b000000000000002e00000000",
            INIT_18 => X"ffffffcaffffffffffffffebffffffff00000018000000000000000c00000000",
            INIT_19 => X"0000000d000000000000002f0000000000000012000000000000000800000000",
            INIT_1A => X"fffffffcfffffffffffffffdfffffffffffffff5ffffffff0000000e00000000",
            INIT_1B => X"fffffffaffffffff0000000e00000000ffffffcfffffffff0000001e00000000",
            INIT_1C => X"000000040000000000000018000000000000000500000000fffffff4ffffffff",
            INIT_1D => X"0000000e00000000000000100000000000000037000000000000003400000000",
            INIT_1E => X"0000001300000000000000080000000000000007000000000000001300000000",
            INIT_1F => X"00000004000000000000000f000000000000000d000000000000001200000000",
            INIT_20 => X"0000001000000000fffffffcffffffff00000009000000000000000900000000",
            INIT_21 => X"0000001000000000000000110000000000000012000000000000000200000000",
            INIT_22 => X"000000020000000000000006000000000000000f000000000000000a00000000",
            INIT_23 => X"ffffffe8ffffffff00000013000000000000002500000000fffffffcffffffff",
            INIT_24 => X"fffffff3ffffffff0000000400000000fffffff7ffffffffffffffdfffffffff",
            INIT_25 => X"0000000100000000fffffffbffffffffffffffe9ffffffffffffffebffffffff",
            INIT_26 => X"fffffffbffffffff00000009000000000000000000000000ffffffe7ffffffff",
            INIT_27 => X"fffffffaffffffff0000000300000000fffffffbffffffffffffffd7ffffffff",
            INIT_28 => X"ffffffddffffffffffffffb9ffffffff00000007000000000000001500000000",
            INIT_29 => X"ffffffe9ffffffffffffffffffffffffffffffd5ffffffffffffffe1ffffffff",
            INIT_2A => X"fffffff2ffffffffffffffe4ffffffff0000000500000000ffffffd7ffffffff",
            INIT_2B => X"fffffffafffffffffffffffaffffffffffffffdfffffffffffffffc8ffffffff",
            INIT_2C => X"ffffffbbffffffff0000002300000000ffffffe9ffffffffffffffe5ffffffff",
            INIT_2D => X"00000013000000000000001300000000ffffffe2ffffffffffffffd8ffffffff",
            INIT_2E => X"0000000200000000000000030000000000000013000000000000001600000000",
            INIT_2F => X"00000045000000000000001f000000000000002b00000000fffffffcffffffff",
            INIT_30 => X"fffffff7fffffffffffffffbffffffff00000000000000000000000400000000",
            INIT_31 => X"0000001f00000000ffffffc0ffffffffffffffdfffffffffffffffefffffffff",
            INIT_32 => X"ffffffeaffffffff0000002a000000000000002e000000000000004800000000",
            INIT_33 => X"0000000e00000000fffffff5ffffffff00000007000000000000001000000000",
            INIT_34 => X"ffffffedffffffffffffffe9ffffffff00000003000000000000000c00000000",
            INIT_35 => X"ffffffeffffffffffffffff2ffffffffffffffe6fffffffffffffff5ffffffff",
            INIT_36 => X"ffffffdbffffffffffffffe1ffffffffffffffb3ffffffffffffffeaffffffff",
            INIT_37 => X"0000001100000000fffffffeffffffff0000000e00000000ffffffd6ffffffff",
            INIT_38 => X"ffffffe3fffffffffffffff5ffffffff0000000e00000000fffffffeffffffff",
            INIT_39 => X"fffffff1ffffffff0000001b00000000ffffffedffffffffffffffe4ffffffff",
            INIT_3A => X"ffffffcaffffffffffffffd9ffffffff0000000f00000000fffffffbffffffff",
            INIT_3B => X"0000001e00000000ffffffdeffffffffffffffbaffffffffffffffc8ffffffff",
            INIT_3C => X"00000014000000000000001500000000fffffffcffffffffffffffc5ffffffff",
            INIT_3D => X"ffffffe5ffffffffffffffceffffffffffffffe8ffffffff0000000500000000",
            INIT_3E => X"0000000c00000000ffffffedffffffffffffffb9fffffffffffffffaffffffff",
            INIT_3F => X"fffffff0ffffffffffffffccffffffffffffffddffffffffffffffd1ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff8ffffffff0000001700000000ffffffeeffffffff0000000000000000",
            INIT_41 => X"00000044000000000000002f000000000000001700000000fffffff0ffffffff",
            INIT_42 => X"0000001100000000fffffffffffffffffffffff8fffffffffffffffaffffffff",
            INIT_43 => X"ffffffcdffffffffffffffd0ffffffff0000000600000000fffffffeffffffff",
            INIT_44 => X"0000000100000000fffffff0ffffffff0000002800000000fffffff0ffffffff",
            INIT_45 => X"00000039000000000000000300000000ffffffecffffffff0000000e00000000",
            INIT_46 => X"0000001b000000000000001d0000000000000028000000000000004b00000000",
            INIT_47 => X"ffffffe6fffffffffffffffdfffffffffffffff6fffffffffffffff0ffffffff",
            INIT_48 => X"000000030000000000000003000000000000000000000000ffffffffffffffff",
            INIT_49 => X"0000000000000000fffffffeffffffff0000001500000000ffffffedffffffff",
            INIT_4A => X"0000002500000000000000190000000000000021000000000000001500000000",
            INIT_4B => X"0000001e000000000000000c00000000ffffffcdffffffff0000001d00000000",
            INIT_4C => X"fffffff7ffffffffffffffd0ffffffff00000018000000000000000400000000",
            INIT_4D => X"ffffffe1ffffffffffffffd7ffffffffffffffe7ffffffffffffffb3ffffffff",
            INIT_4E => X"0000001f00000000ffffffeffffffffffffffffafffffffffffffff9ffffffff",
            INIT_4F => X"000000000000000000000025000000000000000b000000000000000200000000",
            INIT_50 => X"0000001e00000000fffffff8ffffffff0000001a000000000000002200000000",
            INIT_51 => X"0000000000000000fffffff2ffffffff0000002200000000ffffffefffffffff",
            INIT_52 => X"0000000f000000000000000100000000fffffffbffffffff0000001b00000000",
            INIT_53 => X"ffffffe2fffffffffffffff5ffffffffffffffdbffffffff0000000000000000",
            INIT_54 => X"0000001800000000ffffffeeffffffff0000002700000000fffffff5ffffffff",
            INIT_55 => X"ffffffc4ffffffffffffffddffffffff00000031000000000000001200000000",
            INIT_56 => X"ffffff86ffffffffffffffe3ffffffffffffff95ffffffffffffffe2ffffffff",
            INIT_57 => X"000000000000000000000000000000000000001400000000ffffffeaffffffff",
            INIT_58 => X"ffffffffffffffffffffffefffffffff0000000000000000fffffff9ffffffff",
            INIT_59 => X"0000001e00000000fffffff4ffffffff00000004000000000000001d00000000",
            INIT_5A => X"0000000400000000000000270000000000000037000000000000001800000000",
            INIT_5B => X"fffffffbffffffffffffffddffffffff0000000d00000000fffffffdffffffff",
            INIT_5C => X"ffffffe6ffffffffffffffe6ffffffffffffffedffffffff0000001900000000",
            INIT_5D => X"000000380000000000000015000000000000001200000000fffffff8ffffffff",
            INIT_5E => X"0000000200000000fffffffdffffffffffffffe9ffffffff0000004300000000",
            INIT_5F => X"0000001500000000fffffffaffffffff0000001000000000fffffffcffffffff",
            INIT_60 => X"ffffffd7fffffffffffffff0fffffffffffffffaffffffff0000000a00000000",
            INIT_61 => X"ffffffbaffffffffffffffc2ffffffffffffffe5fffffffffffffff1ffffffff",
            INIT_62 => X"ffffffc0ffffffffffffffc5ffffffffffffffcaffffffffffffffb0ffffffff",
            INIT_63 => X"ffffffe2fffffffffffffff5ffffffff0000000800000000ffffffe7ffffffff",
            INIT_64 => X"fffffffcffffffff0000000e00000000ffffffd7ffffffffffffffc2ffffffff",
            INIT_65 => X"ffffffdbfffffffffffffffefffffffffffffffbffffffffffffffeeffffffff",
            INIT_66 => X"fffffff7ffffffffffffffe3ffffffff0000001800000000ffffffeeffffffff",
            INIT_67 => X"fffffff8fffffffffffffff4ffffffffffffffeaffffffff0000003900000000",
            INIT_68 => X"00000008000000000000001600000000fffffff7ffffffffffffffecffffffff",
            INIT_69 => X"0000000900000000ffffffedffffffff0000000800000000fffffffbffffffff",
            INIT_6A => X"fffffff1ffffffffffffffc0ffffffff0000000c00000000ffffffe1ffffffff",
            INIT_6B => X"ffffffe7ffffffffffffffffffffffff0000000500000000ffffffe4ffffffff",
            INIT_6C => X"fffffff8ffffffff0000000000000000ffffffe7ffffffff0000000100000000",
            INIT_6D => X"0000001d00000000fffffff6ffffffff0000002c000000000000000300000000",
            INIT_6E => X"0000000300000000ffffffeffffffffffffffff8ffffffff0000003a00000000",
            INIT_6F => X"00000017000000000000000800000000ffffffe9ffffffff0000001200000000",
            INIT_70 => X"00000017000000000000000c000000000000001000000000fffffff6ffffffff",
            INIT_71 => X"fffffff3ffffffffffffffccffffffff00000016000000000000000000000000",
            INIT_72 => X"0000001900000000fffffffeffffffff00000019000000000000002300000000",
            INIT_73 => X"0000001800000000ffffffeefffffffffffffffefffffffffffffff5ffffffff",
            INIT_74 => X"0000001f00000000ffffffe9ffffffff0000000300000000ffffffe7ffffffff",
            INIT_75 => X"ffffffeaffffffffffffffedffffffff0000001700000000ffffffecffffffff",
            INIT_76 => X"ffffffdcffffffff000000190000000000000003000000000000000800000000",
            INIT_77 => X"ffffffb0ffffffffffffffdbffffffffffffffbaffffffff0000000200000000",
            INIT_78 => X"ffffffcfffffffffffffff84fffffffffffffff3ffffffffffffff86ffffffff",
            INIT_79 => X"0000001100000000ffffffd3ffffffff0000001000000000ffffffe6ffffffff",
            INIT_7A => X"ffffffdaffffffffffffffb6ffffffff0000000700000000ffffffcaffffffff",
            INIT_7B => X"0000001200000000ffffffffffffffffffffffc9ffffffffffffffd9ffffffff",
            INIT_7C => X"ffffffedffffffff00000006000000000000001700000000ffffffecffffffff",
            INIT_7D => X"fffffffeffffffff0000000d0000000000000035000000000000000100000000",
            INIT_7E => X"ffffffe4fffffffffffffff9fffffffffffffff0fffffffffffffff8ffffffff",
            INIT_7F => X"ffffffceffffffff0000002000000000fffffffcfffffffffffffff3ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE8;


    MEM_IWGHT_LAYER2_INSTANCE9 : if BRAM_NAME = "iwght_layer2_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffdeffffffff0000000000000000ffffffdcfffffffffffffff4ffffffff",
            INIT_01 => X"00000000000000000000000000000000fffffffbffffffffffffffdaffffffff",
            INIT_02 => X"ffffffecffffffff000000160000000000000037000000000000002800000000",
            INIT_03 => X"0000002200000000fffffff9ffffffff0000001800000000fffffff6ffffffff",
            INIT_04 => X"ffffffddffffffff0000000a00000000ffffffffffffffff0000002f00000000",
            INIT_05 => X"ffffffe6ffffffff0000000900000000ffffffeffffffffffffffff0ffffffff",
            INIT_06 => X"0000000400000000ffffffeeffffffff00000011000000000000000000000000",
            INIT_07 => X"ffffffd8ffffffffffffffeeffffffff0000001000000000ffffffe0ffffffff",
            INIT_08 => X"0000000900000000ffffffd4fffffffffffffffeffffffff0000000000000000",
            INIT_09 => X"ffffffb5ffffffffffffffeaffffffffffffffaeffffffff0000001800000000",
            INIT_0A => X"ffffffdeffffffffffffffb5ffffffffffffffb5ffffffffffffffadffffffff",
            INIT_0B => X"0000001900000000fffffffffffffffffffffffbfffffffffffffff0ffffffff",
            INIT_0C => X"0000000000000000fffffffaffffffffffffffd3ffffffff0000002100000000",
            INIT_0D => X"0000000f000000000000000b000000000000000200000000ffffffe4ffffffff",
            INIT_0E => X"0000000800000000000000250000000000000003000000000000000900000000",
            INIT_0F => X"000000050000000000000025000000000000002f000000000000000900000000",
            INIT_10 => X"fffffff1ffffffff000000100000000000000004000000000000000900000000",
            INIT_11 => X"fffffff8ffffffffffffffecffffffff0000001600000000fffffff0ffffffff",
            INIT_12 => X"ffffffe1ffffffffffffffe8ffffffff00000050000000000000001500000000",
            INIT_13 => X"0000000900000000ffffffebffffffff0000000f000000000000001a00000000",
            INIT_14 => X"0000000e00000000ffffffecffffffff0000001400000000fffffffaffffffff",
            INIT_15 => X"0000000e00000000ffffffd4ffffffff00000025000000000000000c00000000",
            INIT_16 => X"fffffffaffffffff0000000400000000ffffffe4ffffffffffffffe8ffffffff",
            INIT_17 => X"0000000900000000ffffffe1ffffffff00000014000000000000001c00000000",
            INIT_18 => X"0000003f00000000fffffff5ffffffffffffffd6ffffffff0000003600000000",
            INIT_19 => X"0000000300000000000000050000000000000012000000000000000900000000",
            INIT_1A => X"fffffffdffffffff000000040000000000000017000000000000000800000000",
            INIT_1B => X"00000008000000000000002600000000ffffffdeffffffff0000001e00000000",
            INIT_1C => X"0000002d000000000000001e000000000000001d000000000000000000000000",
            INIT_1D => X"fffffff5ffffffffffffffe4ffffffff00000034000000000000001800000000",
            INIT_1E => X"0000001200000000fffffff1fffffffffffffff2ffffffff0000000800000000",
            INIT_1F => X"0000000c00000000fffffffcffffffffffffffebfffffffffffffff9ffffffff",
            INIT_20 => X"ffffffc4ffffffffffffffd2ffffffff0000001e000000000000000a00000000",
            INIT_21 => X"0000000000000000ffffffbdffffffffffffffcfffffffff0000001700000000",
            INIT_22 => X"ffffffe1ffffffff0000002a000000000000003000000000fffffff2ffffffff",
            INIT_23 => X"ffffffeaffffffffffffffffffffffff00000019000000000000000c00000000",
            INIT_24 => X"0000001600000000ffffffe6ffffffffffffffe9ffffffff0000001c00000000",
            INIT_25 => X"fffffffdffffffff0000000400000000ffffffccfffffffffffffffaffffffff",
            INIT_26 => X"0000002c00000000fffffffffffffffffffffffdffffffff0000000e00000000",
            INIT_27 => X"0000000b0000000000000003000000000000000e000000000000002800000000",
            INIT_28 => X"0000001b00000000000000090000000000000004000000000000000400000000",
            INIT_29 => X"ffffffc8fffffffffffffff8ffffffffffffffecfffffffffffffff4ffffffff",
            INIT_2A => X"ffffffbcffffffffffffff96ffffffffffffffc3ffffffffffffffe9ffffffff",
            INIT_2B => X"fffffff1ffffffffffffffd8ffffffffffffffbeffffffff0000000c00000000",
            INIT_2C => X"ffffffcdffffffffffffffe9ffffffffffffffebffffffffffffffb5ffffffff",
            INIT_2D => X"0000001000000000ffffffd7ffffffffffffffedffffffffffffffc9ffffffff",
            INIT_2E => X"fffffff9fffffffffffffffcffffffffffffffc8ffffffffffffffebffffffff",
            INIT_2F => X"ffffffffffffffff0000001800000000ffffffb7fffffffffffffffeffffffff",
            INIT_30 => X"000000000000000000000001000000000000001100000000ffffffffffffffff",
            INIT_31 => X"00000015000000000000000e000000000000000600000000fffffffbffffffff",
            INIT_32 => X"ffffffc2ffffffffffffffccffffffff0000000000000000ffffffedffffffff",
            INIT_33 => X"ffffffb7ffffffffffffffccffffffffffffffcfffffffffffffffb8ffffffff",
            INIT_34 => X"00000019000000000000000100000000ffffffedffffffff0000000000000000",
            INIT_35 => X"00000025000000000000001700000000ffffffecfffffffffffffffeffffffff",
            INIT_36 => X"fffffff5ffffffff00000019000000000000002c00000000ffffffd7ffffffff",
            INIT_37 => X"0000002200000000ffffffe9ffffffff00000011000000000000001900000000",
            INIT_38 => X"fffffffcffffffff0000000c00000000fffffffeffffffff0000000100000000",
            INIT_39 => X"ffffffcbffffffffffffffc2ffffffffffffffe2ffffffff0000002f00000000",
            INIT_3A => X"0000000400000000ffffffd7ffffffffffffffd8ffffffffffffffaeffffffff",
            INIT_3B => X"fffffffaffffffff000000050000000000000017000000000000000a00000000",
            INIT_3C => X"fffffffdffffffff00000000000000000000003300000000ffffffd9ffffffff",
            INIT_3D => X"0000001200000000ffffffebffffffff0000000a00000000fffffff6ffffffff",
            INIT_3E => X"00000039000000000000001d00000000ffffffefffffffff0000002c00000000",
            INIT_3F => X"00000025000000000000000e0000000000000015000000000000000200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffffffffffff0000000200000000fffffff7ffffffff0000000800000000",
            INIT_41 => X"ffffffc3ffffffff0000001e000000000000002100000000fffffff9ffffffff",
            INIT_42 => X"ffffffe1ffffffffffffffd4ffffffff0000002900000000ffffffceffffffff",
            INIT_43 => X"00000011000000000000000f00000000ffffffd4ffffffff0000001000000000",
            INIT_44 => X"ffffffdefffffffffffffff1ffffffff0000000a00000000ffffffffffffffff",
            INIT_45 => X"fffffff0ffffffff0000001f00000000ffffffe8ffffffffffffffefffffffff",
            INIT_46 => X"0000001a00000000ffffffceffffffff00000001000000000000003000000000",
            INIT_47 => X"00000005000000000000004800000000ffffffd5ffffffff0000000000000000",
            INIT_48 => X"fffffffaffffffff0000000500000000ffffffe6ffffffffffffffc6ffffffff",
            INIT_49 => X"0000001e00000000ffffffffffffffff0000000f00000000fffffff7ffffffff",
            INIT_4A => X"00000022000000000000000c0000000000000005000000000000001600000000",
            INIT_4B => X"0000002600000000ffffffe6ffffffffffffffd8ffffffff0000002c00000000",
            INIT_4C => X"fffffffcffffffff0000000400000000ffffffe5ffffffffffffffe6ffffffff",
            INIT_4D => X"ffffffd2fffffffffffffff7ffffffff00000018000000000000000500000000",
            INIT_4E => X"ffffffd7ffffffffffffffefffffffffffffffdffffffffffffffffaffffffff",
            INIT_4F => X"fffffffdfffffffffffffffeffffffff0000000500000000fffffff2ffffffff",
            INIT_50 => X"fffffff4ffffffffffffffebffffffff00000019000000000000000500000000",
            INIT_51 => X"00000008000000000000001300000000ffffffecffffffff0000001600000000",
            INIT_52 => X"ffffffdfffffffffffffffd0ffffffffffffffbcffffffff0000001000000000",
            INIT_53 => X"ffffffeaffffffffffffffffffffffffffffffd5ffffffffffffff9effffffff",
            INIT_54 => X"ffffffb8ffffffff0000000c000000000000000000000000ffffffeeffffffff",
            INIT_55 => X"0000000d00000000ffffffd6fffffffffffffffbffffffff0000001600000000",
            INIT_56 => X"ffffffa7fffffffffffffff8ffffffff00000025000000000000001300000000",
            INIT_57 => X"0000000d00000000ffffffb1ffffffffffffffbfffffffff0000000200000000",
            INIT_58 => X"0000000c00000000ffffffefffffffffffffffeeffffffff0000000f00000000",
            INIT_59 => X"fffffff9ffffffff0000000e000000000000000300000000ffffffdcffffffff",
            INIT_5A => X"0000000e00000000ffffffccffffffff0000000300000000fffffffcffffffff",
            INIT_5B => X"0000001800000000ffffffe4ffffffff00000003000000000000001900000000",
            INIT_5C => X"0000000c00000000000000000000000000000022000000000000000d00000000",
            INIT_5D => X"ffffffddfffffffffffffff9ffffffffffffffd0ffffffff0000000500000000",
            INIT_5E => X"0000002d0000000000000006000000000000000700000000ffffffe2ffffffff",
            INIT_5F => X"fffffff6ffffffff0000001b00000000fffffffeffffffffffffffd7ffffffff",
            INIT_60 => X"ffffffd1ffffffff0000000800000000fffffff4ffffffffffffffd4ffffffff",
            INIT_61 => X"fffffff8fffffffffffffffeffffffffffffffdfffffffff0000000600000000",
            INIT_62 => X"0000001f000000000000001500000000ffffffe5ffffffff0000000000000000",
            INIT_63 => X"0000003a00000000ffffffebffffffffffffffe2ffffffff0000000200000000",
            INIT_64 => X"ffffffa6ffffffff0000001a000000000000001400000000ffffffceffffffff",
            INIT_65 => X"00000001000000000000001600000000ffffff9affffffff0000001300000000",
            INIT_66 => X"fffffff1ffffffff0000000000000000ffffffe3ffffffff0000000d00000000",
            INIT_67 => X"0000001e00000000fffffffdffffffff0000001500000000ffffffd6ffffffff",
            INIT_68 => X"0000001a000000000000000a00000000fffffff6fffffffffffffff0ffffffff",
            INIT_69 => X"0000000b000000000000001e00000000ffffffc5fffffffffffffffaffffffff",
            INIT_6A => X"0000001900000000fffffff6ffffffffffffffa1ffffffff0000001a00000000",
            INIT_6B => X"0000001f000000000000002f00000000ffffffe7ffffffffffffffd0ffffffff",
            INIT_6C => X"ffffffe7ffffffff0000004b00000000ffffffeaffffffffffffffedffffffff",
            INIT_6D => X"ffffffbaffffffff00000019000000000000002700000000ffffffbbffffffff",
            INIT_6E => X"fffffff5ffffffff00000000000000000000003000000000fffffff3ffffffff",
            INIT_6F => X"000000030000000000000000000000000000002200000000ffffffeaffffffff",
            INIT_70 => X"0000004100000000fffffffdffffffff0000000d000000000000000e00000000",
            INIT_71 => X"000000090000000000000001000000000000002f000000000000002300000000",
            INIT_72 => X"ffffffcfffffffffffffffc2ffffffffffffffabffffffff0000000600000000",
            INIT_73 => X"fffffff3ffffffffffffffffffffffff00000016000000000000002e00000000",
            INIT_74 => X"00000024000000000000000100000000ffffffceffffffffffffffedffffffff",
            INIT_75 => X"ffffffe4ffffffff0000003e00000000ffffffdcffffffff0000004000000000",
            INIT_76 => X"ffffffe3ffffffff0000000200000000fffffffbffffffffffffffd2ffffffff",
            INIT_77 => X"ffffffeffffffffffffffff0ffffffff0000001500000000ffffffb5ffffffff",
            INIT_78 => X"fffffff3fffffffffffffff3ffffffff00000003000000000000001100000000",
            INIT_79 => X"0000002800000000000000030000000000000000000000000000000000000000",
            INIT_7A => X"ffffffecffffffffffffffecffffffff0000002e000000000000001e00000000",
            INIT_7B => X"ffffffeeffffffffffffffcfffffffffffffffc6ffffffff0000001600000000",
            INIT_7C => X"0000001f00000000ffffffebffffffff00000010000000000000000900000000",
            INIT_7D => X"000000180000000000000038000000000000000200000000fffffff9ffffffff",
            INIT_7E => X"0000001a00000000ffffffebffffffffffffffefffffffff0000002700000000",
            INIT_7F => X"fffffff1ffffffff0000001d00000000ffffffeaffffffffffffffd9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE9;


    MEM_IWGHT_LAYER2_INSTANCE10 : if BRAM_NAME = "iwght_layer2_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000ffffffe2fffffffffffffff6ffffffffffffffeaffffffff",
            INIT_01 => X"fffffff6ffffffffffffffd3ffffffffffffffc2ffffffff0000001700000000",
            INIT_02 => X"00000008000000000000001d00000000ffffffdfffffffffffffffddffffffff",
            INIT_03 => X"fffffffeffffffff00000021000000000000002100000000fffffffdffffffff",
            INIT_04 => X"fffffff2ffffffff0000003000000000fffffff9ffffffff0000000100000000",
            INIT_05 => X"ffffffdaffffffff00000011000000000000000c000000000000000c00000000",
            INIT_06 => X"00000009000000000000001a00000000fffffffffffffffffffffff8ffffffff",
            INIT_07 => X"0000001600000000ffffffedffffffff00000028000000000000001500000000",
            INIT_08 => X"fffffff8fffffffffffffff5ffffffffffffffe9ffffffff0000000100000000",
            INIT_09 => X"00000006000000000000000000000000ffffffe4fffffffffffffffcffffffff",
            INIT_0A => X"00000005000000000000003000000000ffffffd7ffffffffffffffeeffffffff",
            INIT_0B => X"0000000700000000fffffff0ffffffffffffffbcffffffffffffffd3ffffffff",
            INIT_0C => X"0000001900000000fffffffdffffffffffffffa3ffffffff0000000f00000000",
            INIT_0D => X"0000002500000000fffffffafffffffffffffff5ffffffff0000000200000000",
            INIT_0E => X"fffffff4ffffffff0000001d00000000ffffffdfffffffffffffffeeffffffff",
            INIT_0F => X"fffffff4fffffffffffffff2ffffffff0000000600000000ffffffe2ffffffff",
            INIT_10 => X"00000033000000000000000d0000000000000006000000000000000100000000",
            INIT_11 => X"ffffffceffffffff0000002c00000000ffffffe0ffffffffffffffc1ffffffff",
            INIT_12 => X"ffffffe4ffffffff0000000200000000ffffffffffffffffffffffdbffffffff",
            INIT_13 => X"000000020000000000000021000000000000001400000000fffffff6ffffffff",
            INIT_14 => X"00000012000000000000001a000000000000001600000000ffffffefffffffff",
            INIT_15 => X"0000001900000000ffffffe3fffffffffffffffafffffffffffffffaffffffff",
            INIT_16 => X"0000003400000000fffffffdfffffffffffffff9ffffffff0000001f00000000",
            INIT_17 => X"0000004d00000000fffffff0ffffffffffffffe9ffffffff0000001200000000",
            INIT_18 => X"fffffffeffffffff0000003500000000fffffff7ffffffff0000000500000000",
            INIT_19 => X"0000000a000000000000000e000000000000003900000000fffffff9ffffffff",
            INIT_1A => X"ffffffd9ffffffffffffffdfffffffffffffffdbffffffffffffffc2ffffffff",
            INIT_1B => X"0000001800000000fffffff1fffffffffffffff7ffffffffffffffdeffffffff",
            INIT_1C => X"0000000000000000fffffff1ffffffff0000002c000000000000001b00000000",
            INIT_1D => X"0000002d00000000fffffff8ffffffffffffffeeffffffff0000001f00000000",
            INIT_1E => X"fffffffdffffffff0000002000000000ffffffd4fffffffffffffff3ffffffff",
            INIT_1F => X"fffffff5ffffffffffffffe4fffffffffffffff4ffffffffffffffe1ffffffff",
            INIT_20 => X"0000000000000000ffffffedfffffffffffffffcfffffffffffffff7ffffffff",
            INIT_21 => X"fffffff4ffffffffffffffe9ffffffffffffffdfffffffff0000000300000000",
            INIT_22 => X"fffffff5ffffffff00000000000000000000000e000000000000000100000000",
            INIT_23 => X"fffffff5fffffffffffffffcffffffffffffffe7fffffffffffffff0ffffffff",
            INIT_24 => X"0000000100000000fffffff5ffffffff0000000b00000000ffffffe7ffffffff",
            INIT_25 => X"0000000700000000fffffff3ffffffff0000000900000000ffffffe9ffffffff",
            INIT_26 => X"0000000c000000000000000400000000ffffffeeffffffff0000000000000000",
            INIT_27 => X"0000000a00000000fffffff6ffffffff0000000800000000ffffffecffffffff",
            INIT_28 => X"fffffff2ffffffff0000000700000000ffffffeffffffffffffffff8ffffffff",
            INIT_29 => X"ffffffe8fffffffffffffffcffffffff0000000400000000fffffff0ffffffff",
            INIT_2A => X"fffffff8fffffffffffffffaffffffff0000000400000000fffffff6ffffffff",
            INIT_2B => X"00000000000000000000000900000000ffffffedffffffff0000000000000000",
            INIT_2C => X"ffffffe7ffffffff0000000300000000fffffff7fffffffffffffffbffffffff",
            INIT_2D => X"00000007000000000000000000000000fffffffdffffffffffffffeaffffffff",
            INIT_2E => X"ffffffdefffffffffffffffcfffffffffffffff6ffffffffffffffecffffffff",
            INIT_2F => X"fffffffbffffffffffffffedffffffffffffffe6fffffffffffffff6ffffffff",
            INIT_30 => X"fffffffbffffffff0000000500000000ffffffffffffffffffffffe4ffffffff",
            INIT_31 => X"ffffffeeffffffff0000000500000000fffffffefffffffffffffff5ffffffff",
            INIT_32 => X"ffffffe7ffffffffffffffe5ffffffff0000000700000000ffffffffffffffff",
            INIT_33 => X"fffffff0fffffffffffffffafffffffffffffff1ffffffff0000000500000000",
            INIT_34 => X"ffffffebffffffff0000000000000000ffffffe4ffffffff0000000400000000",
            INIT_35 => X"0000000500000000ffffffe8fffffffffffffffafffffffffffffffbffffffff",
            INIT_36 => X"ffffffedfffffffffffffff8fffffffffffffff8ffffffffffffffffffffffff",
            INIT_37 => X"fffffffcfffffffffffffff6ffffffff0000000000000000fffffff5ffffffff",
            INIT_38 => X"0000000f00000000ffffffe4fffffffffffffff4ffffffffffffffffffffffff",
            INIT_39 => X"000000020000000000000000000000000000000300000000fffffff6ffffffff",
            INIT_3A => X"fffffff4fffffffffffffff8fffffffffffffffdfffffffffffffff9ffffffff",
            INIT_3B => X"00000001000000000000000200000000ffffffe0fffffffffffffffbffffffff",
            INIT_3C => X"fffffff9fffffffffffffff5ffffffff00000001000000000000001300000000",
            INIT_3D => X"fffffff1ffffffff00000001000000000000001200000000ffffffdaffffffff",
            INIT_3E => X"0000000c000000000000000000000000fffffffcffffffffffffffe9ffffffff",
            INIT_3F => X"ffffffefffffffffffffffebffffffff0000000600000000ffffffe4ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffedffffffffffffffeefffffffffffffff1ffffffff0000000300000000",
            INIT_41 => X"fffffff4ffffffff0000001200000000ffffffebfffffffffffffff2ffffffff",
            INIT_42 => X"fffffff4fffffffffffffff1ffffffffffffffecffffffff0000000300000000",
            INIT_43 => X"ffffffefffffffff0000000300000000ffffffe5ffffffffffffffdfffffffff",
            INIT_44 => X"fffffff5ffffffff000000030000000000000005000000000000000300000000",
            INIT_45 => X"fffffff0ffffffff0000000000000000ffffffe2ffffffff0000000b00000000",
            INIT_46 => X"fffffff6ffffffff000000030000000000000000000000000000000700000000",
            INIT_47 => X"fffffff5fffffffffffffff6fffffffffffffff8ffffffffffffffeaffffffff",
            INIT_48 => X"fffffffeffffffff0000000d0000000000000000000000000000000300000000",
            INIT_49 => X"fffffffcffffffff0000000f00000000fffffff9fffffffffffffff4ffffffff",
            INIT_4A => X"00000015000000000000000300000000fffffff6ffffffff0000000000000000",
            INIT_4B => X"fffffff9ffffffffffffffecfffffffffffffffbffffffff0000000800000000",
            INIT_4C => X"0000000700000000fffffff0ffffffff0000000a00000000fffffff2ffffffff",
            INIT_4D => X"0000000a000000000000000600000000ffffffefffffffff0000000a00000000",
            INIT_4E => X"fffffff5fffffffffffffff1fffffffffffffff4ffffffffffffffe8ffffffff",
            INIT_4F => X"00000004000000000000000900000000ffffffefffffffffffffffe7ffffffff",
            INIT_50 => X"fffffff0ffffffffffffffe9ffffffff0000000300000000fffffff2ffffffff",
            INIT_51 => X"fffffff8ffffffff0000000e00000000fffffff2ffffffffffffffefffffffff",
            INIT_52 => X"0000000400000000fffffffdfffffffffffffff2ffffffffffffffe6ffffffff",
            INIT_53 => X"0000000900000000fffffffaffffffff0000000700000000fffffffaffffffff",
            INIT_54 => X"fffffff5ffffffff000000010000000000000003000000000000000200000000",
            INIT_55 => X"fffffff8ffffffff0000000500000000fffffff6ffffffffffffffe7ffffffff",
            INIT_56 => X"0000000300000000fffffffafffffffffffffff3ffffffffffffffe4ffffffff",
            INIT_57 => X"fffffffcffffffff0000000a0000000000000005000000000000000300000000",
            INIT_58 => X"0000000000000000ffffffe0fffffffffffffff4fffffffffffffff1ffffffff",
            INIT_59 => X"0000000300000000fffffff0ffffffff0000000200000000fffffff8ffffffff",
            INIT_5A => X"0000000500000000ffffffeeffffffffffffffeefffffffffffffff3ffffffff",
            INIT_5B => X"ffffffe9ffffffffffffffedfffffffffffffff8fffffffffffffff0ffffffff",
            INIT_5C => X"fffffffcffffffffffffffecfffffffffffffffafffffffffffffff4ffffffff",
            INIT_5D => X"fffffffcffffffff0000000400000000fffffff2ffffffff0000000900000000",
            INIT_5E => X"ffffffecfffffffffffffff9ffffffffffffffffffffffffffffffebffffffff",
            INIT_5F => X"ffffffecfffffffffffffff9ffffffff0000000000000000ffffffeaffffffff",
            INIT_60 => X"000000080000000000000009000000000000000500000000ffffffefffffffff",
            INIT_61 => X"fffffffcffffffff00000003000000000000000600000000fffffff3ffffffff",
            INIT_62 => X"ffffffe8ffffffffffffffeeffffffff0000000500000000ffffffffffffffff",
            INIT_63 => X"fffffff2fffffffffffffffeffffffff0000000000000000ffffffecffffffff",
            INIT_64 => X"fffffff6ffffffffffffffe8fffffffffffffff4fffffffffffffff4ffffffff",
            INIT_65 => X"fffffff0fffffffffffffff6fffffffffffffff4fffffffffffffff3ffffffff",
            INIT_66 => X"00000008000000000000000100000000fffffff7fffffffffffffff2ffffffff",
            INIT_67 => X"ffffffe2ffffffff0000000700000000ffffffeafffffffffffffffcffffffff",
            INIT_68 => X"0000000e0000000000000005000000000000000800000000ffffffffffffffff",
            INIT_69 => X"0000000000000000ffffffecffffffff0000000d000000000000000000000000",
            INIT_6A => X"ffffffeaffffffffffffffdfffffffffffffffc3ffffffffffffffe7ffffffff",
            INIT_6B => X"fffffff6fffffffffffffff6ffffffffffffffe5fffffffffffffff8ffffffff",
            INIT_6C => X"00000034000000000000003700000000ffffffe1ffffffffffffffc0ffffffff",
            INIT_6D => X"00000028000000000000002f0000000000000037000000000000004800000000",
            INIT_6E => X"0000000a000000000000002000000000fffffffbffffffff0000001700000000",
            INIT_6F => X"ffffffc2fffffffffffffff3ffffffff00000015000000000000000e00000000",
            INIT_70 => X"ffffffceffffffffffffffcfffffffffffffffc3ffffffffffffffddffffffff",
            INIT_71 => X"ffffffd6fffffffffffffff9fffffffffffffff9ffffffff0000000500000000",
            INIT_72 => X"ffffffb2fffffffffffffff2ffffffffffffffddffffffffffffffc2ffffffff",
            INIT_73 => X"ffffffdafffffffffffffffbffffffffffffffd6ffffffffffffffd0ffffffff",
            INIT_74 => X"ffffffdcffffffff0000002100000000ffffffecffffffffffffffe5ffffffff",
            INIT_75 => X"00000014000000000000000900000000ffffffeeffffffffffffffbfffffffff",
            INIT_76 => X"0000000d000000000000000100000000fffffffdffffffff0000000500000000",
            INIT_77 => X"ffffffdbffffffff0000000c0000000000000017000000000000001300000000",
            INIT_78 => X"0000000900000000fffffffaffffffff00000000000000000000000e00000000",
            INIT_79 => X"00000021000000000000002f0000000000000021000000000000000b00000000",
            INIT_7A => X"00000009000000000000000e00000000ffffffe1fffffffffffffffcffffffff",
            INIT_7B => X"0000000b000000000000000600000000fffffffffffffffffffffff9ffffffff",
            INIT_7C => X"000000150000000000000023000000000000002b00000000fffffff8ffffffff",
            INIT_7D => X"ffffffe5fffffffffffffffdffffffff00000005000000000000002300000000",
            INIT_7E => X"0000000a0000000000000000000000000000001100000000ffffffecffffffff",
            INIT_7F => X"00000007000000000000000900000000ffffffeeffffffff0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE10;


    MEM_IWGHT_LAYER2_INSTANCE11 : if BRAM_NAME = "iwght_layer2_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000200000000ffffffdbffffffff00000006000000000000002000000000",
            INIT_01 => X"0000000b00000000000000300000000000000025000000000000001d00000000",
            INIT_02 => X"0000000e0000000000000024000000000000003b000000000000000100000000",
            INIT_03 => X"00000021000000000000002f0000000000000041000000000000005500000000",
            INIT_04 => X"0000000700000000000000100000000000000012000000000000001e00000000",
            INIT_05 => X"ffffffeeffffffffffffffe4fffffffffffffff4ffffffff0000000200000000",
            INIT_06 => X"ffffffe4ffffffffffffffdaffffffff00000010000000000000000300000000",
            INIT_07 => X"0000000d00000000fffffffbffffffffffffffe8fffffffffffffff5ffffffff",
            INIT_08 => X"0000000f000000000000000d000000000000000000000000ffffffffffffffff",
            INIT_09 => X"fffffffaffffffffffffffefffffffff0000000700000000fffffffaffffffff",
            INIT_0A => X"00000009000000000000002e00000000ffffffd5ffffffff0000000b00000000",
            INIT_0B => X"000000200000000000000012000000000000003a000000000000000900000000",
            INIT_0C => X"ffffffd5ffffffff0000000300000000ffffffecffffffff0000000800000000",
            INIT_0D => X"ffffffe0fffffffffffffffdffffffffffffffd5ffffffffffffffebffffffff",
            INIT_0E => X"fffffff4ffffffff0000000a00000000ffffffd9ffffffffffffffe5ffffffff",
            INIT_0F => X"0000000000000000000000290000000000000015000000000000002600000000",
            INIT_10 => X"0000001f00000000fffffff9ffffffff0000000500000000fffffffaffffffff",
            INIT_11 => X"ffffffe3ffffffff0000000800000000ffffffe0ffffffff0000001e00000000",
            INIT_12 => X"fffffffbffffffff0000001a00000000ffffffe4fffffffffffffff5ffffffff",
            INIT_13 => X"fffffff0ffffffff0000000c00000000ffffffd0ffffffffffffffdfffffffff",
            INIT_14 => X"fffffff7ffffffff0000001600000000ffffffc4ffffffffffffffb4ffffffff",
            INIT_15 => X"0000001200000000ffffffe5ffffffffffffffdafffffffffffffffcffffffff",
            INIT_16 => X"ffffffe5ffffffff0000000700000000fffffff1ffffffffffffffe9ffffffff",
            INIT_17 => X"00000005000000000000001900000000fffffffdfffffffffffffff3ffffffff",
            INIT_18 => X"00000017000000000000000600000000ffffffe5fffffffffffffffaffffffff",
            INIT_19 => X"0000002900000000fffffffcffffffff00000027000000000000000e00000000",
            INIT_1A => X"0000002d0000000000000018000000000000001a000000000000005100000000",
            INIT_1B => X"ffffffe3ffffffff0000002d000000000000002c000000000000001b00000000",
            INIT_1C => X"ffffffd7ffffffffffffffdcffffffff00000007000000000000000100000000",
            INIT_1D => X"ffffffc4ffffffff0000000600000000ffffffdeffffffffffffffcaffffffff",
            INIT_1E => X"0000003b00000000ffffffc2ffffffffffffffdcffffffffffffffe5ffffffff",
            INIT_1F => X"00000016000000000000002c0000000000000004000000000000000000000000",
            INIT_20 => X"00000016000000000000000f00000000ffffffefffffffff0000002a00000000",
            INIT_21 => X"ffffffffffffffff000000280000000000000021000000000000001a00000000",
            INIT_22 => X"fffffff2ffffffff000000000000000000000015000000000000000e00000000",
            INIT_23 => X"0000000e000000000000000d00000000ffffffcfffffffff0000000100000000",
            INIT_24 => X"fffffff1ffffffff0000000600000000ffffffffffffffff0000000e00000000",
            INIT_25 => X"fffffff0ffffffff000000020000000000000023000000000000000700000000",
            INIT_26 => X"ffffffd0ffffffffffffffccffffffffffffffe0ffffffffffffffd9ffffffff",
            INIT_27 => X"fffffff5fffffffffffffffcffffffffffffffe9ffffffffffffffffffffffff",
            INIT_28 => X"ffffffecffffffff0000000200000000fffffffcffffffffffffffe4ffffffff",
            INIT_29 => X"000000510000000000000044000000000000001e00000000ffffffeeffffffff",
            INIT_2A => X"00000016000000000000000900000000fffffffdffffffff0000005d00000000",
            INIT_2B => X"ffffffd6ffffffff000000200000000000000021000000000000001b00000000",
            INIT_2C => X"ffffffedfffffffffffffffaffffffff0000002100000000ffffffc0ffffffff",
            INIT_2D => X"0000000000000000ffffffe2ffffffff00000008000000000000001200000000",
            INIT_2E => X"0000001400000000fffffffbffffffffffffffdaffffffffffffffdcffffffff",
            INIT_2F => X"fffffffaffffffff0000000f00000000fffffff2fffffffffffffff5ffffffff",
            INIT_30 => X"ffffffe3ffffffffffffffddffffffffffffffefffffffffffffffb7ffffffff",
            INIT_31 => X"ffffffe4fffffffffffffff4ffffffffffffffcdffffffff0000000000000000",
            INIT_32 => X"fffffffafffffffffffffff1ffffffff0000001a000000000000000800000000",
            INIT_33 => X"0000004800000000fffffffeffffffff0000000a000000000000000000000000",
            INIT_34 => X"0000001900000000ffffffb5ffffffff0000002d000000000000003600000000",
            INIT_35 => X"0000000400000000fffffff1ffffffffffffffcfffffffff0000003600000000",
            INIT_36 => X"000000230000000000000020000000000000003b000000000000003700000000",
            INIT_37 => X"00000004000000000000001800000000ffffffdaffffffff0000002f00000000",
            INIT_38 => X"0000000a00000000000000140000000000000003000000000000000400000000",
            INIT_39 => X"0000002500000000000000110000000000000033000000000000002500000000",
            INIT_3A => X"0000000c00000000ffffffddffffffff0000001c000000000000000200000000",
            INIT_3B => X"fffffffcfffffffffffffffcffffffff00000029000000000000000f00000000",
            INIT_3C => X"000000250000000000000003000000000000000e000000000000001d00000000",
            INIT_3D => X"0000000500000000ffffffeeffffffffffffffe9ffffffff0000000400000000",
            INIT_3E => X"0000001800000000000000040000000000000002000000000000003000000000",
            INIT_3F => X"fffffff2ffffffffffffffe2ffffffff0000001b000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000017000000000000000c00000000fffffffbfffffffffffffff9ffffffff",
            INIT_41 => X"ffffffd5ffffffffffffffefffffffffffffffdfffffffffffffffe8ffffffff",
            INIT_42 => X"ffffffeaffffffff0000000b00000000fffffff2ffffffffffffffd1ffffffff",
            INIT_43 => X"fffffffaffffffffffffffeafffffffffffffff1ffffffffffffffe4ffffffff",
            INIT_44 => X"0000001b000000000000000b0000000000000016000000000000001100000000",
            INIT_45 => X"00000005000000000000003300000000fffffffbfffffffffffffff9ffffffff",
            INIT_46 => X"ffffffd9ffffffffffffffefffffffff0000000500000000fffffffcffffffff",
            INIT_47 => X"0000001400000000fffffffaffffffff0000000d00000000ffffffbfffffffff",
            INIT_48 => X"00000029000000000000000c00000000fffffff7ffffffffffffffd8ffffffff",
            INIT_49 => X"ffffffd3ffffffff0000000700000000ffffffeaffffffff0000001200000000",
            INIT_4A => X"ffffffe0ffffffff0000003f000000000000001800000000ffffffdcffffffff",
            INIT_4B => X"00000021000000000000003f000000000000000600000000fffffff5ffffffff",
            INIT_4C => X"0000002c0000000000000039000000000000001d000000000000002300000000",
            INIT_4D => X"fffffffaffffffff00000012000000000000001a000000000000001600000000",
            INIT_4E => X"ffffffe0fffffffffffffff2ffffffff0000000c00000000ffffffefffffffff",
            INIT_4F => X"fffffff4fffffffffffffff2ffffffffffffffe6ffffffffffffffb2ffffffff",
            INIT_50 => X"00000008000000000000000a000000000000001100000000ffffffeeffffffff",
            INIT_51 => X"ffffffe4ffffffff00000012000000000000001200000000fffffff5ffffffff",
            INIT_52 => X"000000080000000000000000000000000000001d00000000fffffff7ffffffff",
            INIT_53 => X"ffffffe0ffffffff0000000b0000000000000032000000000000000a00000000",
            INIT_54 => X"fffffff9ffffffff0000001300000000ffffffffffffffff0000000e00000000",
            INIT_55 => X"ffffffccffffffffffffffe8ffffffff0000000100000000fffffffbffffffff",
            INIT_56 => X"fffffffcffffffff00000005000000000000000000000000fffffff8ffffffff",
            INIT_57 => X"ffffffd9ffffffffffffffdbffffffffffffffe8ffffffffffffffe8ffffffff",
            INIT_58 => X"0000000000000000ffffffd8ffffffffffffffb8ffffffffffffffc1ffffffff",
            INIT_59 => X"0000001100000000ffffffe4ffffffffffffffe2ffffffff0000000b00000000",
            INIT_5A => X"0000001200000000fffffff3fffffffffffffff0ffffffff0000001900000000",
            INIT_5B => X"000000150000000000000009000000000000000a000000000000000900000000",
            INIT_5C => X"fffffff8ffffffff0000000800000000fffffff7ffffffff0000000600000000",
            INIT_5D => X"0000000f00000000000000240000000000000035000000000000002f00000000",
            INIT_5E => X"ffffffc5ffffffff000000120000000000000017000000000000000e00000000",
            INIT_5F => X"0000000900000000ffffffffffffffffffffffdeffffffffffffffc4ffffffff",
            INIT_60 => X"00000027000000000000000a00000000ffffffe6ffffffff0000000800000000",
            INIT_61 => X"0000000300000000ffffffe8fffffffffffffffdffffffff0000001900000000",
            INIT_62 => X"fffffff3ffffffff000000110000000000000022000000000000000700000000",
            INIT_63 => X"ffffff9fffffffff0000000f0000000000000058000000000000003200000000",
            INIT_64 => X"fffffff4ffffffffffffffb4ffffffffffffffe6ffffffffffffffd1ffffffff",
            INIT_65 => X"0000000c00000000fffffff0fffffffffffffff6ffffffffffffffe8ffffffff",
            INIT_66 => X"0000000d000000000000002d000000000000002c000000000000001a00000000",
            INIT_67 => X"ffffffe1ffffffff000000030000000000000016000000000000000000000000",
            INIT_68 => X"00000008000000000000000c00000000fffffff7ffffffffffffffddffffffff",
            INIT_69 => X"0000001200000000ffffffeaffffffffffffffeeffffffff0000000300000000",
            INIT_6A => X"ffffffc2fffffffffffffff9ffffffffffffffeafffffffffffffffeffffffff",
            INIT_6B => X"ffffffe3ffffffffffffffefffffffffffffffd0fffffffffffffff3ffffffff",
            INIT_6C => X"fffffff7ffffffffffffffdcffffffffffffffd2ffffffff0000000400000000",
            INIT_6D => X"fffffff7fffffffffffffff6ffffffff00000011000000000000000f00000000",
            INIT_6E => X"0000000a00000000fffffff8ffffffffffffffebffffffff0000001700000000",
            INIT_6F => X"0000000600000000000000290000000000000028000000000000001a00000000",
            INIT_70 => X"0000000000000000ffffffe8ffffffff00000014000000000000000b00000000",
            INIT_71 => X"fffffffeffffffff0000001f00000000ffffffc9ffffffffffffffddffffffff",
            INIT_72 => X"00000006000000000000001400000000ffffffd5ffffffffffffffabffffffff",
            INIT_73 => X"000000230000000000000004000000000000001f000000000000000a00000000",
            INIT_74 => X"0000000200000000fffffff2ffffffffffffffeaffffffff0000001600000000",
            INIT_75 => X"ffffffe7ffffffffffffffd2ffffffffffffffddffffffffffffffedffffffff",
            INIT_76 => X"ffffffefffffffffffffffa0ffffffffffffffd1ffffffffffffffddffffffff",
            INIT_77 => X"fffffff0ffffffffffffffe2ffffffffffffffe5ffffffffffffffeaffffffff",
            INIT_78 => X"00000003000000000000001e00000000fffffff2ffffffffffffffedffffffff",
            INIT_79 => X"fffffff7ffffffff0000001000000000fffffffafffffffffffffff0ffffffff",
            INIT_7A => X"ffffffecffffffff0000000d00000000ffffffdafffffffffffffffeffffffff",
            INIT_7B => X"ffffffc4fffffffffffffffefffffffffffffff1ffffffffffffffd5ffffffff",
            INIT_7C => X"ffffffc9ffffffffffffffd6ffffffffffffffd6ffffffffffffffcbffffffff",
            INIT_7D => X"0000000d0000000000000012000000000000000000000000ffffffc4ffffffff",
            INIT_7E => X"fffffff3ffffffff00000024000000000000003c000000000000001e00000000",
            INIT_7F => X"0000002b000000000000001700000000fffffff6ffffffff0000001c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE11;


    MEM_IWGHT_LAYER2_INSTANCE12 : if BRAM_NAME = "iwght_layer2_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000a0000000000000011000000000000002a000000000000000e00000000",
            INIT_01 => X"0000000e00000000fffffffaffffffff00000009000000000000000900000000",
            INIT_02 => X"000000140000000000000004000000000000000d00000000fffffff4ffffffff",
            INIT_03 => X"0000000e0000000000000026000000000000003e000000000000001500000000",
            INIT_04 => X"fffffffafffffffffffffff7fffffffffffffffdffffffff0000000100000000",
            INIT_05 => X"fffffffbfffffffffffffff6fffffffffffffff5ffffffffffffffb4ffffffff",
            INIT_06 => X"00000000000000000000002300000000fffffff1ffffffff0000000d00000000",
            INIT_07 => X"ffffffd9ffffffffffffffe4ffffffffffffff84ffffffffffffffdaffffffff",
            INIT_08 => X"fffffff9ffffffffffffffebffffffff00000031000000000000000700000000",
            INIT_09 => X"ffffffd1fffffffffffffff9ffffffffffffffcfffffffffffffffefffffffff",
            INIT_0A => X"fffffff2ffffffffffffffe9ffffffffffffffd6ffffffffffffffc7ffffffff",
            INIT_0B => X"00000028000000000000003800000000fffffffcffffffffffffffe7ffffffff",
            INIT_0C => X"ffffffe7ffffffff00000002000000000000001c000000000000000d00000000",
            INIT_0D => X"0000000100000000ffffffffffffffff00000009000000000000000b00000000",
            INIT_0E => X"fffffffdfffffffffffffffeffffffff0000000800000000fffffffeffffffff",
            INIT_0F => X"fffffffefffffffffffffffbffffffff00000033000000000000001500000000",
            INIT_10 => X"0000000f00000000000000160000000000000022000000000000002500000000",
            INIT_11 => X"ffffffe1ffffffff0000000900000000ffffffeaffffffffffffffdbffffffff",
            INIT_12 => X"ffffffd2ffffffffffffffe8ffffffff0000000600000000fffffffeffffffff",
            INIT_13 => X"0000002c00000000ffffffa7ffffffffffffffe1ffffffffffffffb7ffffffff",
            INIT_14 => X"fffffff8ffffffffffffffefffffffff0000001d000000000000002f00000000",
            INIT_15 => X"00000004000000000000000d000000000000001f000000000000000800000000",
            INIT_16 => X"0000001700000000000000000000000000000000000000000000001900000000",
            INIT_17 => X"ffffffeafffffffffffffffaffffffff0000000200000000ffffffffffffffff",
            INIT_18 => X"fffffffdffffffff0000000b000000000000000800000000fffffffeffffffff",
            INIT_19 => X"fffffff8ffffffff0000000000000000fffffff8fffffffffffffff6ffffffff",
            INIT_1A => X"0000002000000000ffffffe2ffffffff00000009000000000000000b00000000",
            INIT_1B => X"ffffffc6ffffffffffffffd8ffffffffffffffe1fffffffffffffff1ffffffff",
            INIT_1C => X"fffffff4ffffffff0000000b00000000fffffffeffffffff0000000f00000000",
            INIT_1D => X"0000003d000000000000002d00000000fffffff7fffffffffffffff5ffffffff",
            INIT_1E => X"ffffffe6fffffffffffffff3fffffffffffffff5ffffffff0000003200000000",
            INIT_1F => X"0000005000000000fffffff2ffffffffffffffc3ffffffffffffffddffffffff",
            INIT_20 => X"ffffffe1ffffffffffffffe5ffffffff00000037000000000000003400000000",
            INIT_21 => X"0000001c00000000000000050000000000000015000000000000000000000000",
            INIT_22 => X"0000000b000000000000000b0000000000000024000000000000001d00000000",
            INIT_23 => X"0000000500000000fffffff2fffffffffffffffffffffffffffffff7ffffffff",
            INIT_24 => X"fffffffaffffffff0000000e00000000fffffffbffffffffffffffd5ffffffff",
            INIT_25 => X"fffffff4ffffffff0000001400000000fffffffbfffffffffffffff2ffffffff",
            INIT_26 => X"0000001f000000000000000100000000ffffffecffffffffffffffe9ffffffff",
            INIT_27 => X"0000000e00000000ffffffefffffffffffffffe0ffffffff0000000b00000000",
            INIT_28 => X"fffffff1ffffffffffffffeaffffffffffffffeeffffffffffffffbdffffffff",
            INIT_29 => X"00000008000000000000000000000000ffffffe7ffffffffffffffffffffffff",
            INIT_2A => X"00000013000000000000001d00000000fffffffeffffffff0000001600000000",
            INIT_2B => X"ffffffe9ffffffffffffffcfffffffff0000000200000000ffffffccffffffff",
            INIT_2C => X"fffffff3fffffffffffffff8ffffffffffffffcbffffffffffffffbdffffffff",
            INIT_2D => X"0000001600000000000000180000000000000017000000000000000e00000000",
            INIT_2E => X"ffffffd2ffffffff0000001300000000fffffffdffffffff0000000e00000000",
            INIT_2F => X"ffffffe6ffffffffffffffe1ffffffffffffffffffffffffffffffecffffffff",
            INIT_30 => X"0000002c00000000fffffffdffffffff0000001100000000ffffffedffffffff",
            INIT_31 => X"ffffffd6ffffffffffffffe6ffffffffffffffd4ffffffffffffffcdffffffff",
            INIT_32 => X"0000002d00000000fffffffaffffffffffffffd7fffffffffffffff3ffffffff",
            INIT_33 => X"ffffffefffffffff00000020000000000000000e000000000000004600000000",
            INIT_34 => X"ffffffecffffffffffffffe0ffffffffffffffedffffffffffffffc8ffffffff",
            INIT_35 => X"ffffffeafffffffffffffff8ffffffff0000000900000000ffffffe4ffffffff",
            INIT_36 => X"ffffffeefffffffffffffff4fffffffffffffff4ffffffffffffffd4ffffffff",
            INIT_37 => X"00000033000000000000000300000000fffffffeffffffff0000001700000000",
            INIT_38 => X"00000020000000000000003b0000000000000028000000000000003000000000",
            INIT_39 => X"ffffffb4fffffffffffffff9fffffffffffffffdffffffff0000004000000000",
            INIT_3A => X"0000003d000000000000000c000000000000001900000000fffffff3ffffffff",
            INIT_3B => X"ffffffebffffffff000000010000000000000022000000000000003800000000",
            INIT_3C => X"ffffffe3ffffffffffffffedfffffffffffffff1ffffffff0000001300000000",
            INIT_3D => X"0000000d000000000000000a00000000fffffffcffffffff0000000200000000",
            INIT_3E => X"fffffffaffffffffffffffe8ffffffff00000008000000000000001900000000",
            INIT_3F => X"fffffffbffffffff000000370000000000000002000000000000000600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe0ffffffffffffffe4ffffffff00000006000000000000000100000000",
            INIT_41 => X"0000003400000000fffffff2ffffffff00000004000000000000002400000000",
            INIT_42 => X"fffffff3ffffffff00000032000000000000000f000000000000001200000000",
            INIT_43 => X"0000001000000000fffffff3ffffffffffffffbffffffffffffffff5ffffffff",
            INIT_44 => X"ffffffeafffffffffffffffcffffffffffffff90ffffffffffffffc2ffffffff",
            INIT_45 => X"ffffffcfffffffffffffffe5ffffffff0000003a00000000ffffffd2ffffffff",
            INIT_46 => X"fffffff0ffffffffffffffe7ffffffff0000001c000000000000005300000000",
            INIT_47 => X"0000000600000000ffffffd0ffffffff0000000700000000fffffffeffffffff",
            INIT_48 => X"0000000c000000000000000400000000ffffffffffffffff0000000200000000",
            INIT_49 => X"00000008000000000000000e0000000000000001000000000000000100000000",
            INIT_4A => X"00000001000000000000001d00000000fffffffcffffffffffffffffffffffff",
            INIT_4B => X"0000000b00000000ffffffe5fffffffffffffff5ffffffffffffffd4ffffffff",
            INIT_4C => X"00000028000000000000000300000000fffffff4ffffffff0000001800000000",
            INIT_4D => X"ffffffd8fffffffffffffff8ffffffff0000000f000000000000000800000000",
            INIT_4E => X"fffffff6fffffffffffffffbffffffff0000003a00000000fffffff6ffffffff",
            INIT_4F => X"ffffffe2ffffffffffffffc5ffffffff0000002a000000000000004d00000000",
            INIT_50 => X"00000024000000000000001100000000fffffffbffffffffffffffeaffffffff",
            INIT_51 => X"0000000900000000000000230000000000000000000000000000000900000000",
            INIT_52 => X"0000001000000000ffffffedffffffff00000015000000000000000000000000",
            INIT_53 => X"00000013000000000000001b00000000fffffff0ffffffff0000000900000000",
            INIT_54 => X"00000007000000000000000c000000000000002600000000ffffffffffffffff",
            INIT_55 => X"fffffff9fffffffffffffffbffffffff0000001b000000000000000900000000",
            INIT_56 => X"ffffffe3ffffffffffffffd5ffffffff0000001600000000ffffffdcffffffff",
            INIT_57 => X"0000002100000000fffffff8ffffffffffffffe0ffffffff0000000500000000",
            INIT_58 => X"ffffffefffffffff00000009000000000000001200000000ffffffedffffffff",
            INIT_59 => X"ffffffd7ffffffff0000001c00000000ffffffafffffffffffffffc4ffffffff",
            INIT_5A => X"ffffff96ffffffffffffffdbffffffff0000002e00000000ffffff91ffffffff",
            INIT_5B => X"0000000000000000ffffffd3ffffffffffffffedffffffffffffffe7ffffffff",
            INIT_5C => X"ffffffcbffffffff0000001400000000ffffffecffffffffffffffdfffffffff",
            INIT_5D => X"0000000400000000fffffffeffffffff0000000e00000000ffffffb6ffffffff",
            INIT_5E => X"ffffff9cffffffff0000001000000000ffffffe6ffffffffffffffceffffffff",
            INIT_5F => X"fffffff4fffffffffffffff5ffffffff0000000100000000ffffffdfffffffff",
            INIT_60 => X"0000001000000000000000090000000000000010000000000000001200000000",
            INIT_61 => X"fffffff4fffffffffffffffffffffffffffffffbffffffffffffffeeffffffff",
            INIT_62 => X"fffffff0fffffffffffffff7ffffffffffffffcaffffffffffffffc7ffffffff",
            INIT_63 => X"ffffffdcfffffffffffffff2ffffffff0000003100000000fffffff5ffffffff",
            INIT_64 => X"fffffff0ffffffff0000001f000000000000001000000000ffffffffffffffff",
            INIT_65 => X"ffffffd5ffffffff0000001e000000000000001600000000ffffffecffffffff",
            INIT_66 => X"0000000500000000fffffff8ffffffff0000000000000000fffffff8ffffffff",
            INIT_67 => X"ffffffd8ffffffff0000000a000000000000001300000000fffffffaffffffff",
            INIT_68 => X"ffffffcdffffffffffffffd1ffffffff00000011000000000000000600000000",
            INIT_69 => X"ffffffdcffffffffffffffc9ffffffffffffffe3ffffffffffffffd6ffffffff",
            INIT_6A => X"0000000900000000ffffffd7ffffffffffffffebffffffffffffffe8ffffffff",
            INIT_6B => X"0000000700000000ffffffe4ffffffff0000004e00000000fffffff3ffffffff",
            INIT_6C => X"00000025000000000000003b00000000fffffffeffffffff0000002600000000",
            INIT_6D => X"0000003100000000000000220000000000000014000000000000001200000000",
            INIT_6E => X"00000010000000000000004500000000ffffffffffffffffffffffefffffffff",
            INIT_6F => X"ffffffa0ffffffffffffffb5fffffffffffffff0ffffffff0000001700000000",
            INIT_70 => X"0000004200000000ffffffabffffffffffffffd1ffffffff0000003900000000",
            INIT_71 => X"ffffffdfffffffffffffffc0ffffffffffffffd0fffffffffffffffdffffffff",
            INIT_72 => X"ffffffffffffffffffffffe7ffffffff0000005a00000000ffffffd5ffffffff",
            INIT_73 => X"0000000900000000fffffffaffffffffffffffdfffffffff0000002a00000000",
            INIT_74 => X"fffffffdfffffffffffffffbffffffff0000000e000000000000001c00000000",
            INIT_75 => X"00000017000000000000000a00000000fffffff3ffffffff0000002800000000",
            INIT_76 => X"ffffffddffffffff0000001b00000000fffffff0ffffffffffffffdaffffffff",
            INIT_77 => X"00000006000000000000001400000000fffffffbffffffffffffffe9ffffffff",
            INIT_78 => X"0000001200000000ffffffefffffffff00000012000000000000002f00000000",
            INIT_79 => X"0000002b00000000000000250000000000000003000000000000000800000000",
            INIT_7A => X"0000000100000000000000110000000000000029000000000000002b00000000",
            INIT_7B => X"fffffff5ffffffff00000030000000000000000f00000000ffffffe0ffffffff",
            INIT_7C => X"0000000d0000000000000013000000000000002600000000fffffffaffffffff",
            INIT_7D => X"0000001a00000000000000060000000000000004000000000000000e00000000",
            INIT_7E => X"00000021000000000000002200000000ffffffd4ffffffff0000001600000000",
            INIT_7F => X"fffffff9ffffffff000000270000000000000004000000000000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE12;


    MEM_IWGHT_LAYER2_INSTANCE13 : if BRAM_NAME = "iwght_layer2_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e0000000000000036000000000000001900000000ffffffefffffffff",
            INIT_01 => X"ffffffd7ffffffffffffffc3ffffffffffffffe3ffffffff0000000b00000000",
            INIT_02 => X"0000000f00000000ffffffd1ffffffffffffffbaffffffff0000000900000000",
            INIT_03 => X"00000019000000000000001c00000000ffffffe2fffffffffffffffeffffffff",
            INIT_04 => X"0000002100000000ffffffd0ffffffffffffffd6ffffffff0000001a00000000",
            INIT_05 => X"0000000d00000000fffffff7ffffffffffffffe4ffffffffffffffe5ffffffff",
            INIT_06 => X"0000000700000000ffffffdaffffffffffffffd9ffffffffffffffebffffffff",
            INIT_07 => X"0000001000000000ffffffdbffffffffffffffc9fffffffffffffffaffffffff",
            INIT_08 => X"fffffff5ffffffff0000000100000000ffffffe8ffffffffffffffdcffffffff",
            INIT_09 => X"ffffffdffffffffffffffff2fffffffffffffffcffffffff0000000600000000",
            INIT_0A => X"000000040000000000000014000000000000000e000000000000000800000000",
            INIT_0B => X"0000000400000000fffffff0ffffffff00000004000000000000000b00000000",
            INIT_0C => X"0000001400000000fffffffcffffffff00000009000000000000002800000000",
            INIT_0D => X"0000000e00000000ffffffedffffffffffffffd7fffffffffffffff7ffffffff",
            INIT_0E => X"ffffffe6fffffffffffffff5ffffffffffffffedffffffffffffffefffffffff",
            INIT_0F => X"fffffff1fffffffffffffff2fffffffffffffffdffffffff0000000000000000",
            INIT_10 => X"0000000000000000ffffffe7ffffffffffffffe1ffffffffffffffdcffffffff",
            INIT_11 => X"00000000000000000000000800000000fffffffcfffffffffffffffdffffffff",
            INIT_12 => X"ffffffdcffffffffffffffd5ffffffffffffffd3ffffffffffffffe1ffffffff",
            INIT_13 => X"0000001b00000000ffffffe7ffffffffffffffe9ffffffff0000000700000000",
            INIT_14 => X"ffffffd9fffffffffffffff2ffffffff00000010000000000000000600000000",
            INIT_15 => X"ffffffe2ffffffffffffffe7ffffffff0000000b00000000fffffffeffffffff",
            INIT_16 => X"0000000300000000fffffff4ffffffffffffffeeffffffff0000001400000000",
            INIT_17 => X"ffffffe6ffffffff0000000d00000000fffffffbffffffffffffffecffffffff",
            INIT_18 => X"ffffffebfffffffffffffffffffffffffffffff6fffffffffffffff0ffffffff",
            INIT_19 => X"ffffffe0ffffffffffffffeaffffffffffffffe6ffffffffffffffe9ffffffff",
            INIT_1A => X"fffffff2fffffffffffffff7fffffffffffffffaffffffff0000000b00000000",
            INIT_1B => X"ffffffe0ffffffff0000000800000000fffffffefffffffffffffffcffffffff",
            INIT_1C => X"fffffff2ffffffffffffffe3ffffffffffffffe7ffffffffffffffe2ffffffff",
            INIT_1D => X"fffffffdffffffffffffffe9ffffffffffffffd9fffffffffffffffeffffffff",
            INIT_1E => X"ffffffddffffffffffffffdfffffffff0000000500000000ffffffefffffffff",
            INIT_1F => X"ffffffe2ffffffffffffffe5ffffffffffffffd9ffffffffffffffe7ffffffff",
            INIT_20 => X"00000020000000000000000e00000000ffffffeeffffffffffffffeaffffffff",
            INIT_21 => X"ffffffdcffffffff0000000900000000fffffff2ffffffffffffffe5ffffffff",
            INIT_22 => X"00000002000000000000002100000000fffffff4ffffffffffffffe8ffffffff",
            INIT_23 => X"ffffffeffffffffffffffff3ffffffffffffffe6ffffffff0000000800000000",
            INIT_24 => X"fffffffaffffffff00000002000000000000000600000000fffffff1ffffffff",
            INIT_25 => X"fffffffafffffffffffffffeffffffffffffffdfffffffffffffffe6ffffffff",
            INIT_26 => X"ffffffe0ffffffffffffffecfffffffffffffffeffffffff0000000b00000000",
            INIT_27 => X"00000004000000000000000c00000000ffffffefffffffffffffffddffffffff",
            INIT_28 => X"fffffff2ffffffff0000000e000000000000000900000000fffffff5ffffffff",
            INIT_29 => X"0000000100000000fffffffcffffffff00000010000000000000000700000000",
            INIT_2A => X"ffffffedffffffffffffffe8ffffffff0000000b00000000ffffffdbffffffff",
            INIT_2B => X"00000010000000000000000200000000ffffffe3ffffffff0000000800000000",
            INIT_2C => X"fffffff7ffffffffffffffe5ffffffffffffffe8ffffffffffffffffffffffff",
            INIT_2D => X"ffffffe9fffffffffffffff0ffffffffffffffe5ffffffffffffffd9ffffffff",
            INIT_2E => X"0000001d00000000ffffffefffffffff0000000200000000fffffffbffffffff",
            INIT_2F => X"ffffffe5ffffffffffffffe6fffffffffffffff1fffffffffffffff1ffffffff",
            INIT_30 => X"fffffff4ffffffff00000017000000000000000d00000000fffffffaffffffff",
            INIT_31 => X"00000003000000000000000c000000000000001000000000fffffff8ffffffff",
            INIT_32 => X"fffffffaffffffff00000020000000000000001000000000fffffff3ffffffff",
            INIT_33 => X"000000270000000000000014000000000000001e000000000000001500000000",
            INIT_34 => X"0000000e0000000000000015000000000000000e000000000000000200000000",
            INIT_35 => X"ffffffe2ffffffff0000000300000000ffffffe3ffffffffffffffe9ffffffff",
            INIT_36 => X"fffffff7ffffffff0000000000000000fffffff5ffffffffffffffdeffffffff",
            INIT_37 => X"fffffff3ffffffffffffffddffffffff0000000800000000fffffff8ffffffff",
            INIT_38 => X"ffffffe8ffffffff0000000500000000ffffffe2fffffffffffffffdffffffff",
            INIT_39 => X"fffffff3ffffffff00000029000000000000000c00000000ffffffe8ffffffff",
            INIT_3A => X"00000003000000000000000b000000000000000000000000fffffff2ffffffff",
            INIT_3B => X"fffffffaffffffff0000000d0000000000000002000000000000000a00000000",
            INIT_3C => X"0000001600000000ffffffedffffffffffffffe9ffffffff0000001400000000",
            INIT_3D => X"fffffff0ffffffff000000040000000000000002000000000000001700000000",
            INIT_3E => X"00000000000000000000000300000000ffffffe9ffffffff0000000a00000000",
            INIT_3F => X"fffffffdffffffff0000000a000000000000000300000000ffffffedffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000800000000fffffffeffffffffffffffeefffffffffffffff6ffffffff",
            INIT_41 => X"fffffffbffffffffffffffe8fffffffffffffff6ffffffffffffffdbffffffff",
            INIT_42 => X"00000004000000000000000700000000fffffff6ffffffffffffffe7ffffffff",
            INIT_43 => X"0000000c0000000000000011000000000000001300000000fffffff4ffffffff",
            INIT_44 => X"ffffffdcffffffffffffffeaffffffff0000000900000000fffffffcffffffff",
            INIT_45 => X"ffffffebffffffff00000005000000000000001200000000ffffffebffffffff",
            INIT_46 => X"fffffff5ffffffffffffffe9fffffffffffffffcffffffff0000000200000000",
            INIT_47 => X"fffffffefffffffffffffff5fffffffffffffffffffffffffffffff2ffffffff",
            INIT_48 => X"0000000200000000fffffffeffffffffffffffeaffffffff0000000c00000000",
            INIT_49 => X"fffffffafffffffffffffffbffffffffffffffe8ffffffffffffffdcffffffff",
            INIT_4A => X"ffffffe1ffffffff0000000000000000ffffffe3ffffffffffffffe2ffffffff",
            INIT_4B => X"ffffffebffffffffffffffddfffffffffffffff9fffffffffffffffcffffffff",
            INIT_4C => X"ffffffeeffffffffffffffffffffffff0000000200000000ffffffe8ffffffff",
            INIT_4D => X"fffffffbffffffffffffffd9ffffffffffffffd9ffffffffffffffdcffffffff",
            INIT_4E => X"fffffff6ffffffff0000000700000000ffffffecffffffff0000000600000000",
            INIT_4F => X"fffffffbffffffffffffffe5fffffffffffffff6ffffffffffffffdeffffffff",
            INIT_50 => X"fffffff6fffffffffffffff1fffffffffffffff7ffffffff0000001800000000",
            INIT_51 => X"ffffffc9ffffffff0000000000000000fffffff4fffffffffffffff0ffffffff",
            INIT_52 => X"0000002d000000000000002a000000000000000500000000ffffffbcffffffff",
            INIT_53 => X"ffffffe8ffffffff00000028000000000000002c00000000ffffffddffffffff",
            INIT_54 => X"0000003800000000ffffffebffffffff0000001300000000fffffff2ffffffff",
            INIT_55 => X"0000001100000000000000120000000000000012000000000000001e00000000",
            INIT_56 => X"ffffffeeffffffff000000200000000000000023000000000000001600000000",
            INIT_57 => X"fffffffbfffffffffffffff6fffffffffffffff6fffffffffffffffbffffffff",
            INIT_58 => X"0000002b00000000fffffffafffffffffffffffaffffffff0000000a00000000",
            INIT_59 => X"ffffffd4ffffffff0000000300000000ffffffd2fffffffffffffff0ffffffff",
            INIT_5A => X"ffffffe0ffffffffffffffb2fffffffffffffff5ffffffffffffffedffffffff",
            INIT_5B => X"ffffffcfffffffffffffffb3ffffffffffffffa1ffffffffffffffe7ffffffff",
            INIT_5C => X"ffffffc1ffffffffffffffe3ffffffffffffffbeffffffffffffffbdffffffff",
            INIT_5D => X"0000000e00000000ffffffeeffffffff0000000100000000ffffffd0ffffffff",
            INIT_5E => X"fffffffcfffffffffffffffcffffffffffffffdfffffffff0000001f00000000",
            INIT_5F => X"0000000100000000ffffffe8ffffffffffffffe9ffffffffffffffc8ffffffff",
            INIT_60 => X"fffffff7ffffffff0000000a00000000fffffff8ffffffffffffffeeffffffff",
            INIT_61 => X"0000000200000000ffffffe6ffffffff00000004000000000000000800000000",
            INIT_62 => X"ffffffdaffffffff000000340000000000000007000000000000000700000000",
            INIT_63 => X"ffffffbdffffffffffffffa5fffffffffffffff8ffffffff0000001100000000",
            INIT_64 => X"ffffffc5fffffffffffffff3ffffffffffffffffffffffffffffffebffffffff",
            INIT_65 => X"0000000c00000000ffffffe9ffffffffffffffeeffffffff0000001600000000",
            INIT_66 => X"00000001000000000000000b00000000ffffffd6fffffffffffffffeffffffff",
            INIT_67 => X"ffffffe9ffffffffffffffebffffffffffffffeffffffffffffffff6ffffffff",
            INIT_68 => X"0000000a00000000ffffffd5ffffffffffffffd5ffffffffffffffe8ffffffff",
            INIT_69 => X"0000002500000000fffffff3ffffffff0000001300000000fffffff3ffffffff",
            INIT_6A => X"ffffffdeffffffffffffffdeffffffff00000015000000000000001400000000",
            INIT_6B => X"fffffff4ffffffff00000032000000000000000300000000ffffffeeffffffff",
            INIT_6C => X"0000001b00000000fffffffaffffffff0000003d000000000000000f00000000",
            INIT_6D => X"ffffffa6ffffffffffffffebffffffff00000024000000000000000500000000",
            INIT_6E => X"0000003200000000ffffffd6ffffffffffffffe5ffffffff0000002f00000000",
            INIT_6F => X"fffffff6ffffffffffffffebffffffffffffffedffffffff0000000800000000",
            INIT_70 => X"0000000a00000000fffffffcffffffff0000000300000000fffffff3ffffffff",
            INIT_71 => X"fffffff6ffffffff0000000f00000000ffffffebffffffffffffffeeffffffff",
            INIT_72 => X"0000000c00000000ffffffe1fffffffffffffffbffffffff0000000600000000",
            INIT_73 => X"ffffffd0ffffffffffffffc9ffffffffffffffe5ffffffff0000000800000000",
            INIT_74 => X"0000003200000000fffffffcffffffff00000016000000000000000d00000000",
            INIT_75 => X"00000025000000000000002600000000ffffffebffffffff0000001000000000",
            INIT_76 => X"0000003800000000ffffffecffffffffffffffe1ffffffffffffffdaffffffff",
            INIT_77 => X"fffffff1ffffffffffffffeaffffffff0000000c000000000000002e00000000",
            INIT_78 => X"00000028000000000000001600000000ffffffffffffffff0000000200000000",
            INIT_79 => X"0000000a000000000000000b000000000000002600000000ffffffe1ffffffff",
            INIT_7A => X"0000000f00000000fffffff9ffffffff00000025000000000000002800000000",
            INIT_7B => X"0000000600000000000000080000000000000013000000000000000400000000",
            INIT_7C => X"0000000e00000000fffffffbffffffffffffffe0ffffffff0000000000000000",
            INIT_7D => X"000000130000000000000013000000000000001600000000fffffffbffffffff",
            INIT_7E => X"0000000000000000ffffffb4ffffffff00000001000000000000002d00000000",
            INIT_7F => X"00000007000000000000001200000000fffffff5ffffffffffffffd0ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE13;


    MEM_IWGHT_LAYER2_INSTANCE14 : if BRAM_NAME = "iwght_layer2_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd0fffffffffffffff4ffffffff0000001600000000ffffffebffffffff",
            INIT_01 => X"0000000c000000000000000b00000000ffffffe5ffffffffffffffecffffffff",
            INIT_02 => X"ffffffffffffffff0000000e0000000000000017000000000000000c00000000",
            INIT_03 => X"0000000400000000ffffffe8ffffffffffffffd7ffffffffffffffeaffffffff",
            INIT_04 => X"000000020000000000000002000000000000000100000000ffffffe8ffffffff",
            INIT_05 => X"ffffffeeffffffff00000035000000000000001e000000000000000a00000000",
            INIT_06 => X"000000120000000000000030000000000000003100000000fffffffaffffffff",
            INIT_07 => X"ffffffdfffffffffffffffebfffffffffffffffcffffffff0000001d00000000",
            INIT_08 => X"fffffff8ffffffffffffffddffffffffffffffd3ffffffffffffffe5ffffffff",
            INIT_09 => X"ffffffdcffffffffffffffcaffffffffffffffe3ffffffffffffffd7ffffffff",
            INIT_0A => X"0000000c00000000fffffff7ffffffffffffffc5ffffffffffffff9affffffff",
            INIT_0B => X"0000001e00000000000000290000000000000025000000000000000a00000000",
            INIT_0C => X"ffffffe3ffffffff000000130000000000000005000000000000001700000000",
            INIT_0D => X"fffffffeffffffff0000001700000000ffffffc1ffffffffffffffd6ffffffff",
            INIT_0E => X"ffffffb8ffffffffffffffeeffffffff0000001500000000ffffffecffffffff",
            INIT_0F => X"0000000900000000000000170000000000000024000000000000002d00000000",
            INIT_10 => X"0000000500000000ffffffe7ffffffff00000019000000000000001a00000000",
            INIT_11 => X"00000011000000000000000700000000fffffffaffffffff0000000700000000",
            INIT_12 => X"0000001d000000000000000700000000fffffff1fffffffffffffffeffffffff",
            INIT_13 => X"00000022000000000000002900000000ffffffc2ffffffffffffffd6ffffffff",
            INIT_14 => X"0000000e000000000000001f000000000000003200000000ffffffffffffffff",
            INIT_15 => X"0000002a00000000ffffffb6fffffffffffffff6ffffffff0000001900000000",
            INIT_16 => X"0000001c000000000000002d00000000fffffff2ffffffff0000001b00000000",
            INIT_17 => X"0000001b0000000000000041000000000000003f000000000000002d00000000",
            INIT_18 => X"ffffffeaffffffffffffffe2ffffffffffffffe6fffffffffffffffdffffffff",
            INIT_19 => X"fffffff1ffffffff000000070000000000000000000000000000000700000000",
            INIT_1A => X"fffffff2ffffffff0000000100000000ffffffe0ffffffffffffffecffffffff",
            INIT_1B => X"ffffffffffffffffffffffe7ffffffffffffffe8ffffffffffffffecffffffff",
            INIT_1C => X"0000000c00000000fffffff1ffffffff00000004000000000000000300000000",
            INIT_1D => X"00000004000000000000000500000000fffffffbfffffffffffffffeffffffff",
            INIT_1E => X"0000000700000000fffffff3ffffffff0000000200000000ffffffffffffffff",
            INIT_1F => X"0000000b000000000000000a000000000000000c00000000fffffffaffffffff",
            INIT_20 => X"0000000b00000000000000000000000000000000000000000000000a00000000",
            INIT_21 => X"000000020000000000000002000000000000000400000000fffffff2ffffffff",
            INIT_22 => X"ffffffe1ffffffffffffffe5ffffffffffffffebffffffff0000000000000000",
            INIT_23 => X"fffffff9fffffffffffffff9ffffffff0000000600000000ffffffffffffffff",
            INIT_24 => X"ffffffe4fffffffffffffffbffffffffffffffe6fffffffffffffffaffffffff",
            INIT_25 => X"0000000100000000fffffff9ffffffff00000003000000000000000900000000",
            INIT_26 => X"fffffff7ffffffff00000003000000000000000400000000ffffffeaffffffff",
            INIT_27 => X"ffffffe9fffffffffffffff6ffffffff00000000000000000000000f00000000",
            INIT_28 => X"fffffff3ffffffff0000000d000000000000000300000000ffffffe0ffffffff",
            INIT_29 => X"ffffffdeffffffff0000000000000000ffffffe9ffffffff0000001100000000",
            INIT_2A => X"fffffff6ffffffff00000006000000000000000a000000000000000300000000",
            INIT_2B => X"0000000b00000000ffffffefffffffffffffffedffffffffffffffeeffffffff",
            INIT_2C => X"ffffffeaffffffffffffffebffffffffffffffe5ffffffffffffffefffffffff",
            INIT_2D => X"0000000b00000000ffffffe6ffffffffffffffddfffffffffffffff9ffffffff",
            INIT_2E => X"0000000e000000000000000400000000ffffffe6ffffffffffffffe7ffffffff",
            INIT_2F => X"ffffffe8ffffffff0000000e00000000fffffff0ffffffffffffffefffffffff",
            INIT_30 => X"0000000000000000fffffffbffffffffffffffeafffffffffffffff0ffffffff",
            INIT_31 => X"0000000000000000fffffff3ffffffff0000000200000000fffffff3ffffffff",
            INIT_32 => X"ffffffefffffffffffffffecffffffff0000000000000000fffffff1ffffffff",
            INIT_33 => X"ffffffefffffffff0000000a000000000000001100000000fffffff3ffffffff",
            INIT_34 => X"ffffffe9ffffffff00000000000000000000000200000000fffffffcffffffff",
            INIT_35 => X"ffffffe4ffffffff00000001000000000000000000000000fffffff2ffffffff",
            INIT_36 => X"fffffffaffffffff0000000300000000fffffff8ffffffff0000000700000000",
            INIT_37 => X"000000080000000000000000000000000000000000000000fffffffcffffffff",
            INIT_38 => X"00000013000000000000000000000000fffffffefffffffffffffffbffffffff",
            INIT_39 => X"0000000000000000ffffffffffffffff0000000d000000000000000800000000",
            INIT_3A => X"ffffffe7fffffffffffffffaffffffffffffffe5ffffffffffffffdfffffffff",
            INIT_3B => X"fffffff0fffffffffffffffaffffffffffffffecfffffffffffffffeffffffff",
            INIT_3C => X"ffffffe8ffffffffffffffe6ffffffffffffffe8fffffffffffffffbffffffff",
            INIT_3D => X"fffffffeffffffffffffffe6ffffffffffffffe4ffffffff0000000400000000",
            INIT_3E => X"ffffffffffffffffffffffdbffffffffffffffdfffffffff0000000b00000000",
            INIT_3F => X"fffffffbfffffffffffffffeffffffff00000008000000000000000100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffedffffffff0000000700000000ffffffffffffffffffffffe0ffffffff",
            INIT_41 => X"0000000300000000ffffffd8fffffffffffffff0ffffffffffffffe7ffffffff",
            INIT_42 => X"fffffffdffffffffffffffe5ffffffff00000002000000000000000e00000000",
            INIT_43 => X"0000000200000000ffffffffffffffff00000005000000000000000000000000",
            INIT_44 => X"ffffffedffffffff0000000d00000000ffffffe9ffffffff0000000300000000",
            INIT_45 => X"0000000d00000000ffffffebffffffffffffffdfffffffff0000000000000000",
            INIT_46 => X"ffffffe0ffffffffffffffe2fffffffffffffff4ffffffffffffffdeffffffff",
            INIT_47 => X"fffffff9fffffffffffffff7fffffffffffffff8ffffffff0000000300000000",
            INIT_48 => X"00000001000000000000001100000000ffffffe5fffffffffffffff7ffffffff",
            INIT_49 => X"fffffff3ffffffff0000000400000000ffffffeaffffffff0000000d00000000",
            INIT_4A => X"ffffffdbffffffff0000000000000000fffffffaffffffff0000000c00000000",
            INIT_4B => X"0000000c00000000ffffffeefffffffffffffff1fffffffffffffff4ffffffff",
            INIT_4C => X"ffffffe8fffffffffffffff7ffffffffffffffe9ffffffffffffffffffffffff",
            INIT_4D => X"ffffffe5ffffffff0000000100000000fffffff6ffffffffffffffdeffffffff",
            INIT_4E => X"0000000400000000ffffffebffffffffffffffecffffffffffffffe4ffffffff",
            INIT_4F => X"ffffffe7ffffffff0000000300000000fffffff9ffffffffffffffe2ffffffff",
            INIT_50 => X"ffffffe7ffffffffffffffffffffffffffffffffffffffff0000000400000000",
            INIT_51 => X"0000000a00000000ffffffe6ffffffffffffffe0fffffffffffffff2ffffffff",
            INIT_52 => X"0000000300000000fffffff7fffffffffffffffeffffffff0000000000000000",
            INIT_53 => X"ffffffebffffffff00000004000000000000000a00000000ffffffe7ffffffff",
            INIT_54 => X"0000000200000000fffffffafffffffffffffffaffffffffffffffeeffffffff",
            INIT_55 => X"fffffff6ffffffff0000000300000000fffffff5fffffffffffffff4ffffffff",
            INIT_56 => X"fffffff8fffffffffffffff1ffffffffffffffeeffffffffffffffe3ffffffff",
            INIT_57 => X"ffffffefffffffff0000000200000000ffffffedffffffffffffffeeffffffff",
            INIT_58 => X"000000000000000000000002000000000000000500000000fffffff4ffffffff",
            INIT_59 => X"0000000900000000fffffffbffffffffffffffe1ffffffff0000000c00000000",
            INIT_5A => X"0000000400000000ffffffedffffffffffffffeffffffffffffffff8ffffffff",
            INIT_5B => X"fffffff3ffffffff0000000300000000ffffffdfffffffffffffffe4ffffffff",
            INIT_5C => X"00000005000000000000000600000000ffffffe2ffffffff0000000600000000",
            INIT_5D => X"000000020000000000000002000000000000000100000000fffffffeffffffff",
            INIT_5E => X"00000010000000000000000900000000ffffffebffffffff0000000b00000000",
            INIT_5F => X"fffffffeffffffff0000001500000000ffffffffffffffff0000000600000000",
            INIT_60 => X"0000000b00000000ffffffe9ffffffff0000000200000000fffffffdffffffff",
            INIT_61 => X"fffffffaffffffffffffffe1ffffffffffffffe2ffffffff0000000100000000",
            INIT_62 => X"000000230000000000000025000000000000001d00000000ffffffd5ffffffff",
            INIT_63 => X"0000006200000000fffffff6fffffffffffffff9ffffffff0000002100000000",
            INIT_64 => X"fffffffeffffffff0000000c0000000000000005000000000000002300000000",
            INIT_65 => X"0000000f00000000ffffffa3fffffffffffffffeffffffffffffffcdffffffff",
            INIT_66 => X"0000003500000000ffffffb9ffffffffffffffbaffffffff0000001000000000",
            INIT_67 => X"fffffff3ffffffff0000000a000000000000001e00000000ffffffd2ffffffff",
            INIT_68 => X"ffffffdcffffffffffffffd1ffffffff0000002200000000ffffffffffffffff",
            INIT_69 => X"0000000e00000000ffffffc8ffffffffffffffe5ffffffff0000002e00000000",
            INIT_6A => X"00000001000000000000002a00000000ffffffcfffffffffffffffdbffffffff",
            INIT_6B => X"0000001e00000000ffffffdbffffffff0000004000000000ffffffdaffffffff",
            INIT_6C => X"0000001000000000000000230000000000000000000000000000003c00000000",
            INIT_6D => X"ffffffd8ffffffff000000350000000000000035000000000000001000000000",
            INIT_6E => X"ffffffe4ffffffffffffff9affffffffffffffedffffffff0000001100000000",
            INIT_6F => X"fffffffcfffffffffffffff6ffffffffffffffd9ffffffff0000000600000000",
            INIT_70 => X"000000110000000000000011000000000000000e000000000000000600000000",
            INIT_71 => X"ffffffdcfffffffffffffffbfffffffffffffff3ffffffffffffffefffffffff",
            INIT_72 => X"00000034000000000000000300000000ffffffa2ffffffff0000004b00000000",
            INIT_73 => X"ffffffd4ffffffff0000002500000000ffffffecffffffffffffffd3ffffffff",
            INIT_74 => X"ffffffedffffffff0000001a00000000fffffffaffffffff0000000100000000",
            INIT_75 => X"fffffff0ffffffffffffffeaffffffff0000002f00000000ffffffc8ffffffff",
            INIT_76 => X"fffffffbffffffff0000000f00000000fffffff3ffffffff0000002600000000",
            INIT_77 => X"ffffffe2fffffffffffffff3ffffffff0000000100000000fffffff4ffffffff",
            INIT_78 => X"0000004000000000ffffffdcffffffff0000000200000000ffffffe2ffffffff",
            INIT_79 => X"ffffffddffffffff00000021000000000000000f00000000ffffffe3ffffffff",
            INIT_7A => X"ffffffd0ffffffffffffffb2ffffffff00000030000000000000000700000000",
            INIT_7B => X"ffffffecffffffffffffffdbffffffffffffffdbffffffff0000000900000000",
            INIT_7C => X"ffffffedffffffff0000000e00000000ffffffe3ffffffffffffff8effffffff",
            INIT_7D => X"ffffffdfffffffff0000004b00000000ffffffceffffffffffffffefffffffff",
            INIT_7E => X"ffffffe1ffffffffffffffe6ffffffff0000001500000000fffffff0ffffffff",
            INIT_7F => X"0000000c00000000fffffff2ffffffff00000007000000000000002d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE14;


    MEM_IWGHT_LAYER2_INSTANCE15 : if BRAM_NAME = "iwght_layer2_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff4fffffffffffffffbfffffffffffffffafffffffffffffff8ffffffff",
            INIT_01 => X"0000001c000000000000000800000000ffffffffffffffff0000000100000000",
            INIT_02 => X"fffffff9ffffffffffffffe7ffffffffffffffe9ffffffff0000002100000000",
            INIT_03 => X"ffffffecffffffffffffffedffffffffffffffe4ffffffff0000001000000000",
            INIT_04 => X"ffffffe3ffffffff00000011000000000000001500000000fffffff2ffffffff",
            INIT_05 => X"0000001200000000ffffffdfffffffff0000000d000000000000002100000000",
            INIT_06 => X"0000002700000000fffffff5ffffffff00000006000000000000001c00000000",
            INIT_07 => X"0000003a00000000000000170000000000000015000000000000003200000000",
            INIT_08 => X"fffffff8ffffffff00000037000000000000002b000000000000001a00000000",
            INIT_09 => X"000000180000000000000035000000000000003a000000000000003c00000000",
            INIT_0A => X"0000001c00000000fffffff4ffffffff0000001c000000000000000c00000000",
            INIT_0B => X"0000000600000000ffffffe9ffffffffffffffeaffffffff0000000a00000000",
            INIT_0C => X"000000250000000000000008000000000000002600000000ffffffcaffffffff",
            INIT_0D => X"00000009000000000000003500000000fffffff8fffffffffffffff4ffffffff",
            INIT_0E => X"fffffff8ffffffff0000000e000000000000001b000000000000001600000000",
            INIT_0F => X"fffffff6ffffffffffffffe5ffffffff00000021000000000000001e00000000",
            INIT_10 => X"fffffff3ffffffffffffffe7ffffffffffffffe0ffffffff0000001700000000",
            INIT_11 => X"ffffffedffffffffffffffe6ffffffffffffffe1ffffffffffffffd2ffffffff",
            INIT_12 => X"0000000b00000000ffffffe8ffffffff00000020000000000000000800000000",
            INIT_13 => X"fffffff9ffffffffffffffe8ffffffffffffffdfffffffff0000004100000000",
            INIT_14 => X"fffffffaffffffffffffffc4fffffffffffffffcffffffff0000002500000000",
            INIT_15 => X"ffffffecffffffff0000000900000000ffffffbdffffffff0000001800000000",
            INIT_16 => X"fffffff1ffffffff0000003d0000000000000005000000000000000300000000",
            INIT_17 => X"0000000300000000000000040000000000000038000000000000001b00000000",
            INIT_18 => X"0000001a00000000fffffff1ffffffff00000020000000000000002f00000000",
            INIT_19 => X"0000001700000000fffffff2ffffffffffffffd9ffffffff0000001700000000",
            INIT_1A => X"00000016000000000000000d000000000000001400000000ffffffefffffffff",
            INIT_1B => X"0000000e00000000fffffffeffffffff00000005000000000000002a00000000",
            INIT_1C => X"0000001400000000ffffffe6ffffffffffffffcaffffffffffffffcfffffffff",
            INIT_1D => X"0000000300000000fffffff4ffffffffffffffd4ffffffff0000001700000000",
            INIT_1E => X"0000000500000000ffffffd0ffffffffffffffd7ffffffff0000001f00000000",
            INIT_1F => X"0000000f000000000000000c00000000ffffffe2ffffffff0000001800000000",
            INIT_20 => X"fffffff4ffffffff0000000400000000ffffffdfffffffffffffffd1ffffffff",
            INIT_21 => X"ffffffecffffffff0000000f000000000000000400000000ffffffecffffffff",
            INIT_22 => X"00000015000000000000000000000000ffffffcaffffffff0000002900000000",
            INIT_23 => X"0000001500000000ffffffc8ffffffffffffffb6ffffffffffffffc0ffffffff",
            INIT_24 => X"00000018000000000000001700000000ffffffd1ffffffff0000000400000000",
            INIT_25 => X"000000100000000000000014000000000000000a00000000ffffffd5ffffffff",
            INIT_26 => X"0000000d000000000000001d00000000ffffffe3ffffffff0000001600000000",
            INIT_27 => X"ffffffedffffffff0000000b000000000000001d00000000fffffff1ffffffff",
            INIT_28 => X"fffffff5ffffffffffffffd5ffffffffffffffd8ffffffffffffffe0ffffffff",
            INIT_29 => X"ffffffc4ffffffffffffffdbfffffffffffffff0ffffffffffffffeaffffffff",
            INIT_2A => X"ffffffecffffffff0000001a000000000000001700000000ffffffd4ffffffff",
            INIT_2B => X"00000041000000000000001100000000ffffffc6fffffffffffffff1ffffffff",
            INIT_2C => X"fffffff7ffffffffffffffc6ffffffff0000004d000000000000007400000000",
            INIT_2D => X"fffffff8ffffffffffffff9bffffffffffffffafffffffffffffffdeffffffff",
            INIT_2E => X"ffffffa3ffffffff00000018000000000000003e000000000000001000000000",
            INIT_2F => X"ffffffbbffffffffffffffbbffffffffffffffb6ffffffffffffffe9ffffffff",
            INIT_30 => X"0000003b000000000000003400000000ffffffe6ffffffff0000000b00000000",
            INIT_31 => X"ffffffe9fffffffffffffffcffffffffffffffd8ffffffffffffffc9ffffffff",
            INIT_32 => X"0000000000000000ffffffe6ffffffff0000001800000000ffffffe2ffffffff",
            INIT_33 => X"ffffffe6fffffffffffffff3ffffffff0000002f000000000000002c00000000",
            INIT_34 => X"fffffff5ffffffff00000027000000000000003d000000000000006300000000",
            INIT_35 => X"fffffff5ffffffff0000002200000000ffffffacffffffffffffffcfffffffff",
            INIT_36 => X"ffffffd7ffffffff00000000000000000000000100000000ffffffd9ffffffff",
            INIT_37 => X"0000000600000000ffffffe3ffffffff00000014000000000000001e00000000",
            INIT_38 => X"0000001800000000fffffff6ffffffff0000000b000000000000003c00000000",
            INIT_39 => X"ffffffa5ffffffffffffffe0ffffffffffffffc2ffffffffffffffefffffffff",
            INIT_3A => X"ffffff9affffffffffffffaefffffffffffffffdffffffffffffffcfffffffff",
            INIT_3B => X"00000000000000000000000e00000000ffffffb7ffffffffffffffd1ffffffff",
            INIT_3C => X"00000000000000000000000c000000000000000a000000000000003a00000000",
            INIT_3D => X"0000001900000000000000290000000000000010000000000000000a00000000",
            INIT_3E => X"ffffffeefffffffffffffff8ffffffffffffffebffffffff0000001600000000",
            INIT_3F => X"ffffffc4fffffffffffffffcfffffffffffffff2ffffffffffffffddffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002400000000fffffffcfffffffffffffff5fffffffffffffff5ffffffff",
            INIT_41 => X"ffffffdbffffffffffffffebffffffffffffffbfffffffff0000000700000000",
            INIT_42 => X"ffffffecffffffff0000000a00000000ffffffd6ffffffffffffffeeffffffff",
            INIT_43 => X"0000001400000000fffffff3ffffffffffffffc6ffffffffffffffa1ffffffff",
            INIT_44 => X"000000570000000000000049000000000000002a000000000000001500000000",
            INIT_45 => X"0000002a00000000ffffffd3ffffffff0000001a000000000000005e00000000",
            INIT_46 => X"0000000800000000000000320000000000000022000000000000003900000000",
            INIT_47 => X"0000000500000000fffffffbffffffffffffffdbffffffffffffffd7ffffffff",
            INIT_48 => X"00000015000000000000001100000000fffffff1ffffffff0000000000000000",
            INIT_49 => X"0000000700000000fffffff8ffffffff0000000500000000ffffffffffffffff",
            INIT_4A => X"0000000e000000000000002400000000fffffff9ffffffff0000001f00000000",
            INIT_4B => X"00000001000000000000001d000000000000000b000000000000000800000000",
            INIT_4C => X"ffffffe8fffffffffffffff2ffffffffffffffdaffffffff0000000200000000",
            INIT_4D => X"00000007000000000000002b00000000ffffffe4ffffffffffffffb9ffffffff",
            INIT_4E => X"0000001a000000000000003700000000fffffffaffffffff0000002a00000000",
            INIT_4F => X"ffffffc1ffffffffffffffe7ffffffff0000000c000000000000001300000000",
            INIT_50 => X"00000000000000000000000a00000000fffffffdffffffffffffffd1ffffffff",
            INIT_51 => X"000000040000000000000038000000000000002100000000ffffffffffffffff",
            INIT_52 => X"ffffffebffffffffffffffedffffffff00000007000000000000000d00000000",
            INIT_53 => X"0000000400000000ffffffeaffffffff0000001200000000ffffffedffffffff",
            INIT_54 => X"ffffffdfffffffffffffffe0ffffffffffffffdfffffffffffffffe8ffffffff",
            INIT_55 => X"000000140000000000000018000000000000002a000000000000001c00000000",
            INIT_56 => X"ffffffbbffffffffffffffdefffffffffffffffbffffffffffffffeaffffffff",
            INIT_57 => X"ffffffecffffffff0000000c000000000000001000000000ffffffefffffffff",
            INIT_58 => X"0000000e00000000fffffff2ffffffffffffffeafffffffffffffff2ffffffff",
            INIT_59 => X"0000003b000000000000002a00000000ffffffe5ffffffff0000000700000000",
            INIT_5A => X"00000028000000000000001e0000000000000005000000000000001800000000",
            INIT_5B => X"ffffffc8fffffffffffffff1ffffffff0000001100000000ffffffd7ffffffff",
            INIT_5C => X"ffffffc3ffffffffffffffecffffffffffffffbcffffffffffffffdcffffffff",
            INIT_5D => X"0000001c0000000000000002000000000000001b00000000ffffffbbffffffff",
            INIT_5E => X"ffffffedffffffff00000016000000000000001c000000000000001400000000",
            INIT_5F => X"ffffffebffffffffffffffc1fffffffffffffffaffffffff0000001900000000",
            INIT_60 => X"0000001100000000ffffffffffffffff0000001600000000ffffffe4ffffffff",
            INIT_61 => X"ffffffd6ffffffffffffffecffffffff0000001c000000000000001200000000",
            INIT_62 => X"00000020000000000000000c00000000ffffffe9fffffffffffffffeffffffff",
            INIT_63 => X"0000000000000000ffffffd7ffffffffffffffbdffffffff0000000500000000",
            INIT_64 => X"ffffffdafffffffffffffff5ffffffff0000000000000000ffffffdfffffffff",
            INIT_65 => X"fffffff6ffffffffffffffc0ffffffff0000001800000000ffffffdcffffffff",
            INIT_66 => X"ffffffeffffffffffffffff2fffffffffffffff2ffffffff0000000000000000",
            INIT_67 => X"0000001600000000fffffff3ffffffffffffffe7ffffffff0000002000000000",
            INIT_68 => X"00000013000000000000001d000000000000000200000000ffffffffffffffff",
            INIT_69 => X"000000080000000000000007000000000000001d000000000000002100000000",
            INIT_6A => X"0000000000000000ffffffdcffffffffffffffb7ffffffffffffffb5ffffffff",
            INIT_6B => X"00000010000000000000000c000000000000000e000000000000001a00000000",
            INIT_6C => X"fffffff4ffffffffffffffc4ffffffffffffffe2ffffffff0000001800000000",
            INIT_6D => X"0000001d00000000fffffffaffffffffffffffc5ffffffffffffffddffffffff",
            INIT_6E => X"0000000400000000000000070000000000000001000000000000001300000000",
            INIT_6F => X"ffffffdcffffffffffffffd1ffffffffffffffcfffffffff0000000e00000000",
            INIT_70 => X"ffffffebffffffffffffffe7fffffffffffffff1ffffffffffffffdfffffffff",
            INIT_71 => X"ffffffefffffffffffffffedfffffffffffffff8fffffffffffffff2ffffffff",
            INIT_72 => X"0000001c000000000000002d000000000000002c000000000000002000000000",
            INIT_73 => X"0000002000000000fffffffeffffffff0000000d000000000000000e00000000",
            INIT_74 => X"0000002600000000000000190000000000000011000000000000001200000000",
            INIT_75 => X"0000002e0000000000000017000000000000003f000000000000002400000000",
            INIT_76 => X"ffffffdbffffffff0000000a0000000000000009000000000000000900000000",
            INIT_77 => X"0000001d00000000fffffff3ffffffff0000002200000000ffffffd4ffffffff",
            INIT_78 => X"0000002e00000000000000130000000000000000000000000000003400000000",
            INIT_79 => X"fffffff6ffffffff00000012000000000000000a00000000ffffffd3ffffffff",
            INIT_7A => X"ffffffe6ffffffffffffffd3ffffffff0000002c000000000000001c00000000",
            INIT_7B => X"0000001400000000fffffff2ffffffffffffffd6ffffffffffffffffffffffff",
            INIT_7C => X"0000000f000000000000001e000000000000001600000000fffffff6ffffffff",
            INIT_7D => X"00000009000000000000000f000000000000000d000000000000000f00000000",
            INIT_7E => X"00000011000000000000000e00000000ffffffe9ffffffff0000001c00000000",
            INIT_7F => X"fffffff7ffffffff00000033000000000000001400000000fffffff1ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE15;


    MEM_IWGHT_LAYER2_INSTANCE16 : if BRAM_NAME = "iwght_layer2_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffefffffffff0000001000000000fffffffcffffffffffffffccffffffff",
            INIT_01 => X"0000003c00000000ffffffe6ffffffff0000002700000000fffffffcffffffff",
            INIT_02 => X"0000000c0000000000000022000000000000002300000000fffffff3ffffffff",
            INIT_03 => X"0000001100000000000000000000000000000030000000000000002100000000",
            INIT_04 => X"00000032000000000000001f0000000000000002000000000000001c00000000",
            INIT_05 => X"ffffffc8fffffffffffffff8ffffffffffffffebffffffffffffffccffffffff",
            INIT_06 => X"ffffffe4ffffffffffffffd8fffffffffffffff4ffffffffffffffc9ffffffff",
            INIT_07 => X"ffffffeaffffffffffffffc3ffffffffffffffcffffffffffffffffdffffffff",
            INIT_08 => X"ffffffe9fffffffffffffff9ffffffffffffffceffffffffffffffddffffffff",
            INIT_09 => X"fffffffaffffffffffffffd6ffffffffffffffbffffffffffffffff5ffffffff",
            INIT_0A => X"0000001b000000000000000b00000000ffffffeaffffffff0000001600000000",
            INIT_0B => X"0000001400000000000000470000000000000049000000000000002200000000",
            INIT_0C => X"ffffffe7ffffffffffffffe7fffffffffffffffcffffffff0000002300000000",
            INIT_0D => X"0000000000000000ffffffcbffffffffffffffe6ffffffffffffffefffffffff",
            INIT_0E => X"ffffffc0ffffffffffffff96ffffffffffffff7affffffffffffffd9ffffffff",
            INIT_0F => X"0000000d000000000000000300000000ffffffdfffffffffffffff8effffffff",
            INIT_10 => X"ffffffeffffffffffffffff8fffffffffffffff5fffffffffffffff4ffffffff",
            INIT_11 => X"fffffff8fffffffffffffff6fffffffffffffffbffffffff0000000e00000000",
            INIT_12 => X"00000000000000000000000500000000fffffff9ffffffff0000000500000000",
            INIT_13 => X"0000002200000000ffffffe6ffffffffffffffd8ffffffff0000002700000000",
            INIT_14 => X"0000000d00000000ffffffefffffffff0000001c000000000000000e00000000",
            INIT_15 => X"ffffffdeffffffffffffffd7ffffffffffffffc2ffffffff0000000600000000",
            INIT_16 => X"00000058000000000000001f00000000ffffffedffffffffffffffe6ffffffff",
            INIT_17 => X"ffffffc4ffffffff0000001000000000ffffffeafffffffffffffff9ffffffff",
            INIT_18 => X"ffffffdeffffffff0000002700000000ffffffbbffffffffffffffb4ffffffff",
            INIT_19 => X"ffffffecfffffffffffffff0ffffffff00000009000000000000002f00000000",
            INIT_1A => X"ffffffdcfffffffffffffff7fffffffffffffff5ffffffffffffffecffffffff",
            INIT_1B => X"ffffffe1ffffffff00000000000000000000002c00000000ffffffd0ffffffff",
            INIT_1C => X"ffffffe6ffffffff0000000600000000fffffffaffffffff0000001100000000",
            INIT_1D => X"00000010000000000000002a000000000000001f000000000000001200000000",
            INIT_1E => X"ffffffeeffffffffffffffe4ffffffff00000003000000000000003100000000",
            INIT_1F => X"0000000e0000000000000013000000000000000700000000ffffffcaffffffff",
            INIT_20 => X"ffffffc3fffffffffffffff6ffffffff0000000a00000000fffffffdffffffff",
            INIT_21 => X"fffffff8ffffffffffffffeaffffffff0000001c000000000000000000000000",
            INIT_22 => X"0000001000000000ffffffdefffffffffffffffbffffffffffffffffffffffff",
            INIT_23 => X"000000120000000000000011000000000000000f000000000000000e00000000",
            INIT_24 => X"ffffffdbffffffff000000010000000000000002000000000000000800000000",
            INIT_25 => X"ffffffbeffffffffffffffc2ffffffff0000000e00000000ffffffccffffffff",
            INIT_26 => X"ffffffe5fffffffffffffff9ffffffff00000012000000000000000600000000",
            INIT_27 => X"ffffffe0ffffffffffffffc8fffffffffffffffcfffffffffffffff2ffffffff",
            INIT_28 => X"0000003a0000000000000034000000000000001300000000ffffffedffffffff",
            INIT_29 => X"ffffffd8ffffffff0000002f00000000fffffff4fffffffffffffffdffffffff",
            INIT_2A => X"ffffffdfffffffff0000002e00000000fffffffeffffffff0000001600000000",
            INIT_2B => X"0000000d00000000ffffffd2ffffffff0000001300000000ffffffd3ffffffff",
            INIT_2C => X"fffffffcffffffff0000002800000000ffffffe4ffffffff0000005b00000000",
            INIT_2D => X"ffffffe1ffffffffffffffceffffffffffffffceffffffff0000000f00000000",
            INIT_2E => X"ffffffebffffffffffffffbfffffffffffffffecffffffffffffffebffffffff",
            INIT_2F => X"0000001300000000fffffff1ffffffff0000001b000000000000000c00000000",
            INIT_30 => X"ffffffeafffffffffffffffbffffffff00000006000000000000001300000000",
            INIT_31 => X"0000002b00000000fffffffafffffffffffffff6ffffffffffffffd6ffffffff",
            INIT_32 => X"ffffffdbffffffff00000031000000000000000100000000ffffffcaffffffff",
            INIT_33 => X"fffffff2fffffffffffffffbffffffff00000027000000000000001800000000",
            INIT_34 => X"ffffffe6ffffffff0000001b00000000fffffffbffffffffffffffd8ffffffff",
            INIT_35 => X"ffffffcdffffffff0000000200000000ffffffd6ffffffffffffffe9ffffffff",
            INIT_36 => X"ffffffedffffffff0000001900000000ffffffddffffffffffffffbdffffffff",
            INIT_37 => X"00000018000000000000001a000000000000004200000000ffffffd4ffffffff",
            INIT_38 => X"00000008000000000000002b0000000000000031000000000000002a00000000",
            INIT_39 => X"0000000000000000fffffff3ffffffff00000005000000000000001300000000",
            INIT_3A => X"0000000a00000000fffffff6ffffffff0000001900000000ffffffedffffffff",
            INIT_3B => X"0000001200000000ffffffecffffffffffffffffffffffff0000003400000000",
            INIT_3C => X"ffffffcfffffffffffffffe8ffffffff0000000100000000fffffff7ffffffff",
            INIT_3D => X"fffffff3ffffffffffffffe7ffffffffffffffe2ffffffffffffffc3ffffffff",
            INIT_3E => X"0000001100000000ffffffc1ffffffffffffff9cffffffffffffffa6ffffffff",
            INIT_3F => X"000000090000000000000026000000000000000a000000000000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffd3ffffffff0000001f0000000000000001000000000000000a00000000",
            INIT_41 => X"0000002800000000ffffffdcffffffffffffffe8ffffffffffffffd7ffffffff",
            INIT_42 => X"0000002f000000000000001b00000000ffffffedffffffff0000000e00000000",
            INIT_43 => X"000000090000000000000004000000000000001d000000000000001700000000",
            INIT_44 => X"00000014000000000000001500000000fffffff2ffffffff0000001000000000",
            INIT_45 => X"fffffff5ffffffffffffffeeffffffff0000001400000000fffffff9ffffffff",
            INIT_46 => X"000000010000000000000006000000000000000300000000fffffff1ffffffff",
            INIT_47 => X"0000005100000000fffffff6fffffffffffffff0ffffffffffffffe0ffffffff",
            INIT_48 => X"fffffff2ffffffff000000070000000000000031000000000000003b00000000",
            INIT_49 => X"ffffffedfffffffffffffffdfffffffffffffff2ffffffff0000000d00000000",
            INIT_4A => X"fffffff6ffffffff00000017000000000000000500000000fffffffbffffffff",
            INIT_4B => X"0000000000000000ffffffefffffffff0000000d000000000000001b00000000",
            INIT_4C => X"ffffffc3ffffffffffffffc2fffffffffffffff1ffffffff0000001d00000000",
            INIT_4D => X"00000001000000000000003500000000ffffffe0ffffffff0000000f00000000",
            INIT_4E => X"0000002b000000000000002e00000000ffffffeaffffffffffffffc9ffffffff",
            INIT_4F => X"000000060000000000000003000000000000001f000000000000001d00000000",
            INIT_50 => X"0000000f00000000fffffffcffffffffffffffffffffffff0000001700000000",
            INIT_51 => X"ffffffd6ffffffff0000000a000000000000000900000000fffffffcffffffff",
            INIT_52 => X"ffffffd0ffffffffffffffe6ffffffffffffffe9ffffffff0000001700000000",
            INIT_53 => X"ffffffeeffffffff0000000500000000fffffff4ffffffffffffffe5ffffffff",
            INIT_54 => X"ffffffbdffffffffffffff98ffffffffffffffe4ffffffffffffffd6ffffffff",
            INIT_55 => X"ffffffc2ffffffffffffffdefffffffffffffff6ffffffffffffff6cffffffff",
            INIT_56 => X"0000004100000000000000150000000000000000000000000000002200000000",
            INIT_57 => X"fffffff2fffffffffffffffcffffffff00000039000000000000001e00000000",
            INIT_58 => X"00000000000000000000000300000000fffffffaffffffff0000000e00000000",
            INIT_59 => X"fffffff8ffffffff0000000600000000fffffff4ffffffffffffffefffffffff",
            INIT_5A => X"ffffffe1ffffffff00000006000000000000000000000000fffffffaffffffff",
            INIT_5B => X"ffffffddffffffffffffffd0ffffffffffffffc3ffffffff0000000000000000",
            INIT_5C => X"0000002400000000ffffffe8ffffffffffffffe2ffffffffffffffe8ffffffff",
            INIT_5D => X"000000320000000000000025000000000000002100000000fffffff9ffffffff",
            INIT_5E => X"0000001a00000000ffffffd4ffffffff0000001a000000000000001300000000",
            INIT_5F => X"00000003000000000000000800000000fffffff7ffffffff0000001b00000000",
            INIT_60 => X"00000000000000000000001b000000000000001f000000000000000500000000",
            INIT_61 => X"0000002400000000fffffff0ffffffffffffffdffffffffffffffff1ffffffff",
            INIT_62 => X"ffffffbfffffffff0000000000000000ffffff9dffffffffffffffd4ffffffff",
            INIT_63 => X"ffffffc2fffffffffffffff6ffffffffffffffebffffffffffffffd0ffffffff",
            INIT_64 => X"0000000100000000ffffffe7ffffffffffffffe9ffffffff0000000000000000",
            INIT_65 => X"0000001500000000ffffffe0ffffffffffffffd3ffffffffffffffc9ffffffff",
            INIT_66 => X"0000002a00000000000000290000000000000027000000000000000c00000000",
            INIT_67 => X"0000001400000000000000220000000000000018000000000000005100000000",
            INIT_68 => X"ffffffd6ffffffff000000060000000000000008000000000000000d00000000",
            INIT_69 => X"ffffffe9fffffffffffffffcffffffffffffffcdffffffffffffffd5ffffffff",
            INIT_6A => X"ffffffd3ffffffffffffffe4fffffffffffffffefffffffffffffff5ffffffff",
            INIT_6B => X"0000002600000000ffffffa6ffffffffffffffc4ffffffffffffffc1ffffffff",
            INIT_6C => X"0000000200000000fffffffbffffffff00000023000000000000001500000000",
            INIT_6D => X"0000002900000000fffffff7fffffffffffffffbffffffff0000000600000000",
            INIT_6E => X"ffffffe5fffffffffffffffdffffffffffffffecfffffffffffffffdffffffff",
            INIT_6F => X"0000002e0000000000000018000000000000001700000000fffffffbffffffff",
            INIT_70 => X"ffffffe4ffffffffffffffe1ffffffff00000011000000000000003400000000",
            INIT_71 => X"fffffff4ffffffff0000000300000000fffffffaffffffff0000000400000000",
            INIT_72 => X"00000022000000000000002100000000fffffff7fffffffffffffffeffffffff",
            INIT_73 => X"000000150000000000000011000000000000000d000000000000002600000000",
            INIT_74 => X"0000001d00000000ffffffe2ffffffffffffffe0fffffffffffffff4ffffffff",
            INIT_75 => X"0000001b0000000000000017000000000000000d000000000000001600000000",
            INIT_76 => X"fffffffcffffffff00000034000000000000000400000000ffffffeeffffffff",
            INIT_77 => X"fffffffbffffffffffffffcaffffffffffffffccffffffffffffffbcffffffff",
            INIT_78 => X"ffffffeaffffffffffffffdcffffffffffffffeafffffffffffffff8ffffffff",
            INIT_79 => X"0000002300000000fffffff1ffffffff0000001300000000fffffffaffffffff",
            INIT_7A => X"ffffffc5ffffffffffffffe1ffffffff0000000000000000fffffff9ffffffff",
            INIT_7B => X"ffffffeaffffffffffffffcdffffffffffffffedffffffffffffffc9ffffffff",
            INIT_7C => X"00000015000000000000000c00000000ffffffe9ffffffffffffffcdffffffff",
            INIT_7D => X"000000310000000000000010000000000000001e000000000000000700000000",
            INIT_7E => X"0000000a0000000000000028000000000000001f000000000000001900000000",
            INIT_7F => X"ffffffdfffffffff0000000000000000ffffffecfffffffffffffff1ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE16;


    MEM_IWGHT_LAYER2_INSTANCE17 : if BRAM_NAME = "iwght_layer2_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffcffffffffffffffcdfffffffffffffff4fffffffffffffff5ffffffff",
            INIT_01 => X"00000003000000000000000c00000000fffffff2fffffffffffffff8ffffffff",
            INIT_02 => X"00000005000000000000000c00000000ffffffe4ffffffffffffffebffffffff",
            INIT_03 => X"0000000f00000000fffffff3ffffffff0000000c00000000ffffffe9ffffffff",
            INIT_04 => X"0000000400000000ffffffe7ffffffff00000012000000000000002c00000000",
            INIT_05 => X"0000000b00000000ffffffebffffffffffffffd9ffffffff0000002c00000000",
            INIT_06 => X"0000001700000000ffffffe2ffffffffffffffe5ffffffffffffffeaffffffff",
            INIT_07 => X"00000024000000000000002f000000000000000400000000ffffffd5ffffffff",
            INIT_08 => X"0000001c000000000000002c00000000ffffffd9ffffffff0000001d00000000",
            INIT_09 => X"0000000a00000000fffffffffffffffffffffff8ffffffff0000001700000000",
            INIT_0A => X"0000000200000000ffffffd3ffffffff0000002700000000fffffff7ffffffff",
            INIT_0B => X"fffffffaffffffffffffffa7ffffffffffffffdbffffffff0000002200000000",
            INIT_0C => X"ffffff75ffffffff0000003100000000ffffffc0ffffffffffffffb4ffffffff",
            INIT_0D => X"ffffffd8ffffffffffffffa7ffffffff0000004100000000fffffff2ffffffff",
            INIT_0E => X"ffffffffffffffffffffffd1ffffffffffffffbefffffffffffffffeffffffff",
            INIT_0F => X"ffffffcdffffffff0000000700000000ffffffc8ffffffffffffffbaffffffff",
            INIT_10 => X"fffffffaffffffffffffffe2ffffffff0000000a00000000ffffffe5ffffffff",
            INIT_11 => X"0000001900000000ffffffe5ffffffff00000020000000000000001f00000000",
            INIT_12 => X"0000000000000000ffffffeffffffffffffffffcffffffff0000000d00000000",
            INIT_13 => X"0000001e00000000fffffffefffffffffffffff5ffffffff0000001b00000000",
            INIT_14 => X"0000004000000000fffffff7ffffffffffffffc9ffffffffffffffe5ffffffff",
            INIT_15 => X"00000008000000000000001100000000fffffffcffffffffffffffc3ffffffff",
            INIT_16 => X"ffffffedffffffff0000001900000000ffffffe6fffffffffffffffaffffffff",
            INIT_17 => X"0000000300000000ffffffe5ffffffff0000000e00000000ffffffe3ffffffff",
            INIT_18 => X"fffffffdffffffffffffffecffffffff00000001000000000000000a00000000",
            INIT_19 => X"0000001700000000ffffffc9ffffffff00000010000000000000000400000000",
            INIT_1A => X"0000002d00000000fffffffdffffffffffffffd2ffffffff0000003000000000",
            INIT_1B => X"fffffff5ffffffff0000002a0000000000000002000000000000002300000000",
            INIT_1C => X"ffffffe7fffffffffffffffdffffffff00000028000000000000000800000000",
            INIT_1D => X"0000003400000000fffffffeffffffffffffffcafffffffffffffff0ffffffff",
            INIT_1E => X"0000002000000000ffffffccfffffffffffffffcffffffffffffffe5ffffffff",
            INIT_1F => X"0000001000000000000000040000000000000009000000000000000200000000",
            INIT_20 => X"fffffff3fffffffffffffff3ffffffff0000000700000000fffffff9ffffffff",
            INIT_21 => X"ffffffb8ffffffff000000000000000000000015000000000000000a00000000",
            INIT_22 => X"0000002300000000ffffffe9fffffffffffffffaffffffff0000000700000000",
            INIT_23 => X"0000002500000000ffffffdcffffffff00000027000000000000003700000000",
            INIT_24 => X"0000000d000000000000001200000000fffffffffffffffffffffff5ffffffff",
            INIT_25 => X"00000022000000000000001c00000000ffffffe8ffffffff0000002100000000",
            INIT_26 => X"0000000f00000000fffffffdffffffffffffffe4ffffffffffffffcfffffffff",
            INIT_27 => X"0000000e000000000000003900000000fffffff1ffffffffffffffeaffffffff",
            INIT_28 => X"0000000200000000ffffffcdffffffff0000001c00000000fffffff5ffffffff",
            INIT_29 => X"0000001a000000000000001000000000ffffffcaffffffff0000004200000000",
            INIT_2A => X"0000000800000000fffffff0fffffffffffffff2ffffffffffffffe6ffffffff",
            INIT_2B => X"fffffff0ffffffffffffffe6ffffffffffffffc9ffffffffffffffddffffffff",
            INIT_2C => X"ffffffedffffffff0000003000000000ffffffbeffffffff0000000e00000000",
            INIT_2D => X"ffffffe7ffffffff0000000500000000fffffff8ffffffff0000001600000000",
            INIT_2E => X"ffffffeffffffffffffffff7ffffffff0000000600000000ffffffeeffffffff",
            INIT_2F => X"ffffffe4ffffffffffffffffffffffffffffff89ffffffff0000000100000000",
            INIT_30 => X"fffffffffffffffffffffff7ffffffffffffffeaffffffffffffffc0ffffffff",
            INIT_31 => X"fffffff7fffffffffffffffdfffffffffffffff8ffffffffffffffd2ffffffff",
            INIT_32 => X"0000000700000000ffffffedffffffffffffffd5ffffffff0000002300000000",
            INIT_33 => X"0000001500000000fffffff1ffffffffffffffc7ffffffffffffffd6ffffffff",
            INIT_34 => X"0000001c0000000000000033000000000000003b000000000000001600000000",
            INIT_35 => X"fffffff3fffffffffffffff2ffffffff0000000a00000000fffffff0ffffffff",
            INIT_36 => X"ffffffe3fffffffffffffff7ffffffff0000001100000000fffffff4ffffffff",
            INIT_37 => X"00000006000000000000001e000000000000003200000000fffffff6ffffffff",
            INIT_38 => X"fffffff1ffffffffffffffe7ffffffffffffffccffffffff0000001a00000000",
            INIT_39 => X"ffffffecffffffff0000003f00000000ffffffc7ffffffffffffffe7ffffffff",
            INIT_3A => X"ffffffd9ffffffffffffffe8ffffffff0000003400000000fffffff1ffffffff",
            INIT_3B => X"0000000c00000000ffffffdfffffffffffffffdcfffffffffffffffeffffffff",
            INIT_3C => X"fffffffcffffffff0000000000000000ffffffdaffffffffffffffd4ffffffff",
            INIT_3D => X"ffffffe6ffffffff00000018000000000000001500000000fffffff8ffffffff",
            INIT_3E => X"0000000400000000ffffffddffffffffffffffd5ffffffffffffffd2ffffffff",
            INIT_3F => X"fffffff3ffffffff00000014000000000000000400000000fffffff4ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000090000000000000002000000000000000300000000fffffffcffffffff",
            INIT_41 => X"00000030000000000000000200000000ffffff91ffffffffffffffdfffffffff",
            INIT_42 => X"ffffffc9ffffffff0000001300000000ffffffa8ffffffffffffff9affffffff",
            INIT_43 => X"0000001e0000000000000015000000000000001600000000ffffffd6ffffffff",
            INIT_44 => X"ffffffe1fffffffffffffff4ffffffff0000001700000000fffffffbffffffff",
            INIT_45 => X"ffffffdfffffffff0000000a0000000000000021000000000000001b00000000",
            INIT_46 => X"0000001a000000000000000f00000000fffffff3ffffffff0000001000000000",
            INIT_47 => X"ffffffd3ffffffff0000002b000000000000001300000000ffffffeaffffffff",
            INIT_48 => X"0000000200000000ffffffe4ffffffffffffffe1ffffffffffffffe0ffffffff",
            INIT_49 => X"ffffffe5fffffffffffffff7ffffffffffffffe0fffffffffffffff4ffffffff",
            INIT_4A => X"0000003c0000000000000036000000000000003200000000ffffffbbffffffff",
            INIT_4B => X"000000340000000000000041000000000000004e000000000000001e00000000",
            INIT_4C => X"000000220000000000000016000000000000004f000000000000001600000000",
            INIT_4D => X"ffffffc8ffffffffffffffdaffffffffffffffbeffffffff0000000800000000",
            INIT_4E => X"ffffffd9ffffffff0000000900000000fffffffdffffffffffffffeeffffffff",
            INIT_4F => X"00000009000000000000001b000000000000001200000000fffffff4ffffffff",
            INIT_50 => X"fffffff4ffffffffffffffecfffffffffffffff5fffffffffffffff2ffffffff",
            INIT_51 => X"0000000800000000000000020000000000000010000000000000001b00000000",
            INIT_52 => X"00000007000000000000000500000000fffffff9ffffffff0000000200000000",
            INIT_53 => X"00000024000000000000002f000000000000001300000000ffffffefffffffff",
            INIT_54 => X"00000019000000000000001000000000fffffffaffffffff0000000200000000",
            INIT_55 => X"fffffffcffffffff000000020000000000000007000000000000000e00000000",
            INIT_56 => X"fffffff2ffffffffffffff90ffffffffffffffbfffffffff0000002d00000000",
            INIT_57 => X"ffffffddffffffff0000001200000000ffffffdafffffffffffffff7ffffffff",
            INIT_58 => X"ffffffe7ffffffffffffffe9fffffffffffffffeffffffffffffffe5ffffffff",
            INIT_59 => X"fffffff1ffffffffffffffd3ffffffffffffffd4ffffffff0000000a00000000",
            INIT_5A => X"fffffffdffffffffffffffd5ffffffffffffffecffffffff0000000600000000",
            INIT_5B => X"ffffffc6ffffffffffffffdcffffffffffffffd5ffffffffffffffb0ffffffff",
            INIT_5C => X"00000026000000000000000b000000000000001600000000ffffffc2ffffffff",
            INIT_5D => X"0000001500000000fffffffeffffffff0000000f000000000000000800000000",
            INIT_5E => X"fffffff3ffffffffffffffd3ffffffff0000001c000000000000002100000000",
            INIT_5F => X"fffffff6ffffffff0000001d00000000ffffffeaffffffffffffffafffffffff",
            INIT_60 => X"0000002000000000ffffffd6fffffffffffffffbfffffffffffffff4ffffffff",
            INIT_61 => X"ffffffc5fffffffffffffff6ffffffff00000027000000000000000f00000000",
            INIT_62 => X"ffffffb1ffffffffffffffd9fffffffffffffff1ffffffffffffffd2ffffffff",
            INIT_63 => X"ffffffabffffffff0000000b00000000fffffff4fffffffffffffffdffffffff",
            INIT_64 => X"fffffff2ffffffff0000000400000000ffffffd3ffffffffffffffc6ffffffff",
            INIT_65 => X"00000000000000000000000a000000000000000f00000000ffffffefffffffff",
            INIT_66 => X"fffffff1ffffffff0000000b0000000000000019000000000000001100000000",
            INIT_67 => X"fffffff5ffffffff0000000d000000000000000700000000fffffffaffffffff",
            INIT_68 => X"ffffffedffffffff0000000c00000000ffffffedffffffff0000000100000000",
            INIT_69 => X"fffffff1ffffffffffffffffffffffffffffffefffffffffffffffebffffffff",
            INIT_6A => X"ffffffb2fffffffffffffff4ffffffff0000003b00000000fffffffaffffffff",
            INIT_6B => X"0000000a000000000000001c00000000fffffff5ffffffffffffffe1ffffffff",
            INIT_6C => X"0000000b000000000000000c000000000000000e000000000000001f00000000",
            INIT_6D => X"ffffffecffffffff0000000300000000fffffff8ffffffff0000001400000000",
            INIT_6E => X"0000001100000000ffffffedffffffffffffffdbffffffffffffffcbffffffff",
            INIT_6F => X"00000000000000000000002f00000000fffffff6ffffffff0000000100000000",
            INIT_70 => X"000000250000000000000019000000000000000200000000ffffffdbffffffff",
            INIT_71 => X"00000029000000000000001500000000fffffff7ffffffff0000002500000000",
            INIT_72 => X"ffffffcdffffffff00000043000000000000001d000000000000003100000000",
            INIT_73 => X"ffffffdbffffffff0000001700000000ffffffecffffffffffffffd5ffffffff",
            INIT_74 => X"ffffffd3fffffffffffffffaffffffff0000003800000000fffffff9ffffffff",
            INIT_75 => X"0000001f000000000000002400000000fffffffdffffffff0000001f00000000",
            INIT_76 => X"ffffffe8ffffffff000000000000000000000008000000000000001d00000000",
            INIT_77 => X"00000023000000000000001c000000000000000000000000ffffffe9ffffffff",
            INIT_78 => X"ffffffe6ffffffffffffffdcffffffffffffffb5ffffffffffffffdbffffffff",
            INIT_79 => X"00000020000000000000002900000000ffffffcaffffffffffffffbeffffffff",
            INIT_7A => X"ffffffa6ffffffffffffffbbffffffffffffffdeffffffff0000002300000000",
            INIT_7B => X"fffffff0ffffffffffffffd4fffffffffffffff6ffffffff0000000400000000",
            INIT_7C => X"0000001400000000ffffffdbffffffff0000004800000000fffffff7ffffffff",
            INIT_7D => X"0000002500000000ffffffdfffffffff00000006000000000000001f00000000",
            INIT_7E => X"fffffffffffffffffffffffbfffffffffffffff3fffffffffffffffeffffffff",
            INIT_7F => X"00000008000000000000000000000000ffffffd5fffffffffffffff2ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE17;


    MEM_IWGHT_LAYER2_INSTANCE18 : if BRAM_NAME = "iwght_layer2_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff7ffffffffffffffe8ffffffff0000001e00000000ffffffdeffffffff",
            INIT_01 => X"0000000d00000000fffffff7ffffffffffffffc5ffffffffffffffceffffffff",
            INIT_02 => X"0000000400000000fffffff4ffffffffffffffe5ffffffffffffffdeffffffff",
            INIT_03 => X"0000002d00000000000000040000000000000006000000000000001a00000000",
            INIT_04 => X"00000007000000000000000500000000ffffffceffffffff0000000600000000",
            INIT_05 => X"0000001500000000fffffff8ffffffff0000001f00000000fffffffeffffffff",
            INIT_06 => X"0000002700000000fffffff4ffffffffffffffe2ffffffffffffffffffffffff",
            INIT_07 => X"fffffffcffffffffffffffe3ffffffffffffffe3ffffffffffffffeaffffffff",
            INIT_08 => X"00000000000000000000000c00000000ffffffeeffffffff0000000900000000",
            INIT_09 => X"00000025000000000000000400000000ffffffd9ffffffff0000000500000000",
            INIT_0A => X"fffffffdffffffffffffffe2ffffffffffffffe3fffffffffffffff3ffffffff",
            INIT_0B => X"000000000000000000000012000000000000000d000000000000002800000000",
            INIT_0C => X"ffffffdbffffffff00000018000000000000000900000000ffffffedffffffff",
            INIT_0D => X"ffffffe8ffffffffffffffc3fffffffffffffffefffffffffffffff6ffffffff",
            INIT_0E => X"00000011000000000000001f0000000000000006000000000000000000000000",
            INIT_0F => X"ffffffddffffffff0000000b000000000000000000000000ffffffcfffffffff",
            INIT_10 => X"fffffff1ffffffff00000029000000000000002b000000000000000900000000",
            INIT_11 => X"0000000200000000ffffffefffffffff0000002100000000fffffff6ffffffff",
            INIT_12 => X"00000044000000000000000f000000000000001e00000000fffffffaffffffff",
            INIT_13 => X"fffffff9ffffffff000000540000000000000031000000000000001e00000000",
            INIT_14 => X"ffffffc9fffffffffffffff8ffffffff0000000a000000000000001600000000",
            INIT_15 => X"fffffff1fffffffffffffffafffffffffffffffaffffffffffffffc2ffffffff",
            INIT_16 => X"ffffffdbffffffff00000032000000000000002f000000000000001b00000000",
            INIT_17 => X"0000000b00000000ffffffedffffffff0000000300000000fffffff5ffffffff",
            INIT_18 => X"0000000c00000000000000050000000000000010000000000000000000000000",
            INIT_19 => X"ffffffe9ffffffffffffffe1ffffffffffffffe2ffffffffffffffeeffffffff",
            INIT_1A => X"fffffff1ffffffffffffffe5ffffffffffffffedffffffffffffffdfffffffff",
            INIT_1B => X"ffffffe0ffffffffffffffdfffffffffffffffa6ffffffffffffffeaffffffff",
            INIT_1C => X"fffffffcffffffffffffffc6ffffffffffffff8fffffffffffffffbdffffffff",
            INIT_1D => X"ffffffdafffffffffffffff4ffffffffffffffe3ffffffffffffffdbffffffff",
            INIT_1E => X"fffffff8ffffffffffffffe9ffffffffffffffd5ffffffffffffffecffffffff",
            INIT_1F => X"00000027000000000000000700000000fffffff2ffffffffffffffdaffffffff",
            INIT_20 => X"fffffffcffffffff000000050000000000000039000000000000001000000000",
            INIT_21 => X"fffffff7ffffffff000000030000000000000006000000000000002600000000",
            INIT_22 => X"0000000e00000000000000130000000000000013000000000000001000000000",
            INIT_23 => X"fffffffcfffffffffffffffcfffffffffffffff6ffffffff0000000d00000000",
            INIT_24 => X"ffffffb7ffffffffffffffe2ffffffffffffffb6ffffffffffffffeeffffffff",
            INIT_25 => X"0000000800000000fffffffeffffffffffffffcdfffffffffffffffaffffffff",
            INIT_26 => X"0000002000000000000000110000000000000032000000000000001000000000",
            INIT_27 => X"0000001800000000fffffffcffffffff0000000b000000000000001700000000",
            INIT_28 => X"0000001b0000000000000006000000000000000a00000000fffffff0ffffffff",
            INIT_29 => X"ffffffe2ffffffffffffffe8ffffffff00000010000000000000000800000000",
            INIT_2A => X"ffffffe4ffffffffffffffedffffffffffffffedfffffffffffffff8ffffffff",
            INIT_2B => X"fffffff2ffffffffffffffd3ffffffffffffffc6ffffffffffffffccffffffff",
            INIT_2C => X"0000000d00000000ffffffebffffffffffffffebffffffff0000000500000000",
            INIT_2D => X"ffffff74ffffffffffffffa5ffffffffffffffabffffffff0000000900000000",
            INIT_2E => X"ffffffbdffffffffffffffcfffffffffffffffaaffffffffffffffbdffffffff",
            INIT_2F => X"00000017000000000000000d000000000000003a000000000000001000000000",
            INIT_30 => X"fffffffbfffffffffffffff5fffffffffffffffafffffffffffffffcffffffff",
            INIT_31 => X"fffffff9ffffffff0000001300000000ffffffedfffffffffffffff4ffffffff",
            INIT_32 => X"ffffffc7ffffffffffffffdefffffffffffffff7fffffffffffffffcffffffff",
            INIT_33 => X"0000003600000000fffffff7fffffffffffffff6fffffffffffffff0ffffffff",
            INIT_34 => X"fffffffbffffffffffffffecffffffffffffffefffffffff0000000700000000",
            INIT_35 => X"fffffff9ffffffffffffffeffffffffffffffff4ffffffff0000000f00000000",
            INIT_36 => X"ffffffd5ffffffffffffffdaffffffffffffffeaffffffff0000000c00000000",
            INIT_37 => X"0000000000000000ffffffcbffffffffffffff99ffffffffffffffebffffffff",
            INIT_38 => X"ffffffccffffffffffffffc8ffffffff0000000000000000fffffffbffffffff",
            INIT_39 => X"ffffffeaffffffffffffffd3ffffffff0000000500000000ffffffc9ffffffff",
            INIT_3A => X"fffffff4ffffffff00000022000000000000002c000000000000000900000000",
            INIT_3B => X"0000001200000000ffffffe1ffffffff00000005000000000000001900000000",
            INIT_3C => X"0000003f000000000000001a00000000ffffffd7ffffffff0000001400000000",
            INIT_3D => X"fffffff1fffffffffffffff9fffffffffffffff3ffffffffffffffedffffffff",
            INIT_3E => X"ffffffdbffffffffffffffe3ffffffffffffffe9ffffffffffffffdeffffffff",
            INIT_3F => X"0000001600000000fffffff5ffffffff0000001900000000fffffff7ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000ffffffebfffffffffffffff9ffffffffffffffdcffffffff",
            INIT_41 => X"ffffffefffffffff0000003d000000000000002000000000ffffffd2ffffffff",
            INIT_42 => X"ffffffe9ffffffff0000000a0000000000000011000000000000000f00000000",
            INIT_43 => X"0000001e000000000000003000000000fffffff3fffffffffffffff9ffffffff",
            INIT_44 => X"0000000f0000000000000006000000000000000e000000000000001500000000",
            INIT_45 => X"fffffffcffffffff00000016000000000000000a000000000000000900000000",
            INIT_46 => X"ffffffffffffffffffffffeaffffffffffffffdaffffffffffffffd3ffffffff",
            INIT_47 => X"00000013000000000000001400000000ffffffb4ffffffffffffffc6ffffffff",
            INIT_48 => X"ffffffdaffffffffffffffd4ffffffffffffffaeffffffff0000004600000000",
            INIT_49 => X"fffffffcffffffffffffffccffffffffffffffc8ffffffffffffffccffffffff",
            INIT_4A => X"fffffffafffffffffffffff9ffffffff00000037000000000000002400000000",
            INIT_4B => X"0000000a000000000000000c000000000000000b000000000000000c00000000",
            INIT_4C => X"fffffff6ffffffffffffffcafffffffffffffffcffffffffffffffffffffffff",
            INIT_4D => X"00000001000000000000000100000000fffffff7ffffffff0000000800000000",
            INIT_4E => X"ffffffe8ffffffff00000024000000000000000f000000000000001000000000",
            INIT_4F => X"0000000000000000ffffffebffffffff0000000000000000ffffffffffffffff",
            INIT_50 => X"0000001b000000000000000c00000000fffffffbffffffff0000002700000000",
            INIT_51 => X"ffffffa1ffffffffffffffaaffffffffffffff8dffffffff0000002000000000",
            INIT_52 => X"ffffffffffffffffffffffcbffffffffffffffa0ffffffffffffffc6ffffffff",
            INIT_53 => X"fffffff0ffffffffffffffeaffffffff0000001d000000000000001800000000",
            INIT_54 => X"ffffffdaffffffff0000000e00000000fffffffaffffffffffffffeaffffffff",
            INIT_55 => X"0000002f000000000000002c00000000ffffffeefffffffffffffffcffffffff",
            INIT_56 => X"0000000a00000000000000000000000000000025000000000000001700000000",
            INIT_57 => X"0000001600000000ffffffe7ffffffffffffffeefffffffffffffffdffffffff",
            INIT_58 => X"fffffff0ffffffff0000001600000000ffffffebffffffff0000001500000000",
            INIT_59 => X"fffffffdffffffffffffffeafffffffffffffff7ffffffffffffffddffffffff",
            INIT_5A => X"00000019000000000000001600000000fffffffdfffffffffffffff9ffffffff",
            INIT_5B => X"00000006000000000000001500000000ffffffe8ffffffff0000000000000000",
            INIT_5C => X"ffffffd1ffffffffffffffcaffffffffffffffdfffffffff0000001b00000000",
            INIT_5D => X"00000026000000000000002300000000fffffff5ffffffffffffffc3ffffffff",
            INIT_5E => X"fffffff3ffffffff0000000300000000fffffff4fffffffffffffffbffffffff",
            INIT_5F => X"000000250000000000000019000000000000001e000000000000000500000000",
            INIT_60 => X"ffffffecfffffffffffffff7ffffffffffffffecffffffff0000001400000000",
            INIT_61 => X"0000001c00000000ffffffdfffffffffffffffecffffffffffffffd5ffffffff",
            INIT_62 => X"fffffff4fffffffffffffff7ffffffff00000014000000000000003700000000",
            INIT_63 => X"ffffff9effffffffffffffdfffffffffffffffe5fffffffffffffffeffffffff",
            INIT_64 => X"00000044000000000000000500000000ffffffffffffffff0000002a00000000",
            INIT_65 => X"ffffffe5ffffffffffffffdfffffffff00000045000000000000003900000000",
            INIT_66 => X"ffffffbfffffffffffffffecffffffffffffffd3ffffffffffffffdbffffffff",
            INIT_67 => X"0000003b00000000fffffffdffffffffffffffe6ffffffff0000000400000000",
            INIT_68 => X"0000000f00000000fffffff3ffffffff00000027000000000000000a00000000",
            INIT_69 => X"ffffffe8ffffffffffffffdcffffffffffffffe6fffffffffffffff2ffffffff",
            INIT_6A => X"ffffffd9ffffffff0000001900000000fffffffdfffffffffffffff0ffffffff",
            INIT_6B => X"fffffffaffffffffffffffe1ffffffffffffffe7fffffffffffffffdffffffff",
            INIT_6C => X"ffffff8affffffffffffff9affffffffffffffc5ffffffffffffffe8ffffffff",
            INIT_6D => X"0000003a000000000000000d0000000000000002000000000000001a00000000",
            INIT_6E => X"fffffffbffffffff000000100000000000000034000000000000001f00000000",
            INIT_6F => X"00000001000000000000001800000000fffffff3ffffffff0000002100000000",
            INIT_70 => X"fffffffbfffffffffffffffbffffffff0000000400000000ffffffd4ffffffff",
            INIT_71 => X"ffffffe8ffffffffffffffccffffffffffffffc4ffffffff0000001d00000000",
            INIT_72 => X"0000000d0000000000000007000000000000000000000000ffffffdbffffffff",
            INIT_73 => X"fffffff1ffffffffffffffbaffffffffffffffacffffffffffffffcaffffffff",
            INIT_74 => X"ffffffbdffffffffffffffe3ffffffffffffffe8ffffffff0000000100000000",
            INIT_75 => X"ffffffb2ffffffffffffffaeffffffffffffffd2ffffffffffffff9dffffffff",
            INIT_76 => X"0000001400000000ffffffdaffffffffffffffdcffffffff0000000c00000000",
            INIT_77 => X"fffffffdffffffff000000130000000000000034000000000000002b00000000",
            INIT_78 => X"00000006000000000000001700000000fffffff1ffffffff0000000000000000",
            INIT_79 => X"ffffffbbffffffff0000000000000000ffffffefffffffff0000000c00000000",
            INIT_7A => X"ffffffb6ffffffffffffffc5ffffffffffffffa0ffffffffffffff8cffffffff",
            INIT_7B => X"0000003d00000000ffffffe7ffffffff0000003800000000ffffff9cffffffff",
            INIT_7C => X"000000000000000000000020000000000000000b000000000000000800000000",
            INIT_7D => X"ffffffebffffffff0000000500000000fffffffaffffffff0000000900000000",
            INIT_7E => X"ffffffceffffffffffffffd2ffffffffffffffdaffffffff0000000000000000",
            INIT_7F => X"0000002a0000000000000005000000000000000000000000fffffffaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE18;


    MEM_IWGHT_LAYER2_INSTANCE19 : if BRAM_NAME = "iwght_layer2_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff93fffffffffffffff6ffffffff00000022000000000000000500000000",
            INIT_01 => X"000000350000000000000021000000000000000800000000ffffffc3ffffffff",
            INIT_02 => X"ffffffbeffffffff000000360000000000000012000000000000000200000000",
            INIT_03 => X"00000000000000000000001c00000000ffffffe4ffffffffffffffe8ffffffff",
            INIT_04 => X"fffffff7ffffffff0000003b0000000000000018000000000000000f00000000",
            INIT_05 => X"fffffff1ffffffff0000001a000000000000000d000000000000000a00000000",
            INIT_06 => X"0000001e000000000000001c00000000fffffff7fffffffffffffffbffffffff",
            INIT_07 => X"ffffffd5ffffffffffffffd3ffffffffffffffddffffffff0000000700000000",
            INIT_08 => X"0000001b00000000ffffffaaffffffffffffffb4ffffffffffffffcdffffffff",
            INIT_09 => X"ffffffc0ffffffffffffffd9ffffffff0000000500000000fffffff1ffffffff",
            INIT_0A => X"fffffffbfffffffffffffffdffffffffffffffd3ffffffffffffffbbffffffff",
            INIT_0B => X"000000090000000000000007000000000000000b000000000000000700000000",
            INIT_0C => X"0000002500000000000000290000000000000030000000000000000500000000",
            INIT_0D => X"ffffffcbffffffffffffffe4fffffffffffffff4ffffffff0000000e00000000",
            INIT_0E => X"ffffffe9fffffffffffffff3ffffffff00000007000000000000001500000000",
            INIT_0F => X"0000000b000000000000001200000000fffffff7ffffffffffffffdfffffffff",
            INIT_10 => X"ffffff9fffffffffffffffa7ffffffffffffffbdffffffff0000001800000000",
            INIT_11 => X"000000420000000000000004000000000000000400000000fffffff6ffffffff",
            INIT_12 => X"0000002f00000000000000140000000000000043000000000000002600000000",
            INIT_13 => X"00000004000000000000001000000000fffffffdffffffff0000002c00000000",
            INIT_14 => X"fffffffbffffffffffffffeeffffffff0000000e000000000000001700000000",
            INIT_15 => X"00000007000000000000001f00000000ffffffffffffffff0000002200000000",
            INIT_16 => X"ffffffe0fffffffffffffffeffffffff0000000d000000000000001f00000000",
            INIT_17 => X"0000002100000000000000030000000000000014000000000000000b00000000",
            INIT_18 => X"ffffffd2fffffffffffffff3ffffffff0000000b000000000000001b00000000",
            INIT_19 => X"ffffffb5ffffffffffffffcbffffffffffffff8bffffffffffffffc9ffffffff",
            INIT_1A => X"0000003e000000000000001b00000000ffffffeffffffffffffffff2ffffffff",
            INIT_1B => X"0000000e00000000fffffff8ffffffff0000001d000000000000002c00000000",
            INIT_1C => X"0000000000000000fffffffeffffffffffffffe8fffffffffffffffeffffffff",
            INIT_1D => X"0000003600000000000000130000000000000018000000000000001a00000000",
            INIT_1E => X"0000001500000000ffffffefffffffff0000001c000000000000001100000000",
            INIT_1F => X"0000000100000000ffffffefffffffff00000000000000000000000600000000",
            INIT_20 => X"fffffff8ffffffff00000005000000000000000b00000000fffffff9ffffffff",
            INIT_21 => X"00000000000000000000000b00000000ffffffd7ffffffff0000000100000000",
            INIT_22 => X"ffffffe3ffffffff000000070000000000000014000000000000000f00000000",
            INIT_23 => X"ffffffecffffffffffffffe6ffffffffffffffe0ffffffffffffffc7ffffffff",
            INIT_24 => X"ffffffd6ffffffffffffffbaffffffff00000018000000000000001f00000000",
            INIT_25 => X"0000001b000000000000001c000000000000001400000000ffffffbfffffffff",
            INIT_26 => X"fffffffcffffffff0000002c000000000000001f000000000000000e00000000",
            INIT_27 => X"00000007000000000000001300000000ffffffe3ffffffff0000001b00000000",
            INIT_28 => X"0000000b000000000000000d0000000000000018000000000000000b00000000",
            INIT_29 => X"0000000100000000fffffffbffffffffffffffdbffffffff0000002500000000",
            INIT_2A => X"ffffffd4fffffffffffffffbfffffffffffffff5fffffffffffffffeffffffff",
            INIT_2B => X"0000000c00000000ffffffffffffffff0000000600000000ffffffe5ffffffff",
            INIT_2C => X"ffffffc2ffffffff0000000300000000fffffff3ffffffff0000000e00000000",
            INIT_2D => X"00000002000000000000000600000000ffffffe5ffffffffffffffa0ffffffff",
            INIT_2E => X"0000000800000000000000160000000000000018000000000000001d00000000",
            INIT_2F => X"ffffffe6ffffffffffffffd5ffffffffffffffe4ffffffffffffffd3ffffffff",
            INIT_30 => X"0000003d000000000000002000000000ffffffffffffffff0000002000000000",
            INIT_31 => X"00000017000000000000001e0000000000000000000000000000001500000000",
            INIT_32 => X"ffffffcdffffffff0000000100000000ffffffefffffffff0000001000000000",
            INIT_33 => X"00000001000000000000002a00000000fffffff6ffffffffffffffa8ffffffff",
            INIT_34 => X"fffffff0ffffffffffffffe5ffffffff00000008000000000000003c00000000",
            INIT_35 => X"fffffff4ffffffffffffffffffffffff00000030000000000000000300000000",
            INIT_36 => X"fffffffafffffffffffffff2ffffffffffffffb5ffffffffffffffe1ffffffff",
            INIT_37 => X"ffffffd9ffffffff00000013000000000000001600000000ffffffe9ffffffff",
            INIT_38 => X"0000003200000000ffffffdeffffffff0000000000000000fffffffdffffffff",
            INIT_39 => X"ffffffe0fffffffffffffff2ffffffff0000003d000000000000005200000000",
            INIT_3A => X"fffffff4ffffffffffffffdbffffffffffffffc9ffffffffffffffe4ffffffff",
            INIT_3B => X"0000005300000000ffffffecffffffffffffffeeffffffffffffffcbffffffff",
            INIT_3C => X"0000000f00000000fffffff3ffffffff00000042000000000000005100000000",
            INIT_3D => X"ffffffffffffffffffffffd5ffffffff00000014000000000000000c00000000",
            INIT_3E => X"ffffffeffffffffffffffffeffffffffffffffe8ffffffff0000002000000000",
            INIT_3F => X"fffffffbfffffffffffffff5ffffffffffffffbbfffffffffffffff7ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c00000000fffffff7ffffffffffffffeeffffffff0000000200000000",
            INIT_41 => X"0000001f00000000ffffffeeffffffffffffffefffffffff0000000400000000",
            INIT_42 => X"0000003100000000fffffff2ffffffff0000002c000000000000002800000000",
            INIT_43 => X"00000028000000000000001f00000000fffffffaffffffff0000000a00000000",
            INIT_44 => X"fffffffbffffffff0000000c00000000ffffffb5ffffffffffffffeeffffffff",
            INIT_45 => X"00000009000000000000004800000000ffffffe3ffffffffffffffcaffffffff",
            INIT_46 => X"00000021000000000000001100000000ffffffe4ffffffff0000001300000000",
            INIT_47 => X"fffffff5ffffffff00000012000000000000002700000000ffffffdbffffffff",
            INIT_48 => X"0000001000000000ffffffdaffffffff00000000000000000000000b00000000",
            INIT_49 => X"000000010000000000000013000000000000001900000000fffffff9ffffffff",
            INIT_4A => X"fffffff9ffffffff0000002e000000000000002600000000ffffffe3ffffffff",
            INIT_4B => X"ffffffeaffffffffffffffe9ffffffff00000020000000000000003900000000",
            INIT_4C => X"0000001b00000000fffffff2fffffffffffffffcffffffffffffffedffffffff",
            INIT_4D => X"ffffffd3ffffffff0000000200000000fffffff6ffffffff0000003900000000",
            INIT_4E => X"ffffffeefffffffffffffff0ffffffffffffffeeffffffffffffffc8ffffffff",
            INIT_4F => X"0000000c000000000000001a00000000ffffffe6ffffffff0000000500000000",
            INIT_50 => X"0000000f00000000fffffff0ffffffffffffffdbffffffffffffffe9ffffffff",
            INIT_51 => X"0000007500000000000000170000000000000015000000000000003400000000",
            INIT_52 => X"00000036000000000000002800000000fffffff8ffffffff0000003900000000",
            INIT_53 => X"ffffffd2ffffffff0000000100000000fffffff4ffffffffffffffe7ffffffff",
            INIT_54 => X"00000014000000000000000a00000000ffffffdcffffffff0000001400000000",
            INIT_55 => X"00000006000000000000001a000000000000001a000000000000000400000000",
            INIT_56 => X"ffffffc1ffffffff00000039000000000000002c000000000000003800000000",
            INIT_57 => X"0000000d00000000fffffff8ffffffff0000000700000000fffffffcffffffff",
            INIT_58 => X"0000001200000000000000120000000000000006000000000000000100000000",
            INIT_59 => X"ffffffd1ffffffff0000000600000000ffffffeaffffffffffffffe3ffffffff",
            INIT_5A => X"0000001000000000ffffffeaffffffffffffffe2ffffffffffffffcaffffffff",
            INIT_5B => X"00000017000000000000001d000000000000000d00000000ffffffddffffffff",
            INIT_5C => X"0000000400000000ffffffd8ffffffff0000001200000000ffffffe5ffffffff",
            INIT_5D => X"0000000600000000fffffff6ffffffffffffffeaffffffff0000000b00000000",
            INIT_5E => X"ffffffe8ffffffff0000001400000000ffffffecffffffff0000002e00000000",
            INIT_5F => X"0000002300000000ffffffe9ffffffffffffffe7ffffffff0000002900000000",
            INIT_60 => X"ffffffe4ffffffff0000001900000000ffffffcfffffffffffffffc7ffffffff",
            INIT_61 => X"fffffff9fffffffffffffff2fffffffffffffffffffffffffffffff7ffffffff",
            INIT_62 => X"0000001e0000000000000033000000000000000100000000ffffffeeffffffff",
            INIT_63 => X"000000260000000000000039000000000000002a000000000000004c00000000",
            INIT_64 => X"ffffffdcffffffffffffffb4fffffffffffffff7ffffffff0000002900000000",
            INIT_65 => X"ffffffd8ffffffffffffffe6ffffffffffffffffffffffff0000002e00000000",
            INIT_66 => X"0000000d00000000ffffffdfffffffff0000000f000000000000002000000000",
            INIT_67 => X"ffffffe9fffffffffffffffdffffffffffffffdeffffffff0000000900000000",
            INIT_68 => X"0000002500000000ffffffe4ffffffff0000000000000000fffffff1ffffffff",
            INIT_69 => X"000000010000000000000004000000000000000a000000000000001f00000000",
            INIT_6A => X"ffffffcafffffffffffffff3fffffffffffffffdffffffff0000002200000000",
            INIT_6B => X"0000000700000000ffffffd7ffffffff00000011000000000000002100000000",
            INIT_6C => X"00000031000000000000005b000000000000000700000000fffffff0ffffffff",
            INIT_6D => X"0000001b00000000000000260000000000000015000000000000001a00000000",
            INIT_6E => X"0000003200000000ffffff6cffffffffffffff8fffffffffffffff8bffffffff",
            INIT_6F => X"ffffffdffffffffffffffffdffffffffffffffeeffffffff0000000600000000",
            INIT_70 => X"0000002d00000000ffffffd9ffffffffffffffceffffffff0000000400000000",
            INIT_71 => X"fffffffdffffffffffffffffffffffffffffffeaffffffff0000001400000000",
            INIT_72 => X"fffffff2ffffffff0000000100000000fffffff8ffffffff0000000400000000",
            INIT_73 => X"ffffffe3ffffffffffffffb7fffffffffffffff2ffffffff0000001900000000",
            INIT_74 => X"00000033000000000000000400000000ffffffe0fffffffffffffff1ffffffff",
            INIT_75 => X"0000001600000000000000270000000000000043000000000000001f00000000",
            INIT_76 => X"ffffffe9ffffffffffffffe3ffffffffffffffddffffffff0000001a00000000",
            INIT_77 => X"0000001900000000ffffffdcffffffffffffffdeffffffffffffffffffffffff",
            INIT_78 => X"fffffffdfffffffffffffffbffffffff0000000a00000000fffffff6ffffffff",
            INIT_79 => X"0000000400000000ffffffe9ffffffffffffffd2fffffffffffffffdffffffff",
            INIT_7A => X"0000000000000000fffffffeffffffff00000001000000000000001500000000",
            INIT_7B => X"ffffffefffffffffffffffedfffffffffffffff7ffffffff0000000600000000",
            INIT_7C => X"0000002300000000fffffffefffffffffffffffcfffffffffffffffcffffffff",
            INIT_7D => X"000000210000000000000010000000000000001700000000fffffff2ffffffff",
            INIT_7E => X"0000000e0000000000000000000000000000001b000000000000001d00000000",
            INIT_7F => X"0000000900000000ffffffe7fffffffffffffff0fffffffffffffffbffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE19;


    MEM_IWGHT_LAYER2_INSTANCE20 : if BRAM_NAME = "iwght_layer2_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001f00000000fffffff8ffffffffffffffe0ffffffffffffffb7ffffffff",
            INIT_01 => X"00000025000000000000001b0000000000000001000000000000000000000000",
            INIT_02 => X"ffffffe8ffffffff00000018000000000000001f00000000ffffffe7ffffffff",
            INIT_03 => X"ffffffe1ffffffff000000240000000000000038000000000000005700000000",
            INIT_04 => X"ffffffc5ffffffffffffffaeffffffffffffffdefffffffffffffff1ffffffff",
            INIT_05 => X"0000001c00000000ffffffe2ffffffffffffffefffffffffffffffa0ffffffff",
            INIT_06 => X"00000005000000000000001000000000ffffffe7fffffffffffffffdffffffff",
            INIT_07 => X"fffffffcffffffffffffffecffffffff00000017000000000000001d00000000",
            INIT_08 => X"0000000b00000000fffffff5fffffffffffffffafffffffffffffffaffffffff",
            INIT_09 => X"fffffff1fffffffffffffff0ffffffff00000005000000000000000d00000000",
            INIT_0A => X"0000000900000000fffffff2ffffffffffffffd2ffffffff0000000400000000",
            INIT_0B => X"ffffffefffffffff00000012000000000000001a00000000ffffffebffffffff",
            INIT_0C => X"0000001c000000000000001c000000000000000a000000000000000300000000",
            INIT_0D => X"0000000b00000000fffffff6ffffffff00000007000000000000001900000000",
            INIT_0E => X"ffffffbaffffffffffffffd5ffffffffffffffd6ffffffffffffffe1ffffffff",
            INIT_0F => X"ffffffe6fffffffffffffffaffffffff0000000e000000000000002e00000000",
            INIT_10 => X"ffffffe8fffffffffffffff8ffffffff0000001c00000000ffffffcbffffffff",
            INIT_11 => X"00000016000000000000002b0000000000000030000000000000001200000000",
            INIT_12 => X"ffffffdcffffffffffffffe3ffffffff0000001500000000ffffffe7ffffffff",
            INIT_13 => X"fffffff7fffffffffffffff5ffffffffffffffe3ffffffffffffffc7ffffffff",
            INIT_14 => X"fffffffbffffffff0000000e00000000fffffff0ffffffffffffffe1ffffffff",
            INIT_15 => X"0000001600000000ffffffe9ffffffffffffffe7ffffffffffffffd4ffffffff",
            INIT_16 => X"0000004400000000000000330000000000000033000000000000003100000000",
            INIT_17 => X"0000000d000000000000001600000000fffffff3ffffffff0000003300000000",
            INIT_18 => X"000000060000000000000000000000000000000900000000fffffffeffffffff",
            INIT_19 => X"ffffffecffffffff0000000900000000fffffffdffffffff0000000900000000",
            INIT_1A => X"ffffffc8ffffffff0000000e000000000000000100000000ffffffe8ffffffff",
            INIT_1B => X"ffffffe9ffffffffffffffb1ffffffff0000000400000000ffffffedffffffff",
            INIT_1C => X"000000130000000000000011000000000000003700000000fffffff7ffffffff",
            INIT_1D => X"ffffff8bffffffffffffffa5ffffffffffffff68ffffffff0000002400000000",
            INIT_1E => X"0000002700000000ffffffaeffffffffffffffbcffffffffffffff9effffffff",
            INIT_1F => X"00000020000000000000003600000000ffffffffffffffff0000002300000000",
            INIT_20 => X"ffffffd9ffffffffffffffefffffffff00000009000000000000001000000000",
            INIT_21 => X"0000000b00000000fffffffdffffffff00000012000000000000001600000000",
            INIT_22 => X"0000000a00000000000000180000000000000015000000000000000400000000",
            INIT_23 => X"0000000c00000000ffffffedffffffffffffffc8ffffffff0000000e00000000",
            INIT_24 => X"00000002000000000000000500000000fffffff9ffffffffffffffd8ffffffff",
            INIT_25 => X"0000000f00000000fffffff4ffffffff00000020000000000000001c00000000",
            INIT_26 => X"ffffffbbffffffffffffffa4ffffffffffffffc3ffffffff0000001200000000",
            INIT_27 => X"fffffff4fffffffffffffffbffffffffffffffeafffffffffffffffeffffffff",
            INIT_28 => X"ffffffccffffffffffffffe4fffffffffffffff0ffffffffffffffd9ffffffff",
            INIT_29 => X"00000020000000000000002e000000000000003f00000000ffffffffffffffff",
            INIT_2A => X"0000000000000000000000000000000000000014000000000000005300000000",
            INIT_2B => X"ffffffe0ffffffffffffffd5ffffffffffffffe3ffffffff0000000300000000",
            INIT_2C => X"0000000f0000000000000021000000000000001a00000000ffffffe6ffffffff",
            INIT_2D => X"0000001d00000000000000060000000000000030000000000000001700000000",
            INIT_2E => X"ffffffcdfffffffffffffff7ffffffff0000000f00000000fffffffeffffffff",
            INIT_2F => X"ffffffdeffffffffffffffcdffffffffffffffcffffffffffffffff1ffffffff",
            INIT_30 => X"ffffffecffffffff0000000500000000ffffffcfffffffffffffffcaffffffff",
            INIT_31 => X"ffffffc3fffffffffffffffbffffffffffffffe3ffffffffffffffeaffffffff",
            INIT_32 => X"00000013000000000000002e000000000000003b00000000ffffffcdffffffff",
            INIT_33 => X"ffffffa2ffffffff0000000a00000000ffffffd8ffffffffffffffe3ffffffff",
            INIT_34 => X"00000019000000000000003800000000ffffffc8ffffffffffffff9affffffff",
            INIT_35 => X"0000003400000000ffffffe5ffffffffffffffffffffffff0000001900000000",
            INIT_36 => X"fffffffcffffffff000000380000000000000003000000000000002100000000",
            INIT_37 => X"ffffffdbfffffffffffffffbfffffffffffffff8ffffffff0000000c00000000",
            INIT_38 => X"fffffffcffffffffffffffdcffffffffffffffb2ffffffffffffffe1ffffffff",
            INIT_39 => X"0000001300000000fffffffeffffffff00000000000000000000000b00000000",
            INIT_3A => X"fffffffeffffffffffffffe0ffffffff0000000000000000ffffffe2ffffffff",
            INIT_3B => X"0000000f00000000000000280000000000000001000000000000001900000000",
            INIT_3C => X"00000028000000000000001000000000fffffff4ffffffff0000000100000000",
            INIT_3D => X"0000002f000000000000001500000000fffffff9fffffffffffffff6ffffffff",
            INIT_3E => X"0000002e00000000fffffff9ffffffff00000007000000000000003f00000000",
            INIT_3F => X"ffffffffffffffff000000220000000000000004000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003300000000ffffffebffffffff00000019000000000000000200000000",
            INIT_41 => X"ffffffbbffffffffffffffcfffffffffffffff93ffffffff0000000000000000",
            INIT_42 => X"0000001f000000000000000e0000000000000008000000000000000c00000000",
            INIT_43 => X"ffffffecffffffffffffffe6fffffffffffffff2ffffffffffffffd2ffffffff",
            INIT_44 => X"000000290000000000000009000000000000000100000000ffffffebffffffff",
            INIT_45 => X"000000100000000000000017000000000000001400000000ffffffdaffffffff",
            INIT_46 => X"ffffffd6ffffffffffffffb9ffffffff0000002f000000000000002b00000000",
            INIT_47 => X"ffffffe4ffffffffffffffd2ffffffffffffffceffffffffffffffe2ffffffff",
            INIT_48 => X"0000001800000000ffffffd6ffffffffffffffd9ffffffffffffffe8ffffffff",
            INIT_49 => X"0000000b00000000fffffff1ffffffff0000003600000000fffffffcffffffff",
            INIT_4A => X"0000000700000000000000050000000000000024000000000000002f00000000",
            INIT_4B => X"000000000000000000000014000000000000001b000000000000000800000000",
            INIT_4C => X"fffffff8ffffffffffffffc5ffffffff0000000800000000ffffffdfffffffff",
            INIT_4D => X"ffffffdefffffffffffffff8fffffffffffffffcffffffff0000003e00000000",
            INIT_4E => X"0000001d00000000ffffffe8fffffffffffffffaffffffffffffffd4ffffffff",
            INIT_4F => X"fffffffaffffffff000000070000000000000002000000000000001b00000000",
            INIT_50 => X"fffffff6fffffffffffffff4fffffffffffffffbffffffff0000000000000000",
            INIT_51 => X"0000000700000000ffffffe7fffffffffffffffeffffffff0000001300000000",
            INIT_52 => X"0000001100000000000000080000000000000024000000000000000000000000",
            INIT_53 => X"ffffffe9ffffffff0000000700000000fffffffafffffffffffffff3ffffffff",
            INIT_54 => X"fffffffffffffffffffffff0ffffffff0000001e000000000000002100000000",
            INIT_55 => X"0000001700000000000000120000000000000028000000000000002600000000",
            INIT_56 => X"ffffffdfffffffff00000001000000000000002a000000000000000c00000000",
            INIT_57 => X"ffffffc7ffffffffffffffebffffffffffffffdbfffffffffffffff5ffffffff",
            INIT_58 => X"0000002d000000000000000800000000ffffffe5ffffffffffffffddffffffff",
            INIT_59 => X"fffffff7ffffffffffffffeeffffffffffffffd8ffffffff0000000d00000000",
            INIT_5A => X"00000002000000000000001700000000fffffff2fffffffffffffffdffffffff",
            INIT_5B => X"ffffffefffffffff000000160000000000000003000000000000000c00000000",
            INIT_5C => X"0000001700000000ffffffbfffffffffffffffe4ffffffff0000000d00000000",
            INIT_5D => X"0000000200000000ffffffe8ffffffff00000002000000000000000000000000",
            INIT_5E => X"00000011000000000000001900000000ffffffe1ffffffff0000000500000000",
            INIT_5F => X"0000003700000000000000160000000000000012000000000000000400000000",
            INIT_60 => X"000000100000000000000042000000000000000300000000fffffff9ffffffff",
            INIT_61 => X"00000004000000000000002800000000fffffff9ffffffff0000000400000000",
            INIT_62 => X"00000053000000000000002c0000000000000019000000000000000800000000",
            INIT_63 => X"fffffffaffffffff0000000000000000ffffffe6ffffffff0000003000000000",
            INIT_64 => X"ffffffcfffffffffffffffc6fffffffffffffffcffffffff0000000d00000000",
            INIT_65 => X"ffffffe6ffffffffffffffbafffffffffffffff3ffffffffffffffe1ffffffff",
            INIT_66 => X"ffffffdeffffffff0000000000000000ffffffe3ffffffff0000003c00000000",
            INIT_67 => X"0000000700000000fffffff6ffffffffffffffe3fffffffffffffffbffffffff",
            INIT_68 => X"fffffffbffffffffffffffe6fffffffffffffffeffffffff0000000b00000000",
            INIT_69 => X"00000029000000000000001700000000ffffffedffffffff0000001f00000000",
            INIT_6A => X"0000003e00000000000000040000000000000025000000000000000f00000000",
            INIT_6B => X"0000000300000000fffffffbfffffffffffffff7ffffffff0000004a00000000",
            INIT_6C => X"ffffffe6ffffffffffffffdfffffffff0000000500000000ffffffddffffffff",
            INIT_6D => X"ffffffb6ffffffffffffffb6ffffffff00000010000000000000000f00000000",
            INIT_6E => X"ffffffd1ffffffffffffffb8ffffffffffffffc3ffffffffffffffdaffffffff",
            INIT_6F => X"0000002a00000000fffffff7ffffffff0000003e000000000000001500000000",
            INIT_70 => X"000000100000000000000013000000000000000e000000000000003200000000",
            INIT_71 => X"ffffffdcfffffffffffffff0ffffffff0000000f000000000000001e00000000",
            INIT_72 => X"ffffffdfffffffffffffffe4ffffffffffffffd0ffffffffffffffe7ffffffff",
            INIT_73 => X"ffffffebffffffff0000000f000000000000001b00000000ffffffb7ffffffff",
            INIT_74 => X"ffffffdeffffffff0000002a00000000fffffff8fffffffffffffff0ffffffff",
            INIT_75 => X"0000001100000000fffffffeffffffff00000002000000000000001e00000000",
            INIT_76 => X"0000002e00000000ffffffd2ffffffff0000000d000000000000000f00000000",
            INIT_77 => X"fffffffcffffffffffffffeaffffffffffffffebffffffff0000001a00000000",
            INIT_78 => X"0000000600000000ffffffeaffffffff0000000500000000ffffffefffffffff",
            INIT_79 => X"0000000f000000000000001c00000000fffffff8ffffffffffffffebffffffff",
            INIT_7A => X"ffffffeefffffffffffffff2ffffffffffffffb4ffffffff0000001500000000",
            INIT_7B => X"00000048000000000000003800000000ffffffceffffffffffffffedffffffff",
            INIT_7C => X"0000000800000000ffffffe1ffffffff00000044000000000000003e00000000",
            INIT_7D => X"ffffffedffffffff00000003000000000000002c00000000ffffffeeffffffff",
            INIT_7E => X"0000001800000000000000230000000000000043000000000000004600000000",
            INIT_7F => X"0000002300000000000000200000000000000018000000000000000200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE20;


    MEM_IWGHT_LAYER2_INSTANCE21 : if BRAM_NAME = "iwght_layer2_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe1ffffffffffffff96ffffffffffffffd8ffffffffffffffe7ffffffff",
            INIT_01 => X"0000002500000000000000280000000000000030000000000000000c00000000",
            INIT_02 => X"ffffffe7ffffffffffffffdeffffffff00000016000000000000002a00000000",
            INIT_03 => X"0000001900000000fffffff2ffffffff0000001e000000000000001900000000",
            INIT_04 => X"0000001c00000000ffffffe8ffffffff0000001100000000ffffffffffffffff",
            INIT_05 => X"fffffffdffffffffffffffd7ffffffff00000007000000000000001d00000000",
            INIT_06 => X"ffffffe1fffffffffffffff2ffffffffffffffe7ffffffffffffffd6ffffffff",
            INIT_07 => X"0000000c00000000000000090000000000000030000000000000003300000000",
            INIT_08 => X"ffffffc3ffffffff0000001500000000fffffffbffffffffffffffe6ffffffff",
            INIT_09 => X"fffffff2ffffffffffffffd0ffffffff0000001800000000ffffffeaffffffff",
            INIT_0A => X"fffffff2ffffffff0000001500000000fffffff7ffffffff0000000500000000",
            INIT_0B => X"00000028000000000000000d00000000ffffffeaffffffff0000000100000000",
            INIT_0C => X"000000280000000000000028000000000000003f000000000000000400000000",
            INIT_0D => X"00000011000000000000002e0000000000000023000000000000002200000000",
            INIT_0E => X"ffffffffffffffff00000004000000000000000f000000000000002100000000",
            INIT_0F => X"00000034000000000000000700000000fffffff1ffffffff0000000a00000000",
            INIT_10 => X"ffffffbbffffffffffffffeaffffffffffffffc5fffffffffffffff6ffffffff",
            INIT_11 => X"ffffffd3ffffffff0000000000000000ffffffd0ffffffffffffffacffffffff",
            INIT_12 => X"0000002400000000fffffff0ffffffff0000001100000000ffffffe8ffffffff",
            INIT_13 => X"0000003a000000000000000000000000fffffff3ffffffff0000000200000000",
            INIT_14 => X"00000010000000000000000b000000000000001d000000000000001000000000",
            INIT_15 => X"00000000000000000000000e0000000000000035000000000000000500000000",
            INIT_16 => X"fffffffbffffffff0000000500000000fffffff5ffffffffffffffffffffffff",
            INIT_17 => X"0000000300000000fffffffaffffffff00000018000000000000000f00000000",
            INIT_18 => X"fffffff7fffffffffffffffcffffffff0000000a000000000000000d00000000",
            INIT_19 => X"fffffffaffffffff00000006000000000000000400000000ffffffefffffffff",
            INIT_1A => X"ffffffd8ffffffff0000000800000000ffffffd4ffffffffffffffdaffffffff",
            INIT_1B => X"0000003a0000000000000026000000000000004700000000ffffffd3ffffffff",
            INIT_1C => X"0000000c00000000000000130000000000000029000000000000000700000000",
            INIT_1D => X"00000042000000000000000b000000000000001a000000000000000800000000",
            INIT_1E => X"ffffffdfffffffff00000001000000000000000c000000000000001000000000",
            INIT_1F => X"ffffffe6ffffffffffffffdfffffffffffffffd7ffffffffffffffe6ffffffff",
            INIT_20 => X"ffffffb4ffffffffffffffd3ffffffff0000000200000000ffffffdeffffffff",
            INIT_21 => X"ffffffd9ffffffffffffffdaffffffffffffffcdffffffffffffffdfffffffff",
            INIT_22 => X"fffffff0fffffffffffffff8ffffffffffffffeaffffffff0000002100000000",
            INIT_23 => X"ffffffd8ffffffffffffffd2fffffffffffffffaffffffffffffffeaffffffff",
            INIT_24 => X"ffffffeafffffffffffffff6ffffffff00000016000000000000001600000000",
            INIT_25 => X"fffffff7ffffffff000000070000000000000017000000000000001500000000",
            INIT_26 => X"000000130000000000000000000000000000001e00000000fffffff8ffffffff",
            INIT_27 => X"ffffffe8fffffffffffffff0ffffffffffffffafffffffff0000002000000000",
            INIT_28 => X"0000004f000000000000002100000000ffffffe3fffffffffffffff4ffffffff",
            INIT_29 => X"fffffff1ffffffff00000018000000000000000a000000000000003e00000000",
            INIT_2A => X"0000001f00000000ffffffefffffffff0000000300000000fffffffaffffffff",
            INIT_2B => X"fffffffcffffffff00000026000000000000000d000000000000005500000000",
            INIT_2C => X"ffffffd5ffffffff0000001500000000ffffffecffffffffffffffcdffffffff",
            INIT_2D => X"ffffffd8fffffffffffffff7ffffffff00000019000000000000001100000000",
            INIT_2E => X"0000000000000000fffffff7fffffffffffffff7ffffffff0000002300000000",
            INIT_2F => X"00000004000000000000002f00000000ffffffe7ffffffff0000000800000000",
            INIT_30 => X"0000000a00000000000000220000000000000023000000000000002600000000",
            INIT_31 => X"0000001500000000000000090000000000000002000000000000003800000000",
            INIT_32 => X"ffffffc3fffffffffffffff3ffffffff00000009000000000000000b00000000",
            INIT_33 => X"ffffffebffffffffffffffd5ffffffff00000019000000000000000d00000000",
            INIT_34 => X"fffffff7ffffffff0000001e00000000fffffff6ffffffff0000000f00000000",
            INIT_35 => X"ffffffebffffffff0000003700000000ffffffe9ffffffffffffffd1ffffffff",
            INIT_36 => X"ffffffc9fffffffffffffff3fffffffffffffff1fffffffffffffff6ffffffff",
            INIT_37 => X"ffffffd7ffffffff00000024000000000000004d000000000000000c00000000",
            INIT_38 => X"0000001e00000000ffffffedffffffff00000003000000000000001700000000",
            INIT_39 => X"ffffffd6ffffffffffffffefffffffffffffffe2ffffffff0000001000000000",
            INIT_3A => X"0000002200000000ffffffe5ffffffffffffffceffffffffffffffe5ffffffff",
            INIT_3B => X"0000003e000000000000002d0000000000000023000000000000000e00000000",
            INIT_3C => X"000000090000000000000036000000000000000c00000000ffffffffffffffff",
            INIT_3D => X"00000015000000000000000d0000000000000019000000000000001700000000",
            INIT_3E => X"ffffffc0fffffffffffffff5fffffffffffffff1ffffffffffffffefffffffff",
            INIT_3F => X"000000150000000000000001000000000000000d00000000fffffff4ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdcfffffffffffffff9fffffffffffffff0ffffffffffffffe7ffffffff",
            INIT_41 => X"fffffff6fffffffffffffff1ffffffffffffffdefffffffffffffff7ffffffff",
            INIT_42 => X"0000000600000000000000180000000000000006000000000000000300000000",
            INIT_43 => X"fffffffaffffffffffffffe7ffffffffffffffe2ffffffff0000000d00000000",
            INIT_44 => X"0000000f00000000fffffff8ffffffff0000000200000000fffffff9ffffffff",
            INIT_45 => X"ffffffe6fffffffffffffff7ffffffffffffffe6ffffffff0000001100000000",
            INIT_46 => X"0000000100000000000000070000000000000002000000000000001600000000",
            INIT_47 => X"fffffff6fffffffffffffff2ffffffff0000000f000000000000000900000000",
            INIT_48 => X"fffffffdffffffffffffffe5ffffffff0000001800000000ffffffe9ffffffff",
            INIT_49 => X"ffffffe6fffffffffffffff8ffffffffffffffecfffffffffffffff8ffffffff",
            INIT_4A => X"fffffff1ffffffffffffffe9fffffffffffffffdffffffffffffffddffffffff",
            INIT_4B => X"fffffff4fffffffffffffff4ffffffffffffffdcffffffffffffffefffffffff",
            INIT_4C => X"ffffffeaffffffffffffffefffffffff0000000100000000ffffffdaffffffff",
            INIT_4D => X"fffffff5ffffffff0000001800000000ffffffedffffffffffffffe1ffffffff",
            INIT_4E => X"0000000500000000fffffffdfffffffffffffffbfffffffffffffff4ffffffff",
            INIT_4F => X"ffffffefffffffff0000000a00000000ffffffe5fffffffffffffffcffffffff",
            INIT_50 => X"fffffff3ffffffff00000000000000000000000700000000fffffff5ffffffff",
            INIT_51 => X"000000090000000000000004000000000000000b000000000000000c00000000",
            INIT_52 => X"fffffffbfffffffffffffffeffffffff0000000900000000fffffffbffffffff",
            INIT_53 => X"fffffff9ffffffff0000000900000000ffffffe6fffffffffffffff3ffffffff",
            INIT_54 => X"ffffffd4ffffffffffffffecffffffffffffffd1ffffffff0000000300000000",
            INIT_55 => X"0000000400000000ffffffcbffffffffffffffebfffffffffffffffeffffffff",
            INIT_56 => X"0000000800000000fffffff9ffffffffffffffd0ffffffffffffffdcffffffff",
            INIT_57 => X"fffffffeffffffffffffffdffffffffffffffff0ffffffffffffffe4ffffffff",
            INIT_58 => X"fffffff0ffffffffffffffeefffffffffffffffafffffffffffffffaffffffff",
            INIT_59 => X"fffffff8ffffffff0000000d00000000fffffff6ffffffff0000000500000000",
            INIT_5A => X"fffffff9fffffffffffffff5ffffffffffffffe8ffffffff0000000000000000",
            INIT_5B => X"ffffffffffffffff0000000b00000000fffffff8fffffffffffffffbffffffff",
            INIT_5C => X"00000008000000000000001000000000fffffff5fffffffffffffff0ffffffff",
            INIT_5D => X"ffffffdafffffffffffffff8ffffffffffffffebffffffffffffffdfffffffff",
            INIT_5E => X"0000000a00000000ffffffebffffffffffffffe5ffffffffffffffeeffffffff",
            INIT_5F => X"fffffff8fffffffffffffffbffffffffffffffe6ffffffffffffffdcffffffff",
            INIT_60 => X"fffffff1fffffffffffffff2ffffffffffffffffffffffff0000000e00000000",
            INIT_61 => X"ffffffd8fffffffffffffff3ffffffff00000001000000000000000a00000000",
            INIT_62 => X"ffffffe3ffffffffffffffe8ffffffffffffffe5fffffffffffffff8ffffffff",
            INIT_63 => X"ffffffdbffffffffffffffdeffffffffffffffe0fffffffffffffff1ffffffff",
            INIT_64 => X"ffffffe9fffffffffffffffbfffffffffffffffcffffffff0000000400000000",
            INIT_65 => X"0000000e00000000fffffffdffffffff0000000900000000fffffff9ffffffff",
            INIT_66 => X"0000000400000000ffffffecffffffffffffffdbffffffffffffffffffffffff",
            INIT_67 => X"000000080000000000000010000000000000000a00000000ffffffe8ffffffff",
            INIT_68 => X"ffffffefffffffffffffffecffffffffffffffeaffffffff0000001500000000",
            INIT_69 => X"fffffffbffffffffffffffeeffffffff0000000d00000000fffffff7ffffffff",
            INIT_6A => X"fffffff4ffffffff0000000700000000ffffffddfffffffffffffff6ffffffff",
            INIT_6B => X"fffffffbffffffff0000001300000000fffffffaffffffffffffffd4ffffffff",
            INIT_6C => X"fffffff2ffffffff0000000a0000000000000012000000000000000b00000000",
            INIT_6D => X"ffffffdaffffffff0000000500000000ffffffe6ffffffffffffffe4ffffffff",
            INIT_6E => X"fffffffbfffffffffffffffcffffffff0000000300000000ffffffffffffffff",
            INIT_6F => X"fffffff8ffffffffffffffecffffffff00000003000000000000000200000000",
            INIT_70 => X"ffffffffffffffff0000000f0000000000000000000000000000000e00000000",
            INIT_71 => X"ffffffe9ffffffffffffffdbfffffffffffffff7ffffffffffffffe9ffffffff",
            INIT_72 => X"fffffff6ffffffffffffffffffffffffffffffeaffffffffffffffe9ffffffff",
            INIT_73 => X"ffffffe1fffffffffffffffcfffffffffffffff6ffffffffffffffdfffffffff",
            INIT_74 => X"ffffffe9ffffffffffffffd5ffffffff0000001f000000000000000400000000",
            INIT_75 => X"fffffffeffffffff0000000000000000ffffffe6ffffffff0000000400000000",
            INIT_76 => X"ffffffdfffffffff0000000f000000000000000300000000fffffff0ffffffff",
            INIT_77 => X"0000001500000000ffffffdbffffffff00000013000000000000001100000000",
            INIT_78 => X"ffffffe6ffffffffffffffebffffffffffffffe7ffffffff0000001200000000",
            INIT_79 => X"ffffffd6ffffffff0000001400000000fffffff7ffffffffffffffe4ffffffff",
            INIT_7A => X"ffffffebffffffffffffffeeffffffff0000000000000000ffffffecffffffff",
            INIT_7B => X"fffffff0fffffffffffffff2ffffffffffffffdfffffffff0000000900000000",
            INIT_7C => X"fffffff9fffffffffffffff3ffffffff0000000c000000000000000600000000",
            INIT_7D => X"ffffffc0ffffffffffffffe5fffffffffffffffefffffffffffffff2ffffffff",
            INIT_7E => X"ffffffd6ffffffffffffffe4ffffffffffffffdeffffffff0000001b00000000",
            INIT_7F => X"0000001400000000000000010000000000000003000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE21;


    MEM_IWGHT_LAYER2_INSTANCE22 : if BRAM_NAME = "iwght_layer2_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe3ffffffff0000001400000000ffffffddffffffffffffffe0ffffffff",
            INIT_01 => X"0000000600000000ffffffe8ffffffffffffffe7fffffffffffffff8ffffffff",
            INIT_02 => X"ffffffffffffffff0000000b00000000fffffff5ffffffffffffffe1ffffffff",
            INIT_03 => X"0000000000000000ffffffecfffffffffffffffbffffffff0000000100000000",
            INIT_04 => X"fffffff8ffffffff00000001000000000000000100000000ffffffdeffffffff",
            INIT_05 => X"000000030000000000000006000000000000000800000000fffffffeffffffff",
            INIT_06 => X"fffffff9ffffffff0000000f00000000ffffffe3ffffffffffffffe2ffffffff",
            INIT_07 => X"0000000600000000fffffffaffffffff0000000600000000ffffffe3ffffffff",
            INIT_08 => X"ffffffedffffffff000000090000000000000000000000000000000900000000",
            INIT_09 => X"0000000300000000000000050000000000000007000000000000000e00000000",
            INIT_0A => X"fffffff6ffffffff000000000000000000000008000000000000000200000000",
            INIT_0B => X"fffffffbfffffffffffffff8ffffffff00000005000000000000000e00000000",
            INIT_0C => X"fffffff6ffffffff0000000b000000000000000000000000fffffff7ffffffff",
            INIT_0D => X"ffffffe7fffffffffffffff2fffffffffffffffbffffffff0000000900000000",
            INIT_0E => X"ffffffedffffffff0000000200000000ffffffeaffffffffffffffedffffffff",
            INIT_0F => X"ffffffe8fffffffffffffff1ffffffff0000000a00000000fffffff7ffffffff",
            INIT_10 => X"ffffffeeffffffffffffffe8ffffffff0000000c00000000ffffffebffffffff",
            INIT_11 => X"fffffff1ffffffff00000009000000000000000400000000fffffffdffffffff",
            INIT_12 => X"000000140000000000000003000000000000000700000000ffffffffffffffff",
            INIT_13 => X"00000006000000000000000d00000000fffffff7ffffffff0000000600000000",
            INIT_14 => X"ffffffeafffffffffffffffaffffffff0000000000000000fffffff1ffffffff",
            INIT_15 => X"fffffffbffffffff00000004000000000000000000000000fffffff8ffffffff",
            INIT_16 => X"fffffff7fffffffffffffffefffffffffffffff7ffffffff0000000400000000",
            INIT_17 => X"ffffffe6ffffffff0000000b00000000fffffff3ffffffff0000000500000000",
            INIT_18 => X"00000001000000000000000200000000fffffffbffffffff0000000d00000000",
            INIT_19 => X"0000000a000000000000000300000000fffffff6ffffffff0000000800000000",
            INIT_1A => X"fffffff7fffffffffffffffdffffffffffffffedfffffffffffffff9ffffffff",
            INIT_1B => X"ffffffe9ffffffff0000000800000000ffffffeaffffffff0000000600000000",
            INIT_1C => X"fffffff9ffffffffffffffe2fffffffffffffff8fffffffffffffffeffffffff",
            INIT_1D => X"fffffff9fffffffffffffffaffffffff00000000000000000000000400000000",
            INIT_1E => X"ffffffe8ffffffff0000000300000000fffffff2ffffffff0000000000000000",
            INIT_1F => X"0000000800000000ffffffeeffffffff0000000b00000000ffffffe8ffffffff",
            INIT_20 => X"fffffff7fffffffffffffffeffffffffffffffeeffffffffffffffecffffffff",
            INIT_21 => X"00000009000000000000000700000000fffffff3ffffffffffffffedffffffff",
            INIT_22 => X"ffffffefffffffffffffffebfffffffffffffff6ffffffffffffffeeffffffff",
            INIT_23 => X"fffffff4ffffffffffffffe4ffffffff0000000800000000ffffffedffffffff",
            INIT_24 => X"0000000f000000000000000000000000fffffff6ffffffffffffffe8ffffffff",
            INIT_25 => X"0000001000000000ffffffffffffffff0000000e000000000000000600000000",
            INIT_26 => X"fffffff0fffffffffffffff1ffffffffffffffebfffffffffffffffaffffffff",
            INIT_27 => X"0000000600000000fffffff4ffffffff00000001000000000000000400000000",
            INIT_28 => X"00000011000000000000000a000000000000000400000000fffffff2ffffffff",
            INIT_29 => X"fffffff2fffffffffffffff6fffffffffffffff0ffffffff0000001100000000",
            INIT_2A => X"ffffffebffffffff0000000000000000ffffffffffffffff0000000700000000",
            INIT_2B => X"fffffffbffffffff00000006000000000000000d000000000000000400000000",
            INIT_2C => X"fffffff8fffffffffffffffffffffffffffffff1ffffffff0000000700000000",
            INIT_2D => X"00000010000000000000000f00000000fffffffafffffffffffffff0ffffffff",
            INIT_2E => X"0000000f00000000fffffff1ffffffffffffffefffffffff0000000200000000",
            INIT_2F => X"fffffff1fffffffffffffffbfffffffffffffff0ffffffff0000001400000000",
            INIT_30 => X"ffffffe7ffffffff0000000000000000ffffffedffffffff0000001000000000",
            INIT_31 => X"ffffffeeffffffff0000000900000000ffffffecffffffff0000000800000000",
            INIT_32 => X"fffffff1ffffffff0000000900000000ffffffebfffffffffffffff3ffffffff",
            INIT_33 => X"fffffffbfffffffffffffff6ffffffff0000001500000000fffffff6ffffffff",
            INIT_34 => X"0000001200000000fffffff8fffffffffffffff2ffffffff0000000a00000000",
            INIT_35 => X"0000000500000000fffffff0ffffffffffffffe8fffffffffffffff7ffffffff",
            INIT_36 => X"fffffffcffffffff0000000100000000fffffff5fffffffffffffff6ffffffff",
            INIT_37 => X"fffffffeffffffffffffffedffffffff0000000000000000fffffff2ffffffff",
            INIT_38 => X"fffffff8fffffffffffffff3ffffffffffffffe3ffffffffffffffe6ffffffff",
            INIT_39 => X"ffffffefffffffff0000001300000000fffffffcffffffffffffffffffffffff",
            INIT_3A => X"fffffff0ffffffffffffffebfffffffffffffff8ffffffff0000000b00000000",
            INIT_3B => X"fffffff1ffffffff00000005000000000000000e000000000000000e00000000",
            INIT_3C => X"fffffff1ffffffff00000005000000000000000000000000fffffff2ffffffff",
            INIT_3D => X"000000120000000000000001000000000000000c00000000fffffff3ffffffff",
            INIT_3E => X"ffffffeffffffffffffffff8ffffffffffffffe2ffffffff0000000d00000000",
            INIT_3F => X"fffffff4ffffffffffffffe2fffffffffffffff0ffffffffffffffffffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffafffffffffffffff0fffffffffffffff3ffffffff0000000400000000",
            INIT_41 => X"fffffffdffffffffffffffeeffffffff00000000000000000000000e00000000",
            INIT_42 => X"0000000900000000fffffff8fffffffffffffff7ffffffffffffffffffffffff",
            INIT_43 => X"ffffffeafffffffffffffffaffffffff0000000a000000000000000700000000",
            INIT_44 => X"ffffffeefffffffffffffffefffffffffffffff7fffffffffffffffcffffffff",
            INIT_45 => X"ffffffebffffffffffffffeaffffffff0000000e000000000000000200000000",
            INIT_46 => X"fffffff4ffffffff0000000c00000000fffffff1ffffffff0000000900000000",
            INIT_47 => X"fffffffcffffffff0000000700000000ffffffebffffffffffffffeeffffffff",
            INIT_48 => X"ffffffe6fffffffffffffff9ffffffffffffffeafffffffffffffff8ffffffff",
            INIT_49 => X"fffffffaffffffff0000000e00000000ffffffecffffffffffffffe9ffffffff",
            INIT_4A => X"0000000c00000000fffffffafffffffffffffffefffffffffffffff2ffffffff",
            INIT_4B => X"fffffff9fffffffffffffff6fffffffffffffffaffffffff0000000300000000",
            INIT_4C => X"ffffffebffffffff000000000000000000000006000000000000000100000000",
            INIT_4D => X"ffffffe3fffffffffffffff0fffffffffffffff3fffffffffffffffdffffffff",
            INIT_4E => X"fffffff9ffffffff000000050000000000000003000000000000000b00000000",
            INIT_4F => X"00000008000000000000000b00000000fffffff7ffffffff0000000300000000",
            INIT_50 => X"ffffffd6ffffffffffffffdfffffffffffffffadffffffffffffffb9ffffffff",
            INIT_51 => X"00000020000000000000000900000000fffffff4ffffffffffffffd7ffffffff",
            INIT_52 => X"0000002b000000000000001f000000000000002000000000ffffffecffffffff",
            INIT_53 => X"00000023000000000000002b0000000000000037000000000000002300000000",
            INIT_54 => X"fffffff9ffffffffffffffc7ffffffff00000001000000000000000500000000",
            INIT_55 => X"ffffffe3ffffffffffffffffffffffff00000003000000000000000900000000",
            INIT_56 => X"ffffffe7ffffffffffffffefffffffffffffffefffffffffffffffe8ffffffff",
            INIT_57 => X"0000002d00000000fffffff3ffffffff00000007000000000000001c00000000",
            INIT_58 => X"0000000f0000000000000015000000000000000400000000ffffffc7ffffffff",
            INIT_59 => X"fffffff8fffffffffffffff1ffffffff00000013000000000000000700000000",
            INIT_5A => X"0000001500000000ffffffdfffffffffffffffefffffffff0000001c00000000",
            INIT_5B => X"0000000d0000000000000029000000000000000d00000000ffffffd9ffffffff",
            INIT_5C => X"fffffff9ffffffffffffffd3ffffffff00000021000000000000001a00000000",
            INIT_5D => X"fffffffdffffffffffffffe2ffffffffffffffccffffffffffffffe0ffffffff",
            INIT_5E => X"ffffffd1ffffffffffffffe1fffffffffffffffbffffffffffffffd2ffffffff",
            INIT_5F => X"ffffffe1ffffffffffffffc8ffffffffffffffe8ffffffff0000000e00000000",
            INIT_60 => X"fffffff7fffffffffffffff6ffffffffffffffe1ffffffffffffffcfffffffff",
            INIT_61 => X"0000001200000000ffffffffffffffff00000021000000000000000b00000000",
            INIT_62 => X"ffffffe7ffffffffffffffd7fffffffffffffffbffffffffffffffd8ffffffff",
            INIT_63 => X"0000000c00000000fffffff3ffffffffffffffcdffffffffffffffe8ffffffff",
            INIT_64 => X"0000000b000000000000001c000000000000002500000000ffffffe5ffffffff",
            INIT_65 => X"00000011000000000000001900000000ffffffe5ffffffff0000000000000000",
            INIT_66 => X"ffffffbeffffffffffffffd0ffffffff0000001200000000ffffffd2ffffffff",
            INIT_67 => X"fffffffcffffffff0000000c00000000fffffff5ffffffffffffffe6ffffffff",
            INIT_68 => X"ffffffd1fffffffffffffff3ffffffff0000001400000000ffffffebffffffff",
            INIT_69 => X"ffffffecffffffffffffffe3ffffffff0000002400000000ffffffecffffffff",
            INIT_6A => X"ffffffe0ffffffffffffffe3ffffffffffffffeaffffffffffffffcfffffffff",
            INIT_6B => X"0000001200000000ffffffd9fffffffffffffff8ffffffffffffffe3ffffffff",
            INIT_6C => X"fffffffbffffffff0000001e00000000ffffffe4ffffffff0000000900000000",
            INIT_6D => X"0000000800000000ffffffddffffffff0000002f000000000000001b00000000",
            INIT_6E => X"ffffffedffffffff0000003400000000ffffffedffffffff0000000c00000000",
            INIT_6F => X"00000006000000000000000f0000000000000006000000000000000c00000000",
            INIT_70 => X"000000060000000000000004000000000000000c00000000fffffff9ffffffff",
            INIT_71 => X"ffffffd4fffffffffffffffbfffffffffffffffcfffffffffffffff9ffffffff",
            INIT_72 => X"ffffffdbffffffff0000002300000000fffffff5fffffffffffffff0ffffffff",
            INIT_73 => X"ffffffe2ffffffffffffffcaffffffff0000000a000000000000002400000000",
            INIT_74 => X"ffffffe5ffffffff0000000400000000fffffffbffffffff0000000000000000",
            INIT_75 => X"ffffffdeffffffff00000004000000000000000800000000ffffffd0ffffffff",
            INIT_76 => X"00000033000000000000001b0000000000000026000000000000002f00000000",
            INIT_77 => X"0000001500000000fffffffbfffffffffffffffdffffffff0000000200000000",
            INIT_78 => X"0000002f000000000000001a000000000000002000000000ffffffdfffffffff",
            INIT_79 => X"0000002200000000000000300000000000000004000000000000001700000000",
            INIT_7A => X"ffffffd2fffffffffffffffefffffffffffffff1ffffffff0000000a00000000",
            INIT_7B => X"0000001000000000ffffffd6ffffffff0000002000000000fffffff8ffffffff",
            INIT_7C => X"0000000e000000000000000000000000fffffff2ffffffff0000004c00000000",
            INIT_7D => X"0000001000000000fffffff0ffffffff0000001e000000000000001b00000000",
            INIT_7E => X"fffffff7ffffffff0000000800000000ffffffd8ffffffffffffffddffffffff",
            INIT_7F => X"0000000c00000000ffffffa0ffffffffffffffb8fffffffffffffff2ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE22;


    MEM_IWGHT_LAYER2_INSTANCE23 : if BRAM_NAME = "iwght_layer2_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000a000000000000000c00000000ffffffeafffffffffffffffaffffffff",
            INIT_01 => X"ffffffc3ffffffff0000000d00000000ffffffc9ffffffffffffffe8ffffffff",
            INIT_02 => X"ffffffd1ffffffffffffffccffffffffffffffcbffffffff0000000c00000000",
            INIT_03 => X"fffffff2ffffffff0000000100000000ffffffe9ffffffffffffffd1ffffffff",
            INIT_04 => X"ffffffe5fffffffffffffff2ffffffff0000000000000000ffffffd5ffffffff",
            INIT_05 => X"0000000d00000000000000090000000000000038000000000000000500000000",
            INIT_06 => X"0000000a00000000000000170000000000000000000000000000003a00000000",
            INIT_07 => X"ffffffe8ffffffff0000001a000000000000003800000000ffffffeaffffffff",
            INIT_08 => X"0000001b000000000000001b00000000fffffff9ffffffff0000002500000000",
            INIT_09 => X"ffffffe4fffffffffffffff0ffffffff0000000d000000000000000100000000",
            INIT_0A => X"fffffff6ffffffff0000000100000000fffffffcffffffff0000001200000000",
            INIT_0B => X"000000060000000000000006000000000000000a00000000ffffffe6ffffffff",
            INIT_0C => X"0000000800000000000000240000000000000006000000000000004d00000000",
            INIT_0D => X"0000001300000000fffffffdfffffffffffffff9ffffffffffffffedffffffff",
            INIT_0E => X"00000011000000000000000e0000000000000023000000000000000f00000000",
            INIT_0F => X"0000000000000000fffffff4ffffffff0000001600000000ffffffd1ffffffff",
            INIT_10 => X"ffffffe9fffffffffffffffbffffffffffffffe5ffffffff0000001900000000",
            INIT_11 => X"00000021000000000000002b00000000ffffffe5fffffffffffffff1ffffffff",
            INIT_12 => X"000000070000000000000001000000000000003f000000000000000400000000",
            INIT_13 => X"00000001000000000000000b00000000ffffffffffffffff0000000c00000000",
            INIT_14 => X"0000001100000000fffffffbffffffffffffffeaffffffff0000002000000000",
            INIT_15 => X"fffffff9ffffffff0000002500000000fffffff4fffffffffffffffcffffffff",
            INIT_16 => X"00000005000000000000000600000000ffffffe1ffffffffffffffacffffffff",
            INIT_17 => X"000000090000000000000015000000000000000e00000000fffffff1ffffffff",
            INIT_18 => X"ffffffe9ffffffff0000001a000000000000002400000000ffffffe9ffffffff",
            INIT_19 => X"fffffff8ffffffffffffffebfffffffffffffff6fffffffffffffff6ffffffff",
            INIT_1A => X"ffffffdaffffffff00000007000000000000001400000000fffffff6ffffffff",
            INIT_1B => X"00000046000000000000001600000000ffffffe9ffffffff0000004b00000000",
            INIT_1C => X"ffffffd5ffffffffffffffdffffffffffffffff7fffffffffffffff6ffffffff",
            INIT_1D => X"ffffffecffffffffffffffdefffffffffffffffdffffffffffffffeaffffffff",
            INIT_1E => X"0000001c00000000ffffff82ffffffffffffffacffffffffffffffcbffffffff",
            INIT_1F => X"0000001a000000000000002500000000ffffffc7ffffffff0000001b00000000",
            INIT_20 => X"ffffffc2ffffffff0000003800000000ffffffffffffffffffffffc4ffffffff",
            INIT_21 => X"0000001800000000fffffff5ffffffff00000042000000000000000d00000000",
            INIT_22 => X"00000041000000000000000c00000000ffffffeaffffffff0000002a00000000",
            INIT_23 => X"ffffffddffffffff00000022000000000000000800000000ffffffe6ffffffff",
            INIT_24 => X"0000001200000000ffffffd5ffffffff0000002b000000000000001200000000",
            INIT_25 => X"00000035000000000000001b00000000ffffffe1ffffffff0000002a00000000",
            INIT_26 => X"ffffffdcffffffff0000000400000000ffffffe7fffffffffffffff1ffffffff",
            INIT_27 => X"ffffffe6ffffffffffffffbcffffffff0000000200000000ffffffebffffffff",
            INIT_28 => X"0000001200000000ffffffedffffffff00000005000000000000001a00000000",
            INIT_29 => X"fffffff2ffffffff0000001500000000ffffffefffffffff0000000f00000000",
            INIT_2A => X"0000000000000000ffffffd8ffffffff00000010000000000000001a00000000",
            INIT_2B => X"00000027000000000000001c00000000ffffffc6ffffffff0000000b00000000",
            INIT_2C => X"0000001700000000fffffff3ffffffffffffffe6fffffffffffffff6ffffffff",
            INIT_2D => X"ffffffefffffffff0000002400000000ffffffccfffffffffffffffaffffffff",
            INIT_2E => X"0000002900000000fffffff8ffffffff0000001600000000ffffffe0ffffffff",
            INIT_2F => X"0000001300000000fffffffaffffffff00000012000000000000000d00000000",
            INIT_30 => X"0000004000000000ffffffdffffffffffffffff6ffffffffffffffc6ffffffff",
            INIT_31 => X"ffffffe9ffffffffffffffffffffffff0000000a000000000000002700000000",
            INIT_32 => X"ffffffc8ffffffffffffffcdffffffffffffffd4ffffffffffffffd9ffffffff",
            INIT_33 => X"ffffffe2fffffffffffffff2ffffffffffffffe8fffffffffffffff4ffffffff",
            INIT_34 => X"ffffffd3ffffffffffffffc5fffffffffffffff7ffffffffffffffdcffffffff",
            INIT_35 => X"00000036000000000000004e00000000fffffff9ffffffffffffffceffffffff",
            INIT_36 => X"0000000a000000000000003000000000fffffffeffffffff0000000600000000",
            INIT_37 => X"00000011000000000000000e000000000000004300000000ffffffecffffffff",
            INIT_38 => X"00000014000000000000000d00000000fffffffcfffffffffffffffaffffffff",
            INIT_39 => X"0000001000000000fffffffbffffffff0000000a000000000000000700000000",
            INIT_3A => X"ffffffc9ffffffff000000070000000000000035000000000000000a00000000",
            INIT_3B => X"fffffff7fffffffffffffff4ffffffff0000000c000000000000000300000000",
            INIT_3C => X"ffffffffffffffff0000003f00000000ffffffcdfffffffffffffff3ffffffff",
            INIT_3D => X"0000000400000000fffffff3ffffffff0000003900000000ffffffcfffffffff",
            INIT_3E => X"fffffff8ffffffffffffffcaffffffff00000024000000000000003400000000",
            INIT_3F => X"0000002200000000fffffff6ffffffff0000001f000000000000003800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffb5fffffffffffffff3fffffffffffffff4ffffffff0000001400000000",
            INIT_41 => X"0000002200000000ffffffe3ffffffff0000000600000000fffffff5ffffffff",
            INIT_42 => X"ffffffe3ffffffff000000480000000000000027000000000000000300000000",
            INIT_43 => X"ffffffe8fffffffffffffffdffffffffffffffeffffffffffffffff4ffffffff",
            INIT_44 => X"fffffffaffffffffffffffdaffffffff00000020000000000000000b00000000",
            INIT_45 => X"fffffff5fffffffffffffff2fffffffffffffffcffffffffffffffe0ffffffff",
            INIT_46 => X"fffffffaffffffff0000000000000000ffffffe6ffffffff0000001400000000",
            INIT_47 => X"00000009000000000000000d0000000000000003000000000000000000000000",
            INIT_48 => X"ffffffddffffffffffffffe0fffffffffffffff9fffffffffffffffaffffffff",
            INIT_49 => X"00000015000000000000003d00000000ffffffe0fffffffffffffffdffffffff",
            INIT_4A => X"ffffffe4fffffffffffffffdffffffff0000000a000000000000003000000000",
            INIT_4B => X"0000000500000000ffffffe8ffffffffffffffd0ffffffffffffffeeffffffff",
            INIT_4C => X"0000000700000000fffffff5ffffffff0000000d00000000ffffffe7ffffffff",
            INIT_4D => X"0000002900000000ffffffebffffffffffffffc3ffffffff0000000800000000",
            INIT_4E => X"fffffffbffffffffffffffddffffffffffffffcbffffffff0000003900000000",
            INIT_4F => X"fffffff2ffffffff0000002e000000000000000f00000000fffffff7ffffffff",
            INIT_50 => X"ffffffedffffffff0000001400000000fffffff8ffffffff0000001200000000",
            INIT_51 => X"0000000100000000ffffffe8ffffffff00000013000000000000001b00000000",
            INIT_52 => X"0000002000000000fffffffcffffffffffffffd7ffffffff0000000d00000000",
            INIT_53 => X"fffffffcffffffff0000000500000000fffffffffffffffffffffffeffffffff",
            INIT_54 => X"fffffffdffffffffffffffeeffffffff0000001d00000000ffffffefffffffff",
            INIT_55 => X"00000005000000000000000300000000fffffff4ffffffff0000001000000000",
            INIT_56 => X"0000001600000000fffffff6ffffffff00000007000000000000001c00000000",
            INIT_57 => X"0000000d000000000000000800000000ffffffe8fffffffffffffff9ffffffff",
            INIT_58 => X"fffffffeffffffff0000000300000000ffffffeaffffffff0000000500000000",
            INIT_59 => X"ffffffefffffffffffffffddffffffff0000000300000000fffffff3ffffffff",
            INIT_5A => X"ffffffc0ffffffffffffffd5ffffffffffffffccffffffffffffffe2ffffffff",
            INIT_5B => X"fffffffffffffffffffffffcffffffffffffffb3ffffffffffffffd2ffffffff",
            INIT_5C => X"0000002f00000000fffffff8ffffffffffffffe7ffffffff0000002100000000",
            INIT_5D => X"00000009000000000000003600000000ffffffe1ffffffffffffffd9ffffffff",
            INIT_5E => X"ffffffd0ffffffff0000000e000000000000000300000000ffffffffffffffff",
            INIT_5F => X"0000000c00000000ffffffe3ffffffffffffffd8ffffffff0000002900000000",
            INIT_60 => X"00000015000000000000002800000000ffffffedffffffffffffffe9ffffffff",
            INIT_61 => X"fffffff2ffffffffffffffe6fffffffffffffffdffffffff0000000c00000000",
            INIT_62 => X"00000014000000000000002000000000fffffff6ffffffff0000001000000000",
            INIT_63 => X"0000001d00000000ffffffefffffffffffffffffffffffff0000002e00000000",
            INIT_64 => X"0000000e000000000000001f00000000ffffffddfffffffffffffff5ffffffff",
            INIT_65 => X"0000002e00000000ffffffceffffffffffffffa9ffffffff0000000200000000",
            INIT_66 => X"0000001200000000fffffff1ffffffff0000000c00000000ffffffe6ffffffff",
            INIT_67 => X"fffffffbffffffffffffffd7fffffffffffffff4ffffffff0000001000000000",
            INIT_68 => X"ffffffc9ffffffff0000001600000000fffffff6ffffffffffffffe8ffffffff",
            INIT_69 => X"ffffffe7fffffffffffffffaffffffffffffffcdffffffff0000002600000000",
            INIT_6A => X"0000000a000000000000002700000000ffffffcdffffffffffffffceffffffff",
            INIT_6B => X"0000000300000000ffffffe2ffffffff00000019000000000000001600000000",
            INIT_6C => X"0000001700000000000000090000000000000008000000000000000200000000",
            INIT_6D => X"0000000d0000000000000016000000000000002e000000000000000f00000000",
            INIT_6E => X"0000000800000000ffffffdfffffffffffffffedffffffff0000001900000000",
            INIT_6F => X"ffffffeeffffffff00000005000000000000000a00000000fffffffdffffffff",
            INIT_70 => X"0000000000000000fffffff9ffffffff0000002300000000fffffffdffffffff",
            INIT_71 => X"ffffffeafffffffffffffff2ffffffffffffffeffffffffffffffff2ffffffff",
            INIT_72 => X"0000000700000000ffffffd5ffffffffffffffdcfffffffffffffffeffffffff",
            INIT_73 => X"0000001d00000000ffffffddffffffffffffffdcffffffff0000000200000000",
            INIT_74 => X"00000021000000000000001600000000fffffffdffffffff0000001700000000",
            INIT_75 => X"fffffff7ffffffff0000001500000000ffffffe3ffffffffffffffe6ffffffff",
            INIT_76 => X"ffffffe0ffffffff00000006000000000000000800000000ffffffdcffffffff",
            INIT_77 => X"ffffffe7fffffffffffffffeffffffff0000001600000000fffffffeffffffff",
            INIT_78 => X"00000028000000000000000d0000000000000002000000000000000600000000",
            INIT_79 => X"fffffffcffffffffffffffe7ffffffff0000000d000000000000002400000000",
            INIT_7A => X"fffffffeffffffff0000000a000000000000001100000000ffffffecffffffff",
            INIT_7B => X"ffffffbdffffffffffffffebffffffff00000002000000000000000d00000000",
            INIT_7C => X"0000000a000000000000002800000000ffffffc5ffffffffffffffbcffffffff",
            INIT_7D => X"0000000400000000fffffffafffffffffffffff6ffffffff0000000500000000",
            INIT_7E => X"0000001c000000000000001300000000ffffffd5ffffffff0000002000000000",
            INIT_7F => X"0000000200000000000000020000000000000019000000000000001000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE23;


    MEM_IWGHT_LAYER2_INSTANCE24 : if BRAM_NAME = "iwght_layer2_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000060000000000000001000000000000001100000000ffffffffffffffff",
            INIT_01 => X"00000000000000000000000c00000000fffffffcfffffffffffffffdffffffff",
            INIT_02 => X"fffffffeffffffff000000120000000000000000000000000000001400000000",
            INIT_03 => X"fffffff8ffffffffffffffecfffffffffffffffcffffffff0000000100000000",
            INIT_04 => X"fffffff0ffffffffffffffdcffffffff0000000000000000fffffff7ffffffff",
            INIT_05 => X"00000000000000000000001e00000000ffffffd9ffffffffffffffddffffffff",
            INIT_06 => X"0000001400000000fffffff8ffffffff0000002b000000000000003000000000",
            INIT_07 => X"0000000a0000000000000004000000000000001e00000000fffffffdffffffff",
            INIT_08 => X"fffffffbffffffff00000025000000000000001500000000fffffff6ffffffff",
            INIT_09 => X"00000037000000000000000200000000ffffffffffffffff0000000900000000",
            INIT_0A => X"000000150000000000000034000000000000001300000000fffffffeffffffff",
            INIT_0B => X"ffffffb5ffffffff0000000c00000000ffffffe8ffffffffffffffaeffffffff",
            INIT_0C => X"000000050000000000000003000000000000001b00000000ffffffe7ffffffff",
            INIT_0D => X"0000001500000000fffffff3ffffffffffffffd7fffffffffffffff0ffffffff",
            INIT_0E => X"0000001c000000000000000900000000fffffffeffffffff0000000900000000",
            INIT_0F => X"fffffff0ffffffff00000012000000000000000b000000000000000500000000",
            INIT_10 => X"00000021000000000000002a00000000fffffffdfffffffffffffffdffffffff",
            INIT_11 => X"0000002200000000000000360000000000000026000000000000001600000000",
            INIT_12 => X"ffffffebffffffffffffffb6ffffffffffffffa6ffffffffffffffddffffffff",
            INIT_13 => X"ffffffecffffffffffffffe1ffffffffffffffecfffffffffffffff9ffffffff",
            INIT_14 => X"ffffffd2ffffffffffffffd2ffffffff00000015000000000000000900000000",
            INIT_15 => X"0000001400000000ffffffe0ffffffffffffffd4fffffffffffffff3ffffffff",
            INIT_16 => X"00000051000000000000001900000000ffffffebffffffff0000002e00000000",
            INIT_17 => X"ffffffecffffffff0000000000000000fffffff2ffffffff0000001400000000",
            INIT_18 => X"0000001b000000000000002b000000000000002c00000000ffffffecffffffff",
            INIT_19 => X"ffffffeaffffffff0000000800000000ffffffe5ffffffff0000001700000000",
            INIT_1A => X"0000001200000000ffffffeeffffffffffffffebfffffffffffffffbffffffff",
            INIT_1B => X"fffffffbffffffffffffffe6fffffffffffffff9ffffffff0000000700000000",
            INIT_1C => X"ffffffffffffffffffffffeffffffffffffffffdffffffffffffffdbffffffff",
            INIT_1D => X"ffffffdcffffffffffffffe0fffffffffffffff6ffffffff0000000000000000",
            INIT_1E => X"0000001000000000fffffffafffffffffffffff1ffffffff0000002300000000",
            INIT_1F => X"ffffffe3ffffffffffffffd6ffffffffffffffebffffffff0000001000000000",
            INIT_20 => X"fffffffeffffffff0000002100000000ffffffccffffffffffffffbcffffffff",
            INIT_21 => X"0000000f00000000000000710000000000000051000000000000001500000000",
            INIT_22 => X"0000001e000000000000006a0000000000000018000000000000001e00000000",
            INIT_23 => X"ffffffdfffffffffffffffe7ffffffffffffffddffffffff0000002300000000",
            INIT_24 => X"fffffff2fffffffffffffff3ffffffff0000002a00000000ffffffecffffffff",
            INIT_25 => X"ffffffeeffffffff0000000c000000000000001500000000ffffffe7ffffffff",
            INIT_26 => X"00000021000000000000001f000000000000000800000000ffffffedffffffff",
            INIT_27 => X"ffffffeffffffffffffffffaffffffff0000000b00000000ffffffeeffffffff",
            INIT_28 => X"ffffffcbffffffffffffffe9ffffffff0000000700000000ffffffddffffffff",
            INIT_29 => X"0000000000000000ffffffe3fffffffffffffff9ffffffff0000000c00000000",
            INIT_2A => X"0000000900000000ffffffa8ffffffffffffffd7ffffffffffffffedffffffff",
            INIT_2B => X"ffffffc9ffffffff0000000c000000000000000600000000ffffffe0ffffffff",
            INIT_2C => X"ffffffdafffffffffffffff3ffffffff0000002000000000ffffffffffffffff",
            INIT_2D => X"0000002400000000ffffffabffffffffffffffbdffffffff0000003100000000",
            INIT_2E => X"ffffffafffffffff000000690000000000000014000000000000001b00000000",
            INIT_2F => X"0000001800000000ffffffd5ffffffff00000012000000000000001800000000",
            INIT_30 => X"ffffffffffffffff0000000200000000ffffffeeffffffff0000000400000000",
            INIT_31 => X"00000013000000000000000500000000fffffffbffffffff0000000700000000",
            INIT_32 => X"00000000000000000000001d00000000fffffffdffffffff0000000100000000",
            INIT_33 => X"ffffffa9ffffffff000000420000000000000013000000000000001900000000",
            INIT_34 => X"0000000000000000ffffffa8ffffffffffffffffffffffff0000001c00000000",
            INIT_35 => X"0000000400000000ffffffd5ffffffffffffff4effffffffffffffb3ffffffff",
            INIT_36 => X"ffffffc4ffffffffffffffddffffffffffffffddffffffff0000001700000000",
            INIT_37 => X"ffffffedfffffffffffffff3ffffffff0000000a00000000fffffff6ffffffff",
            INIT_38 => X"00000000000000000000001b0000000000000019000000000000000200000000",
            INIT_39 => X"ffffffe6ffffffff0000000700000000fffffff6fffffffffffffff9ffffffff",
            INIT_3A => X"ffffffd8ffffffff0000001a00000000ffffffffffffffffffffffc8ffffffff",
            INIT_3B => X"0000001700000000ffffffefffffffff0000004000000000fffffffdffffffff",
            INIT_3C => X"00000013000000000000001a000000000000003e000000000000005700000000",
            INIT_3D => X"0000000e00000000ffffffb4fffffffffffffffbffffffff0000003500000000",
            INIT_3E => X"ffffffedffffffffffffffffffffffffffffffd1fffffffffffffff2ffffffff",
            INIT_3F => X"fffffff9fffffffffffffff9ffffffff0000000a00000000ffffffd2ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002600000000ffffffe8fffffffffffffff3ffffffff0000001300000000",
            INIT_41 => X"ffffffddfffffffffffffffbffffffff00000029000000000000001700000000",
            INIT_42 => X"ffffffefffffffffffffffcdffffffffffffffebfffffffffffffff7ffffffff",
            INIT_43 => X"ffffffc2ffffffff0000000f00000000ffffffc6ffffffffffffffcfffffffff",
            INIT_44 => X"000000570000000000000006000000000000003000000000ffffffd2ffffffff",
            INIT_45 => X"fffffffaffffffff0000000e0000000000000013000000000000009700000000",
            INIT_46 => X"0000001e00000000ffffffbbffffffffffffffffffffffff0000002100000000",
            INIT_47 => X"0000000c00000000ffffffedffffffffffffffadffffffffffffffecffffffff",
            INIT_48 => X"ffffffebffffffff0000000100000000fffffffaffffffff0000000100000000",
            INIT_49 => X"fffffffdfffffffffffffff8ffffffffffffffeeffffffff0000000200000000",
            INIT_4A => X"0000000800000000fffffff6ffffffffffffffdaffffffff0000000f00000000",
            INIT_4B => X"ffffffc4ffffffff0000000d00000000fffffffdffffffffffffffd6ffffffff",
            INIT_4C => X"0000000900000000000000320000000000000000000000000000000100000000",
            INIT_4D => X"00000008000000000000001c000000000000001300000000fffffff0ffffffff",
            INIT_4E => X"ffffffcfffffffff0000003c0000000000000005000000000000003600000000",
            INIT_4F => X"0000000d00000000ffffffccffffffff0000001600000000fffffff2ffffffff",
            INIT_50 => X"0000000b0000000000000011000000000000000e000000000000000600000000",
            INIT_51 => X"0000000e00000000ffffffeefffffffffffffffdffffffff0000000800000000",
            INIT_52 => X"ffffffccfffffffffffffff4fffffffffffffffcfffffffffffffff7ffffffff",
            INIT_53 => X"0000000800000000ffffffc0ffffffffffffffb0ffffffffffffffefffffffff",
            INIT_54 => X"ffffffe0ffffffff0000000500000000ffffffdffffffffffffffffdffffffff",
            INIT_55 => X"0000001200000000fffffffcffffffff00000017000000000000001800000000",
            INIT_56 => X"ffffffe9fffffffffffffff2ffffffff0000000400000000ffffffe9ffffffff",
            INIT_57 => X"fffffffdffffffffffffffeffffffffffffffff7fffffffffffffffcffffffff",
            INIT_58 => X"0000000400000000ffffffe7ffffffffffffffd9ffffffffffffffedffffffff",
            INIT_59 => X"000000170000000000000014000000000000000400000000ffffffe4ffffffff",
            INIT_5A => X"ffffffddffffffffffffffd5ffffffffffffffeaffffffff0000002600000000",
            INIT_5B => X"fffffff9ffffffff00000016000000000000002a00000000fffffff3ffffffff",
            INIT_5C => X"ffffffe9ffffffffffffff99ffffffff0000000d00000000ffffffe7ffffffff",
            INIT_5D => X"00000017000000000000000000000000ffffffd3ffffffff0000001100000000",
            INIT_5E => X"ffffffcfffffffffffffffd1ffffffffffffffedffffffff0000000100000000",
            INIT_5F => X"ffffffe0ffffffffffffffe3ffffffff0000000b00000000ffffffeaffffffff",
            INIT_60 => X"ffffffe4ffffffff00000012000000000000001500000000fffffffaffffffff",
            INIT_61 => X"fffffff5ffffffffffffffd5ffffffff00000002000000000000000000000000",
            INIT_62 => X"0000001100000000ffffffd5ffffffffffffffb2ffffffffffffffe5ffffffff",
            INIT_63 => X"00000012000000000000002200000000fffffff3ffffffff0000002800000000",
            INIT_64 => X"fffffff1ffffffff00000017000000000000001700000000fffffff2ffffffff",
            INIT_65 => X"0000000d00000000ffffffeaffffffff00000012000000000000000000000000",
            INIT_66 => X"00000008000000000000000100000000ffffffdefffffffffffffff1ffffffff",
            INIT_67 => X"00000023000000000000003c00000000fffffffcfffffffffffffffaffffffff",
            INIT_68 => X"0000000f0000000000000037000000000000002c000000000000000100000000",
            INIT_69 => X"0000003100000000fffffff4ffffffffffffffd5ffffffff0000003d00000000",
            INIT_6A => X"ffffffdfffffffff0000001100000000fffffff3ffffffffffffffd6ffffffff",
            INIT_6B => X"ffffffd8ffffffff000000160000000000000038000000000000000b00000000",
            INIT_6C => X"0000001500000000fffffff6ffffffff00000011000000000000000900000000",
            INIT_6D => X"ffffffdfffffffff0000000f00000000ffffffd6ffffffff0000001800000000",
            INIT_6E => X"0000000c00000000fffffff8ffffffff0000000d00000000ffffffe3ffffffff",
            INIT_6F => X"00000014000000000000000100000000fffffffeffffffff0000003f00000000",
            INIT_70 => X"ffffffeafffffffffffffff6ffffffffffffffeaffffffffffffffedffffffff",
            INIT_71 => X"fffffff9ffffffffffffffe9fffffffffffffff5fffffffffffffffbffffffff",
            INIT_72 => X"0000000d00000000fffffff6ffffffffffffffe6ffffffffffffffefffffffff",
            INIT_73 => X"fffffff3ffffffff0000000500000000fffffffdfffffffffffffff2ffffffff",
            INIT_74 => X"fffffff5fffffffffffffff3ffffffffffffffe7ffffffffffffffffffffffff",
            INIT_75 => X"0000000b000000000000000300000000fffffffcffffffff0000001200000000",
            INIT_76 => X"fffffffaffffffffffffffeeffffffff00000009000000000000000e00000000",
            INIT_77 => X"00000006000000000000000d0000000000000000000000000000000900000000",
            INIT_78 => X"fffffff2ffffffff0000000f000000000000000d00000000ffffffeaffffffff",
            INIT_79 => X"000000100000000000000008000000000000000700000000fffffff8ffffffff",
            INIT_7A => X"0000000200000000ffffffeefffffffffffffff3fffffffffffffff6ffffffff",
            INIT_7B => X"fffffffdffffffffffffffe3ffffffffffffffffffffffff0000000800000000",
            INIT_7C => X"0000000600000000fffffff9ffffffff0000000400000000ffffffe8ffffffff",
            INIT_7D => X"fffffffffffffffffffffff2ffffffffffffffdfffffffffffffffebffffffff",
            INIT_7E => X"0000000500000000fffffffdffffffff0000000900000000ffffffe4ffffffff",
            INIT_7F => X"00000001000000000000000f00000000fffffffbffffffff0000000c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE24;


    MEM_IWGHT_LAYER2_INSTANCE25 : if BRAM_NAME = "iwght_layer2_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffffffffffffffffffecffffffffffffffe8ffffffff0000000a00000000",
            INIT_01 => X"00000004000000000000000000000000fffffff6fffffffffffffffdffffffff",
            INIT_02 => X"ffffffe9fffffffffffffff8ffffffffffffffeaffffffff0000000b00000000",
            INIT_03 => X"fffffff6fffffffffffffff8ffffffff00000005000000000000000a00000000",
            INIT_04 => X"00000003000000000000001000000000ffffffeafffffffffffffff9ffffffff",
            INIT_05 => X"00000005000000000000000f00000000fffffff1ffffffff0000000a00000000",
            INIT_06 => X"0000000500000000ffffffffffffffff0000000000000000fffffffbffffffff",
            INIT_07 => X"00000003000000000000000d00000000fffffff5fffffffffffffffdffffffff",
            INIT_08 => X"0000000f00000000ffffffeeffffffffffffffeeffffffff0000000400000000",
            INIT_09 => X"0000000d000000000000000c000000000000000a00000000ffffffedffffffff",
            INIT_0A => X"fffffffffffffffffffffffcffffffff00000006000000000000000400000000",
            INIT_0B => X"fffffffffffffffffffffffaffffffff0000000900000000fffffff6ffffffff",
            INIT_0C => X"fffffff6ffffffff0000000200000000ffffffecffffffff0000000300000000",
            INIT_0D => X"ffffffeaffffffff0000000300000000fffffff2ffffffff0000000600000000",
            INIT_0E => X"fffffffbfffffffffffffff6ffffffffffffffe3fffffffffffffff9ffffffff",
            INIT_0F => X"00000013000000000000000d00000000fffffffffffffffffffffff6ffffffff",
            INIT_10 => X"ffffffeffffffffffffffffaffffffff0000000f00000000ffffffedffffffff",
            INIT_11 => X"fffffff7ffffffff0000000700000000ffffffeffffffffffffffffdffffffff",
            INIT_12 => X"ffffffe9fffffffffffffff4ffffffff0000000400000000ffffffedffffffff",
            INIT_13 => X"0000000e00000000fffffff1fffffffffffffffbffffffff0000000200000000",
            INIT_14 => X"00000004000000000000000a00000000ffffffe8ffffffff0000000000000000",
            INIT_15 => X"0000000e000000000000000d00000000fffffffeffffffffffffffe9ffffffff",
            INIT_16 => X"0000000500000000ffffffe5ffffffff0000000a000000000000000600000000",
            INIT_17 => X"ffffffffffffffffffffffedffffffff0000001000000000ffffffe6ffffffff",
            INIT_18 => X"fffffff8fffffffffffffff2ffffffff0000000a00000000fffffff5ffffffff",
            INIT_19 => X"fffffff0fffffffffffffff9ffffffff0000000000000000ffffffe4ffffffff",
            INIT_1A => X"fffffff6ffffffffffffffe1fffffffffffffffaffffffff0000000400000000",
            INIT_1B => X"0000001300000000fffffff5ffffffff00000012000000000000000300000000",
            INIT_1C => X"fffffffdfffffffffffffff8fffffffffffffffcfffffffffffffff6ffffffff",
            INIT_1D => X"ffffffeeffffffffffffffecffffffff0000000e000000000000001100000000",
            INIT_1E => X"00000000000000000000000600000000ffffffedffffffff0000000c00000000",
            INIT_1F => X"ffffffe5ffffffff0000000a000000000000001700000000fffffff0ffffffff",
            INIT_20 => X"fffffff3ffffffff00000014000000000000001000000000fffffff2ffffffff",
            INIT_21 => X"0000000100000000fffffff4ffffffff00000003000000000000000e00000000",
            INIT_22 => X"ffffffedffffffff0000000400000000fffffff4ffffffffffffffedffffffff",
            INIT_23 => X"0000000800000000ffffffeaffffffff0000000600000000ffffffe7ffffffff",
            INIT_24 => X"ffffffedffffffff0000001000000000ffffffedfffffffffffffff0ffffffff",
            INIT_25 => X"0000000d00000000fffffff0ffffffff0000000100000000fffffff9ffffffff",
            INIT_26 => X"0000000400000000ffffffe9fffffffffffffff8fffffffffffffff2ffffffff",
            INIT_27 => X"ffffffecffffffffffffffffffffffff0000000200000000fffffffbffffffff",
            INIT_28 => X"ffffffeefffffffffffffffbffffffff0000000b00000000fffffff1ffffffff",
            INIT_29 => X"fffffff6ffffffff000000020000000000000008000000000000000300000000",
            INIT_2A => X"ffffffeaffffffffffffffedfffffffffffffff9fffffffffffffff7ffffffff",
            INIT_2B => X"00000011000000000000000100000000ffffffe9ffffffff0000000600000000",
            INIT_2C => X"0000000500000000fffffff6ffffffff00000006000000000000000500000000",
            INIT_2D => X"0000000600000000fffffffafffffffffffffffbfffffffffffffff0ffffffff",
            INIT_2E => X"0000001500000000fffffffdffffffff0000000b00000000ffffffffffffffff",
            INIT_2F => X"0000000b000000000000000b000000000000000a00000000ffffffffffffffff",
            INIT_30 => X"0000000200000000fffffff0fffffffffffffff9fffffffffffffff4ffffffff",
            INIT_31 => X"ffffffecfffffffffffffff9fffffffffffffffaffffffff0000000400000000",
            INIT_32 => X"fffffff3ffffffff0000000800000000fffffff1fffffffffffffff4ffffffff",
            INIT_33 => X"fffffff2ffffffffffffffe9fffffffffffffffbffffffff0000000500000000",
            INIT_34 => X"ffffffffffffffff0000000500000000fffffff2fffffffffffffff0ffffffff",
            INIT_35 => X"ffffffeaffffffff0000000600000000fffffff7ffffffffffffffebffffffff",
            INIT_36 => X"ffffffffffffffff0000000500000000fffffffafffffffffffffff6ffffffff",
            INIT_37 => X"fffffff7ffffffff0000000f000000000000000100000000fffffff0ffffffff",
            INIT_38 => X"fffffff5fffffffffffffff3ffffffff0000000c00000000fffffff9ffffffff",
            INIT_39 => X"fffffffefffffffffffffffeffffffff0000000f00000000fffffff6ffffffff",
            INIT_3A => X"000000080000000000000004000000000000000000000000fffffffcffffffff",
            INIT_3B => X"ffffffebffffffffffffffe4ffffffff0000000000000000fffffff5ffffffff",
            INIT_3C => X"0000000400000000fffffff6fffffffffffffffbfffffffffffffff8ffffffff",
            INIT_3D => X"ffffffe7ffffffffffffffecffffffffffffffeefffffffffffffffcffffffff",
            INIT_3E => X"ffffffecffffffff00000003000000000000001400000000fffffff0ffffffff",
            INIT_3F => X"ffffffecfffffffffffffffdfffffffffffffff3fffffffffffffff2ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffedffffffff0000000c000000000000000a000000000000000300000000",
            INIT_41 => X"0000000d00000000fffffff1fffffffffffffff5ffffffffffffffefffffffff",
            INIT_42 => X"fffffff6ffffffff0000000200000000fffffff1ffffffffffffffffffffffff",
            INIT_43 => X"00000000000000000000000900000000ffffffffffffffff0000000200000000",
            INIT_44 => X"ffffffffffffffff0000001300000000fffffff5ffffffff0000000c00000000",
            INIT_45 => X"ffffffefffffffff0000000600000000fffffffeffffffffffffffeeffffffff",
            INIT_46 => X"0000000400000000fffffff2ffffffff0000000000000000ffffffffffffffff",
            INIT_47 => X"0000000200000000fffffffdfffffffffffffff7fffffffffffffff8ffffffff",
            INIT_48 => X"fffffff1fffffffffffffff6fffffffffffffffeffffffffffffffe2ffffffff",
            INIT_49 => X"0000001300000000fffffffcffffffff0000000b000000000000001400000000",
            INIT_4A => X"ffffffeeffffffff000000050000000000000003000000000000000800000000",
            INIT_4B => X"ffffffeaffffffff0000000600000000fffffff5ffffffff0000000300000000",
            INIT_4C => X"fffffff0fffffffffffffffbffffffffffffffffffffffff0000000300000000",
            INIT_4D => X"fffffff7ffffffff0000000000000000ffffffedfffffffffffffffcffffffff",
            INIT_4E => X"0000000800000000ffffffe6ffffffff0000000d00000000ffffffe0ffffffff",
            INIT_4F => X"fffffff2ffffffffffffffeffffffffffffffff4fffffffffffffff9ffffffff",
            INIT_50 => X"0000001400000000fffffffbfffffffffffffff3ffffffff0000001200000000",
            INIT_51 => X"fffffff3ffffffffffffffd0ffffffffffffffebffffffffffffffecffffffff",
            INIT_52 => X"0000000b00000000fffffff0fffffffffffffff3ffffffff0000001000000000",
            INIT_53 => X"0000000000000000fffffffdffffffff00000012000000000000000000000000",
            INIT_54 => X"0000000500000000ffffffdefffffffffffffff3ffffffff0000000200000000",
            INIT_55 => X"0000000d00000000fffffff4ffffffff0000000300000000ffffffeeffffffff",
            INIT_56 => X"ffffffe5fffffffffffffff6ffffffff00000008000000000000001400000000",
            INIT_57 => X"0000000a00000000ffffffefffffffff0000001e00000000ffffffeeffffffff",
            INIT_58 => X"fffffff4ffffffff0000000e00000000fffffff7fffffffffffffffdffffffff",
            INIT_59 => X"0000000500000000fffffffcffffffff00000003000000000000000600000000",
            INIT_5A => X"000000090000000000000003000000000000000500000000ffffffefffffffff",
            INIT_5B => X"ffffffeffffffffffffffffbffffffff00000000000000000000000f00000000",
            INIT_5C => X"fffffff6ffffffff0000000f00000000fffffff5ffffffffffffffedffffffff",
            INIT_5D => X"ffffffdeffffffff0000000500000000fffffff2ffffffffffffffedffffffff",
            INIT_5E => X"fffffff1ffffffff0000000c00000000ffffffecfffffffffffffff1ffffffff",
            INIT_5F => X"ffffffe3ffffffff0000000600000000fffffff7fffffffffffffffeffffffff",
            INIT_60 => X"fffffff9ffffffff0000000c0000000000000001000000000000000e00000000",
            INIT_61 => X"ffffffe6fffffffffffffffefffffffffffffff1ffffffff0000000300000000",
            INIT_62 => X"00000000000000000000001b00000000fffffffeffffffffffffffeaffffffff",
            INIT_63 => X"fffffff0fffffffffffffff7fffffffffffffffcfffffffffffffff9ffffffff",
            INIT_64 => X"fffffffeffffffff00000018000000000000000f00000000ffffffdfffffffff",
            INIT_65 => X"ffffffe2ffffffffffffffe6ffffffff0000000900000000ffffffeaffffffff",
            INIT_66 => X"ffffffeeffffffff000000000000000000000000000000000000000500000000",
            INIT_67 => X"ffffffeeffffffff0000000200000000ffffffeeffffffffffffffefffffffff",
            INIT_68 => X"ffffffe7ffffffff0000000800000000ffffffecfffffffffffffff5ffffffff",
            INIT_69 => X"fffffff8ffffffff00000000000000000000000800000000fffffffbffffffff",
            INIT_6A => X"fffffffcffffffffffffffeeffffffff00000001000000000000000400000000",
            INIT_6B => X"ffffffefffffffff0000000000000000fffffff8ffffffffffffffdaffffffff",
            INIT_6C => X"ffffffe5fffffffffffffff4fffffffffffffff1fffffffffffffffbffffffff",
            INIT_6D => X"000000110000000000000004000000000000000300000000ffffffe5ffffffff",
            INIT_6E => X"fffffff3fffffffffffffff0ffffffffffffffdffffffffffffffff2ffffffff",
            INIT_6F => X"ffffffd7ffffffffffffffe2ffffffff0000000800000000fffffffbffffffff",
            INIT_70 => X"fffffff1fffffffffffffff7fffffffffffffff7ffffffffffffffebffffffff",
            INIT_71 => X"ffffffdcffffffff00000003000000000000000f000000000000000b00000000",
            INIT_72 => X"ffffffe6ffffffffffffffe7ffffffff0000000d000000000000000000000000",
            INIT_73 => X"fffffffbfffffffffffffffbfffffffffffffff1ffffffffffffffebffffffff",
            INIT_74 => X"0000000200000000fffffff1ffffffffffffffffffffffffffffffe7ffffffff",
            INIT_75 => X"fffffff8fffffffffffffffffffffffffffffff9fffffffffffffff5ffffffff",
            INIT_76 => X"ffffffecfffffffffffffff9ffffffffffffffebfffffffffffffff3ffffffff",
            INIT_77 => X"fffffff6ffffffff0000000600000000ffffffe0ffffffff0000000a00000000",
            INIT_78 => X"000000000000000000000006000000000000000700000000fffffffdffffffff",
            INIT_79 => X"00000017000000000000000700000000ffffffe7ffffffffffffffe8ffffffff",
            INIT_7A => X"fffffffdffffffffffffffeaffffffff00000002000000000000000600000000",
            INIT_7B => X"ffffffefffffffff0000001100000000ffffffe5ffffffff0000000100000000",
            INIT_7C => X"000000050000000000000005000000000000000800000000ffffffedffffffff",
            INIT_7D => X"00000003000000000000000200000000ffffffecfffffffffffffff3ffffffff",
            INIT_7E => X"fffffff0ffffffff0000000000000000ffffffdcfffffffffffffff4ffffffff",
            INIT_7F => X"fffffff2ffffffff00000005000000000000000200000000ffffffefffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE25;


    MEM_IWGHT_LAYER2_INSTANCE26 : if BRAM_NAME = "iwght_layer2_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000001c000000000000001f000000000000002200000000",
            INIT_01 => X"fffffffcffffffff00000016000000000000001500000000ffffffffffffffff",
            INIT_02 => X"ffffffc4ffffffffffffffc6ffffffffffffffeaffffffff0000001a00000000",
            INIT_03 => X"ffffffddffffffffffffffcdffffffffffffffc8fffffffffffffff7ffffffff",
            INIT_04 => X"00000014000000000000001e00000000ffffffa5ffffffffffffffa8ffffffff",
            INIT_05 => X"fffffff0ffffffffffffffe2ffffffffffffffd8ffffffff0000000e00000000",
            INIT_06 => X"fffffffeffffffffffffffecfffffffffffffff5fffffffffffffff4ffffffff",
            INIT_07 => X"ffffffeeffffffff0000000a0000000000000003000000000000000a00000000",
            INIT_08 => X"0000001a000000000000001e0000000000000032000000000000000b00000000",
            INIT_09 => X"fffffffbffffffff00000005000000000000001d000000000000000600000000",
            INIT_0A => X"0000001d000000000000000100000000fffffff4ffffffffffffffedffffffff",
            INIT_0B => X"0000000200000000ffffffe8ffffffffffffffcbffffffff0000000100000000",
            INIT_0C => X"000000140000000000000001000000000000000100000000ffffffefffffffff",
            INIT_0D => X"ffffffeaffffffffffffffedffffffff0000000a000000000000000200000000",
            INIT_0E => X"00000014000000000000001f00000000fffffff9ffffffff0000001500000000",
            INIT_0F => X"0000001b00000000ffffffe9ffffffffffffffb5ffffffffffffffe6ffffffff",
            INIT_10 => X"0000001a00000000000000200000000000000016000000000000000700000000",
            INIT_11 => X"00000008000000000000000a000000000000002a000000000000001b00000000",
            INIT_12 => X"0000000700000000000000260000000000000026000000000000002100000000",
            INIT_13 => X"00000026000000000000001f000000000000000e000000000000001200000000",
            INIT_14 => X"fffffffefffffffffffffffcffffffff0000000700000000ffffffecffffffff",
            INIT_15 => X"ffffffeefffffffffffffffbffffffff0000000b00000000ffffffe6ffffffff",
            INIT_16 => X"0000003300000000ffffffffffffffffffffffe0ffffffff0000000e00000000",
            INIT_17 => X"0000001800000000000000120000000000000004000000000000001c00000000",
            INIT_18 => X"fffffff7ffffffff000000240000000000000018000000000000001f00000000",
            INIT_19 => X"0000000e00000000ffffffefffffffff0000001400000000ffffffe5ffffffff",
            INIT_1A => X"0000000e00000000ffffffd8ffffffff00000003000000000000001000000000",
            INIT_1B => X"ffffffb7ffffffff000000000000000000000000000000000000001100000000",
            INIT_1C => X"ffffffdbffffffffffffffd8ffffffffffffffe0ffffffffffffffc1ffffffff",
            INIT_1D => X"ffffffceffffffffffffffeeffffffffffffffd7ffffffffffffffdbffffffff",
            INIT_1E => X"0000000e00000000fffffff0ffffffff00000036000000000000001700000000",
            INIT_1F => X"fffffff3ffffffff0000000600000000fffffffdffffffff0000001100000000",
            INIT_20 => X"000000110000000000000000000000000000000f00000000fffffff7ffffffff",
            INIT_21 => X"fffffff1fffffffffffffff1ffffffff0000000000000000ffffffefffffffff",
            INIT_22 => X"ffffffecffffffffffffffe4ffffffff0000001500000000ffffffeeffffffff",
            INIT_23 => X"ffffffc1ffffffffffffffacffffffffffffffceffffffffffffffe0ffffffff",
            INIT_24 => X"ffffffe0ffffffff000000070000000000000017000000000000000800000000",
            INIT_25 => X"ffffffefffffffffffffffe8fffffffffffffff3ffffffffffffffebffffffff",
            INIT_26 => X"ffffffdbffffffff0000000a0000000000000000000000000000000600000000",
            INIT_27 => X"fffffff6fffffffffffffffbffffffffffffffd2ffffffff0000001400000000",
            INIT_28 => X"fffffffeffffffffffffffc6ffffffffffffffe4ffffffffffffffa3ffffffff",
            INIT_29 => X"ffffffedffffffff0000000400000000ffffffddffffffffffffffc1ffffffff",
            INIT_2A => X"ffffffd5ffffffff0000000b00000000fffffff7ffffffff0000000800000000",
            INIT_2B => X"0000000000000000ffffffdfffffffffffffffeaffffffffffffffe4ffffffff",
            INIT_2C => X"ffffffd9ffffffff0000000100000000ffffffe5ffffffff0000000400000000",
            INIT_2D => X"0000001800000000ffffffeaffffffffffffffedfffffffffffffff1ffffffff",
            INIT_2E => X"00000018000000000000000c0000000000000012000000000000002000000000",
            INIT_2F => X"00000018000000000000000c000000000000001100000000fffffff8ffffffff",
            INIT_30 => X"ffffffccffffffff00000008000000000000000000000000fffffff4ffffffff",
            INIT_31 => X"00000012000000000000000900000000ffffffe6ffffffffffffffacffffffff",
            INIT_32 => X"0000002400000000000000160000000000000011000000000000001d00000000",
            INIT_33 => X"0000000d00000000ffffffe7ffffffffffffffedffffffffffffffbaffffffff",
            INIT_34 => X"fffffffdffffffffffffffebffffffff0000000100000000ffffffffffffffff",
            INIT_35 => X"fffffffeffffffff0000000d00000000ffffffdcffffffffffffffe7ffffffff",
            INIT_36 => X"0000000b00000000fffffff5ffffffffffffffe8ffffffffffffffc9ffffffff",
            INIT_37 => X"ffffffcdfffffffffffffff6ffffffff0000000c00000000ffffffd7ffffffff",
            INIT_38 => X"0000001c000000000000000400000000fffffff0ffffffff0000000100000000",
            INIT_39 => X"fffffffbffffffffffffffe8ffffffffffffffdfffffffff0000001000000000",
            INIT_3A => X"00000001000000000000001900000000ffffffe8ffffffffffffffd9ffffffff",
            INIT_3B => X"0000001800000000fffffff5ffffffff00000011000000000000000d00000000",
            INIT_3C => X"0000000900000000000000340000000000000022000000000000002800000000",
            INIT_3D => X"ffffffeeffffffffffffffefffffffff00000001000000000000000400000000",
            INIT_3E => X"fffffffbffffffffffffffe9fffffffffffffffdffffffff0000000e00000000",
            INIT_3F => X"fffffff7ffffffff0000001c0000000000000006000000000000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001900000000fffffffffffffffffffffffbfffffffffffffffcffffffff",
            INIT_41 => X"0000000c000000000000000a00000000fffffff8ffffffff0000001700000000",
            INIT_42 => X"fffffff5ffffffffffffffebfffffffffffffffcffffffff0000000800000000",
            INIT_43 => X"0000000100000000ffffffecfffffffffffffffaffffffffffffffe2ffffffff",
            INIT_44 => X"0000000500000000ffffffe5ffffffffffffffe3ffffffff0000000d00000000",
            INIT_45 => X"0000002500000000fffffffbffffffffffffffe3ffffffffffffffa9ffffffff",
            INIT_46 => X"0000000c00000000000000250000000000000013000000000000000200000000",
            INIT_47 => X"00000027000000000000003d0000000000000042000000000000002b00000000",
            INIT_48 => X"0000000700000000ffffffe5ffffffffffffffe4ffffffffffffffe6ffffffff",
            INIT_49 => X"fffffff9ffffffff0000000400000000ffffffe6fffffffffffffff5ffffffff",
            INIT_4A => X"0000001b000000000000002f0000000000000014000000000000001100000000",
            INIT_4B => X"ffffffdffffffffffffffff3ffffffffffffffecffffffff0000002600000000",
            INIT_4C => X"0000000b0000000000000007000000000000002d00000000ffffffd9ffffffff",
            INIT_4D => X"00000003000000000000000e000000000000001d00000000ffffffd2ffffffff",
            INIT_4E => X"0000001600000000000000140000000000000016000000000000003b00000000",
            INIT_4F => X"00000004000000000000000500000000fffffff0ffffffff0000000400000000",
            INIT_50 => X"0000001a0000000000000027000000000000000b00000000ffffffeaffffffff",
            INIT_51 => X"00000003000000000000001900000000ffffffebffffffff0000002800000000",
            INIT_52 => X"fffffffbfffffffffffffff5fffffffffffffff4ffffffff0000001300000000",
            INIT_53 => X"fffffffaffffffff00000014000000000000004000000000fffffff0ffffffff",
            INIT_54 => X"fffffffaffffffffffffffe7ffffffff00000000000000000000002500000000",
            INIT_55 => X"ffffffc6fffffffffffffff4fffffffffffffffbffffffffffffffdfffffffff",
            INIT_56 => X"ffffffe4ffffffffffffffd3ffffffff0000000100000000ffffffe2ffffffff",
            INIT_57 => X"ffffffdcffffffff0000000000000000ffffffd8fffffffffffffff0ffffffff",
            INIT_58 => X"ffffffffffffffffffffffc7ffffffffffffffc2ffffffffffffffe1ffffffff",
            INIT_59 => X"0000002000000000ffffffe9fffffffffffffff1ffffffffffffffebffffffff",
            INIT_5A => X"ffffffc8ffffffffffffffa7ffffffffffffffe3ffffffffffffffd9ffffffff",
            INIT_5B => X"ffffffe0fffffffffffffffcffffffffffffffd0ffffffffffffffdeffffffff",
            INIT_5C => X"000000480000000000000009000000000000000300000000ffffffd1ffffffff",
            INIT_5D => X"00000019000000000000000b000000000000000e000000000000000c00000000",
            INIT_5E => X"ffffffecffffffffffffffd6ffffffff00000026000000000000002d00000000",
            INIT_5F => X"0000000300000000fffffff9ffffffff0000000400000000ffffffd0ffffffff",
            INIT_60 => X"ffffffa4ffffffff00000016000000000000000b00000000fffffff6ffffffff",
            INIT_61 => X"ffffffaeffffffffffffffccffffffffffffffafffffffffffffff7cffffffff",
            INIT_62 => X"0000001800000000fffffffefffffffffffffff4ffffffff0000000f00000000",
            INIT_63 => X"0000000c00000000ffffffa0ffffffffffffffd5ffffffffffffffe5ffffffff",
            INIT_64 => X"00000029000000000000002000000000fffffff9ffffffffffffffeeffffffff",
            INIT_65 => X"0000001d00000000ffffffdbfffffffffffffff7fffffffffffffff0ffffffff",
            INIT_66 => X"00000001000000000000000900000000ffffffffffffffffffffffefffffffff",
            INIT_67 => X"fffffff3ffffffff0000000a000000000000003400000000fffffff5ffffffff",
            INIT_68 => X"fffffff0ffffffff0000000c000000000000000b00000000fffffffbffffffff",
            INIT_69 => X"ffffffc0fffffffffffffff0ffffffffffffffefffffffff0000000000000000",
            INIT_6A => X"ffffffc9ffffffffffffffe9fffffffffffffff0ffffffffffffffb9ffffffff",
            INIT_6B => X"0000000000000000ffffffd4ffffffffffffffd8ffffffffffffffecffffffff",
            INIT_6C => X"0000000000000000fffffffdfffffffffffffffeffffffff0000000b00000000",
            INIT_6D => X"fffffffeffffffff000000000000000000000002000000000000001400000000",
            INIT_6E => X"fffffff0ffffffff0000001f000000000000002d000000000000001100000000",
            INIT_6F => X"0000000800000000fffffff0ffffffff00000018000000000000001600000000",
            INIT_70 => X"0000001e000000000000001500000000ffffffffffffffffffffffdaffffffff",
            INIT_71 => X"0000003d00000000ffffffe4ffffffff00000001000000000000001f00000000",
            INIT_72 => X"0000001f00000000fffffffbffffffff00000008000000000000000900000000",
            INIT_73 => X"0000002e000000000000000a00000000fffffff9ffffffff0000000900000000",
            INIT_74 => X"ffffffe5fffffffffffffff5fffffffffffffff5ffffffffffffffdbffffffff",
            INIT_75 => X"00000030000000000000000b00000000fffffffcffffffff0000002a00000000",
            INIT_76 => X"fffffff6ffffffff000000150000000000000010000000000000001200000000",
            INIT_77 => X"ffffffc5ffffffffffffffb7ffffffffffffffddffffffff0000001900000000",
            INIT_78 => X"fffffffcfffffffffffffff8ffffffffffffffdfffffffffffffffe3ffffffff",
            INIT_79 => X"ffffff99ffffffffffffffaeffffffff0000000200000000ffffffc3ffffffff",
            INIT_7A => X"0000000a00000000ffffffb6ffffffffffffffdeffffffffffffffbeffffffff",
            INIT_7B => X"ffffffe2fffffffffffffff7ffffffffffffffd6ffffffff0000000000000000",
            INIT_7C => X"fffffffbffffffff0000001100000000ffffffcdffffffffffffffddffffffff",
            INIT_7D => X"0000000a0000000000000036000000000000002100000000fffffff8ffffffff",
            INIT_7E => X"0000000900000000ffffffefffffffffffffffeaffffffff0000000000000000",
            INIT_7F => X"fffffff4ffffffff0000000900000000fffffff2fffffffffffffffbffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE26;


    MEM_IWGHT_LAYER2_INSTANCE27 : if BRAM_NAME = "iwght_layer2_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff3ffffffff0000000a000000000000000c000000000000000f00000000",
            INIT_01 => X"00000013000000000000000c0000000000000009000000000000002f00000000",
            INIT_02 => X"fffffff1ffffffffffffffe5ffffffff00000016000000000000001f00000000",
            INIT_03 => X"fffffff8ffffffff00000009000000000000001300000000ffffffcdffffffff",
            INIT_04 => X"ffffffd9ffffffff00000015000000000000002b000000000000001500000000",
            INIT_05 => X"fffffff3ffffffffffffffe1ffffffffffffffe1fffffffffffffff6ffffffff",
            INIT_06 => X"00000002000000000000001b000000000000003300000000ffffffedffffffff",
            INIT_07 => X"0000001100000000000000000000000000000017000000000000001800000000",
            INIT_08 => X"0000000a00000000000000110000000000000015000000000000001700000000",
            INIT_09 => X"ffffffe0fffffffffffffffeffffffff00000001000000000000002100000000",
            INIT_0A => X"0000004e00000000fffffffffffffffffffffffdffffffff0000002600000000",
            INIT_0B => X"fffffffcffffffffffffffebffffffff00000017000000000000002c00000000",
            INIT_0C => X"0000000900000000000000000000000000000010000000000000001000000000",
            INIT_0D => X"ffffffbbffffffff0000000700000000fffffffbffffffffffffffefffffffff",
            INIT_0E => X"fffffff6fffffffffffffff3fffffffffffffff4ffffffffffffffd9ffffffff",
            INIT_0F => X"000000350000000000000011000000000000002c00000000fffffff9ffffffff",
            INIT_10 => X"0000001100000000ffffffeaffffffffffffffcfffffffff0000001400000000",
            INIT_11 => X"0000000600000000fffffff0ffffffff0000000000000000fffffff6ffffffff",
            INIT_12 => X"ffffffbdfffffffffffffff4fffffffffffffff9fffffffffffffffaffffffff",
            INIT_13 => X"0000003800000000fffffffbffffffffffffffeefffffffffffffffcffffffff",
            INIT_14 => X"0000001f00000000ffffffebffffffff0000000000000000ffffffaeffffffff",
            INIT_15 => X"0000000e00000000fffffffcffffffff00000001000000000000001b00000000",
            INIT_16 => X"ffffffd3ffffffff0000000600000000ffffffd9ffffffffffffffe1ffffffff",
            INIT_17 => X"fffffff6ffffffffffffffcbffffffff0000002a00000000ffffffecffffffff",
            INIT_18 => X"fffffff4fffffffffffffff8ffffffffffffffeefffffffffffffff5ffffffff",
            INIT_19 => X"ffffffd8ffffffff0000000e00000000ffffffedffffffffffffffeaffffffff",
            INIT_1A => X"00000010000000000000001b00000000ffffffe0fffffffffffffff0ffffffff",
            INIT_1B => X"0000003100000000fffffff1ffffffff0000000500000000ffffffe5ffffffff",
            INIT_1C => X"ffffffedffffffff0000001d00000000fffffffaffffffff0000000000000000",
            INIT_1D => X"fffffff9ffffffffffffffe5ffffffffffffffefffffffff0000002300000000",
            INIT_1E => X"fffffffaffffffff0000000600000000fffffff4ffffffff0000002300000000",
            INIT_1F => X"0000000d00000000ffffffe0ffffffff00000005000000000000000e00000000",
            INIT_20 => X"00000026000000000000000b000000000000002100000000ffffffecffffffff",
            INIT_21 => X"ffffffefffffffffffffffeeffffffff00000014000000000000001f00000000",
            INIT_22 => X"ffffffd1ffffffff0000001000000000ffffffd3ffffffffffffffd8ffffffff",
            INIT_23 => X"ffffffd8fffffffffffffff9ffffffff0000000200000000fffffffbffffffff",
            INIT_24 => X"0000000100000000000000350000000000000028000000000000000a00000000",
            INIT_25 => X"0000004500000000fffffff1ffffffff0000000b000000000000001c00000000",
            INIT_26 => X"ffffffc0ffffffff0000001200000000fffffffbffffffff0000000700000000",
            INIT_27 => X"fffffff8ffffffffffffffddffffffff0000001400000000ffffffe5ffffffff",
            INIT_28 => X"fffffffeffffffff000000070000000000000006000000000000000a00000000",
            INIT_29 => X"00000003000000000000001700000000fffffffdfffffffffffffff7ffffffff",
            INIT_2A => X"ffffffe0fffffffffffffff8ffffffff00000000000000000000000300000000",
            INIT_2B => X"ffffffcffffffffffffffff0ffffffff0000001a00000000ffffffdfffffffff",
            INIT_2C => X"ffffffcaffffffff0000002000000000ffffffbdffffffffffffffb5ffffffff",
            INIT_2D => X"ffffffc3ffffffff000000030000000000000026000000000000000300000000",
            INIT_2E => X"0000002a00000000ffffffeffffffffffffffffcffffffff0000002d00000000",
            INIT_2F => X"fffffffffffffffffffffff1ffffffff00000000000000000000003400000000",
            INIT_30 => X"fffffff1fffffffffffffffcfffffffffffffffbffffffff0000000400000000",
            INIT_31 => X"0000000e000000000000000900000000fffffff3fffffffffffffffaffffffff",
            INIT_32 => X"fffffff5ffffffff0000006200000000ffffffe4ffffffff0000000700000000",
            INIT_33 => X"fffffffeffffffffffffffe8ffffffff00000014000000000000000000000000",
            INIT_34 => X"0000001f00000000ffffffe4ffffffff00000030000000000000001f00000000",
            INIT_35 => X"ffffffffffffffff00000020000000000000001c000000000000000f00000000",
            INIT_36 => X"0000000900000000fffffffcffffffff00000014000000000000003200000000",
            INIT_37 => X"00000020000000000000000800000000fffffffeffffffff0000000b00000000",
            INIT_38 => X"0000004b00000000fffffffeffffffffffffffebffffffffffffffeaffffffff",
            INIT_39 => X"0000001000000000fffffff9ffffffffffffffd3fffffffffffffff7ffffffff",
            INIT_3A => X"ffffffedfffffffffffffff8fffffffffffffffaffffffff0000002c00000000",
            INIT_3B => X"ffffffffffffffff0000001a00000000fffffffaffffffff0000002400000000",
            INIT_3C => X"ffffffd8ffffffff0000001200000000fffffffcffffffff0000000700000000",
            INIT_3D => X"0000000700000000ffffffefffffffffffffffe2ffffffff0000001100000000",
            INIT_3E => X"ffffffffffffffff000000240000000000000002000000000000000000000000",
            INIT_3F => X"0000000f00000000fffffff5ffffffff0000000d000000000000001300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffdffffffff00000012000000000000000a000000000000000600000000",
            INIT_41 => X"0000001100000000fffffff7ffffffffffffffebffffffff0000001100000000",
            INIT_42 => X"ffffffd7ffffffff00000025000000000000000e000000000000001b00000000",
            INIT_43 => X"0000000800000000fffffff6ffffffffffffffd7ffffffffffffffeaffffffff",
            INIT_44 => X"0000000300000000fffffff5ffffffffffffffeafffffffffffffff4ffffffff",
            INIT_45 => X"ffffffdfffffffffffffffd3ffffffff00000012000000000000000100000000",
            INIT_46 => X"0000003300000000fffffff5fffffffffffffff1ffffffff0000002000000000",
            INIT_47 => X"ffffffc6ffffffff00000004000000000000001d00000000ffffffd0ffffffff",
            INIT_48 => X"0000001800000000ffffffecffffffffffffffd0ffffffff0000003100000000",
            INIT_49 => X"ffffffd6ffffffff00000000000000000000000300000000ffffffdbffffffff",
            INIT_4A => X"ffffffe6fffffffffffffff2ffffffffffffffeaffffffff0000001400000000",
            INIT_4B => X"00000015000000000000002c0000000000000002000000000000002500000000",
            INIT_4C => X"fffffff3ffffffffffffffe8ffffffffffffffeefffffffffffffffbffffffff",
            INIT_4D => X"fffffff2ffffffff0000000e000000000000000000000000fffffff0ffffffff",
            INIT_4E => X"ffffffe4fffffffffffffff6ffffffffffffffebffffffff0000001900000000",
            INIT_4F => X"000000070000000000000011000000000000000b000000000000002200000000",
            INIT_50 => X"000000220000000000000028000000000000002500000000fffffff9ffffffff",
            INIT_51 => X"00000017000000000000003600000000ffffffe8ffffffff0000000000000000",
            INIT_52 => X"ffffffd4ffffffff0000001100000000fffffffbffffffff0000001c00000000",
            INIT_53 => X"fffffffeffffffff0000003400000000ffffffe4ffffffffffffffe5ffffffff",
            INIT_54 => X"fffffffaffffffff00000002000000000000002100000000ffffffc4ffffffff",
            INIT_55 => X"0000002d000000000000000300000000fffffffbffffffff0000002100000000",
            INIT_56 => X"ffffffd9ffffffff0000003500000000ffffffbdffffffff0000001700000000",
            INIT_57 => X"0000000400000000ffffffe2ffffffff00000008000000000000001800000000",
            INIT_58 => X"0000001100000000000000230000000000000010000000000000000300000000",
            INIT_59 => X"0000000c0000000000000009000000000000001900000000fffffffcffffffff",
            INIT_5A => X"ffffffe0fffffffffffffffdffffffffffffffeefffffffffffffff3ffffffff",
            INIT_5B => X"0000000800000000ffffffecfffffffffffffff7ffffffffffffffdfffffffff",
            INIT_5C => X"0000000a00000000000000040000000000000012000000000000000c00000000",
            INIT_5D => X"ffffffd0ffffffffffffffccffffffffffffffa9ffffffff0000002a00000000",
            INIT_5E => X"00000002000000000000003e000000000000001300000000fffffffdffffffff",
            INIT_5F => X"00000000000000000000000500000000ffffffe7fffffffffffffffdffffffff",
            INIT_60 => X"ffffffc2ffffffffffffffd6ffffffff0000000b00000000ffffffecffffffff",
            INIT_61 => X"0000001100000000ffffffe3fffffffffffffffaffffffff0000000d00000000",
            INIT_62 => X"ffffffcbffffffffffffffe7ffffffffffffffd3ffffffff0000000b00000000",
            INIT_63 => X"ffffffecffffffff0000000f000000000000001b00000000ffffffb4ffffffff",
            INIT_64 => X"0000001a00000000ffffffdcffffffff0000002d000000000000001b00000000",
            INIT_65 => X"00000029000000000000002b00000000ffffffc7ffffffffffffffdaffffffff",
            INIT_66 => X"fffffff8ffffffffffffffe6ffffffffffffffdbffffffff0000000900000000",
            INIT_67 => X"fffffffaffffffff000000120000000000000019000000000000001e00000000",
            INIT_68 => X"fffffff6ffffffff000000190000000000000034000000000000000000000000",
            INIT_69 => X"0000001300000000fffffffcffffffff00000016000000000000002800000000",
            INIT_6A => X"ffffffd5ffffffffffffffe6ffffffff0000000600000000ffffffdcffffffff",
            INIT_6B => X"0000000f000000000000000600000000ffffffe3ffffffff0000000400000000",
            INIT_6C => X"fffffffefffffffffffffffeffffffff00000025000000000000001b00000000",
            INIT_6D => X"0000000500000000fffffffeffffffff00000016000000000000002300000000",
            INIT_6E => X"00000024000000000000001200000000fffffff5ffffffffffffffdeffffffff",
            INIT_6F => X"0000000e000000000000000f00000000fffffffeffffffff0000000f00000000",
            INIT_70 => X"fffffff0ffffffffffffffe8fffffffffffffffcfffffffffffffffeffffffff",
            INIT_71 => X"ffffffd4ffffffffffffffd1ffffffff0000002e000000000000000400000000",
            INIT_72 => X"000000120000000000000003000000000000000300000000ffffffddffffffff",
            INIT_73 => X"ffffffc7ffffffff0000004c0000000000000018000000000000002200000000",
            INIT_74 => X"0000000000000000fffffffeffffffff00000038000000000000001100000000",
            INIT_75 => X"ffffffe1fffffffffffffff8ffffffff00000002000000000000000d00000000",
            INIT_76 => X"fffffff4fffffffffffffff7ffffffff0000000f000000000000003000000000",
            INIT_77 => X"0000000a000000000000000000000000ffffffc9ffffffffffffffc1ffffffff",
            INIT_78 => X"0000000000000000000000090000000000000008000000000000000c00000000",
            INIT_79 => X"00000002000000000000001100000000ffffffffffffffff0000000700000000",
            INIT_7A => X"ffffffbdffffffffffffffd2ffffffff0000000a000000000000001500000000",
            INIT_7B => X"0000000d000000000000001b000000000000002b00000000ffffffeeffffffff",
            INIT_7C => X"fffffff7ffffffffffffffd0ffffffffffffffd8ffffffffffffffe4ffffffff",
            INIT_7D => X"0000000700000000ffffffc6ffffffffffffffb8fffffffffffffffeffffffff",
            INIT_7E => X"ffffffc0ffffffffffffffc6ffffffffffffffeafffffffffffffffdffffffff",
            INIT_7F => X"ffffffebffffffffffffffdcffffffffffffffccffffffff0000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE27;


    MEM_IWGHT_LAYER2_INSTANCE28 : if BRAM_NAME = "iwght_layer2_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd9fffffffffffffff6ffffffff0000000c00000000ffffffaaffffffff",
            INIT_01 => X"ffffffe0fffffffffffffff0fffffffffffffff7fffffffffffffffeffffffff",
            INIT_02 => X"fffffff4ffffffffffffffccffffffffffffffcbfffffffffffffffcffffffff",
            INIT_03 => X"ffffffebfffffffffffffff9ffffffffffffffeeffffffffffffffd8ffffffff",
            INIT_04 => X"00000004000000000000000a000000000000000e000000000000000d00000000",
            INIT_05 => X"fffffff8ffffffffffffffe4ffffffffffffffeaffffffff0000000300000000",
            INIT_06 => X"ffffffdfffffffffffffffe1ffffffffffffffc6ffffffff0000000a00000000",
            INIT_07 => X"fffffff9ffffffff0000000c000000000000000900000000ffffffe1ffffffff",
            INIT_08 => X"0000002b00000000ffffffe9ffffffffffffffe8ffffffffffffffd5ffffffff",
            INIT_09 => X"0000001600000000fffffff2ffffffff00000023000000000000001f00000000",
            INIT_0A => X"0000000900000000fffffffbffffffffffffffb5ffffffff0000005800000000",
            INIT_0B => X"ffffffdeffffffff0000004d0000000000000016000000000000002800000000",
            INIT_0C => X"0000001600000000ffffffceffffffff0000001f000000000000000500000000",
            INIT_0D => X"ffffffceffffffffffffffe0ffffffffffffffd1ffffffff0000000f00000000",
            INIT_0E => X"ffffffe5fffffffffffffff6ffffffffffffffe8ffffffff0000002400000000",
            INIT_0F => X"0000003d00000000ffffffefffffffffffffffc0ffffffffffffffd5ffffffff",
            INIT_10 => X"0000000500000000000000030000000000000029000000000000002400000000",
            INIT_11 => X"0000001400000000fffffffcffffffff00000000000000000000002200000000",
            INIT_12 => X"ffffffe8ffffffff0000000b000000000000000000000000ffffffe0ffffffff",
            INIT_13 => X"ffffffe9ffffffffffffffdfffffffffffffffe6fffffffffffffffaffffffff",
            INIT_14 => X"0000000900000000fffffffdffffffffffffffe2ffffffff0000001300000000",
            INIT_15 => X"fffffffaffffffff00000005000000000000002a00000000fffffff7ffffffff",
            INIT_16 => X"ffffffdaffffffffffffffe5ffffffff00000010000000000000001800000000",
            INIT_17 => X"ffffffecffffffffffffffc7ffffffffffffffd2ffffffffffffffd2ffffffff",
            INIT_18 => X"ffffffd8ffffffffffffffc6ffffffffffffffedffffffff0000000c00000000",
            INIT_19 => X"0000001e00000000ffffffdfffffffffffffffeaffffffffffffffcdffffffff",
            INIT_1A => X"0000001e00000000ffffffeaffffffffffffffe4ffffffffffffffeeffffffff",
            INIT_1B => X"0000000000000000fffffffaffffffff00000044000000000000001e00000000",
            INIT_1C => X"ffffffe5ffffffffffffffeeffffffffffffffe5ffffffffffffffbaffffffff",
            INIT_1D => X"ffffffcefffffffffffffff1fffffffffffffff2ffffffffffffffcbffffffff",
            INIT_1E => X"ffffffcdffffffffffffffdffffffffffffffff0ffffffffffffffe3ffffffff",
            INIT_1F => X"0000001e000000000000000900000000ffffffccffffffffffffffe8ffffffff",
            INIT_20 => X"0000002200000000ffffffe8fffffffffffffffbffffffff0000001900000000",
            INIT_21 => X"0000000e000000000000003700000000ffffffe2fffffffffffffff3ffffffff",
            INIT_22 => X"00000023000000000000000300000000fffffff2fffffffffffffff0ffffffff",
            INIT_23 => X"0000000b00000000ffffffd5ffffffff00000006000000000000000100000000",
            INIT_24 => X"ffffffe8ffffffffffffffdcfffffffffffffffcffffffffffffffe3ffffffff",
            INIT_25 => X"ffffffedffffffffffffffe6ffffffff00000029000000000000001d00000000",
            INIT_26 => X"0000001100000000fffffff0ffffffffffffffefffffffffffffffccffffffff",
            INIT_27 => X"ffffffb5ffffffff0000002b00000000ffffffedffffffffffffffc1ffffffff",
            INIT_28 => X"ffffffceffffffffffffffb6fffffffffffffffcffffffffffffffeaffffffff",
            INIT_29 => X"0000000b00000000fffffffeffffffffffffffdcfffffffffffffff9ffffffff",
            INIT_2A => X"ffffffe3ffffffffffffffd5ffffffffffffffefffffffffffffffedffffffff",
            INIT_2B => X"ffffffd4ffffffffffffffe1ffffffff0000002000000000ffffffe7ffffffff",
            INIT_2C => X"0000002900000000ffffffc3fffffffffffffffcffffffff0000000500000000",
            INIT_2D => X"fffffff9ffffffff0000001700000000ffffffdcffffffff0000001000000000",
            INIT_2E => X"ffffffd4ffffffffffffffacffffffffffffff99fffffffffffffff9ffffffff",
            INIT_2F => X"00000011000000000000001200000000ffffffccffffffffffffffdeffffffff",
            INIT_30 => X"fffffff7ffffffff0000002300000000ffffffc5fffffffffffffff8ffffffff",
            INIT_31 => X"ffffffb7ffffffff00000004000000000000002800000000ffffffcdffffffff",
            INIT_32 => X"ffffffebffffffff0000000000000000ffffffd1fffffffffffffffeffffffff",
            INIT_33 => X"ffffffc3ffffffffffffffeefffffffffffffff5ffffffffffffffbfffffffff",
            INIT_34 => X"000000540000000000000021000000000000002400000000ffffffd4ffffffff",
            INIT_35 => X"0000000b00000000000000230000000000000006000000000000002400000000",
            INIT_36 => X"fffffff7ffffffff0000001c0000000000000019000000000000001600000000",
            INIT_37 => X"ffffffceffffffffffffffebffffffff0000002c00000000ffffffe5ffffffff",
            INIT_38 => X"ffffffb0ffffffffffffffe8fffffffffffffff0ffffffff0000001a00000000",
            INIT_39 => X"ffffffbaffffffffffffffe4ffffffff0000001c00000000ffffffa6ffffffff",
            INIT_3A => X"fffffff3ffffffffffffffcbffffffffffffffeaffffffffffffff9effffffff",
            INIT_3B => X"ffffffa6ffffffff0000003700000000ffffffcbffffffffffffffdfffffffff",
            INIT_3C => X"ffffffa5ffffffffffffffaaffffffffffffffd1ffffffffffffffd9ffffffff",
            INIT_3D => X"0000001d00000000000000260000000000000025000000000000001200000000",
            INIT_3E => X"0000001e000000000000002500000000fffffffdffffffff0000000600000000",
            INIT_3F => X"fffffffdfffffffffffffff5ffffffff0000001f000000000000002c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000d000000000000000800000000fffffffcffffffff0000001200000000",
            INIT_41 => X"000000060000000000000010000000000000001200000000ffffffecffffffff",
            INIT_42 => X"ffffffadfffffffffffffffaffffffff0000001b00000000ffffffd1ffffffff",
            INIT_43 => X"0000001100000000ffffffdafffffffffffffffeffffffffffffffdaffffffff",
            INIT_44 => X"0000000000000000000000270000000000000041000000000000001700000000",
            INIT_45 => X"0000002600000000000000030000000000000025000000000000001a00000000",
            INIT_46 => X"ffffffeafffffffffffffff3fffffffffffffff7ffffffff0000004200000000",
            INIT_47 => X"0000000900000000ffffffd1ffffffffffffffdfffffffff0000001400000000",
            INIT_48 => X"ffffffadffffffffffffffbeffffffffffffffcdffffffffffffffd8ffffffff",
            INIT_49 => X"ffffffebfffffffffffffff0ffffffffffffffbaffffffff0000002600000000",
            INIT_4A => X"0000002500000000ffffffbcffffffffffffffd5fffffffffffffff6ffffffff",
            INIT_4B => X"ffffffffffffffff0000000a00000000ffffffc5ffffffff0000000000000000",
            INIT_4C => X"fffffffbffffffff0000000e000000000000000000000000ffffffa1ffffffff",
            INIT_4D => X"fffffffdffffffff0000000c0000000000000023000000000000002700000000",
            INIT_4E => X"fffffff5ffffffff00000000000000000000001500000000fffffffbffffffff",
            INIT_4F => X"0000000f00000000fffffffeffffffffffffffd9ffffffff0000001f00000000",
            INIT_50 => X"ffffffe8fffffffffffffff4ffffffffffffffcaffffffffffffffd3ffffffff",
            INIT_51 => X"ffffffbeffffffffffffffbfffffffff0000002300000000ffffffe3ffffffff",
            INIT_52 => X"ffffffc1ffffffffffffff9cffffffff0000001c00000000fffffff5ffffffff",
            INIT_53 => X"0000000700000000ffffffddffffffffffffffe1ffffffffffffffefffffffff",
            INIT_54 => X"fffffffbffffffff0000001200000000fffffffeffffffffffffffe6ffffffff",
            INIT_55 => X"ffffffeafffffffffffffff9ffffffff0000001b00000000fffffff8ffffffff",
            INIT_56 => X"fffffffeffffffff000000050000000000000018000000000000001f00000000",
            INIT_57 => X"ffffffe6fffffffffffffffdffffffffffffffdeffffffffffffffe8ffffffff",
            INIT_58 => X"fffffff0fffffffffffffff7ffffffff0000001e00000000fffffffcffffffff",
            INIT_59 => X"0000001f00000000fffffffbfffffffffffffff8ffffffff0000002100000000",
            INIT_5A => X"ffffffebffffffff00000026000000000000000f00000000fffffffaffffffff",
            INIT_5B => X"ffffffc4fffffffffffffff5ffffffff0000002600000000ffffffc7ffffffff",
            INIT_5C => X"0000001300000000ffffffdeffffffff0000000b000000000000002200000000",
            INIT_5D => X"fffffffaffffffff000000390000000000000003000000000000000900000000",
            INIT_5E => X"ffffffdbffffffff00000018000000000000003200000000fffffffeffffffff",
            INIT_5F => X"fffffff1ffffffff0000002e000000000000001300000000ffffffefffffffff",
            INIT_60 => X"0000001300000000ffffffecffffffff00000018000000000000001f00000000",
            INIT_61 => X"0000002200000000ffffffddfffffffffffffff5ffffffff0000000800000000",
            INIT_62 => X"ffffffb7ffffffffffffffeeffffffffffffff96fffffffffffffff5ffffffff",
            INIT_63 => X"0000001e0000000000000022000000000000000200000000ffffffe1ffffffff",
            INIT_64 => X"000000260000000000000014000000000000000b000000000000001200000000",
            INIT_65 => X"0000002c0000000000000028000000000000001200000000fffffff4ffffffff",
            INIT_66 => X"0000001a000000000000003f00000000fffffffeffffffff0000001000000000",
            INIT_67 => X"00000019000000000000003d000000000000004500000000ffffffe2ffffffff",
            INIT_68 => X"ffffffc3ffffffff0000000400000000ffffffecffffffffffffffe7ffffffff",
            INIT_69 => X"ffffffe2ffffffff0000000100000000ffffffdcffffffffffffffdaffffffff",
            INIT_6A => X"0000002e000000000000001f000000000000002900000000ffffffe6ffffffff",
            INIT_6B => X"00000040000000000000000c0000000000000051000000000000003100000000",
            INIT_6C => X"0000000f000000000000002a0000000000000030000000000000004d00000000",
            INIT_6D => X"00000018000000000000004200000000ffffffecffffffff0000001100000000",
            INIT_6E => X"fffffff5ffffffff000000020000000000000023000000000000000200000000",
            INIT_6F => X"ffffffdcffffffffffffffefffffffffffffffc2ffffffffffffffb3ffffffff",
            INIT_70 => X"fffffff8ffffffffffffffe3ffffffffffffffffffffffffffffffecffffffff",
            INIT_71 => X"0000000200000000ffffffd1ffffffffffffffdfffffffff0000000f00000000",
            INIT_72 => X"000000100000000000000007000000000000000b00000000fffffff3ffffffff",
            INIT_73 => X"ffffffe3ffffffff0000000d000000000000000d000000000000001100000000",
            INIT_74 => X"ffffffdeffffffffffffffe5ffffffffffffffb8fffffffffffffff3ffffffff",
            INIT_75 => X"00000005000000000000001000000000ffffffd6ffffffffffffffccffffffff",
            INIT_76 => X"00000014000000000000000b000000000000000000000000ffffffdbffffffff",
            INIT_77 => X"000000000000000000000011000000000000000400000000fffffff1ffffffff",
            INIT_78 => X"ffffffeaffffffffffffffe6ffffffff00000000000000000000002d00000000",
            INIT_79 => X"ffffffd7ffffffffffffffd6fffffffffffffff8ffffffffffffffd8ffffffff",
            INIT_7A => X"0000003300000000ffffffecffffffffffffffe1ffffffffffffffeeffffffff",
            INIT_7B => X"0000002c000000000000002700000000fffffffffffffffffffffff3ffffffff",
            INIT_7C => X"0000000e00000000ffffffd3fffffffffffffffdffffffff0000002c00000000",
            INIT_7D => X"ffffffccfffffffffffffff1ffffffff0000000100000000ffffffe5ffffffff",
            INIT_7E => X"0000002200000000ffffffe7ffffffffffffffcdffffffffffffffe0ffffffff",
            INIT_7F => X"0000001900000000fffffff9ffffffffffffffceffffffff0000001d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE28;


    MEM_IWGHT_LAYER2_INSTANCE29 : if BRAM_NAME = "iwght_layer2_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffb6ffffffff0000000500000000fffffff5fffffffffffffffcffffffff",
            INIT_01 => X"0000002000000000ffffffbdffffffff0000003700000000ffffffe2ffffffff",
            INIT_02 => X"fffffff3fffffffffffffffdffffffffffffffd8ffffffff0000000000000000",
            INIT_03 => X"0000000900000000ffffffb5ffffffffffffffaeffffffff0000002700000000",
            INIT_04 => X"0000000f00000000000000120000000000000023000000000000003200000000",
            INIT_05 => X"ffffffffffffffffffffffd1ffffffffffffffffffffffff0000000e00000000",
            INIT_06 => X"fffffff4ffffffffffffffffffffffff00000020000000000000000a00000000",
            INIT_07 => X"fffffffeffffffff0000000300000000fffffff1ffffffffffffffd5ffffffff",
            INIT_08 => X"fffffff5ffffffff0000000c000000000000000b000000000000001200000000",
            INIT_09 => X"ffffffe8ffffffff00000000000000000000000f000000000000000500000000",
            INIT_0A => X"00000012000000000000000500000000fffffff2ffffffff0000000300000000",
            INIT_0B => X"00000023000000000000000900000000fffffff8fffffffffffffff4ffffffff",
            INIT_0C => X"0000000700000000fffffff5ffffffffffffffd1fffffffffffffff9ffffffff",
            INIT_0D => X"000000440000000000000026000000000000000b000000000000002d00000000",
            INIT_0E => X"ffffffefffffffff000000210000000000000019000000000000001400000000",
            INIT_0F => X"ffffffd5ffffffffffffffe7ffffffffffffffefffffffffffffffccffffffff",
            INIT_10 => X"0000001a000000000000002d00000000ffffffd8ffffffffffffffddffffffff",
            INIT_11 => X"fffffffeffffffff0000001100000000ffffffeffffffffffffffff6ffffffff",
            INIT_12 => X"ffffffeafffffffffffffff0ffffffff00000026000000000000001300000000",
            INIT_13 => X"0000000900000000fffffffdffffffff00000032000000000000001b00000000",
            INIT_14 => X"fffffff8ffffffff0000001f000000000000001a000000000000002400000000",
            INIT_15 => X"0000000a00000000ffffffe7fffffffffffffffefffffffffffffffaffffffff",
            INIT_16 => X"0000001a00000000000000230000000000000000000000000000000700000000",
            INIT_17 => X"0000001d00000000000000000000000000000004000000000000003800000000",
            INIT_18 => X"0000000000000000ffffffeffffffffffffffffdffffffff0000000700000000",
            INIT_19 => X"fffffff7ffffffffffffffecffffffff00000014000000000000000000000000",
            INIT_1A => X"fffffff8fffffffffffffffbffffffffffffffb4ffffffff0000001100000000",
            INIT_1B => X"ffffffffffffffffffffffe4ffffffffffffffe7ffffffffffffffcfffffffff",
            INIT_1C => X"fffffffcffffffffffffffe4ffffffffffffffddffffffffffffffe6ffffffff",
            INIT_1D => X"0000001300000000000000290000000000000020000000000000000900000000",
            INIT_1E => X"000000140000000000000012000000000000000200000000ffffffffffffffff",
            INIT_1F => X"0000001100000000ffffffecffffffffffffffe0ffffffff0000000000000000",
            INIT_20 => X"ffffffecffffffff000000130000000000000000000000000000000900000000",
            INIT_21 => X"ffffffbfffffffffffffffedffffffffffffffc8ffffffffffffffedffffffff",
            INIT_22 => X"fffffffbffffffffffffffe0ffffffffffffffc5ffffffffffffffd6ffffffff",
            INIT_23 => X"ffffffedffffffff0000000600000000ffffffedffffffffffffffe1ffffffff",
            INIT_24 => X"fffffffaffffffffffffffdfffffffffffffffeeffffffff0000001a00000000",
            INIT_25 => X"0000000000000000fffffff1ffffffff0000000500000000ffffffc7ffffffff",
            INIT_26 => X"0000001c0000000000000009000000000000000700000000ffffffc4ffffffff",
            INIT_27 => X"0000002b00000000ffffffd9ffffffffffffffe7ffffffff0000000500000000",
            INIT_28 => X"0000002f00000000000000250000000000000015000000000000002600000000",
            INIT_29 => X"0000003d0000000000000024000000000000003b000000000000002d00000000",
            INIT_2A => X"0000000b0000000000000002000000000000002c000000000000001b00000000",
            INIT_2B => X"ffffffe7fffffffffffffff1ffffffff00000026000000000000000c00000000",
            INIT_2C => X"0000001100000000fffffffdfffffffffffffff9ffffffffffffffecffffffff",
            INIT_2D => X"ffffffd6ffffffff0000002b0000000000000014000000000000001d00000000",
            INIT_2E => X"ffffffecffffffffffffffc5ffffffff0000001e00000000ffffffecffffffff",
            INIT_2F => X"ffffffe3ffffffffffffffd5ffffffffffffffe3ffffffffffffffd5ffffffff",
            INIT_30 => X"0000001a00000000ffffffeaffffffffffffffebffffffff0000001600000000",
            INIT_31 => X"0000003c00000000000000280000000000000009000000000000002000000000",
            INIT_32 => X"ffffffffffffffff000000130000000000000012000000000000001b00000000",
            INIT_33 => X"ffffffd4ffffffff00000022000000000000001300000000ffffffd9ffffffff",
            INIT_34 => X"0000000800000000ffffffe8ffffffffffffffd7ffffffffffffffe7ffffffff",
            INIT_35 => X"fffffff6ffffffff0000001400000000ffffffefffffffff0000000000000000",
            INIT_36 => X"ffffffdaffffffff00000025000000000000000800000000ffffffe9ffffffff",
            INIT_37 => X"ffffffedfffffffffffffffbffffffff0000000200000000ffffffe6ffffffff",
            INIT_38 => X"0000000000000000ffffffc8ffffffffffffffe8ffffffffffffffd3ffffffff",
            INIT_39 => X"ffffffeeffffffff000000260000000000000016000000000000003000000000",
            INIT_3A => X"ffffffe7ffffffffffffffd6ffffffffffffffd9ffffffffffffffe0ffffffff",
            INIT_3B => X"000000070000000000000009000000000000001b000000000000000500000000",
            INIT_3C => X"fffffffbffffffffffffffbdffffffffffffffcfffffffffffffffbdffffffff",
            INIT_3D => X"0000003200000000ffffffe8ffffffffffffffb6ffffffffffffffdeffffffff",
            INIT_3E => X"0000002600000000ffffffd9ffffffff00000001000000000000000200000000",
            INIT_3F => X"ffffffceffffffff0000000c00000000ffffffeafffffffffffffffdffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffafffffffffffffffdfffffffffffffff8ffffffffffffffddffffffff",
            INIT_41 => X"0000002400000000000000120000000000000015000000000000001200000000",
            INIT_42 => X"000000230000000000000016000000000000001d000000000000000200000000",
            INIT_43 => X"fffffffbfffffffffffffff8ffffffff0000001800000000ffffffd9ffffffff",
            INIT_44 => X"ffffffffffffffff0000003e000000000000003900000000fffffffcffffffff",
            INIT_45 => X"ffffffe9ffffffff000000080000000000000014000000000000001300000000",
            INIT_46 => X"fffffffbfffffffffffffffdffffffffffffffedffffffff0000000900000000",
            INIT_47 => X"00000015000000000000001b000000000000001c000000000000001700000000",
            INIT_48 => X"ffffffdefffffffffffffff8ffffffff0000000d000000000000003000000000",
            INIT_49 => X"ffffffedffffffffffffffd2ffffffff0000000700000000ffffffeaffffffff",
            INIT_4A => X"00000024000000000000001700000000ffffffcbffffffffffffffffffffffff",
            INIT_4B => X"0000000b00000000ffffffe8fffffffffffffffdfffffffffffffffbffffffff",
            INIT_4C => X"ffffffdaffffffffffffffe2ffffffff0000002b00000000fffffff9ffffffff",
            INIT_4D => X"0000001a0000000000000012000000000000004200000000ffffffecffffffff",
            INIT_4E => X"ffffffe0ffffffff00000002000000000000000c00000000fffffff8ffffffff",
            INIT_4F => X"fffffffbffffffff0000000900000000ffffffceffffffff0000000800000000",
            INIT_50 => X"0000000200000000fffffff1ffffffff00000002000000000000001000000000",
            INIT_51 => X"ffffffe7ffffffff000000010000000000000005000000000000000a00000000",
            INIT_52 => X"ffffffd6ffffffffffffffd7fffffffffffffffaffffffffffffffe7ffffffff",
            INIT_53 => X"0000001e00000000fffffff1ffffffffffffffe3ffffffff0000000200000000",
            INIT_54 => X"ffffffceffffffff0000001d0000000000000018000000000000003800000000",
            INIT_55 => X"ffffffe1ffffffffffffffc5ffffffff0000000b000000000000000700000000",
            INIT_56 => X"0000002500000000fffffff1ffffffffffffffd3ffffffff0000002000000000",
            INIT_57 => X"fffffffaffffffffffffffd4ffffffffffffffceffffffffffffffbcffffffff",
            INIT_58 => X"00000015000000000000000a0000000000000008000000000000000c00000000",
            INIT_59 => X"ffffffebffffffff000000170000000000000020000000000000000d00000000",
            INIT_5A => X"ffffffeffffffffffffffffeffffffffffffffe8ffffffffffffffb7ffffffff",
            INIT_5B => X"ffffffecfffffffffffffffeffffffff0000003e000000000000002300000000",
            INIT_5C => X"ffffffebfffffffffffffffbfffffffffffffff9ffffffffffffffcaffffffff",
            INIT_5D => X"fffffff3ffffffff000000240000000000000026000000000000001500000000",
            INIT_5E => X"ffffffe6fffffffffffffff3ffffffff0000002e00000000ffffffe6ffffffff",
            INIT_5F => X"ffffffe9ffffffff0000000200000000fffffff0fffffffffffffffcffffffff",
            INIT_60 => X"00000012000000000000000500000000ffffffdfffffffffffffffb5ffffffff",
            INIT_61 => X"ffffffc1ffffffff000000120000000000000017000000000000000e00000000",
            INIT_62 => X"0000000e000000000000000000000000ffffffdbffffffff0000000d00000000",
            INIT_63 => X"0000001b0000000000000009000000000000000400000000fffffffaffffffff",
            INIT_64 => X"000000020000000000000012000000000000000100000000fffffffbffffffff",
            INIT_65 => X"0000001500000000000000260000000000000015000000000000000200000000",
            INIT_66 => X"ffffffcaffffffff00000017000000000000001600000000ffffffebffffffff",
            INIT_67 => X"ffffffddffffffffffffffd3ffffffffffffffe5ffffffffffffffdfffffffff",
            INIT_68 => X"000000160000000000000029000000000000000a00000000ffffffe4ffffffff",
            INIT_69 => X"fffffffdffffffffffffffe1ffffffffffffffe8ffffffffffffffe0ffffffff",
            INIT_6A => X"0000000700000000ffffffefffffffffffffffd7fffffffffffffff1ffffffff",
            INIT_6B => X"00000007000000000000000f00000000ffffffeeffffffff0000001400000000",
            INIT_6C => X"0000001300000000fffffff3ffffffffffffffe2ffffffff0000001100000000",
            INIT_6D => X"0000000c00000000000000150000000000000010000000000000001c00000000",
            INIT_6E => X"000000010000000000000016000000000000001600000000fffffffaffffffff",
            INIT_6F => X"ffffffb7ffffffff0000003e0000000000000017000000000000000a00000000",
            INIT_70 => X"ffffffd4ffffffffffffff9efffffffffffffff5ffffffffffffffb9ffffffff",
            INIT_71 => X"0000001800000000ffffffedfffffffffffffff6ffffffff0000000200000000",
            INIT_72 => X"fffffff6ffffffffffffffe5ffffffff0000001c00000000ffffffdfffffffff",
            INIT_73 => X"000000240000000000000039000000000000000a000000000000001200000000",
            INIT_74 => X"00000021000000000000000400000000ffffffddffffffff0000002900000000",
            INIT_75 => X"ffffffe2ffffffff0000001200000000fffffff1ffffffff0000000300000000",
            INIT_76 => X"0000000a000000000000000a00000000ffffffefffffffffffffffd6ffffffff",
            INIT_77 => X"0000003300000000000000310000000000000019000000000000003000000000",
            INIT_78 => X"fffffff0ffffffff0000001900000000ffffffdcffffffffffffffebffffffff",
            INIT_79 => X"00000015000000000000001b0000000000000011000000000000001a00000000",
            INIT_7A => X"ffffffebffffffff0000000c0000000000000031000000000000000700000000",
            INIT_7B => X"fffffffeffffffff00000019000000000000000600000000ffffffe2ffffffff",
            INIT_7C => X"0000000e000000000000002400000000fffffff7ffffffffffffffeaffffffff",
            INIT_7D => X"0000000d00000000ffffffcaffffffff0000003100000000ffffffedffffffff",
            INIT_7E => X"fffffff8ffffffff000000040000000000000016000000000000000700000000",
            INIT_7F => X"ffffffe5ffffffff00000003000000000000001c000000000000002600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE29;


    MEM_IWGHT_LAYER2_INSTANCE30 : if BRAM_NAME = "iwght_layer2_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffcffffffffffffffcdffffffffffffffdfffffffff0000001200000000",
            INIT_01 => X"0000000300000000fffffff6ffffffff0000001300000000ffffffedffffffff",
            INIT_02 => X"00000023000000000000000100000000ffffffdbffffffff0000000b00000000",
            INIT_03 => X"ffffffc7ffffffff0000002900000000ffffffdbfffffffffffffff0ffffffff",
            INIT_04 => X"0000002300000000ffffffd1ffffffffffffffe1ffffffff0000001200000000",
            INIT_05 => X"0000000100000000ffffffedfffffffffffffff9ffffffffffffffe6ffffffff",
            INIT_06 => X"fffffffafffffffffffffff2ffffffff0000001700000000ffffffe3ffffffff",
            INIT_07 => X"ffffffc4ffffffff0000000700000000ffffffcfffffffff0000000700000000",
            INIT_08 => X"ffffffedfffffffffffffff0ffffffff0000000900000000ffffffc7ffffffff",
            INIT_09 => X"fffffff1ffffffff0000000700000000fffffff7fffffffffffffff8ffffffff",
            INIT_0A => X"ffffffd4ffffffff00000020000000000000001100000000ffffffd5ffffffff",
            INIT_0B => X"fffffff8ffffffff00000008000000000000000e000000000000000700000000",
            INIT_0C => X"ffffffccffffffff000000090000000000000018000000000000002100000000",
            INIT_0D => X"0000002000000000ffffffe1ffffffffffffffe7ffffffff0000002d00000000",
            INIT_0E => X"ffffffdbffffffffffffffb8ffffffffffffffebffffffff0000002600000000",
            INIT_0F => X"0000000600000000fffffff4ffffffff00000002000000000000000d00000000",
            INIT_10 => X"00000016000000000000000e000000000000001200000000ffffffecffffffff",
            INIT_11 => X"ffffffb8fffffffffffffff1ffffffffffffffebffffffff0000000300000000",
            INIT_12 => X"ffffffb6fffffffffffffff2fffffffffffffffbffffffffffffffdaffffffff",
            INIT_13 => X"0000000900000000ffffffeaffffffff00000000000000000000001b00000000",
            INIT_14 => X"ffffffe3ffffffff00000007000000000000000c00000000ffffffeaffffffff",
            INIT_15 => X"ffffffedffffffffffffffd2ffffffff0000000200000000fffffffeffffffff",
            INIT_16 => X"ffffffe5ffffffffffffffdefffffffffffffffcffffffffffffffddffffffff",
            INIT_17 => X"0000000f000000000000000a0000000000000006000000000000003300000000",
            INIT_18 => X"ffffffedffffffff00000005000000000000000300000000fffffff4ffffffff",
            INIT_19 => X"fffffffdffffffff000000000000000000000005000000000000001200000000",
            INIT_1A => X"00000000000000000000003200000000ffffffeeffffffffffffffe4ffffffff",
            INIT_1B => X"ffffffd8ffffffffffffffd6ffffffffffffffdcffffffffffffffc2ffffffff",
            INIT_1C => X"ffffffd8ffffffff00000012000000000000001e000000000000000400000000",
            INIT_1D => X"0000003100000000fffffff8fffffffffffffffcfffffffffffffffdffffffff",
            INIT_1E => X"ffffffdaffffffff00000048000000000000000d000000000000001a00000000",
            INIT_1F => X"0000000500000000ffffffe2ffffffffffffffdbffffffff0000004600000000",
            INIT_20 => X"00000014000000000000001b00000000ffffffeffffffffffffffffdffffffff",
            INIT_21 => X"ffffff99ffffffffffffffc0ffffffff0000000200000000ffffffe0ffffffff",
            INIT_22 => X"0000000800000000ffffffddfffffffffffffffffffffffffffffff2ffffffff",
            INIT_23 => X"00000000000000000000002b000000000000002b000000000000003400000000",
            INIT_24 => X"ffffffc6ffffffffffffffc7ffffffffffffffd3fffffffffffffff5ffffffff",
            INIT_25 => X"00000009000000000000000d00000000fffffffefffffffffffffff7ffffffff",
            INIT_26 => X"0000002b00000000000000080000000000000012000000000000000100000000",
            INIT_27 => X"ffffffe3ffffffffffffffe0ffffffffffffffedfffffffffffffffcffffffff",
            INIT_28 => X"0000001500000000ffffffdcffffffff0000000a00000000fffffffaffffffff",
            INIT_29 => X"fffffff2fffffffffffffffcffffffffffffffdcffffffffffffffebffffffff",
            INIT_2A => X"ffffffe0ffffffffffffffabffffffffffffffddffffffffffffffd5ffffffff",
            INIT_2B => X"ffffffe1fffffffffffffff4fffffffffffffff0ffffffff0000001800000000",
            INIT_2C => X"ffffffe3fffffffffffffff0fffffffffffffff3ffffffffffffffe6ffffffff",
            INIT_2D => X"fffffffdfffffffffffffff8ffffffffffffffceffffffff0000000e00000000",
            INIT_2E => X"ffffffeafffffffffffffffdffffffff00000016000000000000001000000000",
            INIT_2F => X"fffffff0ffffffff000000050000000000000000000000000000000300000000",
            INIT_30 => X"000000040000000000000029000000000000002200000000ffffffe5ffffffff",
            INIT_31 => X"0000002e00000000ffffffe3ffffffff0000000b000000000000003200000000",
            INIT_32 => X"ffffffeaffffffffffffffd1ffffffff00000010000000000000001000000000",
            INIT_33 => X"0000002c000000000000001a0000000000000009000000000000000a00000000",
            INIT_34 => X"ffffffddfffffffffffffffaffffffff0000000900000000fffffffbffffffff",
            INIT_35 => X"ffffffe6fffffffffffffff2fffffffffffffffaffffffffffffffd0ffffffff",
            INIT_36 => X"ffffffd9fffffffffffffffcfffffffffffffff7ffffffff0000002600000000",
            INIT_37 => X"ffffffe1ffffffff0000001b000000000000000f000000000000001700000000",
            INIT_38 => X"0000000d00000000fffffff9ffffffff00000017000000000000001700000000",
            INIT_39 => X"ffffffe2ffffffff0000005b000000000000002d000000000000003200000000",
            INIT_3A => X"0000001400000000ffffffb9ffffffff00000002000000000000001400000000",
            INIT_3B => X"ffffffe3fffffffffffffff8ffffffffffffffe9ffffffff0000000600000000",
            INIT_3C => X"fffffffdfffffffffffffff9ffffffffffffffcdffffffff0000000c00000000",
            INIT_3D => X"fffffff8ffffffff00000014000000000000002800000000ffffffe2ffffffff",
            INIT_3E => X"0000000400000000ffffffe2ffffffff00000035000000000000000500000000",
            INIT_3F => X"0000001000000000fffffffbfffffffffffffff7ffffffff0000001800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001100000000ffffffebffffffff0000000400000000fffffff8ffffffff",
            INIT_41 => X"fffffff6fffffffffffffffaffffffff0000000d000000000000000d00000000",
            INIT_42 => X"fffffff9fffffffffffffff5fffffffffffffff6ffffffff0000000500000000",
            INIT_43 => X"00000010000000000000000500000000fffffffbffffffff0000001300000000",
            INIT_44 => X"fffffff7fffffffffffffff4ffffffff00000007000000000000001300000000",
            INIT_45 => X"0000000b00000000fffffff6ffffffff0000000d000000000000000400000000",
            INIT_46 => X"00000006000000000000000300000000ffffffe2ffffffffffffffe7ffffffff",
            INIT_47 => X"ffffffe4fffffffffffffff0ffffffffffffffe3ffffffff0000000200000000",
            INIT_48 => X"0000000200000000fffffffcffffffffffffffe4fffffffffffffffdffffffff",
            INIT_49 => X"fffffff5ffffffffffffffe1fffffffffffffff8ffffffff0000001300000000",
            INIT_4A => X"ffffffe8ffffffff0000000000000000ffffffeaffffffff0000000500000000",
            INIT_4B => X"0000001300000000ffffffedfffffffffffffff9fffffffffffffff1ffffffff",
            INIT_4C => X"00000012000000000000001300000000fffffff8ffffffffffffffe9ffffffff",
            INIT_4D => X"0000000200000000fffffffaffffffff0000000e00000000fffffff9ffffffff",
            INIT_4E => X"ffffffe8fffffffffffffff8ffffffffffffffeafffffffffffffffbffffffff",
            INIT_4F => X"ffffffeffffffffffffffff6ffffffff0000000a000000000000001100000000",
            INIT_50 => X"0000000e0000000000000012000000000000000300000000fffffff4ffffffff",
            INIT_51 => X"ffffffeefffffffffffffffbffffffff0000000800000000ffffffe5ffffffff",
            INIT_52 => X"fffffffaffffffff0000000d0000000000000009000000000000000400000000",
            INIT_53 => X"0000000300000000fffffff1ffffffffffffffeeffffffff0000000000000000",
            INIT_54 => X"0000001000000000000000070000000000000006000000000000000500000000",
            INIT_55 => X"0000000c000000000000000000000000ffffffe8fffffffffffffffbffffffff",
            INIT_56 => X"0000000f000000000000000100000000fffffff8ffffffff0000000300000000",
            INIT_57 => X"ffffffe4ffffffffffffffecfffffffffffffff4ffffffffffffffe9ffffffff",
            INIT_58 => X"0000000d00000000ffffffe2ffffffffffffffeeffffffff0000000c00000000",
            INIT_59 => X"fffffffbffffffff0000000b000000000000000000000000ffffffe8ffffffff",
            INIT_5A => X"0000000800000000fffffffbffffffff0000000d00000000ffffffebffffffff",
            INIT_5B => X"0000001800000000fffffff2fffffffffffffffcffffffffffffffefffffffff",
            INIT_5C => X"0000000500000000ffffffedfffffffffffffff7fffffffffffffff8ffffffff",
            INIT_5D => X"0000001100000000fffffff8ffffffffffffffeafffffffffffffff0ffffffff",
            INIT_5E => X"fffffff9ffffffff0000000200000000fffffffffffffffffffffff9ffffffff",
            INIT_5F => X"00000007000000000000000300000000fffffff3fffffffffffffffeffffffff",
            INIT_60 => X"0000000b00000000fffffff6fffffffffffffffeffffffff0000000b00000000",
            INIT_61 => X"0000000c00000000fffffff5fffffffffffffffaffffffff0000000e00000000",
            INIT_62 => X"fffffff0ffffffffffffffffffffffffffffffe5fffffffffffffff9ffffffff",
            INIT_63 => X"ffffffe8fffffffffffffff4fffffffffffffffafffffffffffffff0ffffffff",
            INIT_64 => X"fffffffcfffffffffffffffdfffffffffffffff4fffffffffffffff8ffffffff",
            INIT_65 => X"fffffffdfffffffffffffffefffffffffffffff7ffffffff0000000500000000",
            INIT_66 => X"0000000b00000000ffffffe3fffffffffffffffafffffffffffffff3ffffffff",
            INIT_67 => X"fffffff8ffffffff0000000f00000000fffffff5fffffffffffffffbffffffff",
            INIT_68 => X"ffffffe7ffffffff000000000000000000000009000000000000000800000000",
            INIT_69 => X"fffffffdffffffff000000050000000000000002000000000000000b00000000",
            INIT_6A => X"fffffff0ffffffffffffffe2ffffffffffffffeeffffffffffffffeaffffffff",
            INIT_6B => X"0000000200000000fffffff6fffffffffffffff3fffffffffffffffcffffffff",
            INIT_6C => X"fffffff8fffffffffffffffbfffffffffffffff2ffffffff0000001300000000",
            INIT_6D => X"0000000c00000000fffffff5fffffffffffffffefffffffffffffff1ffffffff",
            INIT_6E => X"ffffffffffffffff0000000e00000000fffffffffffffffffffffff9ffffffff",
            INIT_6F => X"fffffffaffffffff0000000000000000ffffffeeffffffff0000000300000000",
            INIT_70 => X"ffffffe3ffffffffffffffe2ffffffffffffffffffffffffffffffecffffffff",
            INIT_71 => X"fffffff3fffffffffffffff7fffffffffffffff4ffffffffffffffe2ffffffff",
            INIT_72 => X"ffffffeaffffffff0000000b00000000ffffffe6ffffffff0000000000000000",
            INIT_73 => X"ffffffeafffffffffffffff9ffffffff0000000b00000000ffffffebffffffff",
            INIT_74 => X"0000001200000000fffffff6fffffffffffffffaffffffff0000000900000000",
            INIT_75 => X"ffffffecfffffffffffffff8ffffffffffffffedffffffffffffffecffffffff",
            INIT_76 => X"fffffff4ffffffff0000000c0000000000000001000000000000000000000000",
            INIT_77 => X"fffffff2ffffffff0000000200000000fffffffbfffffffffffffff0ffffffff",
            INIT_78 => X"fffffffaffffffff00000003000000000000000800000000fffffffaffffffff",
            INIT_79 => X"0000000f00000000fffffff0ffffffffffffffeefffffffffffffffdffffffff",
            INIT_7A => X"fffffff8ffffffff0000001200000000fffffffefffffffffffffffeffffffff",
            INIT_7B => X"0000000400000000fffffffdfffffffffffffff5ffffffffffffffe8ffffffff",
            INIT_7C => X"fffffff2ffffffffffffffe9fffffffffffffff8fffffffffffffff2ffffffff",
            INIT_7D => X"0000000c00000000fffffffaffffffff0000000d000000000000000f00000000",
            INIT_7E => X"0000000e000000000000000100000000fffffff9ffffffffffffffe9ffffffff",
            INIT_7F => X"fffffff1ffffffff0000000c0000000000000004000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE30;


    MEM_IWGHT_LAYER2_INSTANCE31 : if BRAM_NAME = "iwght_layer2_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffdfffffffffffffffafffffffffffffffafffffffffffffff5ffffffff",
            INIT_01 => X"0000000000000000ffffffeaffffffff0000000000000000fffffff7ffffffff",
            INIT_02 => X"000000030000000000000008000000000000000000000000ffffffeaffffffff",
            INIT_03 => X"fffffffdffffffff000000070000000000000011000000000000000600000000",
            INIT_04 => X"fffffff5fffffffffffffff0ffffffff00000010000000000000000900000000",
            INIT_05 => X"fffffff7ffffffffffffffe7fffffffffffffff0ffffffff0000000a00000000",
            INIT_06 => X"fffffffaffffffff0000000c0000000000000001000000000000000000000000",
            INIT_07 => X"ffffffe1ffffffffffffffecffffffff00000001000000000000000200000000",
            INIT_08 => X"0000002000000000fffffff3ffffffffffffffd4ffffffffffffffc8ffffffff",
            INIT_09 => X"0000001e000000000000002d0000000000000015000000000000000900000000",
            INIT_0A => X"0000000000000000fffffff5fffffffffffffff1ffffffff0000003f00000000",
            INIT_0B => X"fffffff6ffffffff0000002500000000ffffffb9ffffffffffffffc5ffffffff",
            INIT_0C => X"0000002900000000000000260000000000000000000000000000001900000000",
            INIT_0D => X"fffffff7ffffffff000000070000000000000024000000000000000000000000",
            INIT_0E => X"0000001200000000fffffff3ffffffff00000031000000000000001500000000",
            INIT_0F => X"0000000b00000000000000000000000000000010000000000000000700000000",
            INIT_10 => X"00000019000000000000001000000000ffffffe2ffffffff0000003600000000",
            INIT_11 => X"000000000000000000000011000000000000002a000000000000000500000000",
            INIT_12 => X"0000001f00000000ffffffd8ffffffff0000003000000000fffffff0ffffffff",
            INIT_13 => X"fffffffafffffffffffffffdffffffff00000014000000000000000c00000000",
            INIT_14 => X"00000024000000000000001500000000ffffffe0ffffffff0000001c00000000",
            INIT_15 => X"fffffff8ffffffffffffffe8ffffffffffffffecffffffff0000001c00000000",
            INIT_16 => X"ffffffd9ffffffffffffffeeffffffff00000000000000000000000c00000000",
            INIT_17 => X"ffffffa5fffffffffffffffdffffffffffffffd7ffffffff0000004100000000",
            INIT_18 => X"ffffffeaffffffffffffffd7ffffffff0000001500000000ffffffbeffffffff",
            INIT_19 => X"0000001200000000000000090000000000000012000000000000002d00000000",
            INIT_1A => X"00000006000000000000001800000000fffffffffffffffffffffff9ffffffff",
            INIT_1B => X"0000000e00000000fffffff5ffffffff00000003000000000000000300000000",
            INIT_1C => X"000000340000000000000015000000000000003200000000fffffffdffffffff",
            INIT_1D => X"0000001f00000000fffffff5ffffffff00000022000000000000000b00000000",
            INIT_1E => X"ffffffbfffffffffffffffc3ffffffff00000008000000000000002200000000",
            INIT_1F => X"0000002200000000ffffffe3ffffffff00000004000000000000000000000000",
            INIT_20 => X"ffffffedffffffff00000037000000000000001c000000000000000c00000000",
            INIT_21 => X"ffffffbfffffffffffffffd7ffffffff0000000200000000fffffffdffffffff",
            INIT_22 => X"ffffffc2ffffffff00000009000000000000000300000000ffffffd1ffffffff",
            INIT_23 => X"ffffffdcfffffffffffffffdffffffffffffffdeffffffffffffffcfffffffff",
            INIT_24 => X"000000050000000000000015000000000000000000000000ffffffd9ffffffff",
            INIT_25 => X"fffffffdfffffffffffffff4ffffffffffffffeaffffffffffffffe3ffffffff",
            INIT_26 => X"ffffffdfffffffffffffffdbffffffffffffffd9fffffffffffffff2ffffffff",
            INIT_27 => X"fffffff2ffffffff00000001000000000000000600000000ffffffdeffffffff",
            INIT_28 => X"fffffff1ffffffff0000000b00000000ffffffedffffffff0000001000000000",
            INIT_29 => X"ffffffadffffffff00000000000000000000000d000000000000001100000000",
            INIT_2A => X"0000001100000000ffffffe0ffffffffffffffd9ffffffffffffffe4ffffffff",
            INIT_2B => X"0000000300000000ffffff93ffffffff0000003f00000000fffffff4ffffffff",
            INIT_2C => X"00000000000000000000000f0000000000000031000000000000002e00000000",
            INIT_2D => X"0000000900000000fffffff4fffffffffffffffaffffffff0000002800000000",
            INIT_2E => X"0000002700000000fffffffaffffffffffffffe5ffffffff0000000a00000000",
            INIT_2F => X"ffffffe9ffffffff0000001000000000fffffff7fffffffffffffff7ffffffff",
            INIT_30 => X"ffffffdaffffffffffffffdafffffffffffffffdffffffff0000000000000000",
            INIT_31 => X"ffffffc1ffffffffffffffa9ffffffffffffffe3ffffffffffffffe4ffffffff",
            INIT_32 => X"0000002400000000ffffffe4ffffffffffffffe6ffffffffffffffd9ffffffff",
            INIT_33 => X"00000009000000000000001b000000000000000c000000000000000500000000",
            INIT_34 => X"00000025000000000000001700000000ffffffe0ffffffff0000002e00000000",
            INIT_35 => X"0000000b0000000000000030000000000000001f00000000fffffff7ffffffff",
            INIT_36 => X"fffffff4ffffffff0000001e000000000000000100000000fffffff9ffffffff",
            INIT_37 => X"ffffffebfffffffffffffffdffffffffffffffeafffffffffffffff3ffffffff",
            INIT_38 => X"0000003c00000000ffffffe3ffffffff00000011000000000000001200000000",
            INIT_39 => X"ffffffd5ffffffffffffffe6ffffffff0000000f00000000ffffffbbffffffff",
            INIT_3A => X"0000000300000000ffffffdafffffffffffffff9ffffffff0000001400000000",
            INIT_3B => X"ffffffe2fffffffffffffff5ffffffffffffffe7fffffffffffffffdffffffff",
            INIT_3C => X"00000001000000000000000d00000000fffffffcffffffffffffffbfffffffff",
            INIT_3D => X"0000000f000000000000000d000000000000002c000000000000000600000000",
            INIT_3E => X"ffffffc3ffffffff0000002b00000000fffffffafffffffffffffff6ffffffff",
            INIT_3F => X"ffffffdcffffffff00000019000000000000001c00000000fffffff8ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001f000000000000001a00000000fffffffdffffffff0000000900000000",
            INIT_41 => X"0000002c0000000000000022000000000000000f000000000000002700000000",
            INIT_42 => X"0000000000000000ffffffedffffffff0000003d000000000000003500000000",
            INIT_43 => X"0000000c00000000ffffffe6ffffffffffffffffffffffff0000001300000000",
            INIT_44 => X"fffffffbffffffff000000120000000000000000000000000000001d00000000",
            INIT_45 => X"ffffffcefffffffffffffff3ffffffffffffffc9ffffffffffffffc7ffffffff",
            INIT_46 => X"00000000000000000000002a0000000000000021000000000000000c00000000",
            INIT_47 => X"fffffffaffffffff00000000000000000000003e000000000000002e00000000",
            INIT_48 => X"0000000800000000fffffff6ffffffff00000006000000000000001500000000",
            INIT_49 => X"ffffffbeffffffff0000001500000000fffffff2ffffffff0000000800000000",
            INIT_4A => X"ffffffe4ffffffffffffffe1ffffffffffffffd1fffffffffffffffaffffffff",
            INIT_4B => X"00000024000000000000001200000000fffffffeffffffff0000001e00000000",
            INIT_4C => X"00000000000000000000000a00000000ffffffe2ffffffff0000002e00000000",
            INIT_4D => X"ffffffdfffffffff0000000500000000ffffffdfffffffffffffffe0ffffffff",
            INIT_4E => X"fffffff2ffffffff00000008000000000000000400000000fffffff8ffffffff",
            INIT_4F => X"0000002700000000ffffffb5ffffffff00000013000000000000000e00000000",
            INIT_50 => X"0000001300000000fffffffaffffffff0000000e000000000000000600000000",
            INIT_51 => X"fffffff7fffffffffffffff2fffffffffffffffdfffffffffffffff6ffffffff",
            INIT_52 => X"ffffffe9ffffffff0000002d00000000ffffffcbffffffff0000000f00000000",
            INIT_53 => X"ffffffe8ffffffffffffffbeffffffffffffffd4ffffffffffffffa6ffffffff",
            INIT_54 => X"00000018000000000000000000000000ffffffcdffffffffffffffc4ffffffff",
            INIT_55 => X"ffffffcffffffffffffffffbfffffffffffffffaffffffffffffffffffffffff",
            INIT_56 => X"0000000000000000fffffff9ffffffffffffffd9ffffffff0000001d00000000",
            INIT_57 => X"ffffffb1ffffffffffffff99ffffffffffffffdbffffffffffffffd4ffffffff",
            INIT_58 => X"ffffffc6ffffffffffffffbcffffffffffffffcbfffffffffffffffeffffffff",
            INIT_59 => X"ffffffe7ffffffffffffffefffffffffffffffc5ffffffffffffffe8ffffffff",
            INIT_5A => X"ffffffe2ffffffff0000000100000000fffffffeffffffff0000000700000000",
            INIT_5B => X"0000000000000000ffffffe1ffffffffffffffd2ffffffff0000000000000000",
            INIT_5C => X"0000003f00000000ffffffe8fffffffffffffff3ffffffff0000000a00000000",
            INIT_5D => X"0000002c000000000000001800000000ffffffeeffffffff0000001300000000",
            INIT_5E => X"ffffffd1fffffffffffffff2fffffffffffffff1ffffffff0000000e00000000",
            INIT_5F => X"fffffffaffffffff0000000a0000000000000014000000000000000500000000",
            INIT_60 => X"0000000f000000000000000700000000fffffff2ffffffffffffffebffffffff",
            INIT_61 => X"ffffffe9ffffffffffffffdfffffffff0000000a00000000ffffffedffffffff",
            INIT_62 => X"ffffffd9ffffffff0000001600000000ffffffcfffffffff0000000900000000",
            INIT_63 => X"ffffffd0ffffffffffffffceffffffffffffffc1ffffffffffffffd9ffffffff",
            INIT_64 => X"0000000c0000000000000017000000000000000800000000ffffffe3ffffffff",
            INIT_65 => X"00000040000000000000000f0000000000000032000000000000002400000000",
            INIT_66 => X"fffffffbffffffff000000020000000000000025000000000000000200000000",
            INIT_67 => X"00000024000000000000001b000000000000000400000000ffffffffffffffff",
            INIT_68 => X"0000003300000000fffffffcffffffff00000025000000000000000100000000",
            INIT_69 => X"fffffff8ffffffff0000002a0000000000000015000000000000003700000000",
            INIT_6A => X"000000010000000000000002000000000000000e000000000000001600000000",
            INIT_6B => X"ffffffebffffffffffffffaffffffffffffffff2ffffffff0000003600000000",
            INIT_6C => X"0000000900000000fffffff8ffffffffffffffedffffffff0000001600000000",
            INIT_6D => X"ffffffecffffffff0000000c0000000000000027000000000000000400000000",
            INIT_6E => X"0000000c00000000fffffffaffffffff00000022000000000000001500000000",
            INIT_6F => X"fffffff9ffffffff000000120000000000000002000000000000001200000000",
            INIT_70 => X"fffffffbffffffff00000005000000000000000c00000000fffffff6ffffffff",
            INIT_71 => X"0000002100000000fffffff0fffffffffffffff1ffffffffffffffecffffffff",
            INIT_72 => X"ffffffe2fffffffffffffff4fffffffffffffff1ffffffff0000000100000000",
            INIT_73 => X"0000001a000000000000000d000000000000000600000000fffffff3ffffffff",
            INIT_74 => X"0000001100000000fffffff7ffffffff00000015000000000000000900000000",
            INIT_75 => X"00000014000000000000000800000000fffffffeffffffff0000000d00000000",
            INIT_76 => X"0000000f00000000fffffff7ffffffffffffffb4fffffffffffffffcffffffff",
            INIT_77 => X"0000000e000000000000001400000000fffffffefffffffffffffffaffffffff",
            INIT_78 => X"000000080000000000000000000000000000001c000000000000002700000000",
            INIT_79 => X"ffffffecfffffffffffffffafffffffffffffff2ffffffff0000003900000000",
            INIT_7A => X"0000000300000000ffffffd2ffffffffffffffecfffffffffffffffeffffffff",
            INIT_7B => X"fffffff5ffffffffffffffdeffffffff0000002600000000ffffffcbffffffff",
            INIT_7C => X"0000002c000000000000003900000000ffffffd2ffffffffffffffdcffffffff",
            INIT_7D => X"fffffff4ffffffff0000001c000000000000000300000000ffffffd7ffffffff",
            INIT_7E => X"fffffff5ffffffffffffffecffffffff0000002d000000000000000d00000000",
            INIT_7F => X"fffffff8ffffffff000000090000000000000014000000000000001e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE31;


    MEM_IWGHT_LAYER2_INSTANCE32 : if BRAM_NAME = "iwght_layer2_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffffffffffffffffffe2ffffffffffffffe4ffffffff0000002f00000000",
            INIT_01 => X"0000001d0000000000000000000000000000000e00000000ffffffe0ffffffff",
            INIT_02 => X"00000013000000000000001e0000000000000010000000000000001500000000",
            INIT_03 => X"ffffffddffffffff000000020000000000000024000000000000003400000000",
            INIT_04 => X"fffffff2ffffffffffffffcdffffffff0000002d00000000fffffff3ffffffff",
            INIT_05 => X"0000002500000000fffffffcffffffffffffffd3ffffffff0000001800000000",
            INIT_06 => X"ffffffefffffffff0000000d000000000000002500000000fffffff8ffffffff",
            INIT_07 => X"fffffff8fffffffffffffff4ffffffff0000001b00000000fffffff3ffffffff",
            INIT_08 => X"fffffff2ffffffff0000000300000000ffffffe5ffffffff0000001200000000",
            INIT_09 => X"00000026000000000000000d00000000ffffffffffffffffffffffebffffffff",
            INIT_0A => X"fffffff6ffffffffffffffe4ffffffff00000021000000000000001300000000",
            INIT_0B => X"0000000c00000000ffffffd3ffffffffffffffeeffffffff0000002600000000",
            INIT_0C => X"fffffffcffffffffffffffe2ffffffffffffffceffffffffffffffd0ffffffff",
            INIT_0D => X"fffffff6ffffffffffffffdffffffffffffffffbffffffff0000000f00000000",
            INIT_0E => X"0000002f000000000000000000000000ffffffcdffffffff0000002700000000",
            INIT_0F => X"0000000100000000000000030000000000000012000000000000002b00000000",
            INIT_10 => X"fffffffdfffffffffffffff1fffffffffffffffdffffffffffffffe6ffffffff",
            INIT_11 => X"ffffffe7ffffffff000000530000000000000046000000000000000300000000",
            INIT_12 => X"fffffff3ffffffffffffffd1ffffffffffffffe6fffffffffffffffbffffffff",
            INIT_13 => X"00000021000000000000002000000000ffffffefffffffffffffffd5ffffffff",
            INIT_14 => X"0000001200000000fffffff8ffffffff00000000000000000000000e00000000",
            INIT_15 => X"0000003e000000000000000400000000fffffffcfffffffffffffffeffffffff",
            INIT_16 => X"fffffff5ffffffff0000000000000000fffffff4fffffffffffffff7ffffffff",
            INIT_17 => X"fffffff3ffffffffffffffe6ffffffffffffffe0ffffffff0000000a00000000",
            INIT_18 => X"0000000400000000ffffffefffffffffffffffecfffffffffffffffdffffffff",
            INIT_19 => X"00000001000000000000000f000000000000000f000000000000000b00000000",
            INIT_1A => X"ffffffffffffffff00000005000000000000000900000000fffffff6ffffffff",
            INIT_1B => X"0000000500000000ffffffeffffffffffffffffaffffffff0000001200000000",
            INIT_1C => X"0000000500000000000000030000000000000005000000000000000500000000",
            INIT_1D => X"0000000c00000000ffffffebfffffffffffffffcffffffffffffffffffffffff",
            INIT_1E => X"fffffffdffffffff0000000300000000ffffffe8ffffffffffffffefffffffff",
            INIT_1F => X"00000006000000000000000600000000fffffffbffffffffffffffecffffffff",
            INIT_20 => X"000000080000000000000008000000000000000100000000fffffff7ffffffff",
            INIT_21 => X"ffffffedffffffffffffffeaffffffff0000000f00000000fffffff8ffffffff",
            INIT_22 => X"0000000d00000000ffffffedfffffffffffffffcfffffffffffffff5ffffffff",
            INIT_23 => X"0000000700000000fffffffbfffffffffffffffefffffffffffffffaffffffff",
            INIT_24 => X"fffffff5fffffffffffffff7fffffffffffffffefffffffffffffffaffffffff",
            INIT_25 => X"fffffffaffffffff0000000800000000ffffffeaffffffff0000000900000000",
            INIT_26 => X"ffffffecffffffffffffffe4ffffffff0000000700000000fffffff0ffffffff",
            INIT_27 => X"fffffff3fffffffffffffff6fffffffffffffff3ffffffff0000000000000000",
            INIT_28 => X"ffffffffffffffffffffffe9ffffffff0000000b000000000000000700000000",
            INIT_29 => X"fffffff2ffffffffffffffedffffffff0000000b00000000ffffffeaffffffff",
            INIT_2A => X"fffffff6ffffffff0000000c00000000ffffffe3ffffffff0000000a00000000",
            INIT_2B => X"ffffffebfffffffffffffff3ffffffffffffffeeffffffff0000000c00000000",
            INIT_2C => X"000000000000000000000008000000000000000700000000ffffffe9ffffffff",
            INIT_2D => X"00000005000000000000000300000000ffffffe9fffffffffffffffbffffffff",
            INIT_2E => X"ffffffe4fffffffffffffff0ffffffff00000010000000000000000c00000000",
            INIT_2F => X"fffffff1fffffffffffffff0fffffffffffffffdffffffff0000000400000000",
            INIT_30 => X"0000000000000000fffffff0ffffffff0000000900000000ffffffebffffffff",
            INIT_31 => X"fffffffaffffffff0000000a0000000000000005000000000000000300000000",
            INIT_32 => X"0000000300000000fffffffcfffffffffffffff3ffffffffffffffefffffffff",
            INIT_33 => X"000000070000000000000012000000000000001100000000fffffff0ffffffff",
            INIT_34 => X"ffffffffffffffff0000000d00000000ffffffefffffffffffffffecffffffff",
            INIT_35 => X"ffffffeefffffffffffffff2ffffffffffffffe8ffffffff0000000500000000",
            INIT_36 => X"fffffffefffffffffffffff9ffffffff0000000b00000000fffffffeffffffff",
            INIT_37 => X"fffffff6ffffffff0000000900000000ffffffedffffffff0000000f00000000",
            INIT_38 => X"ffffffeffffffffffffffffaffffffff0000000100000000fffffff7ffffffff",
            INIT_39 => X"0000000b000000000000000200000000ffffffecfffffffffffffff4ffffffff",
            INIT_3A => X"fffffff8ffffffff00000007000000000000000300000000fffffff8ffffffff",
            INIT_3B => X"ffffffebffffffff0000000500000000ffffffeefffffffffffffff4ffffffff",
            INIT_3C => X"fffffff0ffffffff00000002000000000000000900000000fffffffcffffffff",
            INIT_3D => X"fffffffaffffffffffffffeefffffffffffffff4ffffffff0000000400000000",
            INIT_3E => X"00000008000000000000000900000000fffffff5ffffffff0000000200000000",
            INIT_3F => X"fffffffdffffffff0000000b000000000000000b000000000000000d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff3fffffffffffffff6fffffffffffffffafffffffffffffffaffffffff",
            INIT_41 => X"fffffffbffffffff00000005000000000000000d000000000000000700000000",
            INIT_42 => X"0000000500000000fffffffffffffffffffffff1ffffffffffffffeaffffffff",
            INIT_43 => X"fffffff3ffffffff0000000000000000fffffffeffffffff0000000300000000",
            INIT_44 => X"0000000800000000fffffff6ffffffff0000000b00000000ffffffffffffffff",
            INIT_45 => X"ffffffebffffffffffffffecffffffff0000000900000000ffffffeeffffffff",
            INIT_46 => X"fffffff1ffffffffffffffebfffffffffffffff0fffffffffffffff3ffffffff",
            INIT_47 => X"0000000100000000000000010000000000000010000000000000000000000000",
            INIT_48 => X"0000001100000000fffffff7fffffffffffffff2ffffffffffffffeeffffffff",
            INIT_49 => X"0000000100000000fffffff1fffffffffffffff6ffffffffffffffe7ffffffff",
            INIT_4A => X"00000001000000000000000b00000000fffffffeffffffff0000000100000000",
            INIT_4B => X"ffffffeefffffffffffffffbfffffffffffffff7ffffffffffffffffffffffff",
            INIT_4C => X"0000000100000000fffffff9ffffffff0000000000000000fffffff3ffffffff",
            INIT_4D => X"ffffffffffffffff0000000300000000fffffff4ffffffff0000001300000000",
            INIT_4E => X"0000000800000000ffffffecffffffff0000000000000000ffffffeaffffffff",
            INIT_4F => X"0000000d000000000000000200000000ffffffe9ffffffffffffffe9ffffffff",
            INIT_50 => X"fffffff1fffffffffffffff8ffffffff00000003000000000000000f00000000",
            INIT_51 => X"fffffff3ffffffffffffffecffffffff0000000200000000ffffffeeffffffff",
            INIT_52 => X"fffffff4fffffffffffffffcffffffff0000000a000000000000000300000000",
            INIT_53 => X"ffffffefffffffffffffffecffffffff00000000000000000000000000000000",
            INIT_54 => X"0000000500000000fffffff3ffffffff0000000900000000fffffff3ffffffff",
            INIT_55 => X"fffffffdfffffffffffffffdffffffffffffffebffffffff0000001100000000",
            INIT_56 => X"00000002000000000000000700000000ffffffedffffffff0000001100000000",
            INIT_57 => X"fffffffdffffffff0000000b000000000000000b00000000ffffffeeffffffff",
            INIT_58 => X"0000000a0000000000000006000000000000000400000000ffffffeeffffffff",
            INIT_59 => X"0000000100000000fffffff9fffffffffffffffcffffffff0000000500000000",
            INIT_5A => X"fffffff4fffffffffffffff7ffffffff0000000f00000000fffffff2ffffffff",
            INIT_5B => X"fffffffbffffffffffffffefffffffffffffffebffffffff0000000400000000",
            INIT_5C => X"fffffff2fffffffffffffff4fffffffffffffff1ffffffff0000000d00000000",
            INIT_5D => X"ffffffebffffffffffffffe5fffffffffffffff5ffffffff0000000700000000",
            INIT_5E => X"ffffffe8ffffffffffffffebffffffff0000000700000000ffffffe1ffffffff",
            INIT_5F => X"0000000a00000000fffffff3fffffffffffffff3ffffffff0000000500000000",
            INIT_60 => X"0000000700000000fffffff0fffffffffffffff8ffffffff0000000100000000",
            INIT_61 => X"fffffff8ffffffffffffffeeffffffff00000018000000000000001500000000",
            INIT_62 => X"00000012000000000000001b000000000000000b00000000ffffffe0ffffffff",
            INIT_63 => X"00000029000000000000004b0000000000000047000000000000006b00000000",
            INIT_64 => X"000000100000000000000017000000000000000a000000000000001e00000000",
            INIT_65 => X"fffffffafffffffffffffff1fffffffffffffff1ffffffff0000000300000000",
            INIT_66 => X"0000000700000000ffffffcdffffffffffffffd4ffffffff0000001700000000",
            INIT_67 => X"ffffffecfffffffffffffff1ffffffff0000000d000000000000001a00000000",
            INIT_68 => X"0000002300000000fffffffbfffffffffffffffafffffffffffffff8ffffffff",
            INIT_69 => X"00000025000000000000001d000000000000000c000000000000001500000000",
            INIT_6A => X"0000000700000000000000140000000000000020000000000000001300000000",
            INIT_6B => X"0000000900000000fffffffbffffffff0000002600000000fffffffeffffffff",
            INIT_6C => X"00000009000000000000000800000000fffffff7ffffffff0000001500000000",
            INIT_6D => X"fffffff2fffffffffffffffbffffffff00000016000000000000000800000000",
            INIT_6E => X"00000015000000000000000b00000000fffffff2fffffffffffffff7ffffffff",
            INIT_6F => X"ffffffe1ffffffff0000000e00000000fffffff5ffffffff0000000200000000",
            INIT_70 => X"fffffff1fffffffffffffff2ffffffffffffffcbffffffffffffffcfffffffff",
            INIT_71 => X"fffffff4ffffffffffffffeeffffffffffffffffffffffff0000000c00000000",
            INIT_72 => X"0000001700000000fffffffbffffffff0000000700000000fffffff9ffffffff",
            INIT_73 => X"ffffffe8ffffffff0000001d0000000000000021000000000000000200000000",
            INIT_74 => X"0000001e00000000ffffffffffffffff0000001800000000fffffff1ffffffff",
            INIT_75 => X"fffffff4fffffffffffffff1fffffffffffffff3fffffffffffffff3ffffffff",
            INIT_76 => X"0000001100000000fffffffaffffffff0000002a000000000000000000000000",
            INIT_77 => X"00000012000000000000000c000000000000000100000000fffffffbffffffff",
            INIT_78 => X"ffffffeefffffffffffffffeffffffffffffffefffffffffffffffe0ffffffff",
            INIT_79 => X"ffffffe8ffffffff0000002600000000ffffffffffffffffffffffe6ffffffff",
            INIT_7A => X"0000001a000000000000001a0000000000000035000000000000001300000000",
            INIT_7B => X"fffffff8ffffffff0000002500000000fffffff3ffffffff0000000300000000",
            INIT_7C => X"ffffffe5ffffffff000000010000000000000023000000000000000d00000000",
            INIT_7D => X"0000000f00000000fffffffeffffffff00000036000000000000002b00000000",
            INIT_7E => X"ffffffe6ffffffff0000001500000000fffffffbffffffff0000000000000000",
            INIT_7F => X"fffffff2fffffffffffffffeffffffffffffffe9ffffffff0000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE32;


    MEM_IWGHT_LAYER2_INSTANCE33 : if BRAM_NAME = "iwght_layer2_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000800000000000000060000000000000009000000000000000600000000",
            INIT_01 => X"0000000000000000fffffff7ffffffff0000000e00000000fffffffdffffffff",
            INIT_02 => X"0000000000000000fffffff3ffffffffffffffebffffffff0000000100000000",
            INIT_03 => X"00000032000000000000002f000000000000002f00000000fffffffeffffffff",
            INIT_04 => X"000000080000000000000006000000000000000800000000ffffffecffffffff",
            INIT_05 => X"fffffff2ffffffffffffffd4fffffffffffffff8ffffffff0000000100000000",
            INIT_06 => X"fffffff3fffffffffffffffbffffffff0000000400000000ffffffedffffffff",
            INIT_07 => X"fffffff6ffffffff00000048000000000000003b000000000000003800000000",
            INIT_08 => X"ffffffd0fffffffffffffff0ffffffff00000010000000000000002f00000000",
            INIT_09 => X"ffffffc6ffffffffffffffe9fffffffffffffff8ffffffff0000000200000000",
            INIT_0A => X"ffffffbcffffffff00000000000000000000001c000000000000000900000000",
            INIT_0B => X"0000000b00000000fffffff4ffffffff0000000c00000000ffffffc4ffffffff",
            INIT_0C => X"00000036000000000000000e0000000000000002000000000000001300000000",
            INIT_0D => X"0000002200000000ffffffe7ffffffffffffffefffffffffffffffe7ffffffff",
            INIT_0E => X"0000001700000000000000190000000000000031000000000000003d00000000",
            INIT_0F => X"fffffff9ffffffff0000000300000000ffffffdbffffffff0000001000000000",
            INIT_10 => X"000000050000000000000038000000000000001a000000000000000800000000",
            INIT_11 => X"00000000000000000000000e00000000fffffffbfffffffffffffffeffffffff",
            INIT_12 => X"0000004d00000000000000300000000000000031000000000000000a00000000",
            INIT_13 => X"ffffffbeffffffff0000001c0000000000000038000000000000003100000000",
            INIT_14 => X"ffffffeeffffffffffffffd6ffffffff0000000300000000ffffffeaffffffff",
            INIT_15 => X"fffffffefffffffffffffff0ffffffff0000000400000000fffffff4ffffffff",
            INIT_16 => X"0000002f00000000fffffff7fffffffffffffffbffffffff0000000f00000000",
            INIT_17 => X"0000001b00000000000000460000000000000038000000000000002400000000",
            INIT_18 => X"0000000300000000000000150000000000000016000000000000002400000000",
            INIT_19 => X"0000001a0000000000000006000000000000001e000000000000002400000000",
            INIT_1A => X"fffffffefffffffffffffff6fffffffffffffff9ffffffff0000000700000000",
            INIT_1B => X"ffffffecffffffff0000000300000000fffffffbffffffff0000000500000000",
            INIT_1C => X"fffffffdffffffff00000006000000000000000100000000ffffffe4ffffffff",
            INIT_1D => X"ffffffecfffffffffffffffeffffffff00000027000000000000000300000000",
            INIT_1E => X"0000000800000000ffffffe8ffffffffffffffd7fffffffffffffffdffffffff",
            INIT_1F => X"ffffffe9ffffffff0000002000000000ffffffffffffffff0000000500000000",
            INIT_20 => X"fffffffbffffffffffffffe0fffffffffffffff4ffffffffffffffe2ffffffff",
            INIT_21 => X"0000003d0000000000000023000000000000002500000000ffffffe1ffffffff",
            INIT_22 => X"ffffffd8ffffffff0000002b00000000fffffff4ffffffffffffffe3ffffffff",
            INIT_23 => X"0000000800000000fffffffcffffffffffffffb5ffffffffffffffdaffffffff",
            INIT_24 => X"0000000b00000000fffffff9ffffffffffffffe4ffffffffffffffe7ffffffff",
            INIT_25 => X"fffffff2ffffffff00000004000000000000001900000000fffffff7ffffffff",
            INIT_26 => X"0000000500000000fffffff3ffffffff0000000500000000ffffffecffffffff",
            INIT_27 => X"0000001a000000000000000100000000ffffffe9ffffffff0000003200000000",
            INIT_28 => X"0000000600000000fffffff2ffffffff0000000d00000000fffffffbffffffff",
            INIT_29 => X"0000000600000000ffffffeaffffffff00000018000000000000000b00000000",
            INIT_2A => X"0000003000000000fffffff5ffffffffffffffe8ffffffff0000000c00000000",
            INIT_2B => X"000000620000000000000007000000000000003a00000000fffffff1ffffffff",
            INIT_2C => X"ffffffdeffffffffffffffc7ffffffff00000058000000000000006200000000",
            INIT_2D => X"ffffffdeffffffffffffffc5ffffffffffffffcaffffffffffffffdcffffffff",
            INIT_2E => X"0000001500000000fffffffcffffffffffffffe2ffffffffffffffddffffffff",
            INIT_2F => X"00000010000000000000000d00000000fffffff1ffffffff0000000200000000",
            INIT_30 => X"00000016000000000000001c00000000fffffff4ffffffff0000001600000000",
            INIT_31 => X"0000000c00000000fffffff3ffffffff0000001b000000000000003100000000",
            INIT_32 => X"fffffff3ffffffffffffffe8ffffffff0000001000000000ffffffebffffffff",
            INIT_33 => X"ffffffaaffffffffffffffc7fffffffffffffff4fffffffffffffff0ffffffff",
            INIT_34 => X"0000001200000000ffffffd2ffffffffffffffd2ffffffff0000000b00000000",
            INIT_35 => X"ffffffd3ffffffff0000000400000000ffffffaaffffffffffffffc4ffffffff",
            INIT_36 => X"ffffffd1ffffffffffffffacffffffffffffffc5ffffffffffffffbcffffffff",
            INIT_37 => X"ffffffeaffffffffffffffe2ffffffffffffffbbffffffffffffffe3ffffffff",
            INIT_38 => X"fffffffeffffffff0000001c000000000000000500000000fffffffbffffffff",
            INIT_39 => X"0000002e0000000000000016000000000000002a000000000000001000000000",
            INIT_3A => X"fffffffaffffffff000000180000000000000009000000000000001900000000",
            INIT_3B => X"fffffffaffffffff00000017000000000000001c000000000000000500000000",
            INIT_3C => X"0000002700000000ffffffd4fffffffffffffff5fffffffffffffffbffffffff",
            INIT_3D => X"0000000000000000ffffffd4ffffffffffffffcffffffffffffffffdffffffff",
            INIT_3E => X"0000000000000000ffffffe7ffffffffffffffeeffffffffffffffd8ffffffff",
            INIT_3F => X"00000000000000000000000600000000fffffff5ffffffff0000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff4ffffffff00000015000000000000001500000000ffffffdcffffffff",
            INIT_41 => X"ffffffc2ffffffffffffffb1ffffffffffffffd4fffffffffffffffeffffffff",
            INIT_42 => X"ffffffb3ffffffffffffff99ffffffffffffffb9ffffffffffffffa0ffffffff",
            INIT_43 => X"ffffffbdffffffff0000000600000000ffffffd5fffffffffffffff8ffffffff",
            INIT_44 => X"0000002c000000000000000000000000ffffffd5ffffffffffffffd3ffffffff",
            INIT_45 => X"ffffffe2ffffffffffffffebffffffff00000005000000000000001e00000000",
            INIT_46 => X"0000001000000000ffffffdcffffffffffffffe3ffffffff0000002c00000000",
            INIT_47 => X"ffffffedfffffffffffffff2ffffffffffffffffffffffffffffffbbffffffff",
            INIT_48 => X"00000010000000000000000700000000ffffffeffffffffffffffffeffffffff",
            INIT_49 => X"0000002600000000000000100000000000000013000000000000000900000000",
            INIT_4A => X"00000000000000000000002100000000fffffff4ffffffff0000000300000000",
            INIT_4B => X"ffffffd3fffffffffffffff8ffffffff0000002200000000ffffffe3ffffffff",
            INIT_4C => X"fffffff5ffffffff0000000c000000000000002c000000000000001600000000",
            INIT_4D => X"0000000d00000000000000040000000000000014000000000000001700000000",
            INIT_4E => X"ffffffdbffffffffffffffd8ffffffff00000003000000000000001f00000000",
            INIT_4F => X"fffffff2ffffffffffffffdbffffffffffffffd3ffffffffffffffffffffffff",
            INIT_50 => X"ffffffe7ffffffff0000001400000000ffffffdffffffffffffffffbffffffff",
            INIT_51 => X"0000000600000000fffffff8ffffffff00000015000000000000001100000000",
            INIT_52 => X"0000000100000000fffffff7ffffffff00000001000000000000002f00000000",
            INIT_53 => X"fffffff8ffffffffffffffffffffffffffffffe1ffffffff0000000000000000",
            INIT_54 => X"ffffffd7ffffffff0000000c00000000fffffffdfffffffffffffff9ffffffff",
            INIT_55 => X"000000030000000000000005000000000000002c000000000000002300000000",
            INIT_56 => X"0000000700000000000000300000000000000014000000000000000d00000000",
            INIT_57 => X"ffffffb8ffffffffffffffd8ffffffffffffffd0ffffffff0000000f00000000",
            INIT_58 => X"fffffffaffffffffffffffb4ffffffffffffffa6ffffffffffffffbaffffffff",
            INIT_59 => X"ffffffcdffffffffffffffe6ffffffffffffffd9ffffffffffffff8fffffffff",
            INIT_5A => X"ffffffe7ffffffffffffffcbffffffffffffffb4fffffffffffffff2ffffffff",
            INIT_5B => X"fffffffdffffffffffffffe1ffffffffffffffeafffffffffffffffdffffffff",
            INIT_5C => X"000000000000000000000015000000000000001400000000fffffffdffffffff",
            INIT_5D => X"0000001a000000000000002300000000ffffffe5ffffffff0000001400000000",
            INIT_5E => X"fffffffcffffffff000000060000000000000019000000000000001100000000",
            INIT_5F => X"ffffffdfffffffffffffffe4fffffffffffffff1ffffffff0000000b00000000",
            INIT_60 => X"ffffffdfffffffffffffffeeffffffff0000000200000000fffffff6ffffffff",
            INIT_61 => X"fffffffeffffffffffffffc2ffffffffffffffb5ffffffff0000002400000000",
            INIT_62 => X"00000005000000000000001100000000ffffffc8ffffffffffffffb3ffffffff",
            INIT_63 => X"0000000100000000fffffffeffffffff0000000200000000ffffffe5ffffffff",
            INIT_64 => X"000000040000000000000017000000000000002a000000000000000800000000",
            INIT_65 => X"fffffff2ffffffff00000016000000000000001200000000ffffffe6ffffffff",
            INIT_66 => X"ffffffe0ffffffff00000006000000000000000d000000000000001500000000",
            INIT_67 => X"0000001900000000000000250000000000000035000000000000001800000000",
            INIT_68 => X"0000001a0000000000000016000000000000001e000000000000001200000000",
            INIT_69 => X"ffffffdfffffffffffffffb2ffffffffffffffaeffffffff0000001300000000",
            INIT_6A => X"ffffffa7ffffffffffffffccffffffffffffff98ffffffffffffffd5ffffffff",
            INIT_6B => X"0000001f000000000000000d00000000ffffffb6ffffffffffffffb0ffffffff",
            INIT_6C => X"00000000000000000000000600000000fffffff8ffffffff0000002400000000",
            INIT_6D => X"fffffffcffffffff00000015000000000000000100000000ffffffe3ffffffff",
            INIT_6E => X"0000001f000000000000000a000000000000000f000000000000001400000000",
            INIT_6F => X"0000000b000000000000001300000000fffffff2fffffffffffffffbffffffff",
            INIT_70 => X"0000000e00000000ffffffe9ffffffffffffffd8ffffffffffffffd0ffffffff",
            INIT_71 => X"0000000e000000000000000e0000000000000000000000000000000800000000",
            INIT_72 => X"fffffff7ffffffffffffffc0ffffffffffffffe2fffffffffffffffcffffffff",
            INIT_73 => X"ffffffe7fffffffffffffffdffffffff0000001400000000fffffff8ffffffff",
            INIT_74 => X"00000015000000000000000200000000ffffffffffffffffffffffceffffffff",
            INIT_75 => X"ffffffe6ffffffffffffffc6ffffffff0000000500000000ffffffdcffffffff",
            INIT_76 => X"0000000200000000ffffffe6ffffffffffffffffffffffff0000000300000000",
            INIT_77 => X"fffffff3ffffffff000000020000000000000016000000000000000000000000",
            INIT_78 => X"00000052000000000000001e000000000000000e000000000000002400000000",
            INIT_79 => X"0000000900000000ffffffe8ffffffff0000000c000000000000001a00000000",
            INIT_7A => X"00000009000000000000000d00000000ffffffe7ffffffff0000000200000000",
            INIT_7B => X"ffffffbcffffffff0000001c000000000000002100000000fffffff2ffffffff",
            INIT_7C => X"ffffffe7ffffffffffffff79ffffffffffffffe1ffffffffffffffe6ffffffff",
            INIT_7D => X"ffffffe1fffffffffffffffbffffffffffffffb6ffffffffffffffc5ffffffff",
            INIT_7E => X"ffffffcbffffffffffffffeaffffffffffffffffffffffffffffffdeffffffff",
            INIT_7F => X"ffffffdffffffffffffffff3ffffffffffffffd7ffffffffffffffd2ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE33;


    MEM_IWGHT_LAYER2_INSTANCE34 : if BRAM_NAME = "iwght_layer2_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd8fffffffffffffff2ffffffff0000000000000000ffffffd7ffffffff",
            INIT_01 => X"0000000800000000ffffffe0fffffffffffffff8ffffffff0000001e00000000",
            INIT_02 => X"0000001500000000fffffff7ffffffff00000016000000000000000800000000",
            INIT_03 => X"00000005000000000000001a0000000000000005000000000000000b00000000",
            INIT_04 => X"000000250000000000000047000000000000001b000000000000002800000000",
            INIT_05 => X"00000016000000000000000c000000000000001600000000ffffffdeffffffff",
            INIT_06 => X"ffffffe6ffffffffffffffeeffffffffffffffdffffffffffffffffeffffffff",
            INIT_07 => X"000000120000000000000002000000000000000400000000fffffff5ffffffff",
            INIT_08 => X"00000006000000000000001700000000ffffffffffffffff0000000000000000",
            INIT_09 => X"0000000800000000fffffff2fffffffffffffff5ffffffffffffffdcffffffff",
            INIT_0A => X"ffffffb5ffffffffffffffebffffffff0000001600000000ffffffc2ffffffff",
            INIT_0B => X"00000005000000000000002000000000fffffff6ffffffff0000000800000000",
            INIT_0C => X"00000032000000000000003b00000000ffffffe8ffffffffffffffedffffffff",
            INIT_0D => X"0000003200000000000000140000000000000017000000000000002b00000000",
            INIT_0E => X"ffffffe7fffffffffffffff9ffffffff0000000300000000ffffffc3ffffffff",
            INIT_0F => X"0000001100000000fffffff0ffffffffffffffc0ffffffff0000001600000000",
            INIT_10 => X"0000001100000000ffffffeeffffffff0000000900000000ffffffeaffffffff",
            INIT_11 => X"ffffffd0fffffffffffffffefffffffffffffffdffffffff0000000400000000",
            INIT_12 => X"ffffffd8ffffffff00000010000000000000000d00000000ffffffd8ffffffff",
            INIT_13 => X"ffffffcefffffffffffffff2ffffffff0000000700000000ffffffe5ffffffff",
            INIT_14 => X"0000000e0000000000000015000000000000000e00000000ffffffedffffffff",
            INIT_15 => X"0000000500000000fffffff4ffffffff0000000e000000000000001c00000000",
            INIT_16 => X"ffffffe1ffffffff0000000f00000000fffffffcfffffffffffffff1ffffffff",
            INIT_17 => X"0000001600000000ffffffd0ffffffffffffffe1ffffffff0000001d00000000",
            INIT_18 => X"ffffffe3ffffffffffffffeefffffffffffffff6ffffffffffffffe0ffffffff",
            INIT_19 => X"ffffffcbffffffffffffffb3ffffffffffffffceffffffff0000000800000000",
            INIT_1A => X"ffffffebfffffffffffffffcfffffffffffffffbffffffff0000000e00000000",
            INIT_1B => X"ffffffedffffffff0000001500000000ffffffedffffffff0000001000000000",
            INIT_1C => X"0000000900000000ffffffccfffffffffffffff3ffffffffffffffdfffffffff",
            INIT_1D => X"0000001400000000ffffffe3ffffffff0000001500000000fffffff7ffffffff",
            INIT_1E => X"ffffffe9fffffffffffffff4fffffffffffffff6ffffffff0000001200000000",
            INIT_1F => X"ffffffeffffffffffffffff4ffffffffffffffecffffffffffffffccffffffff",
            INIT_20 => X"ffffffd4ffffffffffffffc5fffffffffffffffefffffffffffffff5ffffffff",
            INIT_21 => X"ffffffceffffffff0000004200000000ffffffd3ffffffffffffffe7ffffffff",
            INIT_22 => X"ffffffcfffffffff00000000000000000000000e00000000ffffffeeffffffff",
            INIT_23 => X"0000000b00000000ffffffd9ffffffffffffffd8ffffffff0000000700000000",
            INIT_24 => X"0000000200000000ffffffffffffffff0000000e00000000fffffffeffffffff",
            INIT_25 => X"0000001600000000000000000000000000000040000000000000002c00000000",
            INIT_26 => X"0000000300000000000000160000000000000000000000000000001000000000",
            INIT_27 => X"0000000300000000000000050000000000000014000000000000001800000000",
            INIT_28 => X"0000000f00000000000000230000000000000027000000000000001000000000",
            INIT_29 => X"0000001100000000ffffffd3fffffffffffffff8ffffffff0000001a00000000",
            INIT_2A => X"ffffffeafffffffffffffffeffffffffffffffc9ffffffff0000001300000000",
            INIT_2B => X"0000002800000000fffffff1fffffffffffffff3ffffffff0000002300000000",
            INIT_2C => X"00000015000000000000001d00000000ffffffebffffffff0000000a00000000",
            INIT_2D => X"ffffffe4ffffffffffffffedffffffffffffffebffffffffffffffedffffffff",
            INIT_2E => X"ffffffe6ffffffffffffffe4ffffffff00000008000000000000000400000000",
            INIT_2F => X"ffffffeeffffffffffffffe3fffffffffffffff6ffffffffffffffdcffffffff",
            INIT_30 => X"00000005000000000000001400000000ffffffe9fffffffffffffff5ffffffff",
            INIT_31 => X"0000002100000000000000390000000000000011000000000000001d00000000",
            INIT_32 => X"0000001a00000000ffffffd6ffffffffffffffa6ffffffff0000000100000000",
            INIT_33 => X"0000001700000000ffffffcfffffffff0000000900000000fffffff8ffffffff",
            INIT_34 => X"fffffff8ffffffff0000001c00000000fffffff5ffffffff0000000500000000",
            INIT_35 => X"0000000700000000ffffffedffffffff0000001d00000000fffffff8ffffffff",
            INIT_36 => X"000000050000000000000016000000000000001100000000ffffffffffffffff",
            INIT_37 => X"0000002500000000000000220000000000000052000000000000002d00000000",
            INIT_38 => X"0000000e00000000000000200000000000000012000000000000001000000000",
            INIT_39 => X"ffffffe3fffffffffffffff2ffffffff00000024000000000000001b00000000",
            INIT_3A => X"ffffffffffffffff0000000700000000ffffffe9ffffffff0000001600000000",
            INIT_3B => X"0000000000000000000000120000000000000027000000000000002c00000000",
            INIT_3C => X"ffffffd5ffffffff00000014000000000000000d00000000fffffffcffffffff",
            INIT_3D => X"0000002c00000000ffffff92ffffffff00000003000000000000003c00000000",
            INIT_3E => X"0000000c00000000ffffffe2ffffffffffffff8effffffff0000000c00000000",
            INIT_3F => X"fffffff5ffffffff00000002000000000000000c000000000000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff5ffffffffffffffd5ffffffffffffffcdffffffff0000001d00000000",
            INIT_41 => X"0000003200000000ffffffefffffffffffffffdeffffffff0000001d00000000",
            INIT_42 => X"fffffffdffffffff0000001e0000000000000007000000000000000200000000",
            INIT_43 => X"fffffff9ffffffff0000004700000000ffffffb0ffffffff0000002000000000",
            INIT_44 => X"ffffff86ffffffff00000010000000000000003f00000000fffffff1ffffffff",
            INIT_45 => X"fffffff3ffffffffffffffccffffffffffffffecffffffff0000004500000000",
            INIT_46 => X"0000000600000000fffffff5ffffffffffffffe1ffffffff0000000700000000",
            INIT_47 => X"0000001400000000ffffffe3ffffffff0000000500000000ffffffdeffffffff",
            INIT_48 => X"ffffffc7ffffffff0000003600000000fffffffeffffffffffffffdfffffffff",
            INIT_49 => X"ffffffeeffffffffffffffe8ffffffff00000006000000000000001700000000",
            INIT_4A => X"fffffff0ffffffff0000001900000000ffffffffffffffffffffffe2ffffffff",
            INIT_4B => X"ffffffceffffffff0000000c000000000000002200000000ffffffc7ffffffff",
            INIT_4C => X"0000001400000000000000190000000000000023000000000000003100000000",
            INIT_4D => X"fffffff9ffffffffffffffd7ffffffff00000042000000000000000d00000000",
            INIT_4E => X"0000000100000000fffffffeffffffffffffffddffffffff0000002500000000",
            INIT_4F => X"fffffffeffffffff000000060000000000000012000000000000000000000000",
            INIT_50 => X"00000024000000000000000100000000ffffffe1ffffffff0000000b00000000",
            INIT_51 => X"ffffffdeffffffff0000000f000000000000000800000000ffffffd4ffffffff",
            INIT_52 => X"ffffffbbffffffffffffff98ffffffffffffffebfffffffffffffff1ffffffff",
            INIT_53 => X"00000007000000000000003600000000ffffffc9ffffffff0000000300000000",
            INIT_54 => X"ffffffccffffffffffffffe1ffffffff0000001000000000ffffff98ffffffff",
            INIT_55 => X"ffffffdaffffffff00000014000000000000002c00000000ffffffebffffffff",
            INIT_56 => X"0000000400000000ffffffe9ffffffff00000016000000000000000d00000000",
            INIT_57 => X"0000000600000000ffffffeeffffffff00000002000000000000002600000000",
            INIT_58 => X"fffffffdffffffff000000070000000000000000000000000000000000000000",
            INIT_59 => X"000000060000000000000001000000000000000300000000ffffffeaffffffff",
            INIT_5A => X"ffffffdeffffffffffffffcdffffffffffffffe6ffffffff0000002900000000",
            INIT_5B => X"ffffffc3ffffffffffffffe6fffffffffffffff2ffffffffffffffe3ffffffff",
            INIT_5C => X"fffffff5fffffffffffffff8fffffffffffffffbffffffff0000000100000000",
            INIT_5D => X"0000001d000000000000001a00000000fffffff7ffffffff0000001800000000",
            INIT_5E => X"ffffffefffffffff0000003200000000ffffffc8fffffffffffffffeffffffff",
            INIT_5F => X"ffffffceffffffff00000001000000000000003800000000ffffffc9ffffffff",
            INIT_60 => X"0000002c000000000000001200000000ffffffeeffffffff0000003d00000000",
            INIT_61 => X"00000013000000000000001800000000ffffffefffffffff0000001e00000000",
            INIT_62 => X"0000001300000000ffffffc4fffffffffffffff7ffffffffffffffa5ffffffff",
            INIT_63 => X"00000003000000000000001100000000ffffffeafffffffffffffff9ffffffff",
            INIT_64 => X"ffffffe1ffffffff0000000c00000000ffffffffffffffff0000002600000000",
            INIT_65 => X"0000000700000000ffffffe9ffffffff00000011000000000000000c00000000",
            INIT_66 => X"0000000f000000000000001300000000fffffffefffffffffffffff5ffffffff",
            INIT_67 => X"0000001300000000fffffff6fffffffffffffff9ffffffff0000001000000000",
            INIT_68 => X"fffffff4ffffffff0000001900000000ffffffd0ffffffffffffffffffffffff",
            INIT_69 => X"ffffffc5ffffffff0000000c000000000000000c00000000ffffffc0ffffffff",
            INIT_6A => X"ffffffbcffffffffffffffbaffffffffffffffe3ffffffff0000000100000000",
            INIT_6B => X"0000002200000000ffffffc6ffffffffffffffe8ffffffff0000000300000000",
            INIT_6C => X"00000003000000000000000000000000fffffffcffffffffffffffdeffffffff",
            INIT_6D => X"ffffffbffffffffffffffff0ffffffffffffffe5ffffffffffffffcfffffffff",
            INIT_6E => X"ffffffffffffffffffffffedffffffff0000000a00000000ffffffe5ffffffff",
            INIT_6F => X"0000000400000000fffffffeffffffffffffffe3ffffffff0000000500000000",
            INIT_70 => X"0000001f000000000000003200000000ffffffdcffffffffffffffe1ffffffff",
            INIT_71 => X"ffffffd9ffffffff00000032000000000000003400000000fffffffcffffffff",
            INIT_72 => X"ffffffb3ffffffff0000000f0000000000000016000000000000000100000000",
            INIT_73 => X"0000000700000000fffffff6ffffffff00000043000000000000001900000000",
            INIT_74 => X"00000020000000000000001500000000fffffff5ffffffff0000002100000000",
            INIT_75 => X"fffffff4fffffffffffffff7ffffffff0000002500000000ffffffceffffffff",
            INIT_76 => X"ffffffccfffffffffffffff6ffffffffffffffc2ffffffff0000001900000000",
            INIT_77 => X"00000006000000000000001200000000ffffffcfffffffff0000002300000000",
            INIT_78 => X"ffffffddffffffff0000000e00000000ffffffe9ffffffffffffffcdffffffff",
            INIT_79 => X"00000030000000000000000600000000fffffff8ffffffff0000001f00000000",
            INIT_7A => X"00000024000000000000002800000000ffffffdbffffffff0000000100000000",
            INIT_7B => X"00000019000000000000002900000000ffffffddffffffffffffffa0ffffffff",
            INIT_7C => X"ffffffeafffffffffffffff6ffffffff0000001100000000ffffffd7ffffffff",
            INIT_7D => X"0000000b00000000fffffffaffffffff00000005000000000000003600000000",
            INIT_7E => X"ffffffcdffffffff0000001900000000ffffffcbffffffffffffffc8ffffffff",
            INIT_7F => X"0000001100000000ffffffe5ffffffffffffffffffffffff0000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE34;


    MEM_IWGHT_LAYER2_INSTANCE35 : if BRAM_NAME = "iwght_layer2_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffaffffffff0000001000000000fffffff3ffffffff0000000d00000000",
            INIT_01 => X"ffffffcefffffffffffffff9ffffffff0000000100000000ffffffd9ffffffff",
            INIT_02 => X"00000007000000000000000d000000000000001400000000ffffffceffffffff",
            INIT_03 => X"0000000d0000000000000039000000000000001e000000000000003600000000",
            INIT_04 => X"000000200000000000000017000000000000002b000000000000004d00000000",
            INIT_05 => X"000000110000000000000027000000000000001e000000000000000900000000",
            INIT_06 => X"ffffffeeffffffff00000041000000000000003f000000000000002f00000000",
            INIT_07 => X"ffffffd9ffffffff0000000400000000ffffffccffffffff0000003700000000",
            INIT_08 => X"0000005100000000fffffff1ffffffffffffffefffffffffffffffeaffffffff",
            INIT_09 => X"ffffffffffffffffffffffe9fffffffffffffff4fffffffffffffff1ffffffff",
            INIT_0A => X"ffffffd5ffffffffffffffc5ffffffffffffffdcffffffffffffffcfffffffff",
            INIT_0B => X"ffffffeaffffffffffffffeefffffffffffffff2ffffffff0000000b00000000",
            INIT_0C => X"ffffffb4ffffffffffffffc3ffffffffffffffbfffffffffffffffd2ffffffff",
            INIT_0D => X"0000000700000000fffffff4ffffffffffffffffffffffffffffffbdffffffff",
            INIT_0E => X"000000230000000000000019000000000000001d000000000000000400000000",
            INIT_0F => X"ffffffdfffffffffffffffe6ffffffff00000021000000000000002100000000",
            INIT_10 => X"0000000100000000fffffffaffffffff0000000700000000fffffffeffffffff",
            INIT_11 => X"fffffff7ffffffffffffffdeffffffffffffffe2ffffffffffffffeeffffffff",
            INIT_12 => X"ffffffecffffffffffffffe8fffffffffffffff8ffffffff0000000900000000",
            INIT_13 => X"ffffffefffffffffffffffecfffffffffffffff1ffffffff0000001f00000000",
            INIT_14 => X"fffffff9ffffffff000000100000000000000010000000000000000100000000",
            INIT_15 => X"0000003500000000fffffffcfffffffffffffff9ffffffff0000000300000000",
            INIT_16 => X"0000000c00000000ffffffe3ffffffff00000000000000000000001900000000",
            INIT_17 => X"0000001000000000ffffffeaffffffffffffffeeffffffff0000000500000000",
            INIT_18 => X"0000001600000000ffffffdfffffffffffffffafffffffff0000000b00000000",
            INIT_19 => X"fffffff5ffffffff0000002f00000000ffffffffffffffff0000001600000000",
            INIT_1A => X"000000170000000000000003000000000000001100000000ffffffeaffffffff",
            INIT_1B => X"0000003e00000000fffffffdffffffff0000001f000000000000001b00000000",
            INIT_1C => X"0000006000000000000000590000000000000037000000000000002300000000",
            INIT_1D => X"ffffffefffffffffffffffefffffffffffffffdbffffffff0000005e00000000",
            INIT_1E => X"ffffffeeffffffffffffffccffffffffffffffc3ffffffffffffffe7ffffffff",
            INIT_1F => X"00000007000000000000000b00000000ffffff9bffffffffffffffa6ffffffff",
            INIT_20 => X"0000001000000000fffffffdfffffffffffffff9fffffffffffffffaffffffff",
            INIT_21 => X"fffffffeffffffffffffffebffffffffffffffebfffffffffffffff4ffffffff",
            INIT_22 => X"00000020000000000000002000000000ffffffdefffffffffffffffbffffffff",
            INIT_23 => X"0000000a00000000000000410000000000000046000000000000003a00000000",
            INIT_24 => X"ffffffebffffffffffffffcfffffffffffffffdefffffffffffffff8ffffffff",
            INIT_25 => X"ffffffe8ffffffffffffffe3ffffffffffffffd4ffffffffffffffe4ffffffff",
            INIT_26 => X"ffffffe8ffffffffffffffebffffffffffffffd6ffffffffffffffe5ffffffff",
            INIT_27 => X"ffffffb5ffffffff000000000000000000000013000000000000002700000000",
            INIT_28 => X"fffffff8ffffffff00000009000000000000000000000000ffffffffffffffff",
            INIT_29 => X"ffffffc4ffffffffffffffdcffffffff00000014000000000000000800000000",
            INIT_2A => X"0000000300000000000000190000000000000018000000000000001000000000",
            INIT_2B => X"000000300000000000000019000000000000000f000000000000002e00000000",
            INIT_2C => X"ffffffeaffffffffffffffe5fffffffffffffff1ffffffffffffffe7ffffffff",
            INIT_2D => X"0000000800000000fffffff2fffffffffffffff7fffffffffffffff2ffffffff",
            INIT_2E => X"0000000600000000ffffffd3fffffffffffffffcffffffff0000000b00000000",
            INIT_2F => X"0000000c0000000000000005000000000000001200000000ffffffc5ffffffff",
            INIT_30 => X"000000060000000000000023000000000000001400000000fffffffdffffffff",
            INIT_31 => X"00000018000000000000000000000000ffffffc4ffffffff0000001800000000",
            INIT_32 => X"0000004d00000000000000240000000000000031000000000000002000000000",
            INIT_33 => X"ffffffe5ffffffff0000001c0000000000000014000000000000000b00000000",
            INIT_34 => X"00000012000000000000001000000000fffffffcffffffff0000001100000000",
            INIT_35 => X"ffffffffffffffff0000000b000000000000003a00000000ffffffd4ffffffff",
            INIT_36 => X"0000001200000000fffffff2ffffffffffffffe7fffffffffffffff0ffffffff",
            INIT_37 => X"0000003e0000000000000027000000000000003d000000000000003800000000",
            INIT_38 => X"0000001a000000000000000c000000000000000000000000ffffffffffffffff",
            INIT_39 => X"ffffffe4fffffffffffffff3ffffffff00000025000000000000001100000000",
            INIT_3A => X"0000003100000000ffffffe0fffffffffffffff6fffffffffffffffcffffffff",
            INIT_3B => X"fffffff7ffffffff0000001100000000ffffffdeffffffff0000000000000000",
            INIT_3C => X"fffffff1fffffffffffffff4ffffffffffffffbbfffffffffffffff4ffffffff",
            INIT_3D => X"ffffffedffffffff0000000c00000000ffffffdfffffffff0000000b00000000",
            INIT_3E => X"ffffffdaffffffffffffffe3ffffffff0000001000000000ffffffdeffffffff",
            INIT_3F => X"0000000000000000ffffffcbffffffffffffffe7fffffffffffffff4ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000e000000000000000e00000000ffffffd2fffffffffffffff1ffffffff",
            INIT_41 => X"00000002000000000000001d0000000000000034000000000000002a00000000",
            INIT_42 => X"0000001300000000000000040000000000000015000000000000000e00000000",
            INIT_43 => X"ffffffe1ffffffff0000000e0000000000000024000000000000000a00000000",
            INIT_44 => X"fffffff6ffffffffffffffeaffffffff0000000700000000ffffffdcffffffff",
            INIT_45 => X"0000000200000000fffffff4ffffffff00000009000000000000000900000000",
            INIT_46 => X"0000000200000000ffffffdfffffffff0000001300000000fffffff5ffffffff",
            INIT_47 => X"fffffff7fffffffffffffff3ffffffffffffffe5ffffffff0000004e00000000",
            INIT_48 => X"ffffffecffffffff0000000e000000000000000800000000ffffffdeffffffff",
            INIT_49 => X"0000000d00000000fffffffdffffffff00000017000000000000001000000000",
            INIT_4A => X"0000001b000000000000000100000000ffffffe1ffffffff0000000b00000000",
            INIT_4B => X"ffffffc6ffffffff0000003a000000000000001400000000ffffffb1ffffffff",
            INIT_4C => X"000000010000000000000031000000000000001f000000000000003300000000",
            INIT_4D => X"0000000400000000000000040000000000000016000000000000001a00000000",
            INIT_4E => X"0000000c00000000ffffffeeffffffffffffffdeffffffff0000000e00000000",
            INIT_4F => X"00000004000000000000001a00000000fffffffdffffffff0000002900000000",
            INIT_50 => X"ffffffdeffffffffffffffe7fffffffffffffff7ffffffff0000001200000000",
            INIT_51 => X"0000001d00000000fffffffaffffffff00000000000000000000002e00000000",
            INIT_52 => X"00000026000000000000002400000000ffffffffffffffffffffffe9ffffffff",
            INIT_53 => X"0000000300000000fffffffdfffffffffffffffdffffffffffffffccffffffff",
            INIT_54 => X"fffffff9ffffffffffffffebffffffffffffffedffffffffffffffe8ffffffff",
            INIT_55 => X"fffffffcffffffffffffffe6ffffffff0000000900000000fffffff9ffffffff",
            INIT_56 => X"fffffffcffffffffffffffcaffffffffffffffd8ffffffff0000001b00000000",
            INIT_57 => X"ffffffa2ffffffff0000000e000000000000000100000000fffffff2ffffffff",
            INIT_58 => X"0000001000000000ffffffbcffffffff0000001c000000000000000300000000",
            INIT_59 => X"00000042000000000000000e00000000ffffffdcffffffff0000002600000000",
            INIT_5A => X"0000001700000000ffffffe2ffffffff00000011000000000000003f00000000",
            INIT_5B => X"00000002000000000000002500000000ffffffd2ffffffffffffffe0ffffffff",
            INIT_5C => X"00000008000000000000000000000000fffffff1ffffffffffffffbaffffffff",
            INIT_5D => X"0000000700000000fffffff8ffffffffffffffefffffffff0000000200000000",
            INIT_5E => X"0000002000000000ffffffe2ffffffff00000013000000000000001300000000",
            INIT_5F => X"0000002100000000fffffff3ffffffff0000001c00000000fffffffaffffffff",
            INIT_60 => X"fffffff8ffffffff00000018000000000000001e00000000fffffff3ffffffff",
            INIT_61 => X"0000001000000000fffffff2ffffffff0000001e000000000000000f00000000",
            INIT_62 => X"000000100000000000000013000000000000000a000000000000001b00000000",
            INIT_63 => X"ffffffefffffffff0000000100000000ffffffe8ffffffff0000001f00000000",
            INIT_64 => X"fffffff4ffffffff0000000000000000ffffffe9ffffffffffffffeeffffffff",
            INIT_65 => X"fffffff9ffffffffffffffeeffffffff0000000d00000000fffffffcffffffff",
            INIT_66 => X"0000001c00000000ffffffc8fffffffffffffffbffffffff0000002c00000000",
            INIT_67 => X"0000000c000000000000000d000000000000000500000000ffffffe6ffffffff",
            INIT_68 => X"ffffffecffffffff0000000700000000fffffff8fffffffffffffff5ffffffff",
            INIT_69 => X"ffffffb9fffffffffffffff8ffffffff0000000c000000000000000900000000",
            INIT_6A => X"0000000300000000ffffffd9ffffffff00000025000000000000000d00000000",
            INIT_6B => X"0000004500000000fffffffaffffffffffffffdfffffffff0000003b00000000",
            INIT_6C => X"0000002800000000ffffffccffffffff0000000e000000000000004600000000",
            INIT_6D => X"ffffffedffffffff0000003000000000ffffffa7ffffffffffffffefffffffff",
            INIT_6E => X"fffffff1ffffffff0000000f000000000000000700000000ffffffc7ffffffff",
            INIT_6F => X"ffffffc9ffffffffffffffebffffffffffffffdfffffffffffffffe9ffffffff",
            INIT_70 => X"fffffff1ffffffffffffffefffffffffffffffcefffffffffffffff9ffffffff",
            INIT_71 => X"00000013000000000000002900000000ffffffa9ffffffff0000001a00000000",
            INIT_72 => X"fffffffbffffffff0000004300000000fffffff6ffffffffffffffc6ffffffff",
            INIT_73 => X"ffffffecffffffffffffffe3ffffffff0000000b000000000000001300000000",
            INIT_74 => X"fffffff2ffffffff0000002100000000ffffffb2ffffffff0000002800000000",
            INIT_75 => X"0000003700000000ffffffe5ffffffff00000000000000000000003200000000",
            INIT_76 => X"fffffff1ffffffff0000003900000000ffffffd0fffffffffffffff5ffffffff",
            INIT_77 => X"0000000b000000000000000d00000000ffffffe7ffffffffffffffc2ffffffff",
            INIT_78 => X"fffffff5ffffffff000000290000000000000002000000000000000500000000",
            INIT_79 => X"ffffffd7fffffffffffffff2ffffffff0000000f00000000fffffff0ffffffff",
            INIT_7A => X"ffffffccffffffffffffff97fffffffffffffffaffffffff0000001500000000",
            INIT_7B => X"ffffffd3ffffffffffffffd7ffffffffffffffe6ffffffff0000001900000000",
            INIT_7C => X"ffffffe6ffffffffffffffdaffffffff0000002800000000fffffffaffffffff",
            INIT_7D => X"00000022000000000000000c00000000ffffffd5ffffffff0000001b00000000",
            INIT_7E => X"0000000400000000000000020000000000000009000000000000000000000000",
            INIT_7F => X"ffffffe5ffffffff0000000900000000ffffffd6ffffffff0000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE35;


    MEM_IWGHT_LAYER2_INSTANCE36 : if BRAM_NAME = "iwght_layer2_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000c00000000ffffffe5ffffffff0000000a00000000ffffffccffffffff",
            INIT_01 => X"ffffffe4ffffffffffffffe2ffffffffffffffedffffffff0000000700000000",
            INIT_02 => X"0000001900000000ffffffbcffffffff0000000e000000000000000700000000",
            INIT_03 => X"0000001900000000fffffffdffffffffffffffd9fffffffffffffff8ffffffff",
            INIT_04 => X"ffffffd1ffffffff0000002d00000000ffffffedffffffffffffffe4ffffffff",
            INIT_05 => X"0000000300000000ffffffd4ffffffff0000001a00000000fffffff7ffffffff",
            INIT_06 => X"fffffff0fffffffffffffff1ffffffffffffffd4ffffffff0000001800000000",
            INIT_07 => X"0000003c00000000ffffffd2fffffffffffffffdffffffff0000003600000000",
            INIT_08 => X"00000006000000000000002300000000ffffffe5ffffffff0000000200000000",
            INIT_09 => X"0000000c0000000000000008000000000000000800000000ffffffaeffffffff",
            INIT_0A => X"ffffffefffffffff0000000700000000fffffff6ffffffff0000000100000000",
            INIT_0B => X"00000020000000000000002f000000000000000c000000000000001800000000",
            INIT_0C => X"ffffffdafffffffffffffff8ffffffff0000002300000000ffffffd1ffffffff",
            INIT_0D => X"ffffffe1fffffffffffffff0ffffffffffffffd5ffffffff0000003600000000",
            INIT_0E => X"fffffff6fffffffffffffff1ffffffff00000026000000000000001300000000",
            INIT_0F => X"fffffff3ffffffffffffffdbffffffff0000001600000000fffffff9ffffffff",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE36;


    MEM_IFMAP_LAYER0_INSTANCE0 : if BRAM_NAME = "ifmap_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE0;


    MEM_IFMAP_LAYER0_INSTANCE1 : if BRAM_NAME = "ifmap_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE1;


    MEM_IFMAP_LAYER0_INSTANCE2 : if BRAM_NAME = "ifmap_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE2;


    MEM_IFMAP_LAYER0_INSTANCE3 : if BRAM_NAME = "ifmap_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE3;


    MEM_IFMAP_LAYER0_INSTANCE4 : if BRAM_NAME = "ifmap_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE4;


    MEM_IFMAP_LAYER0_INSTANCE5 : if BRAM_NAME = "ifmap_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE0 : if BRAM_NAME = "ifmap_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000009000000000000000a0000000000000010000000000000001000000000",
            INIT_01 => X"0000000d000000000000000c0000000000000008000000000000000600000000",
            INIT_02 => X"0000000f0000000000000014000000000000000b000000000000000500000000",
            INIT_03 => X"0000000000000000000000010000000000000002000000000000000700000000",
            INIT_04 => X"0000000a000000000000000b0000000000000009000000000000000300000000",
            INIT_05 => X"0000002900000000000000050000000000000003000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000001f000000000000000f0000000000000000000000000000000500000000",
            INIT_08 => X"0000004c000000000000000c000000000000000a000000000000000800000000",
            INIT_09 => X"0000000000000000000000000000000000000013000000000000002c00000000",
            INIT_0A => X"0000000000000000000000000000000000000012000000000000002100000000",
            INIT_0B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000030000000000000000000000000000000300000000",
            INIT_0D => X"0000002d00000000000000290000000000000001000000000000000800000000",
            INIT_0E => X"000000000000000000000000000000000000001c000000000000002400000000",
            INIT_0F => X"0000000e00000000000000110000000000000000000000000000002700000000",
            INIT_10 => X"000000130000000000000033000000000000000a000000000000000000000000",
            INIT_11 => X"0000000b00000000000000110000000000000000000000000000000d00000000",
            INIT_12 => X"0000006900000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000007f000000000000003a0000000000000027000000000000002b00000000",
            INIT_14 => X"0000000000000000000000140000000000000025000000000000007c00000000",
            INIT_15 => X"0000000e000000000000003c0000000000000053000000000000000000000000",
            INIT_16 => X"0000002a000000000000005e0000000000000000000000000000000300000000",
            INIT_17 => X"0000001a000000000000001e0000000000000013000000000000002e00000000",
            INIT_18 => X"000000000000000000000017000000000000002c000000000000004f00000000",
            INIT_19 => X"0000000000000000000000010000000000000013000000000000005600000000",
            INIT_1A => X"00000007000000000000003b0000000000000058000000000000000200000000",
            INIT_1B => X"00000080000000000000003b000000000000000b000000000000000000000000",
            INIT_1C => X"0000004d000000000000001e000000000000002c000000000000005000000000",
            INIT_1D => X"000000200000000000000025000000000000000f000000000000002300000000",
            INIT_1E => X"0000000e0000000000000041000000000000004f000000000000005f00000000",
            INIT_1F => X"0000000000000000000000320000000000000069000000000000001300000000",
            INIT_20 => X"0000004800000000000000350000000000000012000000000000000100000000",
            INIT_21 => X"0000007100000000000000000000000000000003000000000000001500000000",
            INIT_22 => X"0000002e000000000000000c0000000000000040000000000000005e00000000",
            INIT_23 => X"000000170000000000000000000000000000001b000000000000002400000000",
            INIT_24 => X"0000000000000000000000000000000000000035000000000000004b00000000",
            INIT_25 => X"000000540000000000000035000000000000000f000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_27 => X"00000000000000000000003c0000000000000072000000000000002200000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000004c00000000000000670000000000000056000000000000000100000000",
            INIT_2A => X"00000047000000000000008700000000000000c4000000000000002100000000",
            INIT_2B => X"0000000c00000000000000110000000000000027000000000000004800000000",
            INIT_2C => X"0000001e00000000000000170000000000000014000000000000001500000000",
            INIT_2D => X"0000006d00000000000000510000000000000044000000000000001000000000",
            INIT_2E => X"000000130000000000000016000000000000001500000000000000a300000000",
            INIT_2F => X"0000000700000000000000060000000000000007000000000000000f00000000",
            INIT_30 => X"00000023000000000000000e000000000000002a000000000000001f00000000",
            INIT_31 => X"000000390000000000000090000000000000004d000000000000000a00000000",
            INIT_32 => X"000000160000000000000010000000000000000f000000000000001500000000",
            INIT_33 => X"00000024000000000000002c000000000000001f000000000000001400000000",
            INIT_34 => X"000000180000000000000029000000000000004a000000000000000b00000000",
            INIT_35 => X"0000002600000000000000240000000000000050000000000000001c00000000",
            INIT_36 => X"0000000b000000000000000c000000000000001c000000000000003100000000",
            INIT_37 => X"0000001b0000000000000003000000000000001a000000000000001b00000000",
            INIT_38 => X"00000080000000000000007c000000000000007a000000000000001f00000000",
            INIT_39 => X"00000081000000000000007c0000000000000080000000000000008000000000",
            INIT_3A => X"0000006100000000000000710000000000000087000000000000008b00000000",
            INIT_3B => X"0000007000000000000000710000000000000069000000000000006400000000",
            INIT_3C => X"0000008200000000000000870000000000000083000000000000008100000000",
            INIT_3D => X"000000740000000000000072000000000000007b000000000000008300000000",
            INIT_3E => X"0000002d0000000000000025000000000000003c000000000000004e00000000",
            INIT_3F => X"00000060000000000000006b000000000000005d000000000000004600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008700000000000000850000000000000082000000000000006700000000",
            INIT_41 => X"000000310000000000000035000000000000003e000000000000007100000000",
            INIT_42 => X"0000001700000000000000190000000000000017000000000000002f00000000",
            INIT_43 => X"0000005c00000000000000140000000000000059000000000000003e00000000",
            INIT_44 => X"0000005900000000000000720000000000000088000000000000007200000000",
            INIT_45 => X"0000003b000000000000001b0000000000000025000000000000003500000000",
            INIT_46 => X"0000001f000000000000000e0000000000000023000000000000001400000000",
            INIT_47 => X"00000059000000000000003d0000000000000000000000000000005500000000",
            INIT_48 => X"0000001a000000000000003d0000000000000043000000000000008700000000",
            INIT_49 => X"00000024000000000000003e0000000000000016000000000000001900000000",
            INIT_4A => X"0000004200000000000000140000000000000022000000000000001800000000",
            INIT_4B => X"0000005f000000000000004d0000000000000022000000000000000400000000",
            INIT_4C => X"0000002000000000000000180000000000000028000000000000003600000000",
            INIT_4D => X"0000000c0000000000000014000000000000005c000000000000000d00000000",
            INIT_4E => X"00000009000000000000001b0000000000000016000000000000002600000000",
            INIT_4F => X"0000005500000000000000500000000000000044000000000000000300000000",
            INIT_50 => X"0000000b00000000000000170000000000000020000000000000004300000000",
            INIT_51 => X"0000001e00000000000000110000000000000001000000000000004600000000",
            INIT_52 => X"00000000000000000000000c0000000000000020000000000000001f00000000",
            INIT_53 => X"0000004500000000000000520000000000000035000000000000002c00000000",
            INIT_54 => X"0000004b0000000000000016000000000000001a000000000000000a00000000",
            INIT_55 => X"000000240000000000000024000000000000000d000000000000001100000000",
            INIT_56 => X"0000000000000000000000050000000000000001000000000000003d00000000",
            INIT_57 => X"0000001c00000000000000200000000000000031000000000000002300000000",
            INIT_58 => X"0000003100000000000000270000000000000033000000000000002000000000",
            INIT_59 => X"00000066000000000000003c0000000000000024000000000000000d00000000",
            INIT_5A => X"000000190000000000000000000000000000000d000000000000000d00000000",
            INIT_5B => X"0000000f00000000000000300000000000000033000000000000001000000000",
            INIT_5C => X"00000014000000000000000a0000000000000028000000000000002c00000000",
            INIT_5D => X"0000000f00000000000000680000000000000062000000000000003400000000",
            INIT_5E => X"0000000000000000000000470000000000000000000000000000000f00000000",
            INIT_5F => X"000000000000000000000000000000000000001f000000000000001600000000",
            INIT_60 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"000000000000000000000000000000000000003b000000000000000200000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000110000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE0;


    MEM_IFMAP_LAYER1_INSTANCE1 : if BRAM_NAME = "ifmap_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_03 => X"0000000000000000000000170000000000000016000000000000000000000000",
            INIT_04 => X"0000000f000000000000000b0000000000000025000000000000000000000000",
            INIT_05 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000021000000000000001200000000",
            INIT_08 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_0A => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_0C => X"000000000000000000000000000000000000000b000000000000002300000000",
            INIT_0D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_0E => X"0000003c00000000000000320000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000005000000000000000700000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_12 => X"00000020000000000000002f000000000000002e000000000000000000000000",
            INIT_13 => X"000000000000000000000000000000000000001c000000000000000b00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000170000000000000022000000000000002c000000000000003500000000",
            INIT_17 => X"0000003600000000000000180000000000000016000000000000002c00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_19 => X"00000041000000000000001b000000000000001b000000000000000600000000",
            INIT_1A => X"0000006200000000000000320000000000000028000000000000003600000000",
            INIT_1B => X"0000002000000000000000290000000000000025000000000000003000000000",
            INIT_1C => X"00000025000000000000001e000000000000001b000000000000001800000000",
            INIT_1D => X"0000002900000000000000260000000000000029000000000000002500000000",
            INIT_1E => X"0000001a00000000000000380000000000000057000000000000002000000000",
            INIT_1F => X"0000001600000000000000140000000000000014000000000000001900000000",
            INIT_20 => X"0000002d000000000000002a0000000000000027000000000000002000000000",
            INIT_21 => X"0000002a00000000000000230000000000000035000000000000003200000000",
            INIT_22 => X"0000001a000000000000001a000000000000001b000000000000005800000000",
            INIT_23 => X"0000002600000000000000200000000000000019000000000000001800000000",
            INIT_24 => X"000000390000000000000037000000000000002c000000000000003100000000",
            INIT_25 => X"0000003c000000000000001e000000000000002a000000000000003000000000",
            INIT_26 => X"00000017000000000000001e0000000000000019000000000000001300000000",
            INIT_27 => X"0000002000000000000000260000000000000023000000000000001a00000000",
            INIT_28 => X"00000011000000000000002e0000000000000042000000000000002d00000000",
            INIT_29 => X"0000001000000000000000150000000000000015000000000000001a00000000",
            INIT_2A => X"0000000a000000000000000a000000000000000f000000000000001900000000",
            INIT_2B => X"0000001800000000000000150000000000000011000000000000000b00000000",
            INIT_2C => X"0000000e000000000000000b0000000000000006000000000000000a00000000",
            INIT_2D => X"0000005000000000000000190000000000000013000000000000001100000000",
            INIT_2E => X"0000003800000000000000110000000000000010000000000000000e00000000",
            INIT_2F => X"0000000f0000000000000014000000000000001c000000000000003700000000",
            INIT_30 => X"0000000f00000000000000160000000000000011000000000000000b00000000",
            INIT_31 => X"000000350000000000000041000000000000000d000000000000001000000000",
            INIT_32 => X"00000070000000000000006b000000000000001c000000000000001900000000",
            INIT_33 => X"0000001d00000000000000050000000000000030000000000000006600000000",
            INIT_34 => X"00000011000000000000000c000000000000001d000000000000002b00000000",
            INIT_35 => X"0000003d000000000000004d0000000000000033000000000000001b00000000",
            INIT_36 => X"000000460000000000000079000000000000005e000000000000004100000000",
            INIT_37 => X"000000840000000000000012000000000000000f000000000000004800000000",
            INIT_38 => X"0000009e000000000000003d0000000000000022000000000000006a00000000",
            INIT_39 => X"000000380000000000000053000000000000007e000000000000007600000000",
            INIT_3A => X"0000004600000000000000460000000000000079000000000000005400000000",
            INIT_3B => X"000000b000000000000000980000000000000000000000000000002a00000000",
            INIT_3C => X"000000a100000000000000c1000000000000002c000000000000003d00000000",
            INIT_3D => X"000000780000000000000038000000000000005b00000000000000a100000000",
            INIT_3E => X"00000049000000000000004c000000000000005d000000000000009b00000000",
            INIT_3F => X"0000003600000000000000a300000000000000a3000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac00000000000000970000000000000059000000000000001c00000000",
            INIT_41 => X"00000095000000000000008f0000000000000051000000000000008700000000",
            INIT_42 => X"0000004000000000000000580000000000000047000000000000005300000000",
            INIT_43 => X"00000036000000000000004400000000000000c900000000000000b800000000",
            INIT_44 => X"0000007800000000000000af00000000000000af000000000000003b00000000",
            INIT_45 => X"000000550000000000000094000000000000007f000000000000005b00000000",
            INIT_46 => X"000000dc00000000000000430000000000000058000000000000004d00000000",
            INIT_47 => X"0000004b0000000000000080000000000000008200000000000000d700000000",
            INIT_48 => X"00000055000000000000005a0000000000000061000000000000006e00000000",
            INIT_49 => X"00000036000000000000004a000000000000004d000000000000004000000000",
            INIT_4A => X"000000d800000000000000e80000000000000021000000000000004300000000",
            INIT_4B => X"0000004e0000000000000067000000000000008f000000000000009f00000000",
            INIT_4C => X"0000005a000000000000004f0000000000000090000000000000007d00000000",
            INIT_4D => X"000000290000000000000026000000000000001a000000000000004000000000",
            INIT_4E => X"0000009f00000000000000c900000000000000d0000000000000001e00000000",
            INIT_4F => X"000000a5000000000000006e00000000000000e100000000000000d400000000",
            INIT_50 => X"000000380000000000000043000000000000007d00000000000000c800000000",
            INIT_51 => X"00000053000000000000005f000000000000005a000000000000004c00000000",
            INIT_52 => X"000000f700000000000000ba00000000000000e200000000000000a600000000",
            INIT_53 => X"00000084000000000000008500000000000000a200000000000000e500000000",
            INIT_54 => X"00000089000000000000007d0000000000000072000000000000007a00000000",
            INIT_55 => X"000000940000000000000099000000000000009a000000000000009900000000",
            INIT_56 => X"000000bb00000000000000f900000000000000d7000000000000009700000000",
            INIT_57 => X"0000007b000000000000007c000000000000007f000000000000008900000000",
            INIT_58 => X"0000009d000000000000009a0000000000000090000000000000008000000000",
            INIT_59 => X"0000008a00000000000000a800000000000000ba00000000000000a400000000",
            INIT_5A => X"0000008e000000000000009100000000000000fa00000000000000a600000000",
            INIT_5B => X"000000910000000000000085000000000000007b000000000000008800000000",
            INIT_5C => X"000000b200000000000000a200000000000000a2000000000000009b00000000",
            INIT_5D => X"00000089000000000000009f00000000000000ac00000000000000af00000000",
            INIT_5E => X"0000008d000000000000007f0000000000000073000000000000009300000000",
            INIT_5F => X"00000092000000000000009f0000000000000091000000000000008e00000000",
            INIT_60 => X"0000009600000000000000c800000000000000ba000000000000009700000000",
            INIT_61 => X"0000006f000000000000006c000000000000006d000000000000007100000000",
            INIT_62 => X"0000007c00000000000000710000000000000062000000000000007100000000",
            INIT_63 => X"000000620000000000000068000000000000006e000000000000007700000000",
            INIT_64 => X"0000006d000000000000006a0000000000000062000000000000005f00000000",
            INIT_65 => X"0000006c0000000000000073000000000000006c000000000000006800000000",
            INIT_66 => X"0000007500000000000000670000000000000061000000000000003c00000000",
            INIT_67 => X"00000046000000000000002a000000000000001d000000000000003a00000000",
            INIT_68 => X"00000076000000000000006d0000000000000062000000000000005c00000000",
            INIT_69 => X"0000008f00000000000000770000000000000076000000000000007200000000",
            INIT_6A => X"0000000d00000000000000260000000000000058000000000000007f00000000",
            INIT_6B => X"0000003a000000000000002c0000000000000028000000000000002900000000",
            INIT_6C => X"0000006800000000000000030000000000000038000000000000005100000000",
            INIT_6D => X"00000026000000000000004c0000000000000067000000000000006e00000000",
            INIT_6E => X"0000004f0000000000000022000000000000002c000000000000002800000000",
            INIT_6F => X"00000037000000000000002f0000000000000048000000000000003d00000000",
            INIT_70 => X"0000003900000000000000650000000000000000000000000000003000000000",
            INIT_71 => X"00000036000000000000003d0000000000000003000000000000000000000000",
            INIT_72 => X"0000002f0000000000000023000000000000000c000000000000003e00000000",
            INIT_73 => X"0000004300000000000000260000000000000028000000000000002400000000",
            INIT_74 => X"000000650000000000000076000000000000006a000000000000002a00000000",
            INIT_75 => X"0000002f0000000000000030000000000000003e000000000000005800000000",
            INIT_76 => X"0000002800000000000000570000000000000051000000000000000000000000",
            INIT_77 => X"0000003a00000000000000310000000000000012000000000000002b00000000",
            INIT_78 => X"000000250000000000000037000000000000007b000000000000006200000000",
            INIT_79 => X"00000000000000000000003e0000000000000040000000000000004900000000",
            INIT_7A => X"0000001b00000000000000270000000000000036000000000000005c00000000",
            INIT_7B => X"0000001c000000000000002f000000000000002b000000000000002900000000",
            INIT_7C => X"0000007800000000000000190000000000000025000000000000004900000000",
            INIT_7D => X"0000005d0000000000000024000000000000004d000000000000005c00000000",
            INIT_7E => X"0000005200000000000000380000000000000023000000000000004700000000",
            INIT_7F => X"0000002000000000000000460000000000000022000000000000003400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE1;


    MEM_IFMAP_LAYER1_INSTANCE2 : if BRAM_NAME = "ifmap_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003000000000000000510000000000000066000000000000003b00000000",
            INIT_01 => X"00000070000000000000004c0000000000000055000000000000001a00000000",
            INIT_02 => X"0000005200000000000000400000000000000035000000000000003800000000",
            INIT_03 => X"0000002d0000000000000004000000000000004c000000000000003100000000",
            INIT_04 => X"0000002400000000000000130000000000000024000000000000003300000000",
            INIT_05 => X"00000002000000000000002b0000000000000065000000000000006000000000",
            INIT_06 => X"000000300000000000000025000000000000006d000000000000003600000000",
            INIT_07 => X"0000000000000000000000030000000000000000000000000000005800000000",
            INIT_08 => X"0000002b000000000000003f000000000000004b000000000000000000000000",
            INIT_09 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000280000000000000037000000000000001e000000000000002800000000",
            INIT_0B => X"000000380000000000000074000000000000009d000000000000000000000000",
            INIT_0C => X"00000002000000000000000c000000000000001f000000000000003700000000",
            INIT_0D => X"0000000400000000000000000000000000000000000000000000000200000000",
            INIT_0E => X"0000004e00000000000000180000000000000016000000000000000000000000",
            INIT_0F => X"0000000700000000000000040000000000000004000000000000008800000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_11 => X"0000000400000000000000000000000000000005000000000000000000000000",
            INIT_12 => X"00000032000000000000008b0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_14 => X"0000000700000000000000090000000000000002000000000000000000000000",
            INIT_15 => X"000000000000000000000005000000000000001c000000000000000000000000",
            INIT_16 => X"0000001400000000000000230000000000000043000000000000000500000000",
            INIT_17 => X"0000000000000000000000000000000000000009000000000000001900000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000001300000000000000030000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_20 => X"000000120000000000000000000000000000000d000000000000000500000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_22 => X"00000000000000000000000a0000000000000005000000000000003e00000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000009000000000000000a00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000001c0000000000000000000000000000000d000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000016000000000000000c00000000",
            INIT_36 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000300000000000000000000000000000000000000000",
            INIT_39 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000007000000000000002600000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000f000000000000002a0000000000000031000000000000000000000000",
            INIT_3E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000007000000000000002e0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001d00000000000000480000000000000004000000000000000700000000",
            INIT_43 => X"00000031000000000000002e0000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000070000000000000019000000000000001c00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000004f00000000000000140000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_4E => X"0000000300000000000000490000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000014000000000000000c00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_52 => X"0000000200000000000000000000000000000000000000000000000600000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000030000000000000009000000000000000000000000",
            INIT_55 => X"0000000600000000000000010000000000000001000000000000000000000000",
            INIT_56 => X"00000000000000000000001d000000000000000d000000000000000000000000",
            INIT_57 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000120000000000000004000000000000000000000000",
            INIT_59 => X"0000000000000000000000030000000000000039000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000007000000000000000900000000",
            INIT_5B => X"0000000000000000000000000000000000000051000000000000000b00000000",
            INIT_5C => X"00000000000000000000001f000000000000000a000000000000000000000000",
            INIT_5D => X"00000000000000000000000c0000000000000000000000000000006500000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000006800000000",
            INIT_60 => X"0000001d00000000000000000000000000000055000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000066000000000000000000000000",
            INIT_62 => X"0000009400000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000080000000000000000000000000000001e00000000",
            INIT_65 => X"0000000000000000000000000000000000000068000000000000001e00000000",
            INIT_66 => X"0000000000000000000001010000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000056000000000000006100000000",
            INIT_6A => X"00000000000000000000000000000000000000cb000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000015000000000000000400000000",
            INIT_6C => X"0000004300000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000005f00000000",
            INIT_6E => X"0000002100000000000000000000000000000000000000000000008000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000090000000000000000000000000000002f000000000000000000000000",
            INIT_71 => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_72 => X"00000020000000000000001f0000000000000000000000000000000e00000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_74 => X"0000003900000000000000080000000000000000000000000000005500000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000002e000000000000002d000000000000000000000000",
            INIT_77 => X"000000dc00000000000000000000000000000000000000000000005e00000000",
            INIT_78 => X"00000000000000000000004b0000000000000000000000000000000000000000",
            INIT_79 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000004e0000000000000000000000000000000a000000000000000d00000000",
            INIT_7B => X"0000000000000000000000960000000000000000000000000000004100000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000500000000000000060000000000000002000000000000000000000000",
            INIT_7E => X"0000005200000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000008500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE2;


    MEM_IFMAP_LAYER1_INSTANCE3 : if BRAM_NAME = "ifmap_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000400000000000000000000000000000005000000000000000800000000",
            INIT_02 => X"000000ac00000000000000000000000000000000000000000000000e00000000",
            INIT_03 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000040000000000000006000000000000000000000000",
            INIT_05 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_06 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000080000000000000016000000000000000000000000",
            INIT_08 => X"0000000400000000000000000000000000000000000000000000000c00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000008000000000000001c00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000001b0000000000000022000000000000000b000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000018000000000000002800000000",
            INIT_15 => X"0000000000000000000000000000000000000007000000000000001b00000000",
            INIT_16 => X"0000001500000000000000050000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000060000000000000000000000000000001700000000",
            INIT_18 => X"000000340000000000000000000000000000000d000000000000000d00000000",
            INIT_19 => X"0000002700000000000000000000000000000000000000000000002900000000",
            INIT_1A => X"0000000f00000000000000160000000000000005000000000000001500000000",
            INIT_1B => X"0000002000000000000000150000000000000017000000000000001100000000",
            INIT_1C => X"00000010000000000000001a0000000000000000000000000000002600000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000024000000000000002a0000000000000016000000000000000a00000000",
            INIT_1F => X"0000002600000000000000140000000000000007000000000000000100000000",
            INIT_20 => X"00000000000000000000000e000000000000002b000000000000002e00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000300000000000000150000000000000018000000000000000f00000000",
            INIT_23 => X"000000170000000000000021000000000000001c000000000000001c00000000",
            INIT_24 => X"0000000000000000000000170000000000000032000000000000002100000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000f00000000000000000000000000000000000000000000000100000000",
            INIT_27 => X"0000002a00000000000000000000000000000000000000000000001500000000",
            INIT_28 => X"00000000000000000000000e0000000000000022000000000000002a00000000",
            INIT_29 => X"0000001600000000000000120000000000000000000000000000000000000000",
            INIT_2A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000001900000000000000090000000000000000000000000000000000000000",
            INIT_2C => X"0000000e0000000000000010000000000000002f000000000000002800000000",
            INIT_2D => X"000000000000000000000011000000000000002e000000000000001900000000",
            INIT_2E => X"00000000000000000000001c000000000000001e000000000000000000000000",
            INIT_2F => X"0000001c0000000000000016000000000000001c000000000000000000000000",
            INIT_30 => X"0000002f00000000000000590000000000000066000000000000004e00000000",
            INIT_31 => X"000000620000000000000041000000000000002c000000000000001700000000",
            INIT_32 => X"0000003b00000000000000420000000000000068000000000000007200000000",
            INIT_33 => X"0000001f000000000000002d0000000000000027000000000000003e00000000",
            INIT_34 => X"00000041000000000000003b0000000000000020000000000000000000000000",
            INIT_35 => X"0000007c0000000000000079000000000000006c000000000000005b00000000",
            INIT_36 => X"0000009500000000000000830000000000000081000000000000008700000000",
            INIT_37 => X"000000320000000000000000000000000000002f000000000000004000000000",
            INIT_38 => X"0000007500000000000000710000000000000073000000000000007600000000",
            INIT_39 => X"000000840000000000000096000000000000008f000000000000008100000000",
            INIT_3A => X"0000008c000000000000009d00000000000000a7000000000000008500000000",
            INIT_3B => X"0000007c0000000000000058000000000000001b000000000000003900000000",
            INIT_3C => X"0000008600000000000000790000000000000076000000000000007e00000000",
            INIT_3D => X"000000a7000000000000008e0000000000000083000000000000008800000000",
            INIT_3E => X"0000006e0000000000000095000000000000009a000000000000007400000000",
            INIT_3F => X"0000006700000000000000650000000000000060000000000000004800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000085000000000000008e0000000000000082000000000000007800000000",
            INIT_41 => X"0000009700000000000000a600000000000000a2000000000000008900000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000005000000000000003f000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE3;


    MEM_IFMAP_LAYER1_INSTANCE4 : if BRAM_NAME = "ifmap_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000130000000000000036000000000000001d000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000001a00000000000000220000000000000022000000000000004800000000",
            INIT_05 => X"0000004300000000000000140000000000000001000000000000000000000000",
            INIT_06 => X"0000001e00000000000000000000000000000002000000000000000100000000",
            INIT_07 => X"00000021000000000000001c0000000000000021000000000000003700000000",
            INIT_08 => X"0000000400000000000000030000000000000007000000000000000b00000000",
            INIT_09 => X"000000030000000000000068000000000000003e000000000000000800000000",
            INIT_0A => X"000000100000000000000057000000000000007d000000000000003d00000000",
            INIT_0B => X"0000003b00000000000000470000000000000000000000000000000e00000000",
            INIT_0C => X"0000000000000000000000190000000000000022000000000000001f00000000",
            INIT_0D => X"000000000000000000000000000000000000002d000000000000001c00000000",
            INIT_0E => X"00000023000000000000002e0000000000000007000000000000000000000000",
            INIT_0F => X"00000000000000000000000d000000000000007f000000000000001300000000",
            INIT_10 => X"000000330000000000000029000000000000001e000000000000001900000000",
            INIT_11 => X"0000001300000000000000000000000000000000000000000000001c00000000",
            INIT_12 => X"000000090000000000000025000000000000001b000000000000004c00000000",
            INIT_13 => X"0000002100000000000000170000000000000009000000000000006000000000",
            INIT_14 => X"00000034000000000000003d000000000000001d000000000000003800000000",
            INIT_15 => X"0000003c000000000000003e000000000000001b000000000000003000000000",
            INIT_16 => X"0000002c00000000000000010000000000000000000000000000000000000000",
            INIT_17 => X"00000009000000000000001d0000000000000003000000000000000f00000000",
            INIT_18 => X"000000120000000000000041000000000000003c000000000000000000000000",
            INIT_19 => X"0000000700000000000000000000000000000021000000000000003600000000",
            INIT_1A => X"00000000000000000000000d0000000000000032000000000000002700000000",
            INIT_1B => X"0000001d00000000000000180000000000000000000000000000000000000000",
            INIT_1C => X"0000005300000000000000140000000000000038000000000000002400000000",
            INIT_1D => X"000000560000000000000038000000000000000b000000000000001500000000",
            INIT_1E => X"0000000900000000000000000000000000000000000000000000001500000000",
            INIT_1F => X"0000004400000000000000000000000000000024000000000000003400000000",
            INIT_20 => X"00000097000000000000009b0000000000000007000000000000003900000000",
            INIT_21 => X"0000000700000000000000040000000000000051000000000000007700000000",
            INIT_22 => X"0000004800000000000000600000000000000045000000000000001d00000000",
            INIT_23 => X"00000028000000000000000e000000000000002c000000000000003000000000",
            INIT_24 => X"000000000000000000000000000000000000008e000000000000004300000000",
            INIT_25 => X"00000034000000000000001e0000000000000004000000000000000100000000",
            INIT_26 => X"00000047000000000000004a000000000000003d000000000000003c00000000",
            INIT_27 => X"0000005100000000000000180000000000000046000000000000004000000000",
            INIT_28 => X"00000035000000000000003a0000000000000000000000000000002400000000",
            INIT_29 => X"0000005100000000000000460000000000000039000000000000003400000000",
            INIT_2A => X"0000006500000000000000420000000000000041000000000000005600000000",
            INIT_2B => X"0000000000000000000000330000000000000044000000000000004100000000",
            INIT_2C => X"0000003900000000000000420000000000000040000000000000002400000000",
            INIT_2D => X"0000003700000000000000400000000000000043000000000000003b00000000",
            INIT_2E => X"0000003d000000000000001d0000000000000062000000000000004000000000",
            INIT_2F => X"0000001e0000000000000000000000000000003a000000000000004400000000",
            INIT_30 => X"0000005100000000000000370000000000000023000000000000002300000000",
            INIT_31 => X"0000007d00000000000000450000000000000041000000000000005400000000",
            INIT_32 => X"0000007b000000000000007d0000000000000037000000000000006000000000",
            INIT_33 => X"0000007900000000000000830000000000000083000000000000008000000000",
            INIT_34 => X"0000006c00000000000000850000000000000091000000000000008900000000",
            INIT_35 => X"000000710000000000000064000000000000005a000000000000005700000000",
            INIT_36 => X"0000008700000000000000880000000000000082000000000000006c00000000",
            INIT_37 => X"0000008b00000000000000750000000000000082000000000000008800000000",
            INIT_38 => X"0000001f0000000000000023000000000000004d000000000000007200000000",
            INIT_39 => X"0000006900000000000000510000000000000036000000000000002900000000",
            INIT_3A => X"0000008a00000000000000860000000000000056000000000000005600000000",
            INIT_3B => X"0000002f00000000000000490000000000000076000000000000008b00000000",
            INIT_3C => X"00000010000000000000001d0000000000000012000000000000001400000000",
            INIT_3D => X"00000030000000000000004c0000000000000029000000000000001800000000",
            INIT_3E => X"0000007700000000000000860000000000000085000000000000003300000000",
            INIT_3F => X"0000000d0000000000000019000000000000003c000000000000004a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000009000000000000001f000000000000002c000000000000001800000000",
            INIT_41 => X"0000003a000000000000001e0000000000000032000000000000000900000000",
            INIT_42 => X"0000005800000000000000570000000000000060000000000000008200000000",
            INIT_43 => X"00000008000000000000000c000000000000001c000000000000003d00000000",
            INIT_44 => X"0000000900000000000000110000000000000029000000000000003700000000",
            INIT_45 => X"0000007e00000000000000290000000000000022000000000000002100000000",
            INIT_46 => X"0000003c0000000000000038000000000000001c000000000000006300000000",
            INIT_47 => X"000000410000000000000007000000000000001a000000000000002f00000000",
            INIT_48 => X"0000000b000000000000000c0000000000000010000000000000001c00000000",
            INIT_49 => X"000000690000000000000055000000000000002c000000000000002200000000",
            INIT_4A => X"0000003000000000000000410000000000000033000000000000002f00000000",
            INIT_4B => X"0000001b00000000000000320000000000000015000000000000002000000000",
            INIT_4C => X"000000290000000000000021000000000000000c000000000000000e00000000",
            INIT_4D => X"0000003600000000000000560000000000000037000000000000002400000000",
            INIT_4E => X"0000001d00000000000000210000000000000039000000000000003300000000",
            INIT_4F => X"00000006000000000000001e0000000000000028000000000000002e00000000",
            INIT_50 => X"000000210000000000000026000000000000003b000000000000002100000000",
            INIT_51 => X"0000002600000000000000430000000000000013000000000000002000000000",
            INIT_52 => X"00000053000000000000001a0000000000000020000000000000002b00000000",
            INIT_53 => X"0000002600000000000000080000000000000011000000000000002100000000",
            INIT_54 => X"0000001e00000000000000250000000000000024000000000000006100000000",
            INIT_55 => X"0000001c000000000000001f0000000000000028000000000000000b00000000",
            INIT_56 => X"0000000a00000000000000190000000000000031000000000000002e00000000",
            INIT_57 => X"00000072000000000000005b0000000000000009000000000000000000000000",
            INIT_58 => X"0000000c0000000000000025000000000000002e000000000000000900000000",
            INIT_59 => X"0000000e000000000000000b0000000000000025000000000000003000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000038000000000000003f000000000000001f000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000044000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"00000000000000000000000b0000000000000011000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_71 => X"0000000a000000000000001b0000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000002f0000000000000014000000000000000000000000",
            INIT_73 => X"0000000200000000000000560000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_75 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000001400000000000000000000000000000035000000000000000000000000",
            INIT_79 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_7E => X"0000000d000000000000006b000000000000001a000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE4;


    MEM_IFMAP_LAYER1_INSTANCE5 : if BRAM_NAME = "ifmap_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_01 => X"0000002100000000000000060000000000000000000000000000000000000000",
            INIT_02 => X"000000030000000000000000000000000000003a000000000000000000000000",
            INIT_03 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000280000000000000012000000000000000f000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000021000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000017000000000000000800000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000003000000000000005c00000000",
            INIT_0B => X"0000002300000000000000240000000000000031000000000000001300000000",
            INIT_0C => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_0E => X"0000002100000000000000060000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000006000000000000001f00000000",
            INIT_10 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_13 => X"0000000300000000000000150000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000025000000000000008800000000",
            INIT_15 => X"00000041000000000000004d000000000000004a000000000000005800000000",
            INIT_16 => X"0000000600000000000000000000000000000001000000000000000e00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000001f000000000000001c0000000000000008000000000000006c00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000700000000000000000000000000000000000000000000000700000000",
            INIT_1C => X"000000000000000000000000000000000000002e000000000000007000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000030000000000000016000000000000000800000000",
            INIT_1F => X"0000001f00000000000000010000000000000000000000000000003f00000000",
            INIT_20 => X"0000001d0000000000000024000000000000001c000000000000005a00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000300000000000000000000000000000000000000000000000300000000",
            INIT_24 => X"0000000200000000000000050000000000000000000000000000000500000000",
            INIT_25 => X"000000000000000000000009000000000000000b000000000000000500000000",
            INIT_26 => X"00000000000000000000000b000000000000000a000000000000000000000000",
            INIT_27 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_28 => X"000000190000000000000014000000000000002e000000000000000000000000",
            INIT_29 => X"000000000000000000000015000000000000000a000000000000000000000000",
            INIT_2A => X"00000000000000000000002e0000000000000006000000000000000000000000",
            INIT_2B => X"0000000000000000000000010000000000000003000000000000000300000000",
            INIT_2C => X"0000000000000000000000000000000000000005000000000000003400000000",
            INIT_2D => X"0000000000000000000000300000000000000000000000000000001c00000000",
            INIT_2E => X"0000000b0000000000000000000000000000005c000000000000000000000000",
            INIT_2F => X"000000090000000000000000000000000000001f000000000000000000000000",
            INIT_30 => X"000000390000000000000000000000000000000e000000000000002400000000",
            INIT_31 => X"00000000000000000000002c0000000000000021000000000000001200000000",
            INIT_32 => X"0000000000000000000000410000000000000000000000000000003e00000000",
            INIT_33 => X"0000003a00000000000000380000000000000026000000000000000000000000",
            INIT_34 => X"0000004d00000000000000000000000000000000000000000000002400000000",
            INIT_35 => X"0000005b00000000000000000000000000000027000000000000000000000000",
            INIT_36 => X"0000000000000000000000500000000000000050000000000000000000000000",
            INIT_37 => X"00000046000000000000001b000000000000002a000000000000001200000000",
            INIT_38 => X"00000000000000000000004a000000000000005c000000000000000000000000",
            INIT_39 => X"0000002d000000000000004d000000000000001e000000000000001100000000",
            INIT_3A => X"0000000000000000000000000000000000000042000000000000000700000000",
            INIT_3B => X"00000000000000000000003b0000000000000030000000000000000100000000",
            INIT_3C => X"0000000000000000000000000000000000000038000000000000005100000000",
            INIT_3D => X"000000300000000000000000000000000000004d000000000000002600000000",
            INIT_3E => X"0000006700000000000000000000000000000000000000000000001100000000",
            INIT_3F => X"0000002c0000000000000000000000000000001e000000000000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000400000000000000030000000000000000000000000000003c00000000",
            INIT_41 => X"0000000000000000000000980000000000000000000000000000004100000000",
            INIT_42 => X"0000000f000000000000000b0000000000000000000000000000005100000000",
            INIT_43 => X"000000440000000000000000000000000000002b000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000003800000000000000000000000000000075000000000000000000000000",
            INIT_46 => X"0000003700000000000000030000000000000000000000000000002200000000",
            INIT_47 => X"0000000000000000000000000000000000000038000000000000001600000000",
            INIT_48 => X"0000000200000000000000000000000000000011000000000000000000000000",
            INIT_49 => X"00000033000000000000005f0000000000000000000000000000006100000000",
            INIT_4A => X"00000024000000000000004c000000000000000f000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000300000000000000000000000000000000000000000000000c00000000",
            INIT_4D => X"00000000000000000000003f00000000000000a3000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_4F => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000003000000000000000000000000000000000000000000000001f00000000",
            INIT_51 => X"0000000000000000000000050000000000000000000000000000007500000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000001f000000000000003e0000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000002000000000000000d000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000002b0000000000000028000000000000000000000000",
            INIT_58 => X"0000000000000000000000110000000000000000000000000000000c00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001200000000000000000000000000000000000000000000000f00000000",
            INIT_5B => X"0000006f00000000000000700000000000000065000000000000003100000000",
            INIT_5C => X"00000074000000000000006b000000000000006b000000000000006f00000000",
            INIT_5D => X"000000460000000000000051000000000000006b000000000000007900000000",
            INIT_5E => X"0000005f0000000000000064000000000000005d000000000000004f00000000",
            INIT_5F => X"0000007100000000000000730000000000000077000000000000006e00000000",
            INIT_60 => X"0000005e000000000000006a000000000000007b000000000000006c00000000",
            INIT_61 => X"000000280000000000000024000000000000002a000000000000003a00000000",
            INIT_62 => X"00000044000000000000005a0000000000000047000000000000003200000000",
            INIT_63 => X"0000006e0000000000000075000000000000006f000000000000004600000000",
            INIT_64 => X"0000001e00000000000000250000000000000041000000000000005400000000",
            INIT_65 => X"0000002000000000000000250000000000000025000000000000002600000000",
            INIT_66 => X"00000038000000000000002d0000000000000050000000000000002000000000",
            INIT_67 => X"0000003e0000000000000063000000000000006e000000000000006800000000",
            INIT_68 => X"0000001900000000000000190000000000000020000000000000003e00000000",
            INIT_69 => X"00000018000000000000001c0000000000000022000000000000003800000000",
            INIT_6A => X"00000064000000000000003e0000000000000023000000000000003700000000",
            INIT_6B => X"00000041000000000000004f0000000000000066000000000000004a00000000",
            INIT_6C => X"0000003a000000000000001d000000000000001b000000000000002e00000000",
            INIT_6D => X"0000001f000000000000001f0000000000000023000000000000002e00000000",
            INIT_6E => X"00000048000000000000006a0000000000000033000000000000000f00000000",
            INIT_6F => X"0000003600000000000000530000000000000041000000000000003300000000",
            INIT_70 => X"0000002300000000000000360000000000000021000000000000002b00000000",
            INIT_71 => X"0000001c0000000000000022000000000000001c000000000000001c00000000",
            INIT_72 => X"0000003500000000000000610000000000000046000000000000003000000000",
            INIT_73 => X"0000002b00000000000000350000000000000039000000000000004000000000",
            INIT_74 => X"0000001a0000000000000024000000000000002d000000000000002000000000",
            INIT_75 => X"000000350000000000000027000000000000002b000000000000001c00000000",
            INIT_76 => X"000000310000000000000026000000000000004a000000000000002600000000",
            INIT_77 => X"00000034000000000000002c0000000000000026000000000000003100000000",
            INIT_78 => X"0000002700000000000000150000000000000024000000000000003100000000",
            INIT_79 => X"0000001c00000000000000270000000000000028000000000000004800000000",
            INIT_7A => X"000000300000000000000021000000000000002f000000000000002b00000000",
            INIT_7B => X"0000001c000000000000003a0000000000000023000000000000002900000000",
            INIT_7C => X"0000005e000000000000003e0000000000000019000000000000001c00000000",
            INIT_7D => X"0000001a00000000000000280000000000000025000000000000002a00000000",
            INIT_7E => X"0000003a000000000000002a0000000000000023000000000000002600000000",
            INIT_7F => X"000000080000000000000014000000000000001f000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE6 : if BRAM_NAME = "ifmap_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001500000000000000570000000000000053000000000000002200000000",
            INIT_01 => X"0000004800000000000000280000000000000026000000000000002800000000",
            INIT_02 => X"0000000f0000000000000014000000000000000f000000000000002000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_04 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000000c0000000000000037000000000000002400000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_19 => X"0000000100000000000000090000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_1C => X"0000000000000000000000030000000000000018000000000000000000000000",
            INIT_1D => X"0000002200000000000000250000000000000031000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_20 => X"00000014000000000000000a000000000000000b000000000000000600000000",
            INIT_21 => X"00000015000000000000001a0000000000000023000000000000003b00000000",
            INIT_22 => X"000000230000000000000021000000000000000c000000000000000000000000",
            INIT_23 => X"0000001800000000000000220000000000000015000000000000000000000000",
            INIT_24 => X"00000032000000000000000e000000000000000e000000000000002000000000",
            INIT_25 => X"0000000000000000000000140000000000000006000000000000002500000000",
            INIT_26 => X"00000000000000000000004b0000000000000037000000000000000000000000",
            INIT_27 => X"0000002f0000000000000044000000000000006b000000000000000500000000",
            INIT_28 => X"00000032000000000000004b0000000000000000000000000000001500000000",
            INIT_29 => X"000000000000000000000013000000000000001f000000000000001800000000",
            INIT_2A => X"00000000000000000000000e000000000000003d000000000000003800000000",
            INIT_2B => X"000000290000000000000047000000000000003f000000000000003100000000",
            INIT_2C => X"000000110000000000000031000000000000005a000000000000000e00000000",
            INIT_2D => X"00000042000000000000000b0000000000000023000000000000001900000000",
            INIT_2E => X"0000001b0000000000000000000000000000000a000000000000004d00000000",
            INIT_2F => X"0000001a0000000000000038000000000000003e000000000000005800000000",
            INIT_30 => X"0000002300000000000000140000000000000039000000000000004700000000",
            INIT_31 => X"0000006300000000000000530000000000000010000000000000002400000000",
            INIT_32 => X"0000003c000000000000000d0000000000000039000000000000001e00000000",
            INIT_33 => X"0000001000000000000000220000000000000019000000000000002100000000",
            INIT_34 => X"0000001600000000000000180000000000000015000000000000002200000000",
            INIT_35 => X"0000002d00000000000000650000000000000069000000000000000000000000",
            INIT_36 => X"000000360000000000000017000000000000001c000000000000004a00000000",
            INIT_37 => X"0000001400000000000000260000000000000013000000000000002d00000000",
            INIT_38 => X"000000000000000000000009000000000000000e000000000000000700000000",
            INIT_39 => X"0000007000000000000000330000000000000058000000000000006f00000000",
            INIT_3A => X"0000005f00000000000000510000000000000016000000000000003c00000000",
            INIT_3B => X"0000001c00000000000000100000000000000011000000000000002700000000",
            INIT_3C => X"00000074000000000000001d000000000000002b000000000000002200000000",
            INIT_3D => X"000000670000000000000082000000000000004c000000000000007a00000000",
            INIT_3E => X"0000003c000000000000004a000000000000004b000000000000005000000000",
            INIT_3F => X"00000052000000000000004a0000000000000043000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000066000000000000004d0000000000000050000000000000005300000000",
            INIT_41 => X"00000044000000000000004c0000000000000071000000000000007600000000",
            INIT_42 => X"0000004500000000000000400000000000000041000000000000004100000000",
            INIT_43 => X"0000005c00000000000000550000000000000050000000000000004e00000000",
            INIT_44 => X"00000073000000000000004b0000000000000058000000000000006000000000",
            INIT_45 => X"00000042000000000000004b0000000000000046000000000000007500000000",
            INIT_46 => X"00000055000000000000004d0000000000000047000000000000003f00000000",
            INIT_47 => X"000000650000000000000061000000000000005a000000000000005d00000000",
            INIT_48 => X"0000005a000000000000004f0000000000000056000000000000005600000000",
            INIT_49 => X"0000004b0000000000000053000000000000004d000000000000003f00000000",
            INIT_4A => X"00000054000000000000004c0000000000000050000000000000004c00000000",
            INIT_4B => X"0000003800000000000000490000000000000062000000000000006600000000",
            INIT_4C => X"000000380000000000000039000000000000003a000000000000003800000000",
            INIT_4D => X"0000003b00000000000000490000000000000042000000000000003500000000",
            INIT_4E => X"0000002b00000000000000270000000000000020000000000000002600000000",
            INIT_4F => X"00000043000000000000003a000000000000002c000000000000003100000000",
            INIT_50 => X"000000170000000000000038000000000000003c000000000000003d00000000",
            INIT_51 => X"00000000000000000000001e000000000000002d000000000000003100000000",
            INIT_52 => X"0000002100000000000000080000000000000000000000000000000000000000",
            INIT_53 => X"0000004100000000000000320000000000000011000000000000002800000000",
            INIT_54 => X"0000001000000000000000230000000000000040000000000000004200000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000003f000000000000003b0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000013000000000000002400000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_5B => X"00000000000000000000001e0000000000000027000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000026000000000000002500000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE6;


    MEM_IFMAP_LAYER1_INSTANCE7 : if BRAM_NAME = "ifmap_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE7;


    MEM_IFMAP_LAYER2_INSTANCE0 : if BRAM_NAME = "ifmap_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000001a00000000000000000000000000000001000000000000000000000000",
            INIT_02 => X"00000000000000000000001e0000000000000021000000000000000000000000",
            INIT_03 => X"0000000000000000000000940000000000000004000000000000004b00000000",
            INIT_04 => X"000000740000000000000000000000000000004f000000000000003800000000",
            INIT_05 => X"00000038000000000000003d00000000000000c0000000000000000000000000",
            INIT_06 => X"0000000000000000000000580000000000000034000000000000007800000000",
            INIT_07 => X"000000350000000000000094000000000000004400000000000000a000000000",
            INIT_08 => X"000000bc000000000000002d0000000000000036000000000000005500000000",
            INIT_09 => X"00000000000000000000008600000000000000a0000000000000002d00000000",
            INIT_0A => X"000000fa000000000000002d0000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_0C => X"00000000000000000000003d0000000000000000000000000000001500000000",
            INIT_0D => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000b20000000000000000000000000000000000000000",
            INIT_15 => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000006800000000",
            INIT_17 => X"0000000a0000000000000008000000000000003e000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_1A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000009000000000000000b0000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_20 => X"0000000b00000000000000000000000000000020000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000400000000000000034000000000000000c000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000007a00000000000000000000000000000000000000000000006000000000",
            INIT_26 => X"0000009a0000000000000011000000000000001c000000000000001900000000",
            INIT_27 => X"0000000000000000000000490000000000000000000000000000005c00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000002200000000000000000000000000000033000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000000e000000000000003b000000000000000500000000",
            INIT_2D => X"000000000000000000000000000000000000006d000000000000002500000000",
            INIT_2E => X"0000012100000000000000cb0000000000000000000000000000000000000000",
            INIT_2F => X"0000003f0000000000000000000000000000002900000000000000f200000000",
            INIT_30 => X"0000009e00000000000000ee00000000000000fd00000000000000b700000000",
            INIT_31 => X"000000000000000000000007000000000000000e000000000000000000000000",
            INIT_32 => X"000000360000000000000000000000000000001a000000000000004400000000",
            INIT_33 => X"0000007000000000000000000000000000000062000000000000005600000000",
            INIT_34 => X"0000001800000000000000000000000000000000000000000000000400000000",
            INIT_35 => X"00000000000000000000009e0000000000000003000000000000006a00000000",
            INIT_36 => X"0000006f000000000000003b0000000000000000000000000000001e00000000",
            INIT_37 => X"000000330000000000000000000000000000006b000000000000000000000000",
            INIT_38 => X"00000029000000000000003b0000000000000079000000000000002300000000",
            INIT_39 => X"00000002000000000000003c0000000000000005000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000007500000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000005700000000000000100000000000000044000000000000000000000000",
            INIT_3E => X"0000004400000000000000360000000000000092000000000000005500000000",
            INIT_3F => X"0000002c000000000000009000000000000000b300000000000000e500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005e00000000000000570000000000000000000000000000010900000000",
            INIT_41 => X"000002090000000000000000000000000000006900000000000000e000000000",
            INIT_42 => X"000000f3000000000000003f000000000000001b000000000000002000000000",
            INIT_43 => X"0000000000000000000000fc000000000000000000000000000000fa00000000",
            INIT_44 => X"000000b40000000000000187000000000000002e000000000000002e00000000",
            INIT_45 => X"0000008500000000000000300000000000000047000000000000004a00000000",
            INIT_46 => X"000000000000000000000004000000000000016c00000000000000b800000000",
            INIT_47 => X"000000a700000000000000000000000000000005000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_49 => X"0000002300000000000000300000000000000034000000000000000700000000",
            INIT_4A => X"00000051000000000000007e000000000000009f000000000000001700000000",
            INIT_4B => X"00000042000000000000006e0000000000000063000000000000007200000000",
            INIT_4C => X"0000006a00000000000000000000000000000034000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000115000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_4F => X"0000003200000000000000000000000000000054000000000000002800000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000008500000000000000990000000000000000000000000000004500000000",
            INIT_52 => X"000000ad00000000000000460000000000000075000000000000007a00000000",
            INIT_53 => X"0000000000000000000000040000000000000000000000000000004900000000",
            INIT_54 => X"00000000000000000000000000000000000000b3000000000000004900000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_5E => X"0000009800000000000000ce0000000000000000000000000000000600000000",
            INIT_5F => X"000000d000000000000000a600000000000000a600000000000000d200000000",
            INIT_60 => X"0000011c00000000000000dd000000000000012b00000000000000bb00000000",
            INIT_61 => X"000001530000000000000123000000000000010700000000000000e400000000",
            INIT_62 => X"0000007a000000000000008500000000000000e300000000000000bd00000000",
            INIT_63 => X"00000000000000000000007f0000000000000038000000000000007700000000",
            INIT_64 => X"0000000300000000000000000000000000000016000000000000009200000000",
            INIT_65 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_67 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000005a00000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"00000000000000000000005a000000000000000c000000000000000000000000",
            INIT_6B => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_6D => X"00000014000000000000001e0000000000000013000000000000000000000000",
            INIT_6E => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002300000000000000590000000000000085000000000000003500000000",
            INIT_70 => X"0000007f0000000000000075000000000000006600000000000000a300000000",
            INIT_71 => X"000000d00000000000000080000000000000009c00000000000000bf00000000",
            INIT_72 => X"00000121000000000000010c00000000000000f500000000000000d500000000",
            INIT_73 => X"000000b400000000000000f6000000000000008d00000000000000eb00000000",
            INIT_74 => X"000000d600000000000000da00000000000000de000000000000005500000000",
            INIT_75 => X"000000bc00000000000001a900000000000000e5000000000000004b00000000",
            INIT_76 => X"0000004000000000000000b000000000000000a0000000000000008300000000",
            INIT_77 => X"0000006d0000000000000186000000000000014000000000000000ba00000000",
            INIT_78 => X"0000006100000000000000450000000000000040000000000000007f00000000",
            INIT_79 => X"000000090000000000000029000000000000005e000000000000007e00000000",
            INIT_7A => X"0000000000000000000000000000000000000022000000000000002a00000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000250000000000000029000000000000000a00000000",
            INIT_7E => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000004e00000000000000000000000000000023000000000000009200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE0;


    MEM_IFMAP_LAYER2_INSTANCE1 : if BRAM_NAME = "ifmap_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000065000000000000001a0000000000000027000000000000000000000000",
            INIT_01 => X"0000006a00000000000000860000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_03 => X"0000000000000000000000840000000000000000000000000000000000000000",
            INIT_04 => X"0000000700000000000000000000000000000000000000000000001900000000",
            INIT_05 => X"000000110000000000000000000000000000002b000000000000004500000000",
            INIT_06 => X"000000420000000000000044000000000000001b000000000000002200000000",
            INIT_07 => X"0000010900000000000000ac0000000000000048000000000000000000000000",
            INIT_08 => X"000000850000000000000095000000000000007200000000000000ae00000000",
            INIT_09 => X"000000000000000000000000000000000000004b00000000000000bd00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_0B => X"0000002000000000000000000000000000000000000000000000000400000000",
            INIT_0C => X"0000000000000000000000000000000000000064000000000000001e00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000044000000000000002a000000000000007f000000000000007000000000",
            INIT_0F => X"00000000000000000000005d000000000000004b00000000000000c900000000",
            INIT_10 => X"00000031000000000000007e0000000000000067000000000000000000000000",
            INIT_11 => X"0000005c000000000000003d000000000000003e000000000000007a00000000",
            INIT_12 => X"000000200000000000000000000000000000000c000000000000001200000000",
            INIT_13 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_14 => X"000000000000000000000000000000000000001c000000000000001900000000",
            INIT_15 => X"0000000000000000000000000000000000000065000000000000000800000000",
            INIT_16 => X"0000000000000000000000000000000000000013000000000000001600000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000008a000000000000000000000000",
            INIT_1C => X"0000009b00000000000000900000000000000000000000000000000000000000",
            INIT_1D => X"00000000000000000000002e000000000000008e000000000000007e00000000",
            INIT_1E => X"00000040000000000000004b000000000000002f000000000000000000000000",
            INIT_1F => X"0000000f000000000000001a0000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000200000000000000000000000000000001100000000",
            INIT_21 => X"00000052000000000000002d0000000000000000000000000000000f00000000",
            INIT_22 => X"00000082000000000000005d000000000000007e000000000000000000000000",
            INIT_23 => X"0000001200000000000000d50000000000000078000000000000001000000000",
            INIT_24 => X"0000006300000000000000c9000000000000005900000000000000a300000000",
            INIT_25 => X"0000007700000000000000210000000000000091000000000000001e00000000",
            INIT_26 => X"0000006f000000000000006c000000000000010f000000000000002300000000",
            INIT_27 => X"00000014000000000000002b000000000000004a000000000000007c00000000",
            INIT_28 => X"00000047000000000000004f0000000000000075000000000000008c00000000",
            INIT_29 => X"0000004800000000000000080000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000000000000000000000c100000000",
            INIT_2B => X"000000000000000000000000000000000000001f000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000007c00000000000000ad0000000000000000000000000000000000000000",
            INIT_39 => X"00000020000000000000005c0000000000000062000000000000004b00000000",
            INIT_3A => X"00000032000000000000001a000000000000000f000000000000004800000000",
            INIT_3B => X"0000002a000000000000007e0000000000000046000000000000004600000000",
            INIT_3C => X"0000000000000000000000680000000000000055000000000000002e00000000",
            INIT_3D => X"0000005300000000000000180000000000000029000000000000003500000000",
            INIT_3E => X"0000002d0000000000000000000000000000005e000000000000003900000000",
            INIT_3F => X"000000a2000000000000001c0000000000000060000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c00000000000000bd0000000000000066000000000000008100000000",
            INIT_41 => X"0000000000000000000000200000000000000077000000000000012400000000",
            INIT_42 => X"0000003600000000000000cd0000000000000040000000000000000000000000",
            INIT_43 => X"0000003a00000000000000170000000000000002000000000000001300000000",
            INIT_44 => X"00000088000000000000008600000000000000bf00000000000000aa00000000",
            INIT_45 => X"000000970000000000000093000000000000006d000000000000004f00000000",
            INIT_46 => X"000000480000000000000097000000000000008b00000000000000ad00000000",
            INIT_47 => X"0000006b0000000000000072000000000000006c000000000000007800000000",
            INIT_48 => X"0000007f0000000000000039000000000000008a000000000000002d00000000",
            INIT_49 => X"0000002e00000000000000ae0000000000000027000000000000005300000000",
            INIT_4A => X"0000008500000000000000670000000000000053000000000000007600000000",
            INIT_4B => X"00000000000000000000003d0000000000000028000000000000000000000000",
            INIT_4C => X"00000000000000000000001d0000000000000000000000000000003600000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000c00000000000000510000000000000014000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000200000000000000000000000000000000000000000000004900000000",
            INIT_53 => X"0000002800000000000000180000000000000013000000000000004800000000",
            INIT_54 => X"000000df00000000000000070000000000000000000000000000003200000000",
            INIT_55 => X"0000000000000000000000000000000000000003000000000000002900000000",
            INIT_56 => X"00000000000000000000003a0000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000620000000000000000000000000000004900000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"000000000000000000000000000000000000003a000000000000000000000000",
            INIT_5F => X"0000004500000000000000040000000000000001000000000000005000000000",
            INIT_60 => X"0000008e00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"00000053000000000000007b000000000000002d000000000000008300000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000006100000000",
            INIT_63 => X"000000fb00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"00000021000000000000000f0000000000000031000000000000002f00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000007100000000000000790000000000000071000000000000000000000000",
            INIT_67 => X"0000002f00000000000000000000000000000000000000000000003d00000000",
            INIT_68 => X"0000000000000000000000660000000000000027000000000000003900000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"000000a500000000000000bb00000000000000a300000000000000b200000000",
            INIT_76 => X"00000050000000000000009e0000000000000044000000000000008800000000",
            INIT_77 => X"00000033000000000000003c000000000000008900000000000000bd00000000",
            INIT_78 => X"0000009700000000000000000000000000000021000000000000000000000000",
            INIT_79 => X"0000000000000000000000320000000000000000000000000000005400000000",
            INIT_7A => X"0000005000000000000000620000000000000000000000000000000000000000",
            INIT_7B => X"0000001300000000000000000000000000000011000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE1;


    MEM_IFMAP_LAYER2_INSTANCE2 : if BRAM_NAME = "ifmap_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000007000000000000001c0000000000000031000000000000000000000000",
            INIT_02 => X"000000250000000000000000000000000000000b000000000000003e00000000",
            INIT_03 => X"00000000000000000000002d000000000000000e000000000000002e00000000",
            INIT_04 => X"000000000000000000000031000000000000001b000000000000005b00000000",
            INIT_05 => X"000000570000000000000000000000000000003900000000000000d300000000",
            INIT_06 => X"0000000800000000000000000000000000000000000000000000000500000000",
            INIT_07 => X"00000031000000000000009e000000000000004d00000000000000af00000000",
            INIT_08 => X"00000022000000000000001d000000000000001d000000000000001700000000",
            INIT_09 => X"0000000000000000000000430000000000000083000000000000000000000000",
            INIT_0A => X"00000071000000000000009d0000000000000070000000000000008b00000000",
            INIT_0B => X"0000006200000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000000000000000000000000000d000000000000013000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_11 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_19 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000034000000000000008600000000",
            INIT_1B => X"0000000600000000000000000000000000000000000000000000003100000000",
            INIT_1C => X"0000006a00000000000000000000000000000052000000000000004500000000",
            INIT_1D => X"0000000000000000000000000000000000000061000000000000000000000000",
            INIT_1E => X"000000210000000000000055000000000000000000000000000000a500000000",
            INIT_1F => X"000000000000000000000000000000000000000000000000000000d500000000",
            INIT_20 => X"0000007b00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000370000000000000023000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000c900000000000000b30000000000000000000000000000000000000000",
            INIT_24 => X"000000720000000000000000000000000000000000000000000000d700000000",
            INIT_25 => X"000000d200000000000000ad00000000000000d900000000000000be00000000",
            INIT_26 => X"00000130000000000000012a0000000000000153000000000000016b00000000",
            INIT_27 => X"0000005e00000000000000eb000000000000004a000000000000006400000000",
            INIT_28 => X"00000000000000000000003f000000000000005a000000000000010b00000000",
            INIT_29 => X"0000010b00000000000000480000000000000059000000000000004b00000000",
            INIT_2A => X"0000005c00000000000000000000000000000018000000000000004300000000",
            INIT_2B => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_2C => X"0000003000000000000000720000000000000016000000000000005400000000",
            INIT_2D => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_2E => X"00000007000000000000001e0000000000000017000000000000005400000000",
            INIT_2F => X"00000008000000000000003300000000000000b7000000000000000000000000",
            INIT_30 => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000028000000000000000c000000000000001c000000000000004100000000",
            INIT_32 => X"0000007a0000000000000046000000000000005d000000000000000200000000",
            INIT_33 => X"00000067000000000000005f000000000000002e000000000000004400000000",
            INIT_34 => X"00000049000000000000008c000000000000006f00000000000000cb00000000",
            INIT_35 => X"000000ab00000000000000680000000000000039000000000000005c00000000",
            INIT_36 => X"000000a7000000000000003900000000000000b200000000000000a100000000",
            INIT_37 => X"000000a700000000000000730000000000000025000000000000004600000000",
            INIT_38 => X"0000001c0000000000000090000000000000000000000000000000c000000000",
            INIT_39 => X"000000ac000000000000007f000000000000003a000000000000003700000000",
            INIT_3A => X"000000ac00000000000000320000000000000076000000000000009e00000000",
            INIT_3B => X"0000002b0000000000000078000000000000011d00000000000000a700000000",
            INIT_3C => X"0000007b00000000000000220000000000000029000000000000000000000000",
            INIT_3D => X"000000060000000000000000000000000000000000000000000000b600000000",
            INIT_3E => X"000000000000000000000000000000000000002f000000000000000700000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000006c00000000000000130000000000000013000000000000000000000000",
            INIT_47 => X"0000007000000000000000000000000000000058000000000000001400000000",
            INIT_48 => X"000001bf00000000000001ba000000000000015b00000000000000df00000000",
            INIT_49 => X"0000019f0000000000000136000000000000007f000000000000017300000000",
            INIT_4A => X"0000000000000000000001da00000000000001e000000000000001c400000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000910000000000000000000000000000005b000000000000000000000000",
            INIT_4F => X"0000002100000000000000000000000000000000000000000000004100000000",
            INIT_50 => X"000000000000000000000000000000000000000000000000000000b300000000",
            INIT_51 => X"000000ef000000000000000c0000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000930000000000000000000000000000007200000000",
            INIT_53 => X"000000000000000000000076000000000000000f000000000000000000000000",
            INIT_54 => X"00000090000000000000007d0000000000000024000000000000000000000000",
            INIT_55 => X"0000005a000000000000008b000000000000000000000000000000af00000000",
            INIT_56 => X"000000ab000000000000008b000000000000009a000000000000008e00000000",
            INIT_57 => X"0000002100000000000000290000000000000001000000000000000f00000000",
            INIT_58 => X"0000001b00000000000000290000000000000032000000000000005000000000",
            INIT_59 => X"0000005d00000000000000600000000000000048000000000000002200000000",
            INIT_5A => X"0000003c00000000000000000000000000000054000000000000003c00000000",
            INIT_5B => X"00000039000000000000004d0000000000000031000000000000003500000000",
            INIT_5C => X"0000004400000000000000500000000000000000000000000000005400000000",
            INIT_5D => X"0000004f0000000000000037000000000000003b000000000000001600000000",
            INIT_5E => X"0000001d000000000000003a000000000000001a000000000000000000000000",
            INIT_5F => X"000000000000000000000034000000000000003c000000000000005000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000002900000000000000000000000000000000000000000000000900000000",
            INIT_67 => X"0000000a00000000000000000000000000000056000000000000002100000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_6C => X"00000000000000000000005c00000000000000ea000000000000000000000000",
            INIT_6D => X"000000000000000000000052000000000000008d000000000000000000000000",
            INIT_6E => X"00000047000000000000001b0000000000000000000000000000000000000000",
            INIT_6F => X"000000a200000000000000b10000000000000049000000000000003e00000000",
            INIT_70 => X"000000d800000000000000c6000000000000011f00000000000000d200000000",
            INIT_71 => X"0000010100000000000000c500000000000000b900000000000000d100000000",
            INIT_72 => X"000000550000000000000079000000000000000800000000000000ce00000000",
            INIT_73 => X"000000c5000000000000003f0000000000000094000000000000009000000000",
            INIT_74 => X"000000a7000000000000002e00000000000000ac000000000000000000000000",
            INIT_75 => X"0000000000000000000000b5000000000000004300000000000000b700000000",
            INIT_76 => X"0000003e000000000000003f0000000000000009000000000000005400000000",
            INIT_77 => X"0000002800000000000000910000000000000038000000000000008d00000000",
            INIT_78 => X"0000004600000000000000000000000000000000000000000000002600000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000004200000000000000020000000000000002000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000032000000000000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE2;


    MEM_IFMAP_LAYER2_INSTANCE3 : if BRAM_NAME = "ifmap_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002600000000000000510000000000000000000000000000000800000000",
            INIT_01 => X"0000009700000000000000000000000000000012000000000000004e00000000",
            INIT_02 => X"0000003b0000000000000013000000000000002f000000000000000000000000",
            INIT_03 => X"0000009000000000000000000000000000000007000000000000000000000000",
            INIT_04 => X"00000000000000000000003a0000000000000000000000000000006600000000",
            INIT_05 => X"0000001c000000000000002f000000000000008c00000000000000ad00000000",
            INIT_06 => X"00000069000000000000005b000000000000003b000000000000002800000000",
            INIT_07 => X"0000002700000000000000750000000000000046000000000000006600000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE3;


    MEM_IFMAP_LAYER3_INSTANCE0 : if BRAM_NAME = "ifmap_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000001240000000000000087000000000000003a000000000000004c00000000",
            INIT_02 => X"00000000000000000000000000000000000000c1000000000000000000000000",
            INIT_03 => X"000000ab00000000000000880000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000000000000000001c9000000000000022b00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000b400000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000000000000000000000000000000000000f1000000000000011500000000",
            INIT_08 => X"000000b6000000000000000000000000000000de000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000005e000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000035b00000000000002250000000000000000000000000000000000000000",
            INIT_0E => X"0000019100000000000001a800000000000003f7000000000000024a00000000",
            INIT_0F => X"000000a800000000000001e700000000000001ae00000000000002de00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000670000000000000121000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000000000006b0000000000000000000000000000000000000000",
            INIT_17 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000023300000000000000000000000000000000000000000000009700000000",
            INIT_19 => X"0000018c000000000000011700000000000001ac00000000000001e100000000",
            INIT_1A => X"000002d9000000000000025100000000000002fc00000000000000b200000000",
            INIT_1B => X"0000000000000000000001300000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000001330000000000000000000000000000000000000000",
            INIT_1D => X"000000d800000000000000540000000000000148000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000013b00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000000000000000000000000000000000009d000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000004c000000000000010b000000000000000000000000",
            INIT_2D => X"000000000000000000000101000000000000002d000000000000008f00000000",
            INIT_2E => X"000000000000000000000000000000000000012f000000000000001d00000000",
            INIT_2F => X"000000b900000000000000260000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000440000000000000040000000000000000000000000",
            INIT_32 => X"0000000800000000000000ac0000000000000000000000000000003d00000000",
            INIT_33 => X"00000000000000000000001f0000000000000018000000000000000d00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000be00000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000016600000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000d9000000000000001d0000000000000000000000000000000000000000",
            INIT_3B => X"0000013f00000000000001310000000000000000000000000000020700000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"000000000000000000000000000000000000000000000000000000a400000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000000000000000000000000000000000000c800000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000a000000000000000000000000000000cf000000000000009f00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000b00000000000000800000000000000082000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_4E => X"00000000000000000000029c0000000000000177000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_51 => X"00000024000000000000019600000000000001a5000000000000014c00000000",
            INIT_52 => X"00000000000000000000000000000000000000bc000000000000018700000000",
            INIT_53 => X"00000181000000000000024d0000000000000324000000000000000000000000",
            INIT_54 => X"0000020600000000000002e000000000000002b900000000000002c800000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000009d00000000000001800000000000000000000000000000000000000000",
            INIT_5C => X"0000005a00000000000000000000000000000000000000000000011b00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000001e00000000000000530000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000a40000000000000000000000000000005d00000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000000000000000000124000000000000013b000000000000005100000000",
            INIT_6A => X"000000f2000000000000004f0000000000000000000000000000000000000000",
            INIT_6B => X"0000003d00000000000000510000000000000000000000000000011400000000",
            INIT_6C => X"0000017f000000000000007c0000000000000088000000000000000f00000000",
            INIT_6D => X"0000005e00000000000001650000000000000061000000000000014000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000a500000000000000220000000000000000000000000000000000000000",
            INIT_71 => X"000000e900000000000001330000000000000232000000000000010c00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000011d00000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000bb00000000000001b40000000000000000000000000000008f00000000",
            INIT_77 => X"000000ba0000000000000000000000000000000000000000000000dd00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000012e00000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000020900000000000001ba000000000000015b000000000000018200000000",
            INIT_7D => X"0000001300000000000000a60000000000000012000000000000016800000000",
            INIT_7E => X"000000b700000000000001c000000000000000ee00000000000000ea00000000",
            INIT_7F => X"00000000000000000000001e0000000000000000000000000000013d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER3_INSTANCE0;


    MEM_IFMAP_LAYER3_INSTANCE1 : if BRAM_NAME = "ifmap_layer3_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000d5000000000000011d0000000000000000000000000000000000000000",
            INIT_03 => X"000001a1000000000000018300000000000000f3000000000000008f00000000",
            INIT_04 => X"0000000000000000000000000000000000000050000000000000010000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000011700000000000000000000000000000034000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000ac00000000000000000000000000000000000000000000016700000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001f0000000000000000000000000000000000000000000000a400000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER3_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE0 : if BRAM_NAME = "gold_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000009000000000000000a0000000000000010000000000000001000000000",
            INIT_01 => X"0000000d000000000000000c0000000000000008000000000000000600000000",
            INIT_02 => X"0000000f0000000000000014000000000000000b000000000000000500000000",
            INIT_03 => X"0000000000000000000000010000000000000002000000000000000700000000",
            INIT_04 => X"0000000a000000000000000b0000000000000009000000000000000300000000",
            INIT_05 => X"0000002900000000000000050000000000000003000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000001f000000000000000f0000000000000000000000000000000500000000",
            INIT_08 => X"0000004c000000000000000c000000000000000a000000000000000800000000",
            INIT_09 => X"0000000000000000000000000000000000000013000000000000002c00000000",
            INIT_0A => X"0000000000000000000000000000000000000012000000000000002100000000",
            INIT_0B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000030000000000000000000000000000000300000000",
            INIT_0D => X"0000002d00000000000000290000000000000001000000000000000800000000",
            INIT_0E => X"000000000000000000000000000000000000001c000000000000002400000000",
            INIT_0F => X"0000000e00000000000000110000000000000000000000000000002700000000",
            INIT_10 => X"000000130000000000000033000000000000000a000000000000000000000000",
            INIT_11 => X"0000000b00000000000000110000000000000000000000000000000d00000000",
            INIT_12 => X"0000006900000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000007f000000000000003a0000000000000027000000000000002b00000000",
            INIT_14 => X"0000000000000000000000140000000000000025000000000000007c00000000",
            INIT_15 => X"0000000e000000000000003c0000000000000053000000000000000000000000",
            INIT_16 => X"0000002a000000000000005e0000000000000000000000000000000300000000",
            INIT_17 => X"0000001a000000000000001e0000000000000013000000000000002e00000000",
            INIT_18 => X"000000000000000000000017000000000000002c000000000000004f00000000",
            INIT_19 => X"0000000000000000000000010000000000000013000000000000005600000000",
            INIT_1A => X"00000007000000000000003b0000000000000058000000000000000200000000",
            INIT_1B => X"00000080000000000000003b000000000000000b000000000000000000000000",
            INIT_1C => X"0000004d000000000000001e000000000000002c000000000000005000000000",
            INIT_1D => X"000000200000000000000025000000000000000f000000000000002300000000",
            INIT_1E => X"0000000e0000000000000041000000000000004f000000000000005f00000000",
            INIT_1F => X"0000000000000000000000320000000000000069000000000000001300000000",
            INIT_20 => X"0000004800000000000000350000000000000012000000000000000100000000",
            INIT_21 => X"0000007100000000000000000000000000000003000000000000001500000000",
            INIT_22 => X"0000002e000000000000000c0000000000000040000000000000005e00000000",
            INIT_23 => X"000000170000000000000000000000000000001b000000000000002400000000",
            INIT_24 => X"0000000000000000000000000000000000000035000000000000004b00000000",
            INIT_25 => X"000000540000000000000035000000000000000f000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_27 => X"00000000000000000000003c0000000000000072000000000000002200000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000004c00000000000000670000000000000056000000000000000100000000",
            INIT_2A => X"00000047000000000000008700000000000000c4000000000000002100000000",
            INIT_2B => X"0000000c00000000000000110000000000000027000000000000004800000000",
            INIT_2C => X"0000001e00000000000000170000000000000014000000000000001500000000",
            INIT_2D => X"0000006d00000000000000510000000000000044000000000000001000000000",
            INIT_2E => X"000000130000000000000016000000000000001500000000000000a300000000",
            INIT_2F => X"0000000700000000000000060000000000000007000000000000000f00000000",
            INIT_30 => X"00000023000000000000000e000000000000002a000000000000001f00000000",
            INIT_31 => X"000000390000000000000090000000000000004d000000000000000a00000000",
            INIT_32 => X"000000160000000000000010000000000000000f000000000000001500000000",
            INIT_33 => X"00000024000000000000002c000000000000001f000000000000001400000000",
            INIT_34 => X"000000180000000000000029000000000000004a000000000000000b00000000",
            INIT_35 => X"0000002600000000000000240000000000000050000000000000001c00000000",
            INIT_36 => X"0000000b000000000000000c000000000000001c000000000000003100000000",
            INIT_37 => X"0000001b0000000000000003000000000000001a000000000000001b00000000",
            INIT_38 => X"00000080000000000000007c000000000000007a000000000000001f00000000",
            INIT_39 => X"00000081000000000000007c0000000000000080000000000000008000000000",
            INIT_3A => X"0000006100000000000000710000000000000087000000000000008b00000000",
            INIT_3B => X"0000007000000000000000710000000000000069000000000000006400000000",
            INIT_3C => X"0000008200000000000000870000000000000083000000000000008100000000",
            INIT_3D => X"000000740000000000000072000000000000007b000000000000008300000000",
            INIT_3E => X"0000002d0000000000000025000000000000003c000000000000004e00000000",
            INIT_3F => X"00000060000000000000006b000000000000005d000000000000004600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008700000000000000850000000000000082000000000000006700000000",
            INIT_41 => X"000000310000000000000035000000000000003e000000000000007100000000",
            INIT_42 => X"0000001700000000000000190000000000000017000000000000002f00000000",
            INIT_43 => X"0000005c00000000000000140000000000000059000000000000003e00000000",
            INIT_44 => X"0000005900000000000000720000000000000088000000000000007200000000",
            INIT_45 => X"0000003b000000000000001b0000000000000025000000000000003500000000",
            INIT_46 => X"0000001f000000000000000e0000000000000023000000000000001400000000",
            INIT_47 => X"00000059000000000000003d0000000000000000000000000000005500000000",
            INIT_48 => X"0000001a000000000000003d0000000000000043000000000000008700000000",
            INIT_49 => X"00000024000000000000003e0000000000000016000000000000001900000000",
            INIT_4A => X"0000004200000000000000140000000000000022000000000000001800000000",
            INIT_4B => X"0000005f000000000000004d0000000000000022000000000000000400000000",
            INIT_4C => X"0000002000000000000000180000000000000028000000000000003600000000",
            INIT_4D => X"0000000c0000000000000014000000000000005c000000000000000d00000000",
            INIT_4E => X"00000009000000000000001b0000000000000016000000000000002600000000",
            INIT_4F => X"0000005500000000000000500000000000000044000000000000000300000000",
            INIT_50 => X"0000000b00000000000000170000000000000020000000000000004300000000",
            INIT_51 => X"0000001e00000000000000110000000000000001000000000000004600000000",
            INIT_52 => X"00000000000000000000000c0000000000000020000000000000001f00000000",
            INIT_53 => X"0000004500000000000000520000000000000035000000000000002c00000000",
            INIT_54 => X"0000004b0000000000000016000000000000001a000000000000000a00000000",
            INIT_55 => X"000000240000000000000024000000000000000d000000000000001100000000",
            INIT_56 => X"0000000000000000000000050000000000000001000000000000003d00000000",
            INIT_57 => X"0000001c00000000000000200000000000000031000000000000002300000000",
            INIT_58 => X"0000003100000000000000270000000000000033000000000000002000000000",
            INIT_59 => X"00000066000000000000003c0000000000000024000000000000000d00000000",
            INIT_5A => X"000000190000000000000000000000000000000d000000000000000d00000000",
            INIT_5B => X"0000000f00000000000000300000000000000033000000000000001000000000",
            INIT_5C => X"00000014000000000000000a0000000000000028000000000000002c00000000",
            INIT_5D => X"0000000f00000000000000680000000000000062000000000000003400000000",
            INIT_5E => X"0000000000000000000000470000000000000000000000000000000f00000000",
            INIT_5F => X"000000000000000000000000000000000000001f000000000000001600000000",
            INIT_60 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"000000000000000000000000000000000000003b000000000000000200000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000110000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE0;


    MEM_GOLD_LAYER0_INSTANCE1 : if BRAM_NAME = "gold_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_03 => X"0000000000000000000000170000000000000016000000000000000000000000",
            INIT_04 => X"0000000f000000000000000b0000000000000025000000000000000000000000",
            INIT_05 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000021000000000000001200000000",
            INIT_08 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_0A => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_0C => X"000000000000000000000000000000000000000b000000000000002300000000",
            INIT_0D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_0E => X"0000003c00000000000000320000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000005000000000000000700000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_12 => X"00000020000000000000002f000000000000002e000000000000000000000000",
            INIT_13 => X"000000000000000000000000000000000000001c000000000000000b00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000170000000000000022000000000000002c000000000000003500000000",
            INIT_17 => X"0000003600000000000000180000000000000016000000000000002c00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_19 => X"00000041000000000000001b000000000000001b000000000000000600000000",
            INIT_1A => X"0000006200000000000000320000000000000028000000000000003600000000",
            INIT_1B => X"0000002000000000000000290000000000000025000000000000003000000000",
            INIT_1C => X"00000025000000000000001e000000000000001b000000000000001800000000",
            INIT_1D => X"0000002900000000000000260000000000000029000000000000002500000000",
            INIT_1E => X"0000001a00000000000000380000000000000057000000000000002000000000",
            INIT_1F => X"0000001600000000000000140000000000000014000000000000001900000000",
            INIT_20 => X"0000002d000000000000002a0000000000000027000000000000002000000000",
            INIT_21 => X"0000002a00000000000000230000000000000035000000000000003200000000",
            INIT_22 => X"0000001a000000000000001a000000000000001b000000000000005800000000",
            INIT_23 => X"0000002600000000000000200000000000000019000000000000001800000000",
            INIT_24 => X"000000390000000000000037000000000000002c000000000000003100000000",
            INIT_25 => X"0000003c000000000000001e000000000000002a000000000000003000000000",
            INIT_26 => X"00000017000000000000001e0000000000000019000000000000001300000000",
            INIT_27 => X"0000002000000000000000260000000000000023000000000000001a00000000",
            INIT_28 => X"00000011000000000000002e0000000000000042000000000000002d00000000",
            INIT_29 => X"0000001000000000000000150000000000000015000000000000001a00000000",
            INIT_2A => X"0000000a000000000000000a000000000000000f000000000000001900000000",
            INIT_2B => X"0000001800000000000000150000000000000011000000000000000b00000000",
            INIT_2C => X"0000000e000000000000000b0000000000000006000000000000000a00000000",
            INIT_2D => X"0000005000000000000000190000000000000013000000000000001100000000",
            INIT_2E => X"0000003800000000000000110000000000000010000000000000000e00000000",
            INIT_2F => X"0000000f0000000000000014000000000000001c000000000000003700000000",
            INIT_30 => X"0000000f00000000000000160000000000000011000000000000000b00000000",
            INIT_31 => X"000000350000000000000041000000000000000d000000000000001000000000",
            INIT_32 => X"00000070000000000000006b000000000000001c000000000000001900000000",
            INIT_33 => X"0000001d00000000000000050000000000000030000000000000006600000000",
            INIT_34 => X"00000011000000000000000c000000000000001d000000000000002b00000000",
            INIT_35 => X"0000003d000000000000004d0000000000000033000000000000001b00000000",
            INIT_36 => X"000000460000000000000079000000000000005e000000000000004100000000",
            INIT_37 => X"000000840000000000000012000000000000000f000000000000004800000000",
            INIT_38 => X"0000009e000000000000003d0000000000000022000000000000006a00000000",
            INIT_39 => X"000000380000000000000053000000000000007e000000000000007600000000",
            INIT_3A => X"0000004600000000000000460000000000000079000000000000005400000000",
            INIT_3B => X"000000b000000000000000980000000000000000000000000000002a00000000",
            INIT_3C => X"000000a100000000000000c1000000000000002c000000000000003d00000000",
            INIT_3D => X"000000780000000000000038000000000000005b00000000000000a100000000",
            INIT_3E => X"00000049000000000000004c000000000000005d000000000000009b00000000",
            INIT_3F => X"0000003600000000000000a300000000000000a3000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac00000000000000970000000000000059000000000000001c00000000",
            INIT_41 => X"00000095000000000000008f0000000000000051000000000000008700000000",
            INIT_42 => X"0000004000000000000000580000000000000047000000000000005300000000",
            INIT_43 => X"00000036000000000000004400000000000000c900000000000000b800000000",
            INIT_44 => X"0000007800000000000000af00000000000000af000000000000003b00000000",
            INIT_45 => X"000000550000000000000094000000000000007f000000000000005b00000000",
            INIT_46 => X"000000dc00000000000000430000000000000058000000000000004d00000000",
            INIT_47 => X"0000004b0000000000000080000000000000008200000000000000d700000000",
            INIT_48 => X"00000055000000000000005a0000000000000061000000000000006e00000000",
            INIT_49 => X"00000036000000000000004a000000000000004d000000000000004000000000",
            INIT_4A => X"000000d800000000000000e80000000000000021000000000000004300000000",
            INIT_4B => X"0000004e0000000000000067000000000000008f000000000000009f00000000",
            INIT_4C => X"0000005a000000000000004f0000000000000090000000000000007d00000000",
            INIT_4D => X"000000290000000000000026000000000000001a000000000000004000000000",
            INIT_4E => X"0000009f00000000000000c900000000000000d0000000000000001e00000000",
            INIT_4F => X"000000a5000000000000006e00000000000000e100000000000000d400000000",
            INIT_50 => X"000000380000000000000043000000000000007d00000000000000c800000000",
            INIT_51 => X"00000053000000000000005f000000000000005a000000000000004c00000000",
            INIT_52 => X"000000f700000000000000ba00000000000000e200000000000000a600000000",
            INIT_53 => X"00000084000000000000008500000000000000a200000000000000e500000000",
            INIT_54 => X"00000089000000000000007d0000000000000072000000000000007a00000000",
            INIT_55 => X"000000940000000000000099000000000000009a000000000000009900000000",
            INIT_56 => X"000000bb00000000000000f900000000000000d7000000000000009700000000",
            INIT_57 => X"0000007b000000000000007c000000000000007f000000000000008900000000",
            INIT_58 => X"0000009d000000000000009a0000000000000090000000000000008000000000",
            INIT_59 => X"0000008a00000000000000a800000000000000ba00000000000000a400000000",
            INIT_5A => X"0000008e000000000000009100000000000000fa00000000000000a600000000",
            INIT_5B => X"000000910000000000000085000000000000007b000000000000008800000000",
            INIT_5C => X"000000b200000000000000a200000000000000a2000000000000009b00000000",
            INIT_5D => X"00000089000000000000009f00000000000000ac00000000000000af00000000",
            INIT_5E => X"0000008d000000000000007f0000000000000073000000000000009300000000",
            INIT_5F => X"00000092000000000000009f0000000000000091000000000000008e00000000",
            INIT_60 => X"0000009600000000000000c800000000000000ba000000000000009700000000",
            INIT_61 => X"0000006f000000000000006c000000000000006d000000000000007100000000",
            INIT_62 => X"0000007c00000000000000710000000000000062000000000000007100000000",
            INIT_63 => X"000000620000000000000068000000000000006e000000000000007700000000",
            INIT_64 => X"0000006d000000000000006a0000000000000062000000000000005f00000000",
            INIT_65 => X"0000006c0000000000000073000000000000006c000000000000006800000000",
            INIT_66 => X"0000007500000000000000670000000000000061000000000000003c00000000",
            INIT_67 => X"00000046000000000000002a000000000000001d000000000000003a00000000",
            INIT_68 => X"00000076000000000000006d0000000000000062000000000000005c00000000",
            INIT_69 => X"0000008f00000000000000770000000000000076000000000000007200000000",
            INIT_6A => X"0000000d00000000000000260000000000000058000000000000007f00000000",
            INIT_6B => X"0000003a000000000000002c0000000000000028000000000000002900000000",
            INIT_6C => X"0000006800000000000000030000000000000038000000000000005100000000",
            INIT_6D => X"00000026000000000000004c0000000000000067000000000000006e00000000",
            INIT_6E => X"0000004f0000000000000022000000000000002c000000000000002800000000",
            INIT_6F => X"00000037000000000000002f0000000000000048000000000000003d00000000",
            INIT_70 => X"0000003900000000000000650000000000000000000000000000003000000000",
            INIT_71 => X"00000036000000000000003d0000000000000003000000000000000000000000",
            INIT_72 => X"0000002f0000000000000023000000000000000c000000000000003e00000000",
            INIT_73 => X"0000004300000000000000260000000000000028000000000000002400000000",
            INIT_74 => X"000000650000000000000076000000000000006a000000000000002a00000000",
            INIT_75 => X"0000002f0000000000000030000000000000003e000000000000005800000000",
            INIT_76 => X"0000002800000000000000570000000000000051000000000000000000000000",
            INIT_77 => X"0000003a00000000000000310000000000000012000000000000002b00000000",
            INIT_78 => X"000000250000000000000037000000000000007b000000000000006200000000",
            INIT_79 => X"00000000000000000000003e0000000000000040000000000000004900000000",
            INIT_7A => X"0000001b00000000000000270000000000000036000000000000005c00000000",
            INIT_7B => X"0000001c000000000000002f000000000000002b000000000000002900000000",
            INIT_7C => X"0000007800000000000000190000000000000025000000000000004900000000",
            INIT_7D => X"0000005d0000000000000024000000000000004d000000000000005c00000000",
            INIT_7E => X"0000005200000000000000380000000000000023000000000000004700000000",
            INIT_7F => X"0000002000000000000000460000000000000022000000000000003400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE2 : if BRAM_NAME = "gold_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003000000000000000510000000000000066000000000000003b00000000",
            INIT_01 => X"00000070000000000000004c0000000000000055000000000000001a00000000",
            INIT_02 => X"0000005200000000000000400000000000000035000000000000003800000000",
            INIT_03 => X"0000002d0000000000000004000000000000004c000000000000003100000000",
            INIT_04 => X"0000002400000000000000130000000000000024000000000000003300000000",
            INIT_05 => X"00000002000000000000002b0000000000000065000000000000006000000000",
            INIT_06 => X"000000300000000000000025000000000000006d000000000000003600000000",
            INIT_07 => X"0000000000000000000000030000000000000000000000000000005800000000",
            INIT_08 => X"0000002b000000000000003f000000000000004b000000000000000000000000",
            INIT_09 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000280000000000000037000000000000001e000000000000002800000000",
            INIT_0B => X"000000380000000000000074000000000000009d000000000000000000000000",
            INIT_0C => X"00000002000000000000000c000000000000001f000000000000003700000000",
            INIT_0D => X"0000000400000000000000000000000000000000000000000000000200000000",
            INIT_0E => X"0000004e00000000000000180000000000000016000000000000000000000000",
            INIT_0F => X"0000000700000000000000040000000000000004000000000000008800000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_11 => X"0000000400000000000000000000000000000005000000000000000000000000",
            INIT_12 => X"00000032000000000000008b0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_14 => X"0000000700000000000000090000000000000002000000000000000000000000",
            INIT_15 => X"000000000000000000000005000000000000001c000000000000000000000000",
            INIT_16 => X"0000001400000000000000230000000000000043000000000000000500000000",
            INIT_17 => X"0000000000000000000000000000000000000009000000000000001900000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000001300000000000000030000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_20 => X"000000120000000000000000000000000000000d000000000000000500000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_22 => X"00000000000000000000000a0000000000000005000000000000003e00000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000009000000000000000a00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000001c0000000000000000000000000000000d000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000016000000000000000c00000000",
            INIT_36 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000300000000000000000000000000000000000000000",
            INIT_39 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000007000000000000002600000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000f000000000000002a0000000000000031000000000000000000000000",
            INIT_3E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000007000000000000002e0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001d00000000000000480000000000000004000000000000000700000000",
            INIT_43 => X"00000031000000000000002e0000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000070000000000000019000000000000001c00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000004f00000000000000140000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_4E => X"0000000300000000000000490000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000014000000000000000c00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_52 => X"0000000200000000000000000000000000000000000000000000000600000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000030000000000000009000000000000000000000000",
            INIT_55 => X"0000000600000000000000010000000000000001000000000000000000000000",
            INIT_56 => X"00000000000000000000001d000000000000000d000000000000000000000000",
            INIT_57 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000120000000000000004000000000000000000000000",
            INIT_59 => X"0000000000000000000000030000000000000039000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000007000000000000000900000000",
            INIT_5B => X"0000000000000000000000000000000000000051000000000000000b00000000",
            INIT_5C => X"00000000000000000000001f000000000000000a000000000000000000000000",
            INIT_5D => X"00000000000000000000000c0000000000000000000000000000006500000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000006800000000",
            INIT_60 => X"0000001d00000000000000000000000000000055000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000066000000000000000000000000",
            INIT_62 => X"0000009400000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000080000000000000000000000000000001e00000000",
            INIT_65 => X"0000000000000000000000000000000000000068000000000000001e00000000",
            INIT_66 => X"0000000000000000000001010000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000056000000000000006100000000",
            INIT_6A => X"00000000000000000000000000000000000000cb000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000015000000000000000400000000",
            INIT_6C => X"0000004300000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000005f00000000",
            INIT_6E => X"0000002100000000000000000000000000000000000000000000008000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000090000000000000000000000000000002f000000000000000000000000",
            INIT_71 => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_72 => X"00000020000000000000001f0000000000000000000000000000000e00000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_74 => X"0000003900000000000000080000000000000000000000000000005500000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000002e000000000000002d000000000000000000000000",
            INIT_77 => X"000000dc00000000000000000000000000000000000000000000005e00000000",
            INIT_78 => X"00000000000000000000004b0000000000000000000000000000000000000000",
            INIT_79 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000004e0000000000000000000000000000000a000000000000000d00000000",
            INIT_7B => X"0000000000000000000000960000000000000000000000000000004100000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000500000000000000060000000000000002000000000000000000000000",
            INIT_7E => X"0000005200000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000008500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE2;


    MEM_GOLD_LAYER0_INSTANCE3 : if BRAM_NAME = "gold_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000400000000000000000000000000000005000000000000000800000000",
            INIT_02 => X"000000ac00000000000000000000000000000000000000000000000e00000000",
            INIT_03 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000040000000000000006000000000000000000000000",
            INIT_05 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_06 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000080000000000000016000000000000000000000000",
            INIT_08 => X"0000000400000000000000000000000000000000000000000000000c00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000008000000000000001c00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000001b0000000000000022000000000000000b000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000018000000000000002800000000",
            INIT_15 => X"0000000000000000000000000000000000000007000000000000001b00000000",
            INIT_16 => X"0000001500000000000000050000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000060000000000000000000000000000001700000000",
            INIT_18 => X"000000340000000000000000000000000000000d000000000000000d00000000",
            INIT_19 => X"0000002700000000000000000000000000000000000000000000002900000000",
            INIT_1A => X"0000000f00000000000000160000000000000005000000000000001500000000",
            INIT_1B => X"0000002000000000000000150000000000000017000000000000001100000000",
            INIT_1C => X"00000010000000000000001a0000000000000000000000000000002600000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000024000000000000002a0000000000000016000000000000000a00000000",
            INIT_1F => X"0000002600000000000000140000000000000007000000000000000100000000",
            INIT_20 => X"00000000000000000000000e000000000000002b000000000000002e00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000300000000000000150000000000000018000000000000000f00000000",
            INIT_23 => X"000000170000000000000021000000000000001c000000000000001c00000000",
            INIT_24 => X"0000000000000000000000170000000000000032000000000000002100000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000f00000000000000000000000000000000000000000000000100000000",
            INIT_27 => X"0000002a00000000000000000000000000000000000000000000001500000000",
            INIT_28 => X"00000000000000000000000e0000000000000022000000000000002a00000000",
            INIT_29 => X"0000001600000000000000120000000000000000000000000000000000000000",
            INIT_2A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000001900000000000000090000000000000000000000000000000000000000",
            INIT_2C => X"0000000e0000000000000010000000000000002f000000000000002800000000",
            INIT_2D => X"000000000000000000000011000000000000002e000000000000001900000000",
            INIT_2E => X"00000000000000000000001c000000000000001e000000000000000000000000",
            INIT_2F => X"0000001c0000000000000016000000000000001c000000000000000000000000",
            INIT_30 => X"0000002f00000000000000590000000000000066000000000000004e00000000",
            INIT_31 => X"000000620000000000000041000000000000002c000000000000001700000000",
            INIT_32 => X"0000003b00000000000000420000000000000068000000000000007200000000",
            INIT_33 => X"0000001f000000000000002d0000000000000027000000000000003e00000000",
            INIT_34 => X"00000041000000000000003b0000000000000020000000000000000000000000",
            INIT_35 => X"0000007c0000000000000079000000000000006c000000000000005b00000000",
            INIT_36 => X"0000009500000000000000830000000000000081000000000000008700000000",
            INIT_37 => X"000000320000000000000000000000000000002f000000000000004000000000",
            INIT_38 => X"0000007500000000000000710000000000000073000000000000007600000000",
            INIT_39 => X"000000840000000000000096000000000000008f000000000000008100000000",
            INIT_3A => X"0000008c000000000000009d00000000000000a7000000000000008500000000",
            INIT_3B => X"0000007c0000000000000058000000000000001b000000000000003900000000",
            INIT_3C => X"0000008600000000000000790000000000000076000000000000007e00000000",
            INIT_3D => X"000000a7000000000000008e0000000000000083000000000000008800000000",
            INIT_3E => X"0000006e0000000000000095000000000000009a000000000000007400000000",
            INIT_3F => X"0000006700000000000000650000000000000060000000000000004800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000085000000000000008e0000000000000082000000000000007800000000",
            INIT_41 => X"0000009700000000000000a600000000000000a2000000000000008900000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000005000000000000003f000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE3;


    MEM_GOLD_LAYER0_INSTANCE4 : if BRAM_NAME = "gold_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000130000000000000036000000000000001d000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000001a00000000000000220000000000000022000000000000004800000000",
            INIT_05 => X"0000004300000000000000140000000000000001000000000000000000000000",
            INIT_06 => X"0000001e00000000000000000000000000000002000000000000000100000000",
            INIT_07 => X"00000021000000000000001c0000000000000021000000000000003700000000",
            INIT_08 => X"0000000400000000000000030000000000000007000000000000000b00000000",
            INIT_09 => X"000000030000000000000068000000000000003e000000000000000800000000",
            INIT_0A => X"000000100000000000000057000000000000007d000000000000003d00000000",
            INIT_0B => X"0000003b00000000000000470000000000000000000000000000000e00000000",
            INIT_0C => X"0000000000000000000000190000000000000022000000000000001f00000000",
            INIT_0D => X"000000000000000000000000000000000000002d000000000000001c00000000",
            INIT_0E => X"00000023000000000000002e0000000000000007000000000000000000000000",
            INIT_0F => X"00000000000000000000000d000000000000007f000000000000001300000000",
            INIT_10 => X"000000330000000000000029000000000000001e000000000000001900000000",
            INIT_11 => X"0000001300000000000000000000000000000000000000000000001c00000000",
            INIT_12 => X"000000090000000000000025000000000000001b000000000000004c00000000",
            INIT_13 => X"0000002100000000000000170000000000000009000000000000006000000000",
            INIT_14 => X"00000034000000000000003d000000000000001d000000000000003800000000",
            INIT_15 => X"0000003c000000000000003e000000000000001b000000000000003000000000",
            INIT_16 => X"0000002c00000000000000010000000000000000000000000000000000000000",
            INIT_17 => X"00000009000000000000001d0000000000000003000000000000000f00000000",
            INIT_18 => X"000000120000000000000041000000000000003c000000000000000000000000",
            INIT_19 => X"0000000700000000000000000000000000000021000000000000003600000000",
            INIT_1A => X"00000000000000000000000d0000000000000032000000000000002700000000",
            INIT_1B => X"0000001d00000000000000180000000000000000000000000000000000000000",
            INIT_1C => X"0000005300000000000000140000000000000038000000000000002400000000",
            INIT_1D => X"000000560000000000000038000000000000000b000000000000001500000000",
            INIT_1E => X"0000000900000000000000000000000000000000000000000000001500000000",
            INIT_1F => X"0000004400000000000000000000000000000024000000000000003400000000",
            INIT_20 => X"00000097000000000000009b0000000000000007000000000000003900000000",
            INIT_21 => X"0000000700000000000000040000000000000051000000000000007700000000",
            INIT_22 => X"0000004800000000000000600000000000000045000000000000001d00000000",
            INIT_23 => X"00000028000000000000000e000000000000002c000000000000003000000000",
            INIT_24 => X"000000000000000000000000000000000000008e000000000000004300000000",
            INIT_25 => X"00000034000000000000001e0000000000000004000000000000000100000000",
            INIT_26 => X"00000047000000000000004a000000000000003d000000000000003c00000000",
            INIT_27 => X"0000005100000000000000180000000000000046000000000000004000000000",
            INIT_28 => X"00000035000000000000003a0000000000000000000000000000002400000000",
            INIT_29 => X"0000005100000000000000460000000000000039000000000000003400000000",
            INIT_2A => X"0000006500000000000000420000000000000041000000000000005600000000",
            INIT_2B => X"0000000000000000000000330000000000000044000000000000004100000000",
            INIT_2C => X"0000003900000000000000420000000000000040000000000000002400000000",
            INIT_2D => X"0000003700000000000000400000000000000043000000000000003b00000000",
            INIT_2E => X"0000003d000000000000001d0000000000000062000000000000004000000000",
            INIT_2F => X"0000001e0000000000000000000000000000003a000000000000004400000000",
            INIT_30 => X"0000005100000000000000370000000000000023000000000000002300000000",
            INIT_31 => X"0000007d00000000000000450000000000000041000000000000005400000000",
            INIT_32 => X"0000007b000000000000007d0000000000000037000000000000006000000000",
            INIT_33 => X"0000007900000000000000830000000000000083000000000000008000000000",
            INIT_34 => X"0000006c00000000000000850000000000000091000000000000008900000000",
            INIT_35 => X"000000710000000000000064000000000000005a000000000000005700000000",
            INIT_36 => X"0000008700000000000000880000000000000082000000000000006c00000000",
            INIT_37 => X"0000008b00000000000000750000000000000082000000000000008800000000",
            INIT_38 => X"0000001f0000000000000023000000000000004d000000000000007200000000",
            INIT_39 => X"0000006900000000000000510000000000000036000000000000002900000000",
            INIT_3A => X"0000008a00000000000000860000000000000056000000000000005600000000",
            INIT_3B => X"0000002f00000000000000490000000000000076000000000000008b00000000",
            INIT_3C => X"00000010000000000000001d0000000000000012000000000000001400000000",
            INIT_3D => X"00000030000000000000004c0000000000000029000000000000001800000000",
            INIT_3E => X"0000007700000000000000860000000000000085000000000000003300000000",
            INIT_3F => X"0000000d0000000000000019000000000000003c000000000000004a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000009000000000000001f000000000000002c000000000000001800000000",
            INIT_41 => X"0000003a000000000000001e0000000000000032000000000000000900000000",
            INIT_42 => X"0000005800000000000000570000000000000060000000000000008200000000",
            INIT_43 => X"00000008000000000000000c000000000000001c000000000000003d00000000",
            INIT_44 => X"0000000900000000000000110000000000000029000000000000003700000000",
            INIT_45 => X"0000007e00000000000000290000000000000022000000000000002100000000",
            INIT_46 => X"0000003c0000000000000038000000000000001c000000000000006300000000",
            INIT_47 => X"000000410000000000000007000000000000001a000000000000002f00000000",
            INIT_48 => X"0000000b000000000000000c0000000000000010000000000000001c00000000",
            INIT_49 => X"000000690000000000000055000000000000002c000000000000002200000000",
            INIT_4A => X"0000003000000000000000410000000000000033000000000000002f00000000",
            INIT_4B => X"0000001b00000000000000320000000000000015000000000000002000000000",
            INIT_4C => X"000000290000000000000021000000000000000c000000000000000e00000000",
            INIT_4D => X"0000003600000000000000560000000000000037000000000000002400000000",
            INIT_4E => X"0000001d00000000000000210000000000000039000000000000003300000000",
            INIT_4F => X"00000006000000000000001e0000000000000028000000000000002e00000000",
            INIT_50 => X"000000210000000000000026000000000000003b000000000000002100000000",
            INIT_51 => X"0000002600000000000000430000000000000013000000000000002000000000",
            INIT_52 => X"00000053000000000000001a0000000000000020000000000000002b00000000",
            INIT_53 => X"0000002600000000000000080000000000000011000000000000002100000000",
            INIT_54 => X"0000001e00000000000000250000000000000024000000000000006100000000",
            INIT_55 => X"0000001c000000000000001f0000000000000028000000000000000b00000000",
            INIT_56 => X"0000000a00000000000000190000000000000031000000000000002e00000000",
            INIT_57 => X"00000072000000000000005b0000000000000009000000000000000000000000",
            INIT_58 => X"0000000c0000000000000025000000000000002e000000000000000900000000",
            INIT_59 => X"0000000e000000000000000b0000000000000025000000000000003000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000038000000000000003f000000000000001f000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000044000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"00000000000000000000000b0000000000000011000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_71 => X"0000000a000000000000001b0000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000002f0000000000000014000000000000000000000000",
            INIT_73 => X"0000000200000000000000560000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_75 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000001400000000000000000000000000000035000000000000000000000000",
            INIT_79 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_7E => X"0000000d000000000000006b000000000000001a000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE4;


    MEM_GOLD_LAYER0_INSTANCE5 : if BRAM_NAME = "gold_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_01 => X"0000002100000000000000060000000000000000000000000000000000000000",
            INIT_02 => X"000000030000000000000000000000000000003a000000000000000000000000",
            INIT_03 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000280000000000000012000000000000000f000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000021000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000017000000000000000800000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000003000000000000005c00000000",
            INIT_0B => X"0000002300000000000000240000000000000031000000000000001300000000",
            INIT_0C => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_0E => X"0000002100000000000000060000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000006000000000000001f00000000",
            INIT_10 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_13 => X"0000000300000000000000150000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000025000000000000008800000000",
            INIT_15 => X"00000041000000000000004d000000000000004a000000000000005800000000",
            INIT_16 => X"0000000600000000000000000000000000000001000000000000000e00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000001f000000000000001c0000000000000008000000000000006c00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000700000000000000000000000000000000000000000000000700000000",
            INIT_1C => X"000000000000000000000000000000000000002e000000000000007000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000030000000000000016000000000000000800000000",
            INIT_1F => X"0000001f00000000000000010000000000000000000000000000003f00000000",
            INIT_20 => X"0000001d0000000000000024000000000000001c000000000000005a00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000300000000000000000000000000000000000000000000000300000000",
            INIT_24 => X"0000000200000000000000050000000000000000000000000000000500000000",
            INIT_25 => X"000000000000000000000009000000000000000b000000000000000500000000",
            INIT_26 => X"00000000000000000000000b000000000000000a000000000000000000000000",
            INIT_27 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_28 => X"000000190000000000000014000000000000002e000000000000000000000000",
            INIT_29 => X"000000000000000000000015000000000000000a000000000000000000000000",
            INIT_2A => X"00000000000000000000002e0000000000000006000000000000000000000000",
            INIT_2B => X"0000000000000000000000010000000000000003000000000000000300000000",
            INIT_2C => X"0000000000000000000000000000000000000005000000000000003400000000",
            INIT_2D => X"0000000000000000000000300000000000000000000000000000001c00000000",
            INIT_2E => X"0000000b0000000000000000000000000000005c000000000000000000000000",
            INIT_2F => X"000000090000000000000000000000000000001f000000000000000000000000",
            INIT_30 => X"000000390000000000000000000000000000000e000000000000002400000000",
            INIT_31 => X"00000000000000000000002c0000000000000021000000000000001200000000",
            INIT_32 => X"0000000000000000000000410000000000000000000000000000003e00000000",
            INIT_33 => X"0000003a00000000000000380000000000000026000000000000000000000000",
            INIT_34 => X"0000004d00000000000000000000000000000000000000000000002400000000",
            INIT_35 => X"0000005b00000000000000000000000000000027000000000000000000000000",
            INIT_36 => X"0000000000000000000000500000000000000050000000000000000000000000",
            INIT_37 => X"00000046000000000000001b000000000000002a000000000000001200000000",
            INIT_38 => X"00000000000000000000004a000000000000005c000000000000000000000000",
            INIT_39 => X"0000002d000000000000004d000000000000001e000000000000001100000000",
            INIT_3A => X"0000000000000000000000000000000000000042000000000000000700000000",
            INIT_3B => X"00000000000000000000003b0000000000000030000000000000000100000000",
            INIT_3C => X"0000000000000000000000000000000000000038000000000000005100000000",
            INIT_3D => X"000000300000000000000000000000000000004d000000000000002600000000",
            INIT_3E => X"0000006700000000000000000000000000000000000000000000001100000000",
            INIT_3F => X"0000002c0000000000000000000000000000001e000000000000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000400000000000000030000000000000000000000000000003c00000000",
            INIT_41 => X"0000000000000000000000980000000000000000000000000000004100000000",
            INIT_42 => X"0000000f000000000000000b0000000000000000000000000000005100000000",
            INIT_43 => X"000000440000000000000000000000000000002b000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000003800000000000000000000000000000075000000000000000000000000",
            INIT_46 => X"0000003700000000000000030000000000000000000000000000002200000000",
            INIT_47 => X"0000000000000000000000000000000000000038000000000000001600000000",
            INIT_48 => X"0000000200000000000000000000000000000011000000000000000000000000",
            INIT_49 => X"00000033000000000000005f0000000000000000000000000000006100000000",
            INIT_4A => X"00000024000000000000004c000000000000000f000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000300000000000000000000000000000000000000000000000c00000000",
            INIT_4D => X"00000000000000000000003f00000000000000a3000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_4F => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000003000000000000000000000000000000000000000000000001f00000000",
            INIT_51 => X"0000000000000000000000050000000000000000000000000000007500000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000001f000000000000003e0000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000002000000000000000d000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000002b0000000000000028000000000000000000000000",
            INIT_58 => X"0000000000000000000000110000000000000000000000000000000c00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001200000000000000000000000000000000000000000000000f00000000",
            INIT_5B => X"0000006f00000000000000700000000000000065000000000000003100000000",
            INIT_5C => X"00000074000000000000006b000000000000006b000000000000006f00000000",
            INIT_5D => X"000000460000000000000051000000000000006b000000000000007900000000",
            INIT_5E => X"0000005f0000000000000064000000000000005d000000000000004f00000000",
            INIT_5F => X"0000007100000000000000730000000000000077000000000000006e00000000",
            INIT_60 => X"0000005e000000000000006a000000000000007b000000000000006c00000000",
            INIT_61 => X"000000280000000000000024000000000000002a000000000000003a00000000",
            INIT_62 => X"00000044000000000000005a0000000000000047000000000000003200000000",
            INIT_63 => X"0000006e0000000000000075000000000000006f000000000000004600000000",
            INIT_64 => X"0000001e00000000000000250000000000000041000000000000005400000000",
            INIT_65 => X"0000002000000000000000250000000000000025000000000000002600000000",
            INIT_66 => X"00000038000000000000002d0000000000000050000000000000002000000000",
            INIT_67 => X"0000003e0000000000000063000000000000006e000000000000006800000000",
            INIT_68 => X"0000001900000000000000190000000000000020000000000000003e00000000",
            INIT_69 => X"00000018000000000000001c0000000000000022000000000000003800000000",
            INIT_6A => X"00000064000000000000003e0000000000000023000000000000003700000000",
            INIT_6B => X"00000041000000000000004f0000000000000066000000000000004a00000000",
            INIT_6C => X"0000003a000000000000001d000000000000001b000000000000002e00000000",
            INIT_6D => X"0000001f000000000000001f0000000000000023000000000000002e00000000",
            INIT_6E => X"00000048000000000000006a0000000000000033000000000000000f00000000",
            INIT_6F => X"0000003600000000000000530000000000000041000000000000003300000000",
            INIT_70 => X"0000002300000000000000360000000000000021000000000000002b00000000",
            INIT_71 => X"0000001c0000000000000022000000000000001c000000000000001c00000000",
            INIT_72 => X"0000003500000000000000610000000000000046000000000000003000000000",
            INIT_73 => X"0000002b00000000000000350000000000000039000000000000004000000000",
            INIT_74 => X"0000001a0000000000000024000000000000002d000000000000002000000000",
            INIT_75 => X"000000350000000000000027000000000000002b000000000000001c00000000",
            INIT_76 => X"000000310000000000000026000000000000004a000000000000002600000000",
            INIT_77 => X"00000034000000000000002c0000000000000026000000000000003100000000",
            INIT_78 => X"0000002700000000000000150000000000000024000000000000003100000000",
            INIT_79 => X"0000001c00000000000000270000000000000028000000000000004800000000",
            INIT_7A => X"000000300000000000000021000000000000002f000000000000002b00000000",
            INIT_7B => X"0000001c000000000000003a0000000000000023000000000000002900000000",
            INIT_7C => X"0000005e000000000000003e0000000000000019000000000000001c00000000",
            INIT_7D => X"0000001a00000000000000280000000000000025000000000000002a00000000",
            INIT_7E => X"0000003a000000000000002a0000000000000023000000000000002600000000",
            INIT_7F => X"000000080000000000000014000000000000001f000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE5;


    MEM_GOLD_LAYER0_INSTANCE6 : if BRAM_NAME = "gold_layer0_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001500000000000000570000000000000053000000000000002200000000",
            INIT_01 => X"0000004800000000000000280000000000000026000000000000002800000000",
            INIT_02 => X"0000000f0000000000000014000000000000000f000000000000002000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_04 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000000c0000000000000037000000000000002400000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_19 => X"0000000100000000000000090000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_1C => X"0000000000000000000000030000000000000018000000000000000000000000",
            INIT_1D => X"0000002200000000000000250000000000000031000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_20 => X"00000014000000000000000a000000000000000b000000000000000600000000",
            INIT_21 => X"00000015000000000000001a0000000000000023000000000000003b00000000",
            INIT_22 => X"000000230000000000000021000000000000000c000000000000000000000000",
            INIT_23 => X"0000001800000000000000220000000000000015000000000000000000000000",
            INIT_24 => X"00000032000000000000000e000000000000000e000000000000002000000000",
            INIT_25 => X"0000000000000000000000140000000000000006000000000000002500000000",
            INIT_26 => X"00000000000000000000004b0000000000000037000000000000000000000000",
            INIT_27 => X"0000002f0000000000000044000000000000006b000000000000000500000000",
            INIT_28 => X"00000032000000000000004b0000000000000000000000000000001500000000",
            INIT_29 => X"000000000000000000000013000000000000001f000000000000001800000000",
            INIT_2A => X"00000000000000000000000e000000000000003d000000000000003800000000",
            INIT_2B => X"000000290000000000000047000000000000003f000000000000003100000000",
            INIT_2C => X"000000110000000000000031000000000000005a000000000000000e00000000",
            INIT_2D => X"00000042000000000000000b0000000000000023000000000000001900000000",
            INIT_2E => X"0000001b0000000000000000000000000000000a000000000000004d00000000",
            INIT_2F => X"0000001a0000000000000038000000000000003e000000000000005800000000",
            INIT_30 => X"0000002300000000000000140000000000000039000000000000004700000000",
            INIT_31 => X"0000006300000000000000530000000000000010000000000000002400000000",
            INIT_32 => X"0000003c000000000000000d0000000000000039000000000000001e00000000",
            INIT_33 => X"0000001000000000000000220000000000000019000000000000002100000000",
            INIT_34 => X"0000001600000000000000180000000000000015000000000000002200000000",
            INIT_35 => X"0000002d00000000000000650000000000000069000000000000000000000000",
            INIT_36 => X"000000360000000000000017000000000000001c000000000000004a00000000",
            INIT_37 => X"0000001400000000000000260000000000000013000000000000002d00000000",
            INIT_38 => X"000000000000000000000009000000000000000e000000000000000700000000",
            INIT_39 => X"0000007000000000000000330000000000000058000000000000006f00000000",
            INIT_3A => X"0000005f00000000000000510000000000000016000000000000003c00000000",
            INIT_3B => X"0000001c00000000000000100000000000000011000000000000002700000000",
            INIT_3C => X"00000074000000000000001d000000000000002b000000000000002200000000",
            INIT_3D => X"000000670000000000000082000000000000004c000000000000007a00000000",
            INIT_3E => X"0000003c000000000000004a000000000000004b000000000000005000000000",
            INIT_3F => X"00000052000000000000004a0000000000000043000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000066000000000000004d0000000000000050000000000000005300000000",
            INIT_41 => X"00000044000000000000004c0000000000000071000000000000007600000000",
            INIT_42 => X"0000004500000000000000400000000000000041000000000000004100000000",
            INIT_43 => X"0000005c00000000000000550000000000000050000000000000004e00000000",
            INIT_44 => X"00000073000000000000004b0000000000000058000000000000006000000000",
            INIT_45 => X"00000042000000000000004b0000000000000046000000000000007500000000",
            INIT_46 => X"00000055000000000000004d0000000000000047000000000000003f00000000",
            INIT_47 => X"000000650000000000000061000000000000005a000000000000005d00000000",
            INIT_48 => X"0000005a000000000000004f0000000000000056000000000000005600000000",
            INIT_49 => X"0000004b0000000000000053000000000000004d000000000000003f00000000",
            INIT_4A => X"00000054000000000000004c0000000000000050000000000000004c00000000",
            INIT_4B => X"0000003800000000000000490000000000000062000000000000006600000000",
            INIT_4C => X"000000380000000000000039000000000000003a000000000000003800000000",
            INIT_4D => X"0000003b00000000000000490000000000000042000000000000003500000000",
            INIT_4E => X"0000002b00000000000000270000000000000020000000000000002600000000",
            INIT_4F => X"00000043000000000000003a000000000000002c000000000000003100000000",
            INIT_50 => X"000000170000000000000038000000000000003c000000000000003d00000000",
            INIT_51 => X"00000000000000000000001e000000000000002d000000000000003100000000",
            INIT_52 => X"0000002100000000000000080000000000000000000000000000000000000000",
            INIT_53 => X"0000004100000000000000320000000000000011000000000000002800000000",
            INIT_54 => X"0000001000000000000000230000000000000040000000000000004200000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000003f000000000000003b0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000013000000000000002400000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_5B => X"00000000000000000000001e0000000000000027000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000026000000000000002500000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE6;


    MEM_GOLD_LAYER0_INSTANCE7 : if BRAM_NAME = "gold_layer0_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE7;


    MEM_GOLD_LAYER1_INSTANCE0 : if BRAM_NAME = "gold_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000001a00000000000000000000000000000001000000000000000000000000",
            INIT_02 => X"00000000000000000000001e0000000000000021000000000000000000000000",
            INIT_03 => X"0000000000000000000000940000000000000004000000000000004b00000000",
            INIT_04 => X"000000740000000000000000000000000000004f000000000000003800000000",
            INIT_05 => X"00000038000000000000003d00000000000000c0000000000000000000000000",
            INIT_06 => X"0000000000000000000000580000000000000034000000000000007800000000",
            INIT_07 => X"000000350000000000000094000000000000004400000000000000a000000000",
            INIT_08 => X"000000bc000000000000002d0000000000000036000000000000005500000000",
            INIT_09 => X"00000000000000000000008600000000000000a0000000000000002d00000000",
            INIT_0A => X"000000fa000000000000002d0000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_0C => X"00000000000000000000003d0000000000000000000000000000001500000000",
            INIT_0D => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000b20000000000000000000000000000000000000000",
            INIT_15 => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000006800000000",
            INIT_17 => X"0000000a0000000000000008000000000000003e000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_1A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000009000000000000000b0000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_20 => X"0000000b00000000000000000000000000000020000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"000000400000000000000034000000000000000c000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000007a00000000000000000000000000000000000000000000006000000000",
            INIT_26 => X"0000009a0000000000000011000000000000001c000000000000001900000000",
            INIT_27 => X"0000000000000000000000490000000000000000000000000000005c00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000002200000000000000000000000000000033000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000000e000000000000003b000000000000000500000000",
            INIT_2D => X"000000000000000000000000000000000000006d000000000000002500000000",
            INIT_2E => X"0000012100000000000000cb0000000000000000000000000000000000000000",
            INIT_2F => X"0000003f0000000000000000000000000000002900000000000000f200000000",
            INIT_30 => X"0000009e00000000000000ee00000000000000fd00000000000000b700000000",
            INIT_31 => X"000000000000000000000007000000000000000e000000000000000000000000",
            INIT_32 => X"000000360000000000000000000000000000001a000000000000004400000000",
            INIT_33 => X"0000007000000000000000000000000000000062000000000000005600000000",
            INIT_34 => X"0000001800000000000000000000000000000000000000000000000400000000",
            INIT_35 => X"00000000000000000000009e0000000000000003000000000000006a00000000",
            INIT_36 => X"0000006f000000000000003b0000000000000000000000000000001e00000000",
            INIT_37 => X"000000330000000000000000000000000000006b000000000000000000000000",
            INIT_38 => X"00000029000000000000003b0000000000000079000000000000002300000000",
            INIT_39 => X"00000002000000000000003c0000000000000005000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000007500000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000005700000000000000100000000000000044000000000000000000000000",
            INIT_3E => X"0000004400000000000000360000000000000092000000000000005500000000",
            INIT_3F => X"0000002c000000000000009000000000000000b300000000000000e500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005e00000000000000570000000000000000000000000000010900000000",
            INIT_41 => X"000002090000000000000000000000000000006900000000000000e000000000",
            INIT_42 => X"000000f3000000000000003f000000000000001b000000000000002000000000",
            INIT_43 => X"0000000000000000000000fc000000000000000000000000000000fa00000000",
            INIT_44 => X"000000b40000000000000187000000000000002e000000000000002e00000000",
            INIT_45 => X"0000008500000000000000300000000000000047000000000000004a00000000",
            INIT_46 => X"000000000000000000000004000000000000016c00000000000000b800000000",
            INIT_47 => X"000000a700000000000000000000000000000005000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000005200000000",
            INIT_49 => X"0000002300000000000000300000000000000034000000000000000700000000",
            INIT_4A => X"00000051000000000000007e000000000000009f000000000000001700000000",
            INIT_4B => X"00000042000000000000006e0000000000000063000000000000007200000000",
            INIT_4C => X"0000006a00000000000000000000000000000034000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000115000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_4F => X"0000003200000000000000000000000000000054000000000000002800000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000008500000000000000990000000000000000000000000000004500000000",
            INIT_52 => X"000000ad00000000000000460000000000000075000000000000007a00000000",
            INIT_53 => X"0000000000000000000000040000000000000000000000000000004900000000",
            INIT_54 => X"00000000000000000000000000000000000000b3000000000000004900000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_5E => X"0000009800000000000000ce0000000000000000000000000000000600000000",
            INIT_5F => X"000000d000000000000000a600000000000000a600000000000000d200000000",
            INIT_60 => X"0000011c00000000000000dd000000000000012b00000000000000bb00000000",
            INIT_61 => X"000001530000000000000123000000000000010700000000000000e400000000",
            INIT_62 => X"0000007a000000000000008500000000000000e300000000000000bd00000000",
            INIT_63 => X"00000000000000000000007f0000000000000038000000000000007700000000",
            INIT_64 => X"0000000300000000000000000000000000000016000000000000009200000000",
            INIT_65 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_67 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000005a00000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"00000000000000000000005a000000000000000c000000000000000000000000",
            INIT_6B => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_6D => X"00000014000000000000001e0000000000000013000000000000000000000000",
            INIT_6E => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000002300000000000000590000000000000085000000000000003500000000",
            INIT_70 => X"0000007f0000000000000075000000000000006600000000000000a300000000",
            INIT_71 => X"000000d00000000000000080000000000000009c00000000000000bf00000000",
            INIT_72 => X"00000121000000000000010c00000000000000f500000000000000d500000000",
            INIT_73 => X"000000b400000000000000f6000000000000008d00000000000000eb00000000",
            INIT_74 => X"000000d600000000000000da00000000000000de000000000000005500000000",
            INIT_75 => X"000000bc00000000000001a900000000000000e5000000000000004b00000000",
            INIT_76 => X"0000004000000000000000b000000000000000a0000000000000008300000000",
            INIT_77 => X"0000006d0000000000000186000000000000014000000000000000ba00000000",
            INIT_78 => X"0000006100000000000000450000000000000040000000000000007f00000000",
            INIT_79 => X"000000090000000000000029000000000000005e000000000000007e00000000",
            INIT_7A => X"0000000000000000000000000000000000000022000000000000002a00000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000250000000000000029000000000000000a00000000",
            INIT_7E => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000004e00000000000000000000000000000023000000000000009200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE0;


    MEM_GOLD_LAYER1_INSTANCE1 : if BRAM_NAME = "gold_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000065000000000000001a0000000000000027000000000000000000000000",
            INIT_01 => X"0000006a00000000000000860000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_03 => X"0000000000000000000000840000000000000000000000000000000000000000",
            INIT_04 => X"0000000700000000000000000000000000000000000000000000001900000000",
            INIT_05 => X"000000110000000000000000000000000000002b000000000000004500000000",
            INIT_06 => X"000000420000000000000044000000000000001b000000000000002200000000",
            INIT_07 => X"0000010900000000000000ac0000000000000048000000000000000000000000",
            INIT_08 => X"000000850000000000000095000000000000007200000000000000ae00000000",
            INIT_09 => X"000000000000000000000000000000000000004b00000000000000bd00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_0B => X"0000002000000000000000000000000000000000000000000000000400000000",
            INIT_0C => X"0000000000000000000000000000000000000064000000000000001e00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000044000000000000002a000000000000007f000000000000007000000000",
            INIT_0F => X"00000000000000000000005d000000000000004b00000000000000c900000000",
            INIT_10 => X"00000031000000000000007e0000000000000067000000000000000000000000",
            INIT_11 => X"0000005c000000000000003d000000000000003e000000000000007a00000000",
            INIT_12 => X"000000200000000000000000000000000000000c000000000000001200000000",
            INIT_13 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_14 => X"000000000000000000000000000000000000001c000000000000001900000000",
            INIT_15 => X"0000000000000000000000000000000000000065000000000000000800000000",
            INIT_16 => X"0000000000000000000000000000000000000013000000000000001600000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"000000000000000000000000000000000000008a000000000000000000000000",
            INIT_1C => X"0000009b00000000000000900000000000000000000000000000000000000000",
            INIT_1D => X"00000000000000000000002e000000000000008e000000000000007e00000000",
            INIT_1E => X"00000040000000000000004b000000000000002f000000000000000000000000",
            INIT_1F => X"0000000f000000000000001a0000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000200000000000000000000000000000001100000000",
            INIT_21 => X"00000052000000000000002d0000000000000000000000000000000f00000000",
            INIT_22 => X"00000082000000000000005d000000000000007e000000000000000000000000",
            INIT_23 => X"0000001200000000000000d50000000000000078000000000000001000000000",
            INIT_24 => X"0000006300000000000000c9000000000000005900000000000000a300000000",
            INIT_25 => X"0000007700000000000000210000000000000091000000000000001e00000000",
            INIT_26 => X"0000006f000000000000006c000000000000010f000000000000002300000000",
            INIT_27 => X"00000014000000000000002b000000000000004a000000000000007c00000000",
            INIT_28 => X"00000047000000000000004f0000000000000075000000000000008c00000000",
            INIT_29 => X"0000004800000000000000080000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000000000000000000000c100000000",
            INIT_2B => X"000000000000000000000000000000000000001f000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000007c00000000000000ad0000000000000000000000000000000000000000",
            INIT_39 => X"00000020000000000000005c0000000000000062000000000000004b00000000",
            INIT_3A => X"00000032000000000000001a000000000000000f000000000000004800000000",
            INIT_3B => X"0000002a000000000000007e0000000000000046000000000000004600000000",
            INIT_3C => X"0000000000000000000000680000000000000055000000000000002e00000000",
            INIT_3D => X"0000005300000000000000180000000000000029000000000000003500000000",
            INIT_3E => X"0000002d0000000000000000000000000000005e000000000000003900000000",
            INIT_3F => X"000000a2000000000000001c0000000000000060000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c00000000000000bd0000000000000066000000000000008100000000",
            INIT_41 => X"0000000000000000000000200000000000000077000000000000012400000000",
            INIT_42 => X"0000003600000000000000cd0000000000000040000000000000000000000000",
            INIT_43 => X"0000003a00000000000000170000000000000002000000000000001300000000",
            INIT_44 => X"00000088000000000000008600000000000000bf00000000000000aa00000000",
            INIT_45 => X"000000970000000000000093000000000000006d000000000000004f00000000",
            INIT_46 => X"000000480000000000000097000000000000008b00000000000000ad00000000",
            INIT_47 => X"0000006b0000000000000072000000000000006c000000000000007800000000",
            INIT_48 => X"0000007f0000000000000039000000000000008a000000000000002d00000000",
            INIT_49 => X"0000002e00000000000000ae0000000000000027000000000000005300000000",
            INIT_4A => X"0000008500000000000000670000000000000053000000000000007600000000",
            INIT_4B => X"00000000000000000000003d0000000000000028000000000000000000000000",
            INIT_4C => X"00000000000000000000001d0000000000000000000000000000003600000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000c00000000000000510000000000000014000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000200000000000000000000000000000000000000000000004900000000",
            INIT_53 => X"0000002800000000000000180000000000000013000000000000004800000000",
            INIT_54 => X"000000df00000000000000070000000000000000000000000000003200000000",
            INIT_55 => X"0000000000000000000000000000000000000003000000000000002900000000",
            INIT_56 => X"00000000000000000000003a0000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000620000000000000000000000000000004900000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"000000000000000000000000000000000000003a000000000000000000000000",
            INIT_5F => X"0000004500000000000000040000000000000001000000000000005000000000",
            INIT_60 => X"0000008e00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"00000053000000000000007b000000000000002d000000000000008300000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000006100000000",
            INIT_63 => X"000000fb00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"00000021000000000000000f0000000000000031000000000000002f00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000007100000000000000790000000000000071000000000000000000000000",
            INIT_67 => X"0000002f00000000000000000000000000000000000000000000003d00000000",
            INIT_68 => X"0000000000000000000000660000000000000027000000000000003900000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"000000a500000000000000bb00000000000000a300000000000000b200000000",
            INIT_76 => X"00000050000000000000009e0000000000000044000000000000008800000000",
            INIT_77 => X"00000033000000000000003c000000000000008900000000000000bd00000000",
            INIT_78 => X"0000009700000000000000000000000000000021000000000000000000000000",
            INIT_79 => X"0000000000000000000000320000000000000000000000000000005400000000",
            INIT_7A => X"0000005000000000000000620000000000000000000000000000000000000000",
            INIT_7B => X"0000001300000000000000000000000000000011000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE1;


    MEM_GOLD_LAYER1_INSTANCE2 : if BRAM_NAME = "gold_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000007000000000000001c0000000000000031000000000000000000000000",
            INIT_02 => X"000000250000000000000000000000000000000b000000000000003e00000000",
            INIT_03 => X"00000000000000000000002d000000000000000e000000000000002e00000000",
            INIT_04 => X"000000000000000000000031000000000000001b000000000000005b00000000",
            INIT_05 => X"000000570000000000000000000000000000003900000000000000d300000000",
            INIT_06 => X"0000000800000000000000000000000000000000000000000000000500000000",
            INIT_07 => X"00000031000000000000009e000000000000004d00000000000000af00000000",
            INIT_08 => X"00000022000000000000001d000000000000001d000000000000001700000000",
            INIT_09 => X"0000000000000000000000430000000000000083000000000000000000000000",
            INIT_0A => X"00000071000000000000009d0000000000000070000000000000008b00000000",
            INIT_0B => X"0000006200000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000000000000000000000000000d000000000000013000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_11 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000034000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_19 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000034000000000000008600000000",
            INIT_1B => X"0000000600000000000000000000000000000000000000000000003100000000",
            INIT_1C => X"0000006a00000000000000000000000000000052000000000000004500000000",
            INIT_1D => X"0000000000000000000000000000000000000061000000000000000000000000",
            INIT_1E => X"000000210000000000000055000000000000000000000000000000a500000000",
            INIT_1F => X"000000000000000000000000000000000000000000000000000000d500000000",
            INIT_20 => X"0000007b00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000370000000000000023000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000c900000000000000b30000000000000000000000000000000000000000",
            INIT_24 => X"000000720000000000000000000000000000000000000000000000d700000000",
            INIT_25 => X"000000d200000000000000ad00000000000000d900000000000000be00000000",
            INIT_26 => X"00000130000000000000012a0000000000000153000000000000016b00000000",
            INIT_27 => X"0000005e00000000000000eb000000000000004a000000000000006400000000",
            INIT_28 => X"00000000000000000000003f000000000000005a000000000000010b00000000",
            INIT_29 => X"0000010b00000000000000480000000000000059000000000000004b00000000",
            INIT_2A => X"0000005c00000000000000000000000000000018000000000000004300000000",
            INIT_2B => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_2C => X"0000003000000000000000720000000000000016000000000000005400000000",
            INIT_2D => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_2E => X"00000007000000000000001e0000000000000017000000000000005400000000",
            INIT_2F => X"00000008000000000000003300000000000000b7000000000000000000000000",
            INIT_30 => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000028000000000000000c000000000000001c000000000000004100000000",
            INIT_32 => X"0000007a0000000000000046000000000000005d000000000000000200000000",
            INIT_33 => X"00000067000000000000005f000000000000002e000000000000004400000000",
            INIT_34 => X"00000049000000000000008c000000000000006f00000000000000cb00000000",
            INIT_35 => X"000000ab00000000000000680000000000000039000000000000005c00000000",
            INIT_36 => X"000000a7000000000000003900000000000000b200000000000000a100000000",
            INIT_37 => X"000000a700000000000000730000000000000025000000000000004600000000",
            INIT_38 => X"0000001c0000000000000090000000000000000000000000000000c000000000",
            INIT_39 => X"000000ac000000000000007f000000000000003a000000000000003700000000",
            INIT_3A => X"000000ac00000000000000320000000000000076000000000000009e00000000",
            INIT_3B => X"0000002b0000000000000078000000000000011d00000000000000a700000000",
            INIT_3C => X"0000007b00000000000000220000000000000029000000000000000000000000",
            INIT_3D => X"000000060000000000000000000000000000000000000000000000b600000000",
            INIT_3E => X"000000000000000000000000000000000000002f000000000000000700000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000006c00000000000000130000000000000013000000000000000000000000",
            INIT_47 => X"0000007000000000000000000000000000000058000000000000001400000000",
            INIT_48 => X"000001bf00000000000001ba000000000000015b00000000000000df00000000",
            INIT_49 => X"0000019f0000000000000136000000000000007f000000000000017300000000",
            INIT_4A => X"0000000000000000000001da00000000000001e000000000000001c400000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000910000000000000000000000000000005b000000000000000000000000",
            INIT_4F => X"0000002100000000000000000000000000000000000000000000004100000000",
            INIT_50 => X"000000000000000000000000000000000000000000000000000000b300000000",
            INIT_51 => X"000000ef000000000000000c0000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000930000000000000000000000000000007200000000",
            INIT_53 => X"000000000000000000000076000000000000000f000000000000000000000000",
            INIT_54 => X"00000090000000000000007d0000000000000024000000000000000000000000",
            INIT_55 => X"0000005a000000000000008b000000000000000000000000000000af00000000",
            INIT_56 => X"000000ab000000000000008b000000000000009a000000000000008e00000000",
            INIT_57 => X"0000002100000000000000290000000000000001000000000000000f00000000",
            INIT_58 => X"0000001b00000000000000290000000000000032000000000000005000000000",
            INIT_59 => X"0000005d00000000000000600000000000000048000000000000002200000000",
            INIT_5A => X"0000003c00000000000000000000000000000054000000000000003c00000000",
            INIT_5B => X"00000039000000000000004d0000000000000031000000000000003500000000",
            INIT_5C => X"0000004400000000000000500000000000000000000000000000005400000000",
            INIT_5D => X"0000004f0000000000000037000000000000003b000000000000001600000000",
            INIT_5E => X"0000001d000000000000003a000000000000001a000000000000000000000000",
            INIT_5F => X"000000000000000000000034000000000000003c000000000000005000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000002900000000000000000000000000000000000000000000000900000000",
            INIT_67 => X"0000000a00000000000000000000000000000056000000000000002100000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_6C => X"00000000000000000000005c00000000000000ea000000000000000000000000",
            INIT_6D => X"000000000000000000000052000000000000008d000000000000000000000000",
            INIT_6E => X"00000047000000000000001b0000000000000000000000000000000000000000",
            INIT_6F => X"000000a200000000000000b10000000000000049000000000000003e00000000",
            INIT_70 => X"000000d800000000000000c6000000000000011f00000000000000d200000000",
            INIT_71 => X"0000010100000000000000c500000000000000b900000000000000d100000000",
            INIT_72 => X"000000550000000000000079000000000000000800000000000000ce00000000",
            INIT_73 => X"000000c5000000000000003f0000000000000094000000000000009000000000",
            INIT_74 => X"000000a7000000000000002e00000000000000ac000000000000000000000000",
            INIT_75 => X"0000000000000000000000b5000000000000004300000000000000b700000000",
            INIT_76 => X"0000003e000000000000003f0000000000000009000000000000005400000000",
            INIT_77 => X"0000002800000000000000910000000000000038000000000000008d00000000",
            INIT_78 => X"0000004600000000000000000000000000000000000000000000002600000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000004200000000000000020000000000000002000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000032000000000000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE2;


    MEM_GOLD_LAYER1_INSTANCE3 : if BRAM_NAME = "gold_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002600000000000000510000000000000000000000000000000800000000",
            INIT_01 => X"0000009700000000000000000000000000000012000000000000004e00000000",
            INIT_02 => X"0000003b0000000000000013000000000000002f000000000000000000000000",
            INIT_03 => X"0000009000000000000000000000000000000007000000000000000000000000",
            INIT_04 => X"00000000000000000000003a0000000000000000000000000000006600000000",
            INIT_05 => X"0000001c000000000000002f000000000000008c00000000000000ad00000000",
            INIT_06 => X"00000069000000000000005b000000000000003b000000000000002800000000",
            INIT_07 => X"0000002700000000000000750000000000000046000000000000006600000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE3;


    MEM_GOLD_LAYER2_INSTANCE0 : if BRAM_NAME = "gold_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000001240000000000000087000000000000003a000000000000004c00000000",
            INIT_02 => X"00000000000000000000000000000000000000c1000000000000000000000000",
            INIT_03 => X"000000ab00000000000000880000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000000000000000001c9000000000000022b00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000b400000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000000000000000000000000000000000000f1000000000000011500000000",
            INIT_08 => X"000000b6000000000000000000000000000000de000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000005e000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000035b00000000000002250000000000000000000000000000000000000000",
            INIT_0E => X"0000019100000000000001a800000000000003f7000000000000024a00000000",
            INIT_0F => X"000000a800000000000001e700000000000001ae00000000000002de00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000670000000000000121000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"00000000000000000000006b0000000000000000000000000000000000000000",
            INIT_17 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000023300000000000000000000000000000000000000000000009700000000",
            INIT_19 => X"0000018c000000000000011700000000000001ac00000000000001e100000000",
            INIT_1A => X"000002d9000000000000025100000000000002fc00000000000000b200000000",
            INIT_1B => X"0000000000000000000001300000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000001330000000000000000000000000000000000000000",
            INIT_1D => X"000000d800000000000000540000000000000148000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000013b00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"000000000000000000000000000000000000009d000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000004c000000000000010b000000000000000000000000",
            INIT_2D => X"000000000000000000000101000000000000002d000000000000008f00000000",
            INIT_2E => X"000000000000000000000000000000000000012f000000000000001d00000000",
            INIT_2F => X"000000b900000000000000260000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000440000000000000040000000000000000000000000",
            INIT_32 => X"0000000800000000000000ac0000000000000000000000000000003d00000000",
            INIT_33 => X"00000000000000000000001f0000000000000018000000000000000d00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000be00000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000016600000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000d9000000000000001d0000000000000000000000000000000000000000",
            INIT_3B => X"0000013f00000000000001310000000000000000000000000000020700000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"000000000000000000000000000000000000000000000000000000a400000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000000000000000000000000000000000000c800000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000a000000000000000000000000000000cf000000000000009f00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000b00000000000000800000000000000082000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_4E => X"00000000000000000000029c0000000000000177000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_51 => X"00000024000000000000019600000000000001a5000000000000014c00000000",
            INIT_52 => X"00000000000000000000000000000000000000bc000000000000018700000000",
            INIT_53 => X"00000181000000000000024d0000000000000324000000000000000000000000",
            INIT_54 => X"0000020600000000000002e000000000000002b900000000000002c800000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000009d00000000000001800000000000000000000000000000000000000000",
            INIT_5C => X"0000005a00000000000000000000000000000000000000000000011b00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000001e00000000000000530000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000a40000000000000000000000000000005d00000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000000000000000000124000000000000013b000000000000005100000000",
            INIT_6A => X"000000f2000000000000004f0000000000000000000000000000000000000000",
            INIT_6B => X"0000003d00000000000000510000000000000000000000000000011400000000",
            INIT_6C => X"0000017f000000000000007c0000000000000088000000000000000f00000000",
            INIT_6D => X"0000005e00000000000001650000000000000061000000000000014000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000a500000000000000220000000000000000000000000000000000000000",
            INIT_71 => X"000000e900000000000001330000000000000232000000000000010c00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000011d00000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000bb00000000000001b40000000000000000000000000000008f00000000",
            INIT_77 => X"000000ba0000000000000000000000000000000000000000000000dd00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000012e00000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000020900000000000001ba000000000000015b000000000000018200000000",
            INIT_7D => X"0000001300000000000000a60000000000000012000000000000016800000000",
            INIT_7E => X"000000b700000000000001c000000000000000ee00000000000000ea00000000",
            INIT_7F => X"00000000000000000000001e0000000000000000000000000000013d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE0;


    MEM_GOLD_LAYER2_INSTANCE1 : if BRAM_NAME = "gold_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000d5000000000000011d0000000000000000000000000000000000000000",
            INIT_03 => X"000001a1000000000000018300000000000000f3000000000000008f00000000",
            INIT_04 => X"0000000000000000000000000000000000000050000000000000010000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000011700000000000000000000000000000034000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000ac00000000000000000000000000000000000000000000016700000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001f0000000000000000000000000000000000000000000000a400000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE1;


    MEM_GOLD_LAYER3_INSTANCE0 : if BRAM_NAME = "gold_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000001150000000000000000000000000000022b000000000000012400000000",
            INIT_01 => X"0000012100000000000003f7000000000000005e000000000000000000000000",
            INIT_02 => X"000002fc00000000000000970000000000000000000000000000000000000000",
            INIT_03 => X"00000000000000000000013b0000000000000148000000000000013300000000",
            INIT_04 => X"0000010b0000000000000000000000000000009d000000000000004f00000000",
            INIT_05 => X"0000000000000000000000ac00000000000000b9000000000000012f00000000",
            INIT_06 => X"000000a400000000000002070000000000000000000000000000016600000000",
            INIT_07 => X"000000cf0000000000000035000000000000000000000000000000c800000000",
            INIT_08 => X"00000041000000000000029c0000000000000082000000000000000000000000",
            INIT_09 => X"000000000000000000000000000000000000032400000000000001a500000000",
            INIT_0A => X"000000a40000000000000053000000000000005a000000000000018000000000",
            INIT_0B => X"00000114000000000000013b0000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000000000232000000000000000d000000000000017f00000000",
            INIT_0D => X"00000209000000000000000000000000000000ba00000000000001b400000000",
            INIT_0E => X"0000001000000000000001a1000000000000000000000000000001c000000000",
            INIT_0F => X"000000a400000000000000000000000000000167000000000000011700000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER3_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "sampleifmap_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "sampleifmap_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "sampleifmap_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "sampleifmap_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "sampleifmap_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "sampleifmap_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "sampleifmap_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e600000000000000e700000000000000e800000000000000e900000000",
            INIT_05 => X"000000e900000000000000e800000000000000e800000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e800000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ec00000000000000ec00000000000000ed00000000",
            INIT_0D => X"000000ec00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ea00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_15 => X"000000ea00000000000000e700000000000000e700000000000000e300000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000df00000000000000e400000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000cf00000000000000d100000000000000ba00000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000ec00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000cb00000000000000db00000000000000e900000000000000ec00000000",
            INIT_25 => X"000000e600000000000000d600000000000000c300000000000000a300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_28 => X"000000ec00000000000000ec00000000000000ec00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_2A => X"000000ed00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e500000000000000eb00000000000000e800000000000000ea00000000",
            INIT_2C => X"000000ae00000000000000b900000000000000c200000000000000d000000000",
            INIT_2D => X"000000e200000000000000cf00000000000000b800000000000000a500000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e700000000000000e800000000000000e400000000000000e400000000",
            INIT_31 => X"000000ec00000000000000ed00000000000000ed00000000000000ea00000000",
            INIT_32 => X"000000ef00000000000000ef00000000000000ed00000000000000ed00000000",
            INIT_33 => X"000000dd00000000000000e900000000000000e000000000000000e100000000",
            INIT_34 => X"0000009a000000000000009f00000000000000a100000000000000b700000000",
            INIT_35 => X"000000c6000000000000009c000000000000008f000000000000009000000000",
            INIT_36 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_37 => X"000000ef00000000000000ed00000000000000ec00000000000000eb00000000",
            INIT_38 => X"000000e300000000000000e600000000000000e000000000000000d400000000",
            INIT_39 => X"000000ee00000000000000ed00000000000000ea00000000000000e500000000",
            INIT_3A => X"000000f000000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_3B => X"000000d600000000000000e900000000000000db00000000000000c900000000",
            INIT_3C => X"000000ad00000000000000b800000000000000b900000000000000c100000000",
            INIT_3D => X"000000ba00000000000000a2000000000000009f00000000000000a500000000",
            INIT_3E => X"000000e900000000000000e900000000000000ea00000000000000e500000000",
            INIT_3F => X"000000ee00000000000000ed00000000000000ec00000000000000ea00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000e100000000000000e100000000000000dd00000000000000d800000000",
            INIT_41 => X"000000ee00000000000000ec00000000000000e700000000000000e300000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_43 => X"000000e600000000000000e900000000000000dc00000000000000c500000000",
            INIT_44 => X"000000d000000000000000db00000000000000d100000000000000d100000000",
            INIT_45 => X"000000da00000000000000d900000000000000d200000000000000d100000000",
            INIT_46 => X"000000e600000000000000e400000000000000e400000000000000e100000000",
            INIT_47 => X"000000ee00000000000000ed00000000000000eb00000000000000e600000000",
            INIT_48 => X"00000088000000000000007c0000000000000077000000000000007600000000",
            INIT_49 => X"000000ed00000000000000eb00000000000000e100000000000000ac00000000",
            INIT_4A => X"000000e900000000000000eb00000000000000eb00000000000000ec00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000e100000000000000e700000000000000e300000000000000e400000000",
            INIT_4D => X"000000b900000000000000c900000000000000d900000000000000e100000000",
            INIT_4E => X"000000ba00000000000000a700000000000000a700000000000000ac00000000",
            INIT_4F => X"000000ee00000000000000ec00000000000000eb00000000000000df00000000",
            INIT_50 => X"0000006f000000000000006c0000000000000067000000000000006d00000000",
            INIT_51 => X"000000e500000000000000e300000000000000de000000000000009200000000",
            INIT_52 => X"000000e600000000000000e700000000000000ea00000000000000ec00000000",
            INIT_53 => X"000000e600000000000000e800000000000000e700000000000000e500000000",
            INIT_54 => X"000000df00000000000000e500000000000000e700000000000000e700000000",
            INIT_55 => X"00000089000000000000009200000000000000a400000000000000bf00000000",
            INIT_56 => X"0000009500000000000000790000000000000080000000000000008600000000",
            INIT_57 => X"000000ed00000000000000eb00000000000000ea00000000000000d800000000",
            INIT_58 => X"000000c800000000000000c700000000000000bc00000000000000c300000000",
            INIT_59 => X"000000d300000000000000d500000000000000df00000000000000d100000000",
            INIT_5A => X"000000d200000000000000db00000000000000dc00000000000000d800000000",
            INIT_5B => X"000000dc00000000000000d800000000000000d300000000000000d100000000",
            INIT_5C => X"000000da00000000000000e100000000000000e200000000000000e100000000",
            INIT_5D => X"000000b200000000000000b500000000000000af00000000000000b700000000",
            INIT_5E => X"000000b9000000000000008e00000000000000aa00000000000000ba00000000",
            INIT_5F => X"000000ec00000000000000ea00000000000000e700000000000000db00000000",
            INIT_60 => X"000000d600000000000000ca00000000000000bf00000000000000c100000000",
            INIT_61 => X"000000ab00000000000000cb00000000000000d600000000000000df00000000",
            INIT_62 => X"0000006200000000000000ae00000000000000cf00000000000000b100000000",
            INIT_63 => X"0000007a000000000000006f0000000000000065000000000000005d00000000",
            INIT_64 => X"000000df00000000000000ca0000000000000099000000000000008900000000",
            INIT_65 => X"000000d900000000000000df00000000000000dc00000000000000da00000000",
            INIT_66 => X"000000de00000000000000c400000000000000d400000000000000dd00000000",
            INIT_67 => X"000000eb00000000000000e800000000000000dd00000000000000db00000000",
            INIT_68 => X"0000007d0000000000000071000000000000006f000000000000007100000000",
            INIT_69 => X"000000be00000000000000bf00000000000000aa000000000000008a00000000",
            INIT_6A => X"00000036000000000000009e00000000000000d800000000000000d000000000",
            INIT_6B => X"0000004200000000000000350000000000000031000000000000002d00000000",
            INIT_6C => X"000000ea00000000000000dd000000000000009f000000000000006600000000",
            INIT_6D => X"000000cf00000000000000df00000000000000e300000000000000e900000000",
            INIT_6E => X"000000c700000000000000d400000000000000d300000000000000ca00000000",
            INIT_6F => X"000000dd00000000000000d300000000000000bc00000000000000b300000000",
            INIT_70 => X"00000044000000000000003f0000000000000045000000000000003d00000000",
            INIT_71 => X"000000c30000000000000097000000000000008b000000000000007b00000000",
            INIT_72 => X"0000006700000000000000a300000000000000ce00000000000000d600000000",
            INIT_73 => X"000000b5000000000000008a0000000000000065000000000000005f00000000",
            INIT_74 => X"000000cd00000000000000db00000000000000dd00000000000000cf00000000",
            INIT_75 => X"000000830000000000000093000000000000009e00000000000000b700000000",
            INIT_76 => X"0000008500000000000000880000000000000082000000000000007d00000000",
            INIT_77 => X"000000c500000000000000b6000000000000008a000000000000008000000000",
            INIT_78 => X"0000007f0000000000000055000000000000003a000000000000002800000000",
            INIT_79 => X"000000a300000000000000770000000000000060000000000000008400000000",
            INIT_7A => X"000000b500000000000000b600000000000000b800000000000000ad00000000",
            INIT_7B => X"000000c800000000000000da00000000000000c600000000000000b700000000",
            INIT_7C => X"000000840000000000000091000000000000009f00000000000000ae00000000",
            INIT_7D => X"00000063000000000000005e0000000000000062000000000000007400000000",
            INIT_7E => X"0000008a000000000000007a000000000000006b000000000000006900000000",
            INIT_7F => X"000000b900000000000000bc000000000000009d000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "sampleifmap_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ce0000000000000086000000000000001a000000000000000d00000000",
            INIT_01 => X"000000ac000000000000008d0000000000000076000000000000008a00000000",
            INIT_02 => X"000000e400000000000000dc00000000000000cf00000000000000b500000000",
            INIT_03 => X"000000b000000000000000e200000000000000e600000000000000e000000000",
            INIT_04 => X"00000091000000000000008e000000000000008a000000000000009000000000",
            INIT_05 => X"0000009a00000000000000950000000000000095000000000000009a00000000",
            INIT_06 => X"000000bb00000000000000ad00000000000000a0000000000000009d00000000",
            INIT_07 => X"0000009d00000000000000a500000000000000b200000000000000be00000000",
            INIT_08 => X"000000e100000000000000c8000000000000003a000000000000000500000000",
            INIT_09 => X"000000e200000000000000d400000000000000c700000000000000c500000000",
            INIT_0A => X"000000e600000000000000e800000000000000e900000000000000e500000000",
            INIT_0B => X"000000d200000000000000dd00000000000000df00000000000000d100000000",
            INIT_0C => X"000000bc00000000000000c100000000000000b400000000000000c600000000",
            INIT_0D => X"000000b800000000000000c000000000000000c200000000000000bd00000000",
            INIT_0E => X"0000009000000000000000a100000000000000ab00000000000000ac00000000",
            INIT_0F => X"0000008a00000000000000800000000000000083000000000000008800000000",
            INIT_10 => X"000000ba00000000000000be0000000000000091000000000000002700000000",
            INIT_11 => X"000000c200000000000000c200000000000000c000000000000000b800000000",
            INIT_12 => X"000000be00000000000000c000000000000000bf00000000000000c200000000",
            INIT_13 => X"00000093000000000000009a00000000000000b400000000000000b100000000",
            INIT_14 => X"000000710000000000000092000000000000009c000000000000009100000000",
            INIT_15 => X"0000006f000000000000007e0000000000000084000000000000007200000000",
            INIT_16 => X"0000005e000000000000005d000000000000005b000000000000005c00000000",
            INIT_17 => X"0000008100000000000000810000000000000079000000000000006900000000",
            INIT_18 => X"00000089000000000000008f00000000000000a2000000000000007a00000000",
            INIT_19 => X"00000082000000000000007f0000000000000080000000000000008300000000",
            INIT_1A => X"00000081000000000000007f0000000000000080000000000000008300000000",
            INIT_1B => X"000000640000000000000068000000000000007c000000000000008100000000",
            INIT_1C => X"0000005e00000000000000700000000000000076000000000000006600000000",
            INIT_1D => X"000000530000000000000057000000000000005e000000000000005e00000000",
            INIT_1E => X"00000065000000000000005d0000000000000053000000000000005000000000",
            INIT_1F => X"0000008200000000000000790000000000000073000000000000006c00000000",
            INIT_20 => X"00000050000000000000004d000000000000004c000000000000004900000000",
            INIT_21 => X"0000005a00000000000000570000000000000057000000000000005400000000",
            INIT_22 => X"00000071000000000000006b0000000000000066000000000000005e00000000",
            INIT_23 => X"0000007800000000000000760000000000000076000000000000007300000000",
            INIT_24 => X"00000064000000000000006a000000000000006e000000000000007300000000",
            INIT_25 => X"00000050000000000000004f0000000000000055000000000000005f00000000",
            INIT_26 => X"000000520000000000000050000000000000004d000000000000005000000000",
            INIT_27 => X"00000088000000000000007d0000000000000071000000000000005c00000000",
            INIT_28 => X"0000001200000000000000090000000000000003000000000000000d00000000",
            INIT_29 => X"0000001600000000000000140000000000000015000000000000001200000000",
            INIT_2A => X"00000030000000000000002a0000000000000022000000000000001a00000000",
            INIT_2B => X"000000460000000000000042000000000000003c000000000000003400000000",
            INIT_2C => X"0000003c00000000000000430000000000000048000000000000004700000000",
            INIT_2D => X"0000003900000000000000350000000000000035000000000000003700000000",
            INIT_2E => X"0000005700000000000000480000000000000039000000000000003900000000",
            INIT_2F => X"0000008900000000000000820000000000000078000000000000006800000000",
            INIT_30 => X"000000200000000000000008000000000000000b000000000000002400000000",
            INIT_31 => X"0000000300000000000000080000000000000016000000000000002400000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_33 => X"0000000300000000000000010000000000000005000000000000000600000000",
            INIT_34 => X"0000001500000000000000150000000000000018000000000000000d00000000",
            INIT_35 => X"00000027000000000000001e0000000000000016000000000000001500000000",
            INIT_36 => X"0000007b00000000000000710000000000000055000000000000003900000000",
            INIT_37 => X"000000990000000000000086000000000000007a000000000000007400000000",
            INIT_38 => X"0000001b000000000000000d000000000000001a000000000000002300000000",
            INIT_39 => X"0000001b00000000000000310000000000000046000000000000004700000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000000a000000000000001f0000000000000039000000000000001100000000",
            INIT_3C => X"0000000e00000000000000070000000000000004000000000000000400000000",
            INIT_3D => X"00000056000000000000003e0000000000000029000000000000001900000000",
            INIT_3E => X"0000007200000000000000840000000000000090000000000000007a00000000",
            INIT_3F => X"000000ac00000000000000920000000000000084000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000030000000000000004000000000000000d000000000000001000000000",
            INIT_41 => X"0000002400000000000000360000000000000041000000000000002d00000000",
            INIT_42 => X"0000000000000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"0000008300000000000000a10000000000000076000000000000000700000000",
            INIT_44 => X"0000006d00000000000000690000000000000069000000000000007000000000",
            INIT_45 => X"00000097000000000000009a000000000000008a000000000000007600000000",
            INIT_46 => X"00000078000000000000006a0000000000000069000000000000007f00000000",
            INIT_47 => X"000000b800000000000000a4000000000000008e000000000000008100000000",
            INIT_48 => X"000000000000000000000000000000000000000c000000000000002800000000",
            INIT_49 => X"000000150000000000000020000000000000001e000000000000000c00000000",
            INIT_4A => X"0000000300000000000000020000000000000002000000000000000700000000",
            INIT_4B => X"000000cd00000000000000b60000000000000044000000000000000000000000",
            INIT_4C => X"000000bb00000000000000c300000000000000c200000000000000c400000000",
            INIT_4D => X"00000067000000000000007b000000000000009600000000000000ac00000000",
            INIT_4E => X"00000081000000000000007a0000000000000068000000000000005f00000000",
            INIT_4F => X"000000b900000000000000ab0000000000000098000000000000008400000000",
            INIT_50 => X"000000010000000000000001000000000000001a000000000000004500000000",
            INIT_51 => X"0000000c0000000000000012000000000000000c000000000000000400000000",
            INIT_52 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_53 => X"000000cb00000000000000990000000000000020000000000000000100000000",
            INIT_54 => X"0000009b00000000000000b300000000000000bf00000000000000c300000000",
            INIT_55 => X"0000005e0000000000000051000000000000005b000000000000007700000000",
            INIT_56 => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_57 => X"000000b800000000000000ad00000000000000a2000000000000009000000000",
            INIT_58 => X"000000020000000000000001000000000000002f000000000000005300000000",
            INIT_59 => X"0000000400000000000000070000000000000005000000000000000200000000",
            INIT_5A => X"0000000300000000000000010000000000000001000000000000000100000000",
            INIT_5B => X"000000cd000000000000008e000000000000001b000000000000000100000000",
            INIT_5C => X"00000055000000000000007900000000000000a900000000000000c600000000",
            INIT_5D => X"0000007900000000000000660000000000000055000000000000004a00000000",
            INIT_5E => X"000000840000000000000079000000000000007a000000000000008000000000",
            INIT_5F => X"000000ba00000000000000b000000000000000a5000000000000009300000000",
            INIT_60 => X"0000000300000000000000060000000000000036000000000000005c00000000",
            INIT_61 => X"0000000100000000000000010000000000000001000000000000000200000000",
            INIT_62 => X"0000000100000000000000010000000000000001000000000000000100000000",
            INIT_63 => X"0000009d0000000000000066000000000000000f000000000000000000000000",
            INIT_64 => X"0000004a0000000000000038000000000000004a000000000000007500000000",
            INIT_65 => X"0000007c000000000000007a0000000000000073000000000000006300000000",
            INIT_66 => X"000000880000000000000080000000000000007d000000000000007b00000000",
            INIT_67 => X"000000bc00000000000000b100000000000000a2000000000000009400000000",
            INIT_68 => X"0000000b0000000000000013000000000000002b000000000000005700000000",
            INIT_69 => X"0000000200000000000000020000000000000005000000000000000800000000",
            INIT_6A => X"0000000200000000000000030000000000000003000000000000000300000000",
            INIT_6B => X"00000047000000000000002a0000000000000004000000000000000000000000",
            INIT_6C => X"0000007100000000000000500000000000000039000000000000003500000000",
            INIT_6D => X"00000074000000000000007b0000000000000086000000000000008400000000",
            INIT_6E => X"0000008f000000000000008b0000000000000083000000000000007800000000",
            INIT_6F => X"000000bc00000000000000b600000000000000a9000000000000009c00000000",
            INIT_70 => X"0000001f0000000000000024000000000000002e000000000000005200000000",
            INIT_71 => X"0000001000000000000000110000000000000016000000000000001b00000000",
            INIT_72 => X"0000001300000000000000140000000000000013000000000000001200000000",
            INIT_73 => X"0000004000000000000000250000000000000017000000000000001300000000",
            INIT_74 => X"0000008000000000000000740000000000000068000000000000005700000000",
            INIT_75 => X"0000007300000000000000750000000000000083000000000000008b00000000",
            INIT_76 => X"00000094000000000000008b0000000000000083000000000000007b00000000",
            INIT_77 => X"000000bb00000000000000b900000000000000ae000000000000009f00000000",
            INIT_78 => X"00000037000000000000003a000000000000003e000000000000005500000000",
            INIT_79 => X"00000030000000000000002e000000000000002f000000000000003300000000",
            INIT_7A => X"0000003700000000000000350000000000000033000000000000003100000000",
            INIT_7B => X"0000006800000000000000510000000000000044000000000000003b00000000",
            INIT_7C => X"0000007f0000000000000085000000000000007f000000000000007400000000",
            INIT_7D => X"0000007a00000000000000720000000000000076000000000000007f00000000",
            INIT_7E => X"00000095000000000000008d0000000000000088000000000000008100000000",
            INIT_7F => X"000000ba00000000000000b400000000000000a8000000000000009e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "sampleifmap_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e900000000000000e900000000000000e700000000000000e700000000",
            INIT_05 => X"000000e900000000000000e800000000000000e700000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e900000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000ea00000000000000ea00000000",
            INIT_0D => X"000000ec00000000000000ec00000000000000ea00000000000000eb00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000eb00000000000000eb00000000000000ea00000000000000e900000000",
            INIT_15 => X"000000ea00000000000000e900000000000000eb00000000000000e600000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e200000000000000e600000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000d200000000000000d800000000000000c000000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000d200000000000000e100000000000000ed00000000000000ee00000000",
            INIT_25 => X"000000e500000000000000da00000000000000cd00000000000000ac00000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e700000000000000ed00000000000000e900000000000000eb00000000",
            INIT_2C => X"000000bc00000000000000c600000000000000cd00000000000000d800000000",
            INIT_2D => X"000000e400000000000000d700000000000000c400000000000000b300000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e400000000000000e600000000000000e300000000000000e500000000",
            INIT_31 => X"000000ed00000000000000ed00000000000000ec00000000000000e800000000",
            INIT_32 => X"000000ed00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_33 => X"000000e200000000000000ed00000000000000e400000000000000e500000000",
            INIT_34 => X"000000b000000000000000b400000000000000b400000000000000c500000000",
            INIT_35 => X"000000ce00000000000000a9000000000000009f00000000000000a300000000",
            INIT_36 => X"000000eb00000000000000ec00000000000000ed00000000000000ee00000000",
            INIT_37 => X"000000ed00000000000000ed00000000000000ee00000000000000ec00000000",
            INIT_38 => X"000000e800000000000000ea00000000000000e600000000000000dc00000000",
            INIT_39 => X"000000ed00000000000000ee00000000000000ed00000000000000ea00000000",
            INIT_3A => X"000000ee00000000000000ec00000000000000ed00000000000000ed00000000",
            INIT_3B => X"000000da00000000000000ec00000000000000de00000000000000cc00000000",
            INIT_3C => X"000000bf00000000000000c900000000000000c900000000000000cc00000000",
            INIT_3D => X"000000c700000000000000b000000000000000ae00000000000000b600000000",
            INIT_3E => X"000000ee00000000000000ee00000000000000ef00000000000000ef00000000",
            INIT_3F => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ef00000000000000ee00000000000000ec00000000000000ea00000000",
            INIT_41 => X"000000ec00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_43 => X"000000e700000000000000ea00000000000000dd00000000000000c600000000",
            INIT_44 => X"000000da00000000000000e400000000000000d800000000000000d500000000",
            INIT_45 => X"000000eb00000000000000e900000000000000e000000000000000dd00000000",
            INIT_46 => X"000000f000000000000000ef00000000000000ee00000000000000f000000000",
            INIT_47 => X"000000ee00000000000000f000000000000000f000000000000000f000000000",
            INIT_48 => X"0000009b000000000000008e000000000000008a000000000000008c00000000",
            INIT_49 => X"000000ea00000000000000ec00000000000000ea00000000000000bc00000000",
            INIT_4A => X"000000ed00000000000000ed00000000000000eb00000000000000e900000000",
            INIT_4B => X"000000ed00000000000000ea00000000000000e400000000000000d800000000",
            INIT_4C => X"000000e800000000000000ec00000000000000e600000000000000e600000000",
            INIT_4D => X"000000cc00000000000000db00000000000000e900000000000000ed00000000",
            INIT_4E => X"000000c700000000000000b400000000000000b300000000000000bd00000000",
            INIT_4F => X"000000f000000000000000f000000000000000f100000000000000eb00000000",
            INIT_50 => X"0000007f000000000000007d0000000000000079000000000000008200000000",
            INIT_51 => X"000000e200000000000000e400000000000000e5000000000000009f00000000",
            INIT_52 => X"000000ed00000000000000ec00000000000000ea00000000000000e800000000",
            INIT_53 => X"000000eb00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_54 => X"000000e800000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_55 => X"0000009c00000000000000a500000000000000b800000000000000ce00000000",
            INIT_56 => X"000000a20000000000000085000000000000008c000000000000009500000000",
            INIT_57 => X"000000f000000000000000f000000000000000f100000000000000e400000000",
            INIT_58 => X"000000d300000000000000d300000000000000ca00000000000000d400000000",
            INIT_59 => X"000000d100000000000000d500000000000000e300000000000000d900000000",
            INIT_5A => X"000000dd00000000000000e200000000000000de00000000000000d500000000",
            INIT_5B => X"000000e500000000000000e100000000000000dd00000000000000db00000000",
            INIT_5C => X"000000e700000000000000ed00000000000000ec00000000000000ea00000000",
            INIT_5D => X"000000c200000000000000c800000000000000c600000000000000cc00000000",
            INIT_5E => X"000000c3000000000000009700000000000000b200000000000000c500000000",
            INIT_5F => X"000000f000000000000000f100000000000000f000000000000000e600000000",
            INIT_60 => X"000000d900000000000000d300000000000000ca00000000000000cf00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000db00000000000000e100000000",
            INIT_62 => X"0000007000000000000000b800000000000000d500000000000000b400000000",
            INIT_63 => X"0000008a00000000000000810000000000000079000000000000007200000000",
            INIT_64 => X"000000ec00000000000000d800000000000000a7000000000000009800000000",
            INIT_65 => X"000000e200000000000000ea00000000000000e900000000000000e800000000",
            INIT_66 => X"000000e600000000000000cb00000000000000db00000000000000e400000000",
            INIT_67 => X"000000f100000000000000ef00000000000000e600000000000000e300000000",
            INIT_68 => X"00000083000000000000007d000000000000007d000000000000008200000000",
            INIT_69 => X"000000c700000000000000c900000000000000b6000000000000009100000000",
            INIT_6A => X"0000004700000000000000ac00000000000000e600000000000000db00000000",
            INIT_6B => X"0000005400000000000000490000000000000049000000000000004600000000",
            INIT_6C => X"000000ef00000000000000e300000000000000a8000000000000007200000000",
            INIT_6D => X"000000d300000000000000e400000000000000e700000000000000ed00000000",
            INIT_6E => X"000000ce00000000000000db00000000000000da00000000000000d000000000",
            INIT_6F => X"000000e700000000000000dd00000000000000c500000000000000ba00000000",
            INIT_70 => X"00000055000000000000004f0000000000000056000000000000005100000000",
            INIT_71 => X"000000c8000000000000009d000000000000009b000000000000008d00000000",
            INIT_72 => X"0000007900000000000000b400000000000000df00000000000000e400000000",
            INIT_73 => X"000000c000000000000000970000000000000075000000000000007000000000",
            INIT_74 => X"000000cb00000000000000db00000000000000de00000000000000d400000000",
            INIT_75 => X"0000008a000000000000009a00000000000000a600000000000000ba00000000",
            INIT_76 => X"0000008e0000000000000092000000000000008b000000000000008500000000",
            INIT_77 => X"000000d400000000000000c50000000000000099000000000000008900000000",
            INIT_78 => X"0000009000000000000000620000000000000046000000000000003500000000",
            INIT_79 => X"0000009e0000000000000073000000000000006b000000000000009700000000",
            INIT_7A => X"000000c100000000000000c200000000000000c200000000000000b400000000",
            INIT_7B => X"000000d200000000000000e400000000000000d100000000000000c200000000",
            INIT_7C => X"00000088000000000000009600000000000000a500000000000000b500000000",
            INIT_7D => X"0000006f000000000000006a000000000000006f000000000000007d00000000",
            INIT_7E => X"0000009700000000000000870000000000000079000000000000007600000000",
            INIT_7F => X"000000cb00000000000000ce00000000000000ae00000000000000a400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "sampleifmap_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d8000000000000008c000000000000001d000000000000000f00000000",
            INIT_01 => X"000000a20000000000000085000000000000007b000000000000009600000000",
            INIT_02 => X"000000ea00000000000000e000000000000000d100000000000000b500000000",
            INIT_03 => X"000000bd00000000000000ee00000000000000f100000000000000ea00000000",
            INIT_04 => X"000000a3000000000000009e000000000000009a000000000000009f00000000",
            INIT_05 => X"000000ab00000000000000a500000000000000a500000000000000ab00000000",
            INIT_06 => X"000000cc00000000000000be00000000000000b100000000000000ae00000000",
            INIT_07 => X"000000af00000000000000b700000000000000c400000000000000cf00000000",
            INIT_08 => X"000000e800000000000000cf000000000000003e000000000000000500000000",
            INIT_09 => X"000000e000000000000000d400000000000000cf00000000000000cd00000000",
            INIT_0A => X"000000ee00000000000000ee00000000000000ec00000000000000e600000000",
            INIT_0B => X"000000e400000000000000ee00000000000000ee00000000000000dd00000000",
            INIT_0C => X"000000d500000000000000d800000000000000c800000000000000d900000000",
            INIT_0D => X"000000cc00000000000000d400000000000000d600000000000000d400000000",
            INIT_0E => X"000000a500000000000000b500000000000000bf00000000000000c100000000",
            INIT_0F => X"0000009a000000000000008f0000000000000092000000000000009c00000000",
            INIT_10 => X"000000c400000000000000cc000000000000009b000000000000002d00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000c500000000",
            INIT_12 => X"000000cf00000000000000cf00000000000000cb00000000000000ce00000000",
            INIT_13 => X"000000a900000000000000b000000000000000c600000000000000c100000000",
            INIT_14 => X"0000008500000000000000a300000000000000ab00000000000000a100000000",
            INIT_15 => X"000000870000000000000096000000000000009d000000000000008900000000",
            INIT_16 => X"0000007400000000000000720000000000000070000000000000007300000000",
            INIT_17 => X"0000008e000000000000008d0000000000000085000000000000007d00000000",
            INIT_18 => X"0000009a00000000000000a000000000000000b3000000000000008700000000",
            INIT_19 => X"0000009600000000000000960000000000000098000000000000009800000000",
            INIT_1A => X"0000009500000000000000930000000000000093000000000000009600000000",
            INIT_1B => X"0000007a000000000000007e0000000000000091000000000000009500000000",
            INIT_1C => X"0000006d00000000000000800000000000000086000000000000007800000000",
            INIT_1D => X"0000006700000000000000700000000000000075000000000000007000000000",
            INIT_1E => X"00000075000000000000006f0000000000000067000000000000006100000000",
            INIT_1F => X"000000900000000000000085000000000000007d000000000000007900000000",
            INIT_20 => X"0000005d000000000000005a000000000000005a000000000000005700000000",
            INIT_21 => X"0000006900000000000000660000000000000066000000000000006200000000",
            INIT_22 => X"00000083000000000000007c0000000000000077000000000000006f00000000",
            INIT_23 => X"0000008500000000000000840000000000000088000000000000008900000000",
            INIT_24 => X"00000077000000000000007f0000000000000085000000000000008800000000",
            INIT_25 => X"0000005c00000000000000610000000000000065000000000000006d00000000",
            INIT_26 => X"0000006200000000000000640000000000000064000000000000005e00000000",
            INIT_27 => X"0000009500000000000000870000000000000077000000000000006800000000",
            INIT_28 => X"0000001a0000000000000010000000000000000b000000000000001900000000",
            INIT_29 => X"0000001e00000000000000190000000000000019000000000000001a00000000",
            INIT_2A => X"0000003b0000000000000033000000000000002b000000000000002400000000",
            INIT_2B => X"0000004f000000000000004d000000000000004b000000000000004500000000",
            INIT_2C => X"0000004800000000000000510000000000000058000000000000005700000000",
            INIT_2D => X"0000004500000000000000450000000000000044000000000000004300000000",
            INIT_2E => X"000000640000000000000059000000000000004e000000000000004700000000",
            INIT_2F => X"000000920000000000000088000000000000007c000000000000007100000000",
            INIT_30 => X"0000002c000000000000000d0000000000000010000000000000002e00000000",
            INIT_31 => X"00000008000000000000000b0000000000000019000000000000002d00000000",
            INIT_32 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_33 => X"0000001700000000000000130000000000000012000000000000000d00000000",
            INIT_34 => X"0000001f00000000000000210000000000000026000000000000001d00000000",
            INIT_35 => X"0000003a0000000000000032000000000000002c000000000000002600000000",
            INIT_36 => X"0000007b0000000000000073000000000000005a000000000000004600000000",
            INIT_37 => X"000000a0000000000000008b000000000000007b000000000000007300000000",
            INIT_38 => X"000000290000000000000013000000000000001b000000000000002900000000",
            INIT_39 => X"0000001f00000000000000320000000000000046000000000000005100000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000002400000000000000320000000000000040000000000000001100000000",
            INIT_3C => X"00000023000000000000001e000000000000001e000000000000001e00000000",
            INIT_3D => X"0000006100000000000000470000000000000037000000000000002b00000000",
            INIT_3E => X"0000006900000000000000780000000000000083000000000000007c00000000",
            INIT_3F => X"000000b300000000000000980000000000000086000000000000006f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000000a000000000000000a000000000000000f00000000",
            INIT_41 => X"00000021000000000000002b0000000000000034000000000000002c00000000",
            INIT_42 => X"0000000100000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"00000080000000000000009e0000000000000075000000000000000800000000",
            INIT_44 => X"0000006900000000000000670000000000000069000000000000007000000000",
            INIT_45 => X"0000007e000000000000007e0000000000000073000000000000006b00000000",
            INIT_46 => X"00000074000000000000005e0000000000000056000000000000006a00000000",
            INIT_47 => X"000000c200000000000000ac0000000000000093000000000000008200000000",
            INIT_48 => X"000000040000000000000003000000000000000a000000000000002800000000",
            INIT_49 => X"0000000a000000000000000c000000000000000c000000000000000600000000",
            INIT_4A => X"0000000200000000000000010000000000000001000000000000000600000000",
            INIT_4B => X"000000820000000000000080000000000000003a000000000000000000000000",
            INIT_4C => X"000000710000000000000077000000000000007b000000000000007f00000000",
            INIT_4D => X"00000042000000000000004b0000000000000060000000000000006e00000000",
            INIT_4E => X"000000840000000000000076000000000000005d000000000000004700000000",
            INIT_4F => X"000000c500000000000000b600000000000000a2000000000000008d00000000",
            INIT_50 => X"000000010000000000000001000000000000001d000000000000004d00000000",
            INIT_51 => X"0000000200000000000000030000000000000002000000000000000100000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_53 => X"0000002f000000000000002d000000000000000c000000000000000100000000",
            INIT_54 => X"0000003100000000000000320000000000000030000000000000002e00000000",
            INIT_55 => X"0000004d00000000000000300000000000000026000000000000002a00000000",
            INIT_56 => X"000000870000000000000080000000000000007e000000000000006e00000000",
            INIT_57 => X"000000c600000000000000bb00000000000000b0000000000000009900000000",
            INIT_58 => X"0000000100000000000000010000000000000034000000000000005e00000000",
            INIT_59 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000002000000000000000190000000000000003000000000000000200000000",
            INIT_5C => X"0000001d00000000000000190000000000000019000000000000001900000000",
            INIT_5D => X"00000071000000000000005c0000000000000042000000000000002900000000",
            INIT_5E => X"0000008b000000000000007f000000000000007e000000000000007c00000000",
            INIT_5F => X"000000c900000000000000bf00000000000000b3000000000000009d00000000",
            INIT_60 => X"000000020000000000000007000000000000003c000000000000006600000000",
            INIT_61 => X"0000000200000000000000030000000000000003000000000000000200000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000001f00000000000000130000000000000001000000000000000300000000",
            INIT_64 => X"0000003a000000000000001b000000000000000d000000000000001100000000",
            INIT_65 => X"0000007c000000000000007e0000000000000073000000000000005a00000000",
            INIT_66 => X"0000009100000000000000870000000000000082000000000000007b00000000",
            INIT_67 => X"000000ca00000000000000c000000000000000b0000000000000009f00000000",
            INIT_68 => X"0000000c00000000000000170000000000000033000000000000006300000000",
            INIT_69 => X"00000007000000000000000a000000000000000b000000000000000a00000000",
            INIT_6A => X"0000000300000000000000040000000000000004000000000000000400000000",
            INIT_6B => X"00000015000000000000000d0000000000000005000000000000000600000000",
            INIT_6C => X"00000062000000000000004d0000000000000032000000000000001b00000000",
            INIT_6D => X"0000007d000000000000007e000000000000007e000000000000007100000000",
            INIT_6E => X"0000009a0000000000000094000000000000008a000000000000008000000000",
            INIT_6F => X"000000ca00000000000000c500000000000000b800000000000000a800000000",
            INIT_70 => X"00000023000000000000002c0000000000000039000000000000006000000000",
            INIT_71 => X"00000017000000000000001a000000000000001c000000000000001e00000000",
            INIT_72 => X"0000001700000000000000160000000000000015000000000000001500000000",
            INIT_73 => X"000000370000000000000028000000000000001f000000000000001b00000000",
            INIT_74 => X"0000007000000000000000660000000000000058000000000000004600000000",
            INIT_75 => X"0000007f000000000000007a000000000000007a000000000000007900000000",
            INIT_76 => X"000000a00000000000000095000000000000008b000000000000008500000000",
            INIT_77 => X"000000ca00000000000000c800000000000000bd00000000000000ac00000000",
            INIT_78 => X"0000003d0000000000000043000000000000004b000000000000006500000000",
            INIT_79 => X"0000003700000000000000350000000000000035000000000000003800000000",
            INIT_7A => X"0000003e000000000000003a0000000000000038000000000000003700000000",
            INIT_7B => X"0000006000000000000000540000000000000047000000000000004300000000",
            INIT_7C => X"000000790000000000000074000000000000006d000000000000006700000000",
            INIT_7D => X"00000083000000000000007d000000000000007c000000000000007f00000000",
            INIT_7E => X"000000a200000000000000980000000000000091000000000000008800000000",
            INIT_7F => X"000000c800000000000000c300000000000000b700000000000000ab00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "sampleifmap_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_05 => X"000000e600000000000000e800000000000000ea00000000000000ea00000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e700000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ea00000000000000e900000000000000e900000000",
            INIT_0D => X"000000eb00000000000000ed00000000000000ee00000000000000ed00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ec00000000000000ea00000000000000e700000000000000e700000000",
            INIT_15 => X"000000ea00000000000000eb00000000000000ee00000000000000e900000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e700000000000000e800000000000000e700000000000000e600000000",
            INIT_1D => X"000000e600000000000000d500000000000000db00000000000000c500000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000db00000000000000e600000000000000ed00000000000000ec00000000",
            INIT_25 => X"000000e800000000000000dd00000000000000d000000000000000b300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e800000000000000ed00000000000000ea00000000000000ec00000000",
            INIT_2C => X"000000c800000000000000cf00000000000000d200000000000000da00000000",
            INIT_2D => X"000000e800000000000000dc00000000000000ca00000000000000bd00000000",
            INIT_2E => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e600000000000000e700000000000000e400000000000000e500000000",
            INIT_31 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_32 => X"000000ee00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_33 => X"000000e400000000000000ee00000000000000e500000000000000e600000000",
            INIT_34 => X"000000be00000000000000bf00000000000000be00000000000000cc00000000",
            INIT_35 => X"000000d300000000000000b100000000000000ab00000000000000b100000000",
            INIT_36 => X"000000eb00000000000000e900000000000000ea00000000000000ef00000000",
            INIT_37 => X"000000ee00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_38 => X"000000ea00000000000000ee00000000000000e900000000000000de00000000",
            INIT_39 => X"000000ec00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_3A => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_3B => X"000000da00000000000000eb00000000000000dd00000000000000cb00000000",
            INIT_3C => X"000000cb00000000000000d300000000000000d200000000000000d200000000",
            INIT_3D => X"000000cc00000000000000b900000000000000bb00000000000000c400000000",
            INIT_3E => X"000000ee00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_3F => X"000000ee00000000000000ee00000000000000ee00000000000000ee00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f300000000000000f600000000000000f300000000000000f100000000",
            INIT_41 => X"000000eb00000000000000eb00000000000000ed00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ed00000000000000ed00000000",
            INIT_43 => X"000000e500000000000000e700000000000000da00000000000000c400000000",
            INIT_44 => X"000000e300000000000000eb00000000000000de00000000000000d900000000",
            INIT_45 => X"000000f100000000000000f000000000000000eb00000000000000ea00000000",
            INIT_46 => X"000000f000000000000000f000000000000000f000000000000000f300000000",
            INIT_47 => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_48 => X"000000a100000000000000990000000000000094000000000000009500000000",
            INIT_49 => X"000000e800000000000000e900000000000000e900000000000000bf00000000",
            INIT_4A => X"000000eb00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000ef00000000000000f100000000000000eb00000000000000e800000000",
            INIT_4D => X"000000d300000000000000e200000000000000f300000000000000f700000000",
            INIT_4E => X"000000c900000000000000b900000000000000ba00000000000000c300000000",
            INIT_4F => X"000000ef00000000000000ef00000000000000ef00000000000000eb00000000",
            INIT_50 => X"0000008900000000000000890000000000000085000000000000008d00000000",
            INIT_51 => X"000000e000000000000000e100000000000000e700000000000000a500000000",
            INIT_52 => X"000000eb00000000000000ea00000000000000ea00000000000000e900000000",
            INIT_53 => X"000000ec00000000000000ee00000000000000ec00000000000000eb00000000",
            INIT_54 => X"000000ee00000000000000f100000000000000f000000000000000ee00000000",
            INIT_55 => X"000000a300000000000000ac00000000000000bf00000000000000d500000000",
            INIT_56 => X"000000a6000000000000008f0000000000000099000000000000009f00000000",
            INIT_57 => X"000000ef00000000000000ee00000000000000ef00000000000000e500000000",
            INIT_58 => X"000000df00000000000000e000000000000000d700000000000000e000000000",
            INIT_59 => X"000000ce00000000000000d300000000000000e700000000000000e300000000",
            INIT_5A => X"000000db00000000000000e100000000000000de00000000000000d600000000",
            INIT_5B => X"000000e900000000000000e600000000000000e100000000000000df00000000",
            INIT_5C => X"000000ed00000000000000f100000000000000ef00000000000000ed00000000",
            INIT_5D => X"000000ca00000000000000cf00000000000000cb00000000000000d000000000",
            INIT_5E => X"000000ca00000000000000a400000000000000c400000000000000d300000000",
            INIT_5F => X"000000ef00000000000000ef00000000000000ee00000000000000e900000000",
            INIT_60 => X"000000ea00000000000000e000000000000000d900000000000000de00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000e300000000000000f100000000",
            INIT_62 => X"0000007900000000000000bc00000000000000d600000000000000b700000000",
            INIT_63 => X"00000093000000000000008b0000000000000084000000000000007e00000000",
            INIT_64 => X"000000ed00000000000000dc00000000000000ae00000000000000a100000000",
            INIT_65 => X"000000e900000000000000f000000000000000ee00000000000000eb00000000",
            INIT_66 => X"000000ed00000000000000d400000000000000e500000000000000ed00000000",
            INIT_67 => X"000000f200000000000000f200000000000000e900000000000000ea00000000",
            INIT_68 => X"00000097000000000000008d0000000000000093000000000000009800000000",
            INIT_69 => X"000000cc00000000000000cd00000000000000c100000000000000a500000000",
            INIT_6A => X"0000005c00000000000000b700000000000000ea00000000000000e200000000",
            INIT_6B => X"00000062000000000000005a000000000000005b000000000000005b00000000",
            INIT_6C => X"000000f100000000000000e900000000000000b3000000000000008100000000",
            INIT_6D => X"000000d900000000000000e900000000000000ed00000000000000f100000000",
            INIT_6E => X"000000d600000000000000df00000000000000dc00000000000000d400000000",
            INIT_6F => X"000000ea00000000000000e300000000000000cd00000000000000c400000000",
            INIT_70 => X"0000006600000000000000640000000000000072000000000000006c00000000",
            INIT_71 => X"000000cf00000000000000a400000000000000a4000000000000009b00000000",
            INIT_72 => X"0000008a00000000000000be00000000000000e400000000000000ea00000000",
            INIT_73 => X"000000cf00000000000000a80000000000000087000000000000008300000000",
            INIT_74 => X"000000d400000000000000e300000000000000e800000000000000df00000000",
            INIT_75 => X"0000009300000000000000a300000000000000ae00000000000000c300000000",
            INIT_76 => X"0000009700000000000000980000000000000090000000000000008c00000000",
            INIT_77 => X"000000d800000000000000cb00000000000000a0000000000000009300000000",
            INIT_78 => X"000000990000000000000074000000000000005e000000000000004d00000000",
            INIT_79 => X"000000a10000000000000076000000000000006e000000000000009c00000000",
            INIT_7A => X"000000c800000000000000c600000000000000c500000000000000b600000000",
            INIT_7B => X"000000d900000000000000ec00000000000000d900000000000000ca00000000",
            INIT_7C => X"00000095000000000000009f00000000000000ac00000000000000ba00000000",
            INIT_7D => X"0000007b0000000000000076000000000000007b000000000000008a00000000",
            INIT_7E => X"000000a100000000000000910000000000000082000000000000008000000000",
            INIT_7F => X"000000d000000000000000d500000000000000b800000000000000ae00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "sampleifmap_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000dc0000000000000097000000000000002f000000000000002300000000",
            INIT_01 => X"000000a20000000000000086000000000000007b000000000000009600000000",
            INIT_02 => X"000000e900000000000000e100000000000000d300000000000000b400000000",
            INIT_03 => X"000000be00000000000000ee00000000000000f000000000000000e800000000",
            INIT_04 => X"000000b100000000000000aa00000000000000a200000000000000a300000000",
            INIT_05 => X"000000bb00000000000000b600000000000000b600000000000000bb00000000",
            INIT_06 => X"000000d900000000000000cc00000000000000bf00000000000000bd00000000",
            INIT_07 => X"000000b700000000000000c100000000000000d000000000000000da00000000",
            INIT_08 => X"000000ef00000000000000d9000000000000004f000000000000001800000000",
            INIT_09 => X"000000e500000000000000da00000000000000d300000000000000d400000000",
            INIT_0A => X"000000ef00000000000000f500000000000000f600000000000000ed00000000",
            INIT_0B => X"000000ea00000000000000f100000000000000ef00000000000000dc00000000",
            INIT_0C => X"000000e500000000000000e600000000000000d600000000000000e400000000",
            INIT_0D => X"000000e000000000000000e800000000000000ea00000000000000e700000000",
            INIT_0E => X"000000b300000000000000c500000000000000d100000000000000d400000000",
            INIT_0F => X"000000a5000000000000009e00000000000000a100000000000000a900000000",
            INIT_10 => X"000000d800000000000000de00000000000000b3000000000000004700000000",
            INIT_11 => X"000000e300000000000000e600000000000000e500000000000000d900000000",
            INIT_12 => X"000000dd00000000000000e400000000000000e400000000000000e300000000",
            INIT_13 => X"000000bc00000000000000c100000000000000d700000000000000cf00000000",
            INIT_14 => X"0000009c00000000000000ba00000000000000c300000000000000b800000000",
            INIT_15 => X"0000009e00000000000000ad00000000000000b400000000000000a100000000",
            INIT_16 => X"0000008300000000000000850000000000000087000000000000008a00000000",
            INIT_17 => X"0000009c000000000000009e0000000000000097000000000000008c00000000",
            INIT_18 => X"000000bd00000000000000c200000000000000cf00000000000000a100000000",
            INIT_19 => X"000000c100000000000000c000000000000000be00000000000000bb00000000",
            INIT_1A => X"000000bd00000000000000bd00000000000000be00000000000000c000000000",
            INIT_1B => X"0000009a00000000000000a300000000000000ba00000000000000bc00000000",
            INIT_1C => X"0000009100000000000000a300000000000000aa000000000000009a00000000",
            INIT_1D => X"0000008800000000000000900000000000000099000000000000009400000000",
            INIT_1E => X"0000008d000000000000008b0000000000000086000000000000008200000000",
            INIT_1F => X"0000009c00000000000000940000000000000092000000000000009000000000",
            INIT_20 => X"0000007f000000000000007a0000000000000071000000000000006d00000000",
            INIT_21 => X"000000960000000000000093000000000000008e000000000000008600000000",
            INIT_22 => X"000000ac00000000000000a500000000000000a0000000000000009800000000",
            INIT_23 => X"000000af00000000000000b400000000000000ba00000000000000b500000000",
            INIT_24 => X"0000009b00000000000000a300000000000000a800000000000000ac00000000",
            INIT_25 => X"0000007f0000000000000084000000000000008b000000000000009400000000",
            INIT_26 => X"0000007a00000000000000810000000000000085000000000000008100000000",
            INIT_27 => X"0000009c0000000000000092000000000000008a000000000000007e00000000",
            INIT_28 => X"0000003000000000000000230000000000000019000000000000002900000000",
            INIT_29 => X"0000003d000000000000003a0000000000000038000000000000003400000000",
            INIT_2A => X"00000057000000000000004d0000000000000046000000000000003e00000000",
            INIT_2B => X"0000007e000000000000007e0000000000000079000000000000006a00000000",
            INIT_2C => X"000000700000000000000078000000000000007e000000000000007f00000000",
            INIT_2D => X"0000006600000000000000670000000000000068000000000000006a00000000",
            INIT_2E => X"000000770000000000000073000000000000006e000000000000006900000000",
            INIT_2F => X"00000095000000000000008d0000000000000088000000000000008000000000",
            INIT_30 => X"0000003500000000000000130000000000000014000000000000003700000000",
            INIT_31 => X"00000018000000000000001e0000000000000029000000000000003a00000000",
            INIT_32 => X"00000014000000000000000f000000000000000f000000000000001100000000",
            INIT_33 => X"0000003e000000000000003c0000000000000038000000000000002a00000000",
            INIT_34 => X"0000004c000000000000004d0000000000000051000000000000004700000000",
            INIT_35 => X"0000005a0000000000000053000000000000004f000000000000004e00000000",
            INIT_36 => X"0000008a000000000000008a0000000000000076000000000000006500000000",
            INIT_37 => X"0000009e00000000000000890000000000000080000000000000007d00000000",
            INIT_38 => X"000000290000000000000012000000000000001a000000000000002d00000000",
            INIT_39 => X"000000250000000000000039000000000000004c000000000000005400000000",
            INIT_3A => X"000000070000000000000007000000000000000b000000000000001500000000",
            INIT_3B => X"0000003e000000000000004e000000000000005b000000000000002300000000",
            INIT_3C => X"00000045000000000000003f000000000000003e000000000000003c00000000",
            INIT_3D => X"0000007b00000000000000630000000000000053000000000000004a00000000",
            INIT_3E => X"0000007200000000000000870000000000000095000000000000009200000000",
            INIT_3F => X"000000af00000000000000920000000000000085000000000000007400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000b00000000000000080000000000000009000000000000001100000000",
            INIT_41 => X"00000023000000000000002f0000000000000039000000000000002e00000000",
            INIT_42 => X"0000000300000000000000040000000000000007000000000000001400000000",
            INIT_43 => X"0000009400000000000000b30000000000000086000000000000000f00000000",
            INIT_44 => X"0000007f000000000000007c000000000000007d000000000000008300000000",
            INIT_45 => X"0000008d00000000000000900000000000000085000000000000007e00000000",
            INIT_46 => X"000000740000000000000061000000000000005b000000000000007400000000",
            INIT_47 => X"000000be00000000000000a50000000000000090000000000000008100000000",
            INIT_48 => X"0000000400000000000000030000000000000007000000000000002300000000",
            INIT_49 => X"0000000c00000000000000110000000000000011000000000000000700000000",
            INIT_4A => X"0000000300000000000000020000000000000003000000000000000700000000",
            INIT_4B => X"0000009400000000000000920000000000000040000000000000000200000000",
            INIT_4C => X"000000810000000000000089000000000000008d000000000000009000000000",
            INIT_4D => X"000000450000000000000053000000000000006a000000000000007a00000000",
            INIT_4E => X"0000007e00000000000000710000000000000058000000000000004600000000",
            INIT_4F => X"000000c200000000000000b0000000000000009e000000000000008700000000",
            INIT_50 => X"0000000200000000000000010000000000000015000000000000004000000000",
            INIT_51 => X"0000000500000000000000090000000000000005000000000000000000000000",
            INIT_52 => X"0000000100000000000000000000000000000000000000000000000200000000",
            INIT_53 => X"00000044000000000000003b000000000000000b000000000000000100000000",
            INIT_54 => X"0000003b00000000000000430000000000000045000000000000004300000000",
            INIT_55 => X"00000047000000000000002e000000000000002a000000000000003100000000",
            INIT_56 => X"0000008000000000000000780000000000000074000000000000006600000000",
            INIT_57 => X"000000c400000000000000b700000000000000ab000000000000009300000000",
            INIT_58 => X"000000020000000000000001000000000000002b000000000000005200000000",
            INIT_59 => X"0000000200000000000000050000000000000002000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000003600000000000000260000000000000002000000000000000000000000",
            INIT_5C => X"000000220000000000000024000000000000002b000000000000002e00000000",
            INIT_5D => X"0000006900000000000000520000000000000038000000000000002700000000",
            INIT_5E => X"0000008300000000000000760000000000000073000000000000007300000000",
            INIT_5F => X"000000c700000000000000bb00000000000000ae000000000000009600000000",
            INIT_60 => X"0000000100000000000000030000000000000032000000000000005d00000000",
            INIT_61 => X"0000000200000000000000030000000000000001000000000000000000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000002f000000000000001c0000000000000000000000000000000200000000",
            INIT_64 => X"000000370000000000000016000000000000000c000000000000001700000000",
            INIT_65 => X"00000070000000000000006f0000000000000063000000000000005100000000",
            INIT_66 => X"00000089000000000000007e0000000000000077000000000000007100000000",
            INIT_67 => X"000000c900000000000000bc00000000000000ab000000000000009700000000",
            INIT_68 => X"00000004000000000000000b0000000000000025000000000000005900000000",
            INIT_69 => X"0000000200000000000000040000000000000004000000000000000200000000",
            INIT_6A => X"0000000200000000000000010000000000000001000000000000000100000000",
            INIT_6B => X"00000018000000000000000d0000000000000002000000000000000600000000",
            INIT_6C => X"00000052000000000000003e0000000000000029000000000000001900000000",
            INIT_6D => X"0000006f00000000000000700000000000000071000000000000006500000000",
            INIT_6E => X"000000910000000000000089000000000000007e000000000000007300000000",
            INIT_6F => X"000000c900000000000000c100000000000000b300000000000000a100000000",
            INIT_70 => X"0000001100000000000000160000000000000024000000000000005200000000",
            INIT_71 => X"0000000c000000000000000d000000000000000f000000000000000f00000000",
            INIT_72 => X"0000000f000000000000000e000000000000000d000000000000000c00000000",
            INIT_73 => X"0000002d000000000000001b0000000000000015000000000000001400000000",
            INIT_74 => X"0000005800000000000000550000000000000051000000000000004300000000",
            INIT_75 => X"00000070000000000000006b000000000000006e000000000000006900000000",
            INIT_76 => X"00000097000000000000008a000000000000007f000000000000007700000000",
            INIT_77 => X"000000c800000000000000c400000000000000b700000000000000a400000000",
            INIT_78 => X"0000002500000000000000260000000000000030000000000000005300000000",
            INIT_79 => X"0000002600000000000000220000000000000021000000000000002300000000",
            INIT_7A => X"0000002e000000000000002c0000000000000029000000000000002800000000",
            INIT_7B => X"0000004a000000000000003b0000000000000030000000000000002d00000000",
            INIT_7C => X"000000610000000000000061000000000000005c000000000000005300000000",
            INIT_7D => X"00000075000000000000006c000000000000006a000000000000006b00000000",
            INIT_7E => X"00000099000000000000008d0000000000000085000000000000007b00000000",
            INIT_7F => X"000000c700000000000000bf00000000000000b200000000000000a300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "sampleifmap_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000084000000000000008b000000000000009e000000000000009e00000000",
            INIT_01 => X"000000c100000000000000bb00000000000000b600000000000000a600000000",
            INIT_02 => X"000000ce00000000000000d100000000000000cd00000000000000c700000000",
            INIT_03 => X"000000e600000000000000e300000000000000df00000000000000da00000000",
            INIT_04 => X"000000eb00000000000000e700000000000000e200000000000000d500000000",
            INIT_05 => X"000000ea00000000000000ea00000000000000e800000000000000ec00000000",
            INIT_06 => X"000000ee00000000000000e600000000000000e200000000000000ec00000000",
            INIT_07 => X"000000ee00000000000000ed00000000000000e400000000000000e800000000",
            INIT_08 => X"00000089000000000000009700000000000000ac00000000000000aa00000000",
            INIT_09 => X"000000c700000000000000c500000000000000c100000000000000ae00000000",
            INIT_0A => X"000000d200000000000000d900000000000000d700000000000000ce00000000",
            INIT_0B => X"000000ed00000000000000e900000000000000e700000000000000e100000000",
            INIT_0C => X"000000f200000000000000e800000000000000e400000000000000db00000000",
            INIT_0D => X"000000f200000000000000ec00000000000000ea00000000000000f500000000",
            INIT_0E => X"000000f300000000000000eb00000000000000e400000000000000f100000000",
            INIT_0F => X"000000f600000000000000f600000000000000e800000000000000e900000000",
            INIT_10 => X"0000008e000000000000009d00000000000000b000000000000000ae00000000",
            INIT_11 => X"000000c700000000000000ce00000000000000c900000000000000b500000000",
            INIT_12 => X"000000d400000000000000da00000000000000df00000000000000d100000000",
            INIT_13 => X"000000ef00000000000000e600000000000000e600000000000000e000000000",
            INIT_14 => X"000000ef00000000000000e900000000000000e400000000000000dd00000000",
            INIT_15 => X"000000f300000000000000ec00000000000000d500000000000000e800000000",
            INIT_16 => X"000000f800000000000000ee00000000000000e700000000000000f500000000",
            INIT_17 => X"000000f500000000000000fa00000000000000e600000000000000ed00000000",
            INIT_18 => X"0000009300000000000000a000000000000000b200000000000000b400000000",
            INIT_19 => X"000000cf00000000000000d400000000000000cb00000000000000ba00000000",
            INIT_1A => X"000000d600000000000000dd00000000000000e400000000000000d600000000",
            INIT_1B => X"000000f000000000000000df00000000000000e700000000000000dc00000000",
            INIT_1C => X"000000e400000000000000e900000000000000e400000000000000e000000000",
            INIT_1D => X"000000f300000000000000e600000000000000ac00000000000000b100000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f400000000000000f900000000000000e400000000000000ee00000000",
            INIT_20 => X"0000009300000000000000a500000000000000b900000000000000ba00000000",
            INIT_21 => X"000000cf00000000000000d900000000000000cc00000000000000bd00000000",
            INIT_22 => X"000000d600000000000000de00000000000000e700000000000000d300000000",
            INIT_23 => X"000000eb00000000000000d300000000000000e700000000000000da00000000",
            INIT_24 => X"000000d400000000000000e800000000000000e000000000000000e200000000",
            INIT_25 => X"000000ed00000000000000e000000000000000a8000000000000009f00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f200000000000000f800000000000000ea00000000000000e800000000",
            INIT_28 => X"0000008e00000000000000aa00000000000000be00000000000000c100000000",
            INIT_29 => X"000000d300000000000000db00000000000000cb00000000000000bf00000000",
            INIT_2A => X"000000d600000000000000dd00000000000000ea00000000000000d700000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e400000000000000d600000000",
            INIT_2C => X"000000c100000000000000eb00000000000000ce00000000000000cf00000000",
            INIT_2D => X"000000e600000000000000de000000000000009e000000000000007000000000",
            INIT_2E => X"000000f100000000000000e200000000000000e500000000000000f500000000",
            INIT_2F => X"000000eb00000000000000f300000000000000e700000000000000e400000000",
            INIT_30 => X"0000008500000000000000ac00000000000000bf00000000000000c400000000",
            INIT_31 => X"000000d900000000000000de00000000000000ca00000000000000bf00000000",
            INIT_32 => X"000000d600000000000000da00000000000000eb00000000000000df00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e300000000000000d700000000",
            INIT_34 => X"000000bb00000000000000cd00000000000000ba00000000000000bb00000000",
            INIT_35 => X"000000b700000000000000ac0000000000000089000000000000007800000000",
            INIT_36 => X"000000eb00000000000000d800000000000000df00000000000000db00000000",
            INIT_37 => X"000000eb00000000000000f000000000000000e100000000000000e200000000",
            INIT_38 => X"0000008c00000000000000ae00000000000000c500000000000000cc00000000",
            INIT_39 => X"000000e000000000000000e000000000000000da00000000000000cb00000000",
            INIT_3A => X"000000dc00000000000000dc00000000000000ed00000000000000e800000000",
            INIT_3B => X"000000cd00000000000000c900000000000000dd00000000000000dc00000000",
            INIT_3C => X"000000530000000000000064000000000000008a00000000000000ac00000000",
            INIT_3D => X"0000003c0000000000000041000000000000003e000000000000004700000000",
            INIT_3E => X"000000e400000000000000d100000000000000b6000000000000006800000000",
            INIT_3F => X"000000ec00000000000000ef00000000000000d400000000000000da00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000089000000000000009d00000000000000aa00000000000000af00000000",
            INIT_41 => X"000000c500000000000000af00000000000000ba00000000000000b000000000",
            INIT_42 => X"000000d200000000000000ce00000000000000d400000000000000d100000000",
            INIT_43 => X"000000c100000000000000c100000000000000c900000000000000d400000000",
            INIT_44 => X"0000005b00000000000000590000000000000069000000000000008e00000000",
            INIT_45 => X"00000045000000000000005e0000000000000053000000000000005400000000",
            INIT_46 => X"000000b700000000000000a20000000000000079000000000000004e00000000",
            INIT_47 => X"000000c300000000000000cf00000000000000a300000000000000ae00000000",
            INIT_48 => X"0000006800000000000000710000000000000073000000000000007200000000",
            INIT_49 => X"00000080000000000000006f000000000000006b000000000000006900000000",
            INIT_4A => X"0000009b00000000000000970000000000000092000000000000008b00000000",
            INIT_4B => X"0000009600000000000000970000000000000093000000000000009d00000000",
            INIT_4C => X"0000006300000000000000630000000000000064000000000000007600000000",
            INIT_4D => X"0000005300000000000000560000000000000056000000000000005500000000",
            INIT_4E => X"00000099000000000000009a0000000000000080000000000000008b00000000",
            INIT_4F => X"0000007b0000000000000084000000000000006d000000000000007600000000",
            INIT_50 => X"00000044000000000000004b000000000000004c000000000000004200000000",
            INIT_51 => X"0000005a0000000000000054000000000000005a000000000000005300000000",
            INIT_52 => X"000000670000000000000066000000000000006a000000000000005d00000000",
            INIT_53 => X"0000006c0000000000000072000000000000006b000000000000006a00000000",
            INIT_54 => X"00000055000000000000005b000000000000005a000000000000005a00000000",
            INIT_55 => X"00000072000000000000005f0000000000000042000000000000004800000000",
            INIT_56 => X"000000c70000000000000093000000000000006e000000000000008000000000",
            INIT_57 => X"0000005e000000000000005c0000000000000067000000000000007d00000000",
            INIT_58 => X"0000004d000000000000004b0000000000000041000000000000003500000000",
            INIT_59 => X"000000460000000000000055000000000000006a000000000000006f00000000",
            INIT_5A => X"0000005d000000000000005f0000000000000071000000000000005d00000000",
            INIT_5B => X"00000061000000000000006b0000000000000073000000000000006c00000000",
            INIT_5C => X"000000610000000000000062000000000000005f000000000000006200000000",
            INIT_5D => X"000000bb00000000000000950000000000000055000000000000005a00000000",
            INIT_5E => X"000000cc0000000000000070000000000000009200000000000000b300000000",
            INIT_5F => X"000000550000000000000057000000000000005f000000000000009a00000000",
            INIT_60 => X"0000004a000000000000005e0000000000000056000000000000003a00000000",
            INIT_61 => X"00000055000000000000004d0000000000000064000000000000006400000000",
            INIT_62 => X"0000006c000000000000007f0000000000000085000000000000007800000000",
            INIT_63 => X"000000570000000000000062000000000000006e000000000000006900000000",
            INIT_64 => X"0000005f00000000000000570000000000000051000000000000005100000000",
            INIT_65 => X"000000c300000000000000aa0000000000000070000000000000005f00000000",
            INIT_66 => X"000000ad000000000000007f00000000000000c100000000000000d000000000",
            INIT_67 => X"0000004f0000000000000055000000000000005000000000000000b200000000",
            INIT_68 => X"0000004b00000000000000570000000000000059000000000000004a00000000",
            INIT_69 => X"0000005000000000000000470000000000000044000000000000005200000000",
            INIT_6A => X"0000006f00000000000000760000000000000067000000000000005900000000",
            INIT_6B => X"000000620000000000000069000000000000006a000000000000006500000000",
            INIT_6C => X"0000006d00000000000000620000000000000062000000000000006000000000",
            INIT_6D => X"000000b800000000000000b4000000000000008e000000000000007200000000",
            INIT_6E => X"0000008400000000000000a000000000000000c000000000000000bf00000000",
            INIT_6F => X"00000043000000000000003c000000000000005000000000000000aa00000000",
            INIT_70 => X"0000004e0000000000000052000000000000004f000000000000004d00000000",
            INIT_71 => X"0000005600000000000000460000000000000048000000000000004f00000000",
            INIT_72 => X"0000008500000000000000810000000000000079000000000000006d00000000",
            INIT_73 => X"0000008300000000000000870000000000000088000000000000008900000000",
            INIT_74 => X"0000009600000000000000920000000000000094000000000000009200000000",
            INIT_75 => X"000000b500000000000000b300000000000000a3000000000000009400000000",
            INIT_76 => X"0000006500000000000000aa00000000000000b000000000000000b900000000",
            INIT_77 => X"0000003b00000000000000370000000000000049000000000000005a00000000",
            INIT_78 => X"00000068000000000000006a000000000000005e000000000000006000000000",
            INIT_79 => X"0000008a00000000000000840000000000000083000000000000006d00000000",
            INIT_7A => X"0000009a000000000000009b0000000000000098000000000000009000000000",
            INIT_7B => X"00000094000000000000009e000000000000009b000000000000009b00000000",
            INIT_7C => X"00000092000000000000009c000000000000009d000000000000009600000000",
            INIT_7D => X"000000a900000000000000920000000000000082000000000000007700000000",
            INIT_7E => X"0000006900000000000000a700000000000000a800000000000000b100000000",
            INIT_7F => X"0000004800000000000000560000000000000062000000000000004500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "sampleifmap_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008300000000000000730000000000000065000000000000006a00000000",
            INIT_01 => X"0000008f00000000000000900000000000000087000000000000008100000000",
            INIT_02 => X"0000009a000000000000009a0000000000000096000000000000009200000000",
            INIT_03 => X"0000009000000000000000970000000000000099000000000000009a00000000",
            INIT_04 => X"0000007f000000000000008b0000000000000086000000000000008200000000",
            INIT_05 => X"0000009f00000000000000920000000000000075000000000000005e00000000",
            INIT_06 => X"0000008400000000000000a200000000000000a300000000000000a700000000",
            INIT_07 => X"00000069000000000000009a00000000000000c0000000000000009000000000",
            INIT_08 => X"0000006d0000000000000076000000000000006c000000000000005f00000000",
            INIT_09 => X"000000910000000000000081000000000000005d000000000000005f00000000",
            INIT_0A => X"0000009000000000000000960000000000000097000000000000009500000000",
            INIT_0B => X"0000007b000000000000007a000000000000007e000000000000008600000000",
            INIT_0C => X"00000094000000000000009b0000000000000085000000000000007a00000000",
            INIT_0D => X"0000009c00000000000000a20000000000000093000000000000008300000000",
            INIT_0E => X"0000009500000000000000990000000000000097000000000000009d00000000",
            INIT_0F => X"00000094000000000000009d00000000000000a4000000000000009f00000000",
            INIT_10 => X"0000004600000000000000490000000000000059000000000000006600000000",
            INIT_11 => X"0000008c000000000000007b000000000000006f000000000000005600000000",
            INIT_12 => X"0000007500000000000000780000000000000081000000000000008f00000000",
            INIT_13 => X"0000008d0000000000000085000000000000007e000000000000007800000000",
            INIT_14 => X"0000009f0000000000000099000000000000008e000000000000009600000000",
            INIT_15 => X"000000a100000000000000a5000000000000009d000000000000009700000000",
            INIT_16 => X"00000090000000000000009a0000000000000098000000000000009900000000",
            INIT_17 => X"00000095000000000000007d0000000000000079000000000000008300000000",
            INIT_18 => X"0000006e0000000000000047000000000000003d000000000000005600000000",
            INIT_19 => X"0000007b0000000000000082000000000000008a000000000000008000000000",
            INIT_1A => X"000000840000000000000076000000000000006c000000000000007600000000",
            INIT_1B => X"00000099000000000000009c0000000000000098000000000000008f00000000",
            INIT_1C => X"0000009a00000000000000910000000000000089000000000000009500000000",
            INIT_1D => X"000000a400000000000000a0000000000000009a000000000000009900000000",
            INIT_1E => X"00000069000000000000007d0000000000000090000000000000009800000000",
            INIT_1F => X"000000840000000000000056000000000000004b000000000000005c00000000",
            INIT_20 => X"00000072000000000000006b0000000000000067000000000000006800000000",
            INIT_21 => X"00000076000000000000007b0000000000000074000000000000007300000000",
            INIT_22 => X"00000090000000000000008d0000000000000086000000000000007400000000",
            INIT_23 => X"000000750000000000000085000000000000008d000000000000008f00000000",
            INIT_24 => X"0000009600000000000000820000000000000059000000000000006200000000",
            INIT_25 => X"000000910000000000000098000000000000009a000000000000009700000000",
            INIT_26 => X"00000050000000000000005a0000000000000060000000000000007500000000",
            INIT_27 => X"0000004100000000000000490000000000000047000000000000004100000000",
            INIT_28 => X"0000006f000000000000006f000000000000006b000000000000006300000000",
            INIT_29 => X"0000007e000000000000007d0000000000000077000000000000007200000000",
            INIT_2A => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_2B => X"0000003d000000000000005b0000000000000082000000000000008300000000",
            INIT_2C => X"0000009400000000000000730000000000000038000000000000003900000000",
            INIT_2D => X"0000005f00000000000000720000000000000082000000000000008b00000000",
            INIT_2E => X"0000003a00000000000000490000000000000053000000000000005600000000",
            INIT_2F => X"0000001b0000000000000033000000000000004b000000000000003c00000000",
            INIT_30 => X"0000007200000000000000740000000000000068000000000000003e00000000",
            INIT_31 => X"0000005b00000000000000660000000000000075000000000000007400000000",
            INIT_32 => X"00000070000000000000004e0000000000000051000000000000005400000000",
            INIT_33 => X"0000004c00000000000000600000000000000082000000000000008500000000",
            INIT_34 => X"0000006c000000000000006b0000000000000056000000000000005300000000",
            INIT_35 => X"0000005100000000000000530000000000000058000000000000006000000000",
            INIT_36 => X"0000002d0000000000000033000000000000003d000000000000004600000000",
            INIT_37 => X"00000018000000000000001e000000000000002e000000000000003400000000",
            INIT_38 => X"00000069000000000000006a0000000000000060000000000000003900000000",
            INIT_39 => X"0000003500000000000000410000000000000068000000000000006b00000000",
            INIT_3A => X"0000006e00000000000000440000000000000040000000000000003b00000000",
            INIT_3B => X"0000006200000000000000730000000000000085000000000000008700000000",
            INIT_3C => X"00000050000000000000004e000000000000004f000000000000005800000000",
            INIT_3D => X"0000003700000000000000460000000000000050000000000000005100000000",
            INIT_3E => X"00000029000000000000002d0000000000000031000000000000002c00000000",
            INIT_3F => X"00000018000000000000001b000000000000001e000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000068000000000000005a000000000000004100000000",
            INIT_41 => X"00000049000000000000004f000000000000006d000000000000006d00000000",
            INIT_42 => X"0000006a00000000000000620000000000000058000000000000005500000000",
            INIT_43 => X"0000004100000000000000440000000000000053000000000000006200000000",
            INIT_44 => X"000000520000000000000051000000000000004a000000000000004600000000",
            INIT_45 => X"0000002c00000000000000290000000000000033000000000000004800000000",
            INIT_46 => X"0000002300000000000000270000000000000037000000000000003d00000000",
            INIT_47 => X"00000019000000000000001b000000000000001e000000000000002000000000",
            INIT_48 => X"0000006700000000000000690000000000000057000000000000004300000000",
            INIT_49 => X"0000005100000000000000580000000000000063000000000000006600000000",
            INIT_4A => X"00000039000000000000003b0000000000000045000000000000004c00000000",
            INIT_4B => X"000000460000000000000042000000000000003f000000000000003a00000000",
            INIT_4C => X"00000036000000000000003e0000000000000044000000000000004800000000",
            INIT_4D => X"0000002c0000000000000031000000000000002f000000000000002e00000000",
            INIT_4E => X"0000001c000000000000001e000000000000002e000000000000003800000000",
            INIT_4F => X"0000001e00000000000000180000000000000019000000000000001d00000000",
            INIT_50 => X"0000003a0000000000000041000000000000003a000000000000003600000000",
            INIT_51 => X"0000002c000000000000002d0000000000000032000000000000003700000000",
            INIT_52 => X"0000003a00000000000000370000000000000033000000000000002e00000000",
            INIT_53 => X"0000003a000000000000003e0000000000000040000000000000003e00000000",
            INIT_54 => X"0000003000000000000000250000000000000026000000000000003300000000",
            INIT_55 => X"00000026000000000000002a0000000000000030000000000000003100000000",
            INIT_56 => X"0000001c000000000000001b0000000000000020000000000000002900000000",
            INIT_57 => X"0000001f000000000000001c0000000000000019000000000000001b00000000",
            INIT_58 => X"0000001b000000000000001a000000000000001d000000000000001e00000000",
            INIT_59 => X"0000002700000000000000210000000000000020000000000000001f00000000",
            INIT_5A => X"0000003300000000000000350000000000000034000000000000003100000000",
            INIT_5B => X"0000002800000000000000260000000000000028000000000000002e00000000",
            INIT_5C => X"000000370000000000000042000000000000002c000000000000002600000000",
            INIT_5D => X"0000002500000000000000240000000000000025000000000000002900000000",
            INIT_5E => X"0000001b000000000000001a000000000000001b000000000000001f00000000",
            INIT_5F => X"000000170000000000000021000000000000001e000000000000001c00000000",
            INIT_60 => X"0000001c000000000000001b000000000000001f000000000000002100000000",
            INIT_61 => X"00000020000000000000001f000000000000001e000000000000001c00000000",
            INIT_62 => X"0000001e000000000000001e0000000000000021000000000000002300000000",
            INIT_63 => X"0000002d00000000000000290000000000000027000000000000002200000000",
            INIT_64 => X"0000003100000000000000490000000000000034000000000000002a00000000",
            INIT_65 => X"0000002000000000000000260000000000000023000000000000001e00000000",
            INIT_66 => X"0000001d000000000000001b000000000000001a000000000000001b00000000",
            INIT_67 => X"0000000d000000000000001a0000000000000026000000000000001e00000000",
            INIT_68 => X"0000001a000000000000001a000000000000001e000000000000001f00000000",
            INIT_69 => X"0000001b000000000000001a0000000000000019000000000000001900000000",
            INIT_6A => X"0000002800000000000000250000000000000020000000000000001d00000000",
            INIT_6B => X"0000002a00000000000000280000000000000029000000000000002a00000000",
            INIT_6C => X"000000260000000000000040000000000000002e000000000000002700000000",
            INIT_6D => X"0000001d000000000000001e0000000000000024000000000000001c00000000",
            INIT_6E => X"0000001c000000000000001b0000000000000019000000000000001a00000000",
            INIT_6F => X"0000000400000000000000090000000000000025000000000000002100000000",
            INIT_70 => X"0000001c0000000000000019000000000000001b000000000000001700000000",
            INIT_71 => X"0000002500000000000000220000000000000020000000000000001e00000000",
            INIT_72 => X"0000002700000000000000280000000000000027000000000000002700000000",
            INIT_73 => X"00000021000000000000001e0000000000000023000000000000002600000000",
            INIT_74 => X"0000002400000000000000390000000000000024000000000000001c00000000",
            INIT_75 => X"0000001d000000000000001d000000000000001d000000000000001e00000000",
            INIT_76 => X"0000001b00000000000000170000000000000018000000000000001800000000",
            INIT_77 => X"0000000500000000000000040000000000000013000000000000002400000000",
            INIT_78 => X"000000220000000000000020000000000000001e000000000000001c00000000",
            INIT_79 => X"0000002500000000000000230000000000000022000000000000002100000000",
            INIT_7A => X"0000002200000000000000240000000000000026000000000000002600000000",
            INIT_7B => X"0000000c000000000000000f0000000000000018000000000000001e00000000",
            INIT_7C => X"00000020000000000000002d0000000000000013000000000000000800000000",
            INIT_7D => X"0000001c000000000000001b000000000000001b000000000000001900000000",
            INIT_7E => X"0000002200000000000000140000000000000015000000000000001800000000",
            INIT_7F => X"0000000700000000000000040000000000000005000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "sampleifmap_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009e00000000000000a600000000000000bb00000000000000be00000000",
            INIT_01 => X"000000d800000000000000d300000000000000d000000000000000c100000000",
            INIT_02 => X"000000da00000000000000de00000000000000dd00000000000000db00000000",
            INIT_03 => X"000000ed00000000000000eb00000000000000e800000000000000e500000000",
            INIT_04 => X"000000ef00000000000000ee00000000000000e900000000000000dc00000000",
            INIT_05 => X"000000f100000000000000f100000000000000ef00000000000000f100000000",
            INIT_06 => X"000000f300000000000000eb00000000000000e700000000000000f200000000",
            INIT_07 => X"000000f100000000000000ef00000000000000e700000000000000ed00000000",
            INIT_08 => X"000000a000000000000000b000000000000000c700000000000000c800000000",
            INIT_09 => X"000000da00000000000000da00000000000000d900000000000000c700000000",
            INIT_0A => X"000000db00000000000000e500000000000000e500000000000000df00000000",
            INIT_0B => X"000000f300000000000000ef00000000000000ee00000000000000e900000000",
            INIT_0C => X"000000f500000000000000ee00000000000000ea00000000000000e100000000",
            INIT_0D => X"000000f500000000000000ef00000000000000ed00000000000000f700000000",
            INIT_0E => X"000000f800000000000000ef00000000000000e900000000000000f500000000",
            INIT_0F => X"000000f700000000000000f600000000000000e800000000000000ec00000000",
            INIT_10 => X"000000a200000000000000b300000000000000c800000000000000c900000000",
            INIT_11 => X"000000d600000000000000df00000000000000dc00000000000000c900000000",
            INIT_12 => X"000000db00000000000000e200000000000000e900000000000000dd00000000",
            INIT_13 => X"000000f400000000000000ea00000000000000ea00000000000000e500000000",
            INIT_14 => X"000000f300000000000000ee00000000000000e900000000000000e200000000",
            INIT_15 => X"000000f100000000000000ea00000000000000d600000000000000eb00000000",
            INIT_16 => X"000000fa00000000000000f000000000000000e900000000000000f700000000",
            INIT_17 => X"000000f400000000000000f900000000000000e500000000000000ee00000000",
            INIT_18 => X"000000a400000000000000b300000000000000c700000000000000cb00000000",
            INIT_19 => X"000000d900000000000000e100000000000000d900000000000000c900000000",
            INIT_1A => X"000000d900000000000000e300000000000000eb00000000000000df00000000",
            INIT_1B => X"000000f400000000000000e200000000000000e800000000000000dd00000000",
            INIT_1C => X"000000eb00000000000000ed00000000000000e700000000000000e400000000",
            INIT_1D => X"000000f100000000000000e400000000000000af00000000000000b800000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f200000000000000f700000000000000e300000000000000ed00000000",
            INIT_20 => X"000000a100000000000000b500000000000000cc00000000000000cf00000000",
            INIT_21 => X"000000d500000000000000e100000000000000d600000000000000c900000000",
            INIT_22 => X"000000d700000000000000e200000000000000ed00000000000000d700000000",
            INIT_23 => X"000000ec00000000000000d400000000000000e500000000000000d900000000",
            INIT_24 => X"000000e100000000000000ec00000000000000e100000000000000e300000000",
            INIT_25 => X"000000ec00000000000000e000000000000000ae00000000000000aa00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000ef00000000000000f500000000000000e700000000000000e700000000",
            INIT_28 => X"0000009a00000000000000b700000000000000cd00000000000000d000000000",
            INIT_29 => X"000000d700000000000000e200000000000000d400000000000000c900000000",
            INIT_2A => X"000000d700000000000000df00000000000000ee00000000000000da00000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e500000000000000d700000000",
            INIT_2C => X"000000cc00000000000000ef00000000000000d000000000000000d100000000",
            INIT_2D => X"000000e900000000000000e300000000000000a7000000000000007c00000000",
            INIT_2E => X"000000ef00000000000000e100000000000000e500000000000000f600000000",
            INIT_2F => X"000000e800000000000000f100000000000000e600000000000000e200000000",
            INIT_30 => X"0000008b00000000000000b300000000000000c700000000000000cc00000000",
            INIT_31 => X"000000d500000000000000dd00000000000000cb00000000000000c200000000",
            INIT_32 => X"000000d400000000000000d800000000000000e900000000000000db00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e600000000000000d800000000",
            INIT_34 => X"000000c000000000000000d400000000000000c000000000000000be00000000",
            INIT_35 => X"000000be00000000000000b70000000000000097000000000000008100000000",
            INIT_36 => X"000000e500000000000000d600000000000000e000000000000000e000000000",
            INIT_37 => X"000000e000000000000000eb00000000000000de00000000000000db00000000",
            INIT_38 => X"0000008a00000000000000af00000000000000c600000000000000cd00000000",
            INIT_39 => X"000000cc00000000000000ce00000000000000cb00000000000000c000000000",
            INIT_3A => X"000000d200000000000000d000000000000000df00000000000000d400000000",
            INIT_3B => X"000000ce00000000000000c700000000000000d800000000000000d500000000",
            INIT_3C => X"0000005d0000000000000071000000000000009500000000000000b200000000",
            INIT_3D => X"0000004500000000000000500000000000000050000000000000005500000000",
            INIT_3E => X"000000de00000000000000ce00000000000000b7000000000000006c00000000",
            INIT_3F => X"000000d400000000000000dd00000000000000c500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000085000000000000009a00000000000000a800000000000000ad00000000",
            INIT_41 => X"000000b300000000000000a000000000000000ac00000000000000a500000000",
            INIT_42 => X"000000c300000000000000bd00000000000000c200000000000000be00000000",
            INIT_43 => X"000000c600000000000000c100000000000000bf00000000000000c700000000",
            INIT_44 => X"0000006c000000000000006b0000000000000079000000000000009800000000",
            INIT_45 => X"0000004f000000000000006e0000000000000068000000000000006800000000",
            INIT_46 => X"000000af000000000000009f000000000000007a000000000000005200000000",
            INIT_47 => X"000000af00000000000000be000000000000009500000000000000a300000000",
            INIT_48 => X"0000006900000000000000720000000000000074000000000000007300000000",
            INIT_49 => X"0000007f0000000000000070000000000000006e000000000000006d00000000",
            INIT_4A => X"00000093000000000000008c0000000000000088000000000000008700000000",
            INIT_4B => X"000000a1000000000000009e000000000000008f000000000000009700000000",
            INIT_4C => X"0000007800000000000000780000000000000077000000000000008600000000",
            INIT_4D => X"0000005c0000000000000066000000000000006c000000000000006c00000000",
            INIT_4E => X"0000009100000000000000970000000000000080000000000000008f00000000",
            INIT_4F => X"000000780000000000000082000000000000006a000000000000006e00000000",
            INIT_50 => X"0000005200000000000000560000000000000057000000000000004e00000000",
            INIT_51 => X"0000006400000000000000610000000000000069000000000000006300000000",
            INIT_52 => X"0000006f000000000000006a000000000000006d000000000000006500000000",
            INIT_53 => X"0000007f00000000000000840000000000000076000000000000007200000000",
            INIT_54 => X"0000006b000000000000006e000000000000006d000000000000006d00000000",
            INIT_55 => X"00000077000000000000006c0000000000000057000000000000006000000000",
            INIT_56 => X"000000bf0000000000000090000000000000006f000000000000008400000000",
            INIT_57 => X"000000680000000000000066000000000000006f000000000000007800000000",
            INIT_58 => X"00000062000000000000005f0000000000000055000000000000004a00000000",
            INIT_59 => X"000000510000000000000062000000000000007a000000000000008000000000",
            INIT_5A => X"0000007300000000000000710000000000000081000000000000006800000000",
            INIT_5B => X"0000007b0000000000000086000000000000008b000000000000008400000000",
            INIT_5C => X"0000007700000000000000740000000000000073000000000000007800000000",
            INIT_5D => X"000000bd000000000000009e0000000000000068000000000000007100000000",
            INIT_5E => X"000000c5000000000000006d000000000000009400000000000000b700000000",
            INIT_5F => X"0000006300000000000000630000000000000067000000000000009500000000",
            INIT_60 => X"0000005d0000000000000071000000000000006b000000000000005100000000",
            INIT_61 => X"00000066000000000000005d0000000000000073000000000000007500000000",
            INIT_62 => X"0000008300000000000000950000000000000098000000000000008900000000",
            INIT_63 => X"00000071000000000000007d0000000000000088000000000000008200000000",
            INIT_64 => X"0000007b0000000000000072000000000000006c000000000000006c00000000",
            INIT_65 => X"000000c200000000000000af000000000000007f000000000000007600000000",
            INIT_66 => X"000000a2000000000000007600000000000000bd00000000000000ce00000000",
            INIT_67 => X"000000650000000000000062000000000000005000000000000000a700000000",
            INIT_68 => X"0000005d000000000000006a000000000000006e000000000000006100000000",
            INIT_69 => X"0000006400000000000000590000000000000054000000000000006200000000",
            INIT_6A => X"00000086000000000000008a000000000000007b000000000000006e00000000",
            INIT_6B => X"0000007c00000000000000820000000000000083000000000000007e00000000",
            INIT_6C => X"00000087000000000000007e000000000000007f000000000000007b00000000",
            INIT_6D => X"000000b400000000000000b50000000000000099000000000000008600000000",
            INIT_6E => X"0000007a000000000000009700000000000000b700000000000000b800000000",
            INIT_6F => X"000000590000000000000048000000000000004d00000000000000a000000000",
            INIT_70 => X"0000006100000000000000660000000000000065000000000000006600000000",
            INIT_71 => X"0000006b00000000000000580000000000000058000000000000005f00000000",
            INIT_72 => X"0000009e0000000000000097000000000000008e000000000000008200000000",
            INIT_73 => X"0000009d00000000000000a100000000000000a400000000000000a300000000",
            INIT_74 => X"000000a900000000000000aa00000000000000ad00000000000000ab00000000",
            INIT_75 => X"000000ae00000000000000b100000000000000a900000000000000a200000000",
            INIT_76 => X"0000006200000000000000a400000000000000a800000000000000b000000000",
            INIT_77 => X"0000004b000000000000003f0000000000000046000000000000005700000000",
            INIT_78 => X"0000007c000000000000007f0000000000000076000000000000007b00000000",
            INIT_79 => X"000000a000000000000000980000000000000094000000000000007e00000000",
            INIT_7A => X"000000b400000000000000b300000000000000af00000000000000a700000000",
            INIT_7B => X"000000ae00000000000000b900000000000000b800000000000000b700000000",
            INIT_7C => X"000000a000000000000000af00000000000000b200000000000000ad00000000",
            INIT_7D => X"000000a1000000000000008e0000000000000085000000000000008000000000",
            INIT_7E => X"0000006c00000000000000a600000000000000a200000000000000a900000000",
            INIT_7F => X"000000520000000000000059000000000000005f000000000000004600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "sampleifmap_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000098000000000000008a000000000000007d000000000000008500000000",
            INIT_01 => X"000000a700000000000000a6000000000000009a000000000000009400000000",
            INIT_02 => X"000000b600000000000000b300000000000000ae00000000000000aa00000000",
            INIT_03 => X"000000ab00000000000000b500000000000000b900000000000000b900000000",
            INIT_04 => X"0000008b000000000000009a0000000000000098000000000000009800000000",
            INIT_05 => X"0000009b00000000000000900000000000000078000000000000006600000000",
            INIT_06 => X"0000008800000000000000a300000000000000a200000000000000a500000000",
            INIT_07 => X"0000006c000000000000009900000000000000bb000000000000009100000000",
            INIT_08 => X"00000083000000000000008d0000000000000085000000000000007c00000000",
            INIT_09 => X"000000aa00000000000000980000000000000072000000000000007400000000",
            INIT_0A => X"000000ad00000000000000b000000000000000af00000000000000af00000000",
            INIT_0B => X"00000097000000000000009a00000000000000a000000000000000a700000000",
            INIT_0C => X"000000a000000000000000a80000000000000096000000000000009000000000",
            INIT_0D => X"0000009e00000000000000a50000000000000098000000000000008c00000000",
            INIT_0E => X"00000097000000000000009c000000000000009b00000000000000a300000000",
            INIT_0F => X"000000930000000000000098000000000000009e000000000000009e00000000",
            INIT_10 => X"0000005d00000000000000600000000000000071000000000000008100000000",
            INIT_11 => X"000000a400000000000000940000000000000087000000000000006e00000000",
            INIT_12 => X"000000920000000000000096000000000000009f00000000000000a900000000",
            INIT_13 => X"000000a5000000000000009f0000000000000099000000000000009400000000",
            INIT_14 => X"000000ac00000000000000a800000000000000a000000000000000aa00000000",
            INIT_15 => X"000000a400000000000000a800000000000000a400000000000000a100000000",
            INIT_16 => X"00000092000000000000009e000000000000009e00000000000000a000000000",
            INIT_17 => X"00000096000000000000007d0000000000000079000000000000008400000000",
            INIT_18 => X"0000008700000000000000600000000000000055000000000000007000000000",
            INIT_19 => X"00000093000000000000009c00000000000000a5000000000000009b00000000",
            INIT_1A => X"000000a00000000000000097000000000000008d000000000000008e00000000",
            INIT_1B => X"000000ab00000000000000ae00000000000000ad00000000000000a700000000",
            INIT_1C => X"000000a800000000000000a2000000000000009b00000000000000a700000000",
            INIT_1D => X"000000a600000000000000a300000000000000a100000000000000a300000000",
            INIT_1E => X"0000006f00000000000000820000000000000097000000000000009e00000000",
            INIT_1F => X"0000008a000000000000005c0000000000000052000000000000006200000000",
            INIT_20 => X"0000008f00000000000000870000000000000084000000000000008500000000",
            INIT_21 => X"0000008e0000000000000096000000000000008f000000000000008f00000000",
            INIT_22 => X"000000ab00000000000000a900000000000000a1000000000000008a00000000",
            INIT_23 => X"00000086000000000000009700000000000000a500000000000000a900000000",
            INIT_24 => X"000000a40000000000000094000000000000006b000000000000007400000000",
            INIT_25 => X"00000098000000000000009f00000000000000a300000000000000a300000000",
            INIT_26 => X"0000005b0000000000000066000000000000006c000000000000008000000000",
            INIT_27 => X"000000480000000000000050000000000000004e000000000000004b00000000",
            INIT_28 => X"0000008f0000000000000090000000000000008c000000000000008400000000",
            INIT_29 => X"0000009600000000000000970000000000000093000000000000009000000000",
            INIT_2A => X"0000009a00000000000000940000000000000092000000000000008b00000000",
            INIT_2B => X"0000004e000000000000006e000000000000009c000000000000009f00000000",
            INIT_2C => X"000000a30000000000000084000000000000004a000000000000004b00000000",
            INIT_2D => X"0000006d000000000000007e000000000000008f000000000000009900000000",
            INIT_2E => X"0000004c000000000000005a0000000000000064000000000000006700000000",
            INIT_2F => X"0000002100000000000000390000000000000052000000000000004b00000000",
            INIT_30 => X"0000009200000000000000940000000000000089000000000000005e00000000",
            INIT_31 => X"0000007300000000000000810000000000000091000000000000009200000000",
            INIT_32 => X"0000008700000000000000630000000000000066000000000000006a00000000",
            INIT_33 => X"0000005d0000000000000072000000000000009a000000000000009d00000000",
            INIT_34 => X"0000007c000000000000007d0000000000000068000000000000006500000000",
            INIT_35 => X"000000650000000000000066000000000000006a000000000000007100000000",
            INIT_36 => X"0000003f0000000000000045000000000000004f000000000000005800000000",
            INIT_37 => X"0000001f00000000000000250000000000000035000000000000004300000000",
            INIT_38 => X"000000860000000000000086000000000000007d000000000000005600000000",
            INIT_39 => X"0000004d000000000000005c0000000000000085000000000000008900000000",
            INIT_3A => X"00000083000000000000005c0000000000000059000000000000005200000000",
            INIT_3B => X"0000007300000000000000840000000000000096000000000000009900000000",
            INIT_3C => X"0000006100000000000000600000000000000061000000000000006a00000000",
            INIT_3D => X"0000004f000000000000005f0000000000000065000000000000006300000000",
            INIT_3E => X"00000039000000000000003c0000000000000040000000000000003c00000000",
            INIT_3F => X"0000001f00000000000000220000000000000026000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008300000000000000810000000000000074000000000000005a00000000",
            INIT_41 => X"00000061000000000000006a000000000000008a000000000000008900000000",
            INIT_42 => X"0000007e000000000000007c0000000000000074000000000000006c00000000",
            INIT_43 => X"000000530000000000000054000000000000005f000000000000007100000000",
            INIT_44 => X"000000640000000000000062000000000000005c000000000000005900000000",
            INIT_45 => X"000000450000000000000043000000000000004a000000000000005c00000000",
            INIT_46 => X"0000002e00000000000000330000000000000042000000000000004a00000000",
            INIT_47 => X"0000002000000000000000230000000000000026000000000000002b00000000",
            INIT_48 => X"0000007f00000000000000820000000000000070000000000000005c00000000",
            INIT_49 => X"00000066000000000000006e0000000000000078000000000000007c00000000",
            INIT_4A => X"0000004c0000000000000050000000000000005a000000000000006100000000",
            INIT_4B => X"0000005b00000000000000540000000000000050000000000000004b00000000",
            INIT_4C => X"0000004900000000000000510000000000000059000000000000005f00000000",
            INIT_4D => X"0000003d00000000000000430000000000000041000000000000004100000000",
            INIT_4E => X"00000028000000000000002a000000000000003a000000000000004500000000",
            INIT_4F => X"0000002500000000000000230000000000000028000000000000002a00000000",
            INIT_50 => X"0000004e0000000000000056000000000000004f000000000000004c00000000",
            INIT_51 => X"0000003f00000000000000400000000000000045000000000000004a00000000",
            INIT_52 => X"0000004d000000000000004a0000000000000046000000000000004100000000",
            INIT_53 => X"0000005000000000000000510000000000000052000000000000005100000000",
            INIT_54 => X"000000440000000000000037000000000000003b000000000000004900000000",
            INIT_55 => X"000000320000000000000036000000000000003f000000000000004300000000",
            INIT_56 => X"000000280000000000000028000000000000002d000000000000003600000000",
            INIT_57 => X"0000002500000000000000270000000000000028000000000000002900000000",
            INIT_58 => X"0000002a0000000000000028000000000000002b000000000000002d00000000",
            INIT_59 => X"0000003a00000000000000350000000000000034000000000000003100000000",
            INIT_5A => X"0000004600000000000000480000000000000047000000000000004400000000",
            INIT_5B => X"0000003b000000000000003a000000000000003b000000000000004100000000",
            INIT_5C => X"000000490000000000000055000000000000003f000000000000003800000000",
            INIT_5D => X"0000002f000000000000002f0000000000000033000000000000003900000000",
            INIT_5E => X"0000002800000000000000270000000000000028000000000000002c00000000",
            INIT_5F => X"0000001d000000000000002a000000000000002a000000000000002900000000",
            INIT_60 => X"0000002600000000000000240000000000000028000000000000002b00000000",
            INIT_61 => X"0000003200000000000000310000000000000030000000000000002c00000000",
            INIT_62 => X"0000003100000000000000310000000000000034000000000000003500000000",
            INIT_63 => X"0000003d000000000000003e000000000000003b000000000000003500000000",
            INIT_64 => X"00000042000000000000005e0000000000000045000000000000003700000000",
            INIT_65 => X"00000028000000000000002f000000000000002e000000000000002c00000000",
            INIT_66 => X"0000002a00000000000000280000000000000027000000000000002700000000",
            INIT_67 => X"000000120000000000000020000000000000002e000000000000002900000000",
            INIT_68 => X"0000002400000000000000230000000000000027000000000000002800000000",
            INIT_69 => X"0000002b00000000000000290000000000000029000000000000002700000000",
            INIT_6A => X"0000003a00000000000000380000000000000033000000000000002e00000000",
            INIT_6B => X"00000037000000000000003c000000000000003d000000000000003d00000000",
            INIT_6C => X"000000360000000000000055000000000000003c000000000000002e00000000",
            INIT_6D => X"000000240000000000000025000000000000002e000000000000002800000000",
            INIT_6E => X"0000002a00000000000000280000000000000026000000000000002600000000",
            INIT_6F => X"00000007000000000000000d0000000000000028000000000000002b00000000",
            INIT_70 => X"0000002800000000000000240000000000000026000000000000002200000000",
            INIT_71 => X"000000330000000000000031000000000000002f000000000000002c00000000",
            INIT_72 => X"00000039000000000000003b0000000000000039000000000000003600000000",
            INIT_73 => X"0000002b00000000000000330000000000000037000000000000003900000000",
            INIT_74 => X"00000032000000000000004e0000000000000030000000000000001f00000000",
            INIT_75 => X"0000002300000000000000230000000000000025000000000000002900000000",
            INIT_76 => X"0000002900000000000000240000000000000025000000000000002500000000",
            INIT_77 => X"0000000700000000000000060000000000000014000000000000002d00000000",
            INIT_78 => X"0000002f000000000000002d000000000000002b000000000000002900000000",
            INIT_79 => X"0000003100000000000000300000000000000030000000000000003000000000",
            INIT_7A => X"0000002d00000000000000310000000000000033000000000000003200000000",
            INIT_7B => X"00000011000000000000001a0000000000000022000000000000002800000000",
            INIT_7C => X"0000002c000000000000003f000000000000001b000000000000000800000000",
            INIT_7D => X"0000002300000000000000220000000000000022000000000000002100000000",
            INIT_7E => X"0000002c00000000000000220000000000000022000000000000002300000000",
            INIT_7F => X"0000000800000000000000050000000000000006000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "sampleifmap_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ba00000000000000c200000000000000da00000000000000de00000000",
            INIT_01 => X"000000f100000000000000ee00000000000000ec00000000000000de00000000",
            INIT_02 => X"000000eb00000000000000f400000000000000f500000000000000f300000000",
            INIT_03 => X"000000f500000000000000f200000000000000f100000000000000f000000000",
            INIT_04 => X"000000f800000000000000f500000000000000f000000000000000e300000000",
            INIT_05 => X"000000f300000000000000f300000000000000f300000000000000f900000000",
            INIT_06 => X"000000f700000000000000ef00000000000000eb00000000000000f500000000",
            INIT_07 => X"000000f600000000000000f300000000000000ea00000000000000f100000000",
            INIT_08 => X"000000b800000000000000c900000000000000e200000000000000e500000000",
            INIT_09 => X"000000ee00000000000000f000000000000000f000000000000000df00000000",
            INIT_0A => X"000000e800000000000000f500000000000000f700000000000000f300000000",
            INIT_0B => X"000000f800000000000000f500000000000000f500000000000000f300000000",
            INIT_0C => X"000000fb00000000000000f300000000000000ef00000000000000e600000000",
            INIT_0D => X"000000f400000000000000ee00000000000000ee00000000000000fb00000000",
            INIT_0E => X"000000fc00000000000000f300000000000000ec00000000000000f800000000",
            INIT_0F => X"000000fb00000000000000fa00000000000000ec00000000000000f000000000",
            INIT_10 => X"000000b500000000000000c700000000000000de00000000000000e100000000",
            INIT_11 => X"000000e400000000000000ef00000000000000ee00000000000000db00000000",
            INIT_12 => X"000000e400000000000000ec00000000000000f400000000000000eb00000000",
            INIT_13 => X"000000f700000000000000ee00000000000000ef00000000000000eb00000000",
            INIT_14 => X"000000f600000000000000f100000000000000ec00000000000000e500000000",
            INIT_15 => X"000000ef00000000000000e800000000000000d700000000000000ec00000000",
            INIT_16 => X"000000fc00000000000000f200000000000000eb00000000000000f800000000",
            INIT_17 => X"000000f700000000000000fb00000000000000e800000000000000f100000000",
            INIT_18 => X"000000b300000000000000c200000000000000d800000000000000de00000000",
            INIT_19 => X"000000e100000000000000eb00000000000000e400000000000000d600000000",
            INIT_1A => X"000000dd00000000000000e600000000000000ef00000000000000e500000000",
            INIT_1B => X"000000f700000000000000e600000000000000ec00000000000000e100000000",
            INIT_1C => X"000000ee00000000000000f000000000000000ea00000000000000e600000000",
            INIT_1D => X"000000f100000000000000e500000000000000b000000000000000ba00000000",
            INIT_1E => X"000000fb00000000000000ef00000000000000e900000000000000f800000000",
            INIT_1F => X"000000f300000000000000f800000000000000e400000000000000ee00000000",
            INIT_20 => X"000000ac00000000000000c100000000000000d900000000000000df00000000",
            INIT_21 => X"000000d900000000000000e700000000000000dd00000000000000d200000000",
            INIT_22 => X"000000d700000000000000e100000000000000eb00000000000000da00000000",
            INIT_23 => X"000000ee00000000000000d600000000000000e800000000000000db00000000",
            INIT_24 => X"000000e400000000000000ee00000000000000e300000000000000e500000000",
            INIT_25 => X"000000ef00000000000000e500000000000000b200000000000000b000000000",
            INIT_26 => X"000000f500000000000000ea00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f000000000000000f600000000000000e800000000000000e700000000",
            INIT_28 => X"000000a400000000000000bf00000000000000d500000000000000dc00000000",
            INIT_29 => X"000000d500000000000000e100000000000000d500000000000000ce00000000",
            INIT_2A => X"000000d600000000000000da00000000000000e600000000000000d600000000",
            INIT_2B => X"000000ce00000000000000c800000000000000e300000000000000d600000000",
            INIT_2C => X"000000cf00000000000000ed00000000000000ce00000000000000d000000000",
            INIT_2D => X"000000e900000000000000e600000000000000ad000000000000008200000000",
            INIT_2E => X"000000e800000000000000db00000000000000e100000000000000f400000000",
            INIT_2F => X"000000e600000000000000f200000000000000e700000000000000dd00000000",
            INIT_30 => X"0000009600000000000000b900000000000000ca00000000000000d400000000",
            INIT_31 => X"000000d000000000000000d900000000000000c900000000000000c400000000",
            INIT_32 => X"000000d300000000000000d000000000000000db00000000000000d300000000",
            INIT_33 => X"000000af00000000000000b900000000000000dd00000000000000d400000000",
            INIT_34 => X"000000c500000000000000d200000000000000bd00000000000000bb00000000",
            INIT_35 => X"000000bb00000000000000b8000000000000009d000000000000008900000000",
            INIT_36 => X"000000da00000000000000ce00000000000000dc00000000000000dd00000000",
            INIT_37 => X"000000d800000000000000e700000000000000db00000000000000d100000000",
            INIT_38 => X"0000009300000000000000b300000000000000c900000000000000d300000000",
            INIT_39 => X"000000cb00000000000000ce00000000000000cc00000000000000c500000000",
            INIT_3A => X"000000cd00000000000000c600000000000000d200000000000000d000000000",
            INIT_3B => X"000000cb00000000000000c000000000000000ce00000000000000ce00000000",
            INIT_3C => X"0000006a000000000000007a000000000000009b00000000000000b300000000",
            INIT_3D => X"000000490000000000000058000000000000005e000000000000006400000000",
            INIT_3E => X"000000d700000000000000ca00000000000000b7000000000000006f00000000",
            INIT_3F => X"000000c100000000000000ce00000000000000b900000000000000c600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c00000000000000a000000000000000ad00000000000000b300000000",
            INIT_41 => X"000000b300000000000000a100000000000000af00000000000000aa00000000",
            INIT_42 => X"000000bd00000000000000b400000000000000b800000000000000bb00000000",
            INIT_43 => X"000000c400000000000000ba00000000000000b900000000000000c300000000",
            INIT_44 => X"0000008000000000000000800000000000000089000000000000009f00000000",
            INIT_45 => X"0000005a0000000000000080000000000000007e000000000000007e00000000",
            INIT_46 => X"000000ac000000000000009e000000000000007c000000000000005800000000",
            INIT_47 => X"0000009f00000000000000b00000000000000089000000000000009c00000000",
            INIT_48 => X"00000070000000000000007b000000000000007e000000000000007b00000000",
            INIT_49 => X"0000008000000000000000720000000000000072000000000000007200000000",
            INIT_4A => X"0000009000000000000000890000000000000086000000000000008600000000",
            INIT_4B => X"000000a700000000000000a00000000000000092000000000000009800000000",
            INIT_4C => X"0000008c0000000000000090000000000000008b000000000000009300000000",
            INIT_4D => X"0000006800000000000000780000000000000083000000000000008200000000",
            INIT_4E => X"0000008d00000000000000960000000000000083000000000000009500000000",
            INIT_4F => X"0000007500000000000000800000000000000069000000000000006a00000000",
            INIT_50 => X"0000005800000000000000620000000000000066000000000000005900000000",
            INIT_51 => X"0000006a00000000000000680000000000000073000000000000006b00000000",
            INIT_52 => X"0000007300000000000000710000000000000076000000000000006b00000000",
            INIT_53 => X"0000009200000000000000970000000000000086000000000000007b00000000",
            INIT_54 => X"00000078000000000000007f000000000000007f000000000000008000000000",
            INIT_55 => X"00000080000000000000007a0000000000000068000000000000006f00000000",
            INIT_56 => X"000000b6000000000000008b000000000000006e000000000000008600000000",
            INIT_57 => X"00000070000000000000006d0000000000000075000000000000007200000000",
            INIT_58 => X"0000006a000000000000006e0000000000000068000000000000005800000000",
            INIT_59 => X"0000005e00000000000000710000000000000089000000000000008e00000000",
            INIT_5A => X"0000007d000000000000007f0000000000000092000000000000007400000000",
            INIT_5B => X"0000009700000000000000a500000000000000a5000000000000009400000000",
            INIT_5C => X"0000007f000000000000007f0000000000000082000000000000008e00000000",
            INIT_5D => X"000000bf00000000000000a50000000000000072000000000000007b00000000",
            INIT_5E => X"000000b80000000000000064000000000000008e00000000000000b400000000",
            INIT_5F => X"0000006c000000000000006c000000000000006d000000000000008c00000000",
            INIT_60 => X"0000006800000000000000840000000000000082000000000000006400000000",
            INIT_61 => X"00000076000000000000006d0000000000000082000000000000008100000000",
            INIT_62 => X"0000009700000000000000a800000000000000ab000000000000009a00000000",
            INIT_63 => X"0000008b000000000000009a00000000000000a5000000000000009b00000000",
            INIT_64 => X"0000008c0000000000000081000000000000007d000000000000008200000000",
            INIT_65 => X"000000c100000000000000b30000000000000089000000000000008600000000",
            INIT_66 => X"00000098000000000000007000000000000000b900000000000000cb00000000",
            INIT_67 => X"0000006d0000000000000069000000000000005400000000000000a000000000",
            INIT_68 => X"0000006a000000000000007e0000000000000086000000000000007800000000",
            INIT_69 => X"00000079000000000000006c0000000000000065000000000000007100000000",
            INIT_6A => X"0000009f00000000000000a10000000000000091000000000000008300000000",
            INIT_6B => X"00000095000000000000009e00000000000000a1000000000000009900000000",
            INIT_6C => X"0000009b00000000000000910000000000000093000000000000009200000000",
            INIT_6D => X"000000b100000000000000b600000000000000a1000000000000009600000000",
            INIT_6E => X"00000076000000000000009400000000000000b500000000000000b500000000",
            INIT_6F => X"00000060000000000000004e0000000000000050000000000000009d00000000",
            INIT_70 => X"00000072000000000000007d0000000000000080000000000000007f00000000",
            INIT_71 => X"0000008600000000000000730000000000000071000000000000007400000000",
            INIT_72 => X"000000b800000000000000b000000000000000a8000000000000009f00000000",
            INIT_73 => X"000000b900000000000000be00000000000000bf00000000000000be00000000",
            INIT_74 => X"000000b800000000000000be00000000000000c400000000000000c500000000",
            INIT_75 => X"000000a800000000000000af00000000000000ad00000000000000ac00000000",
            INIT_76 => X"0000006300000000000000a300000000000000a500000000000000ab00000000",
            INIT_77 => X"0000005100000000000000430000000000000047000000000000005700000000",
            INIT_78 => X"00000091000000000000009a0000000000000095000000000000009700000000",
            INIT_79 => X"000000c100000000000000b800000000000000b3000000000000009900000000",
            INIT_7A => X"000000d000000000000000cf00000000000000cd00000000000000c900000000",
            INIT_7B => X"000000c800000000000000d400000000000000d200000000000000d100000000",
            INIT_7C => X"000000ab00000000000000c300000000000000c900000000000000c600000000",
            INIT_7D => X"0000009b000000000000008b0000000000000087000000000000008600000000",
            INIT_7E => X"0000007100000000000000a800000000000000a100000000000000a500000000",
            INIT_7F => X"00000056000000000000005a000000000000005c000000000000004900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "sampleifmap_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b000000000000000a7000000000000009f00000000000000a500000000",
            INIT_01 => X"000000c900000000000000c600000000000000b900000000000000af00000000",
            INIT_02 => X"000000d200000000000000d200000000000000d000000000000000cd00000000",
            INIT_03 => X"000000be00000000000000c900000000000000d000000000000000d200000000",
            INIT_04 => X"0000009400000000000000a900000000000000aa00000000000000aa00000000",
            INIT_05 => X"00000099000000000000008e000000000000007a000000000000006c00000000",
            INIT_06 => X"0000008e00000000000000a700000000000000a500000000000000a700000000",
            INIT_07 => X"0000006f000000000000009800000000000000b5000000000000009300000000",
            INIT_08 => X"0000009d00000000000000ae00000000000000aa000000000000009d00000000",
            INIT_09 => X"000000ca00000000000000b6000000000000008f000000000000008d00000000",
            INIT_0A => X"000000ca00000000000000d100000000000000d300000000000000d000000000",
            INIT_0B => X"000000a200000000000000a700000000000000b500000000000000bf00000000",
            INIT_0C => X"000000a900000000000000b200000000000000a0000000000000009b00000000",
            INIT_0D => X"000000a000000000000000a7000000000000009d000000000000009300000000",
            INIT_0E => X"0000009c00000000000000a100000000000000a200000000000000a900000000",
            INIT_0F => X"0000009400000000000000960000000000000096000000000000009e00000000",
            INIT_10 => X"000000790000000000000080000000000000009400000000000000a200000000",
            INIT_11 => X"000000c200000000000000b100000000000000a4000000000000008a00000000",
            INIT_12 => X"000000ab00000000000000b200000000000000bc00000000000000c700000000",
            INIT_13 => X"000000b000000000000000ac00000000000000ac00000000000000aa00000000",
            INIT_14 => X"000000b500000000000000b000000000000000a800000000000000b400000000",
            INIT_15 => X"000000ac00000000000000af00000000000000ad00000000000000aa00000000",
            INIT_16 => X"0000009600000000000000a300000000000000a500000000000000a800000000",
            INIT_17 => X"00000099000000000000007d0000000000000076000000000000008500000000",
            INIT_18 => X"000000a6000000000000007f0000000000000075000000000000008f00000000",
            INIT_19 => X"000000b000000000000000ba00000000000000c500000000000000bc00000000",
            INIT_1A => X"000000b200000000000000ab00000000000000a300000000000000a900000000",
            INIT_1B => X"000000ba00000000000000bf00000000000000be00000000000000b900000000",
            INIT_1C => X"000000b100000000000000ac00000000000000a500000000000000b400000000",
            INIT_1D => X"000000b200000000000000af00000000000000ac00000000000000ad00000000",
            INIT_1E => X"000000740000000000000088000000000000009c00000000000000a400000000",
            INIT_1F => X"0000009000000000000000620000000000000057000000000000006700000000",
            INIT_20 => X"000000b000000000000000a800000000000000a500000000000000a600000000",
            INIT_21 => X"000000aa00000000000000b300000000000000ae00000000000000b000000000",
            INIT_22 => X"000000bd00000000000000be00000000000000b800000000000000a400000000",
            INIT_23 => X"0000009600000000000000a800000000000000b500000000000000b900000000",
            INIT_24 => X"000000ad000000000000009d0000000000000076000000000000008100000000",
            INIT_25 => X"000000a200000000000000ab00000000000000ad00000000000000ad00000000",
            INIT_26 => X"0000005f000000000000006a0000000000000070000000000000008500000000",
            INIT_27 => X"0000004e00000000000000560000000000000054000000000000005000000000",
            INIT_28 => X"000000af00000000000000b100000000000000ac00000000000000a500000000",
            INIT_29 => X"000000b000000000000000b300000000000000b000000000000000ae00000000",
            INIT_2A => X"000000ad00000000000000ab00000000000000ab00000000000000a400000000",
            INIT_2B => X"0000005e000000000000007e00000000000000ab00000000000000af00000000",
            INIT_2C => X"000000ac000000000000008e0000000000000055000000000000005800000000",
            INIT_2D => X"000000750000000000000088000000000000009800000000000000a200000000",
            INIT_2E => X"00000050000000000000005e0000000000000068000000000000006c00000000",
            INIT_2F => X"00000027000000000000003f0000000000000058000000000000004f00000000",
            INIT_30 => X"000000af00000000000000b200000000000000a6000000000000007c00000000",
            INIT_31 => X"0000008b000000000000009a00000000000000ad00000000000000af00000000",
            INIT_32 => X"0000009a000000000000007a000000000000007e000000000000008200000000",
            INIT_33 => X"0000006c000000000000008300000000000000a900000000000000ae00000000",
            INIT_34 => X"0000008500000000000000860000000000000072000000000000007200000000",
            INIT_35 => X"0000006c000000000000006d0000000000000071000000000000007900000000",
            INIT_36 => X"00000045000000000000004b0000000000000056000000000000005f00000000",
            INIT_37 => X"00000026000000000000002b000000000000003b000000000000004900000000",
            INIT_38 => X"0000009f00000000000000a00000000000000096000000000000006f00000000",
            INIT_39 => X"000000640000000000000074000000000000009e00000000000000a300000000",
            INIT_3A => X"0000009700000000000000730000000000000070000000000000006800000000",
            INIT_3B => X"00000083000000000000009500000000000000a800000000000000ac00000000",
            INIT_3C => X"0000006a000000000000006a000000000000006b000000000000007700000000",
            INIT_3D => X"000000540000000000000064000000000000006c000000000000006a00000000",
            INIT_3E => X"0000004100000000000000440000000000000049000000000000004500000000",
            INIT_3F => X"000000250000000000000028000000000000002c000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009a0000000000000097000000000000008a000000000000007100000000",
            INIT_41 => X"00000077000000000000008000000000000000a200000000000000a100000000",
            INIT_42 => X"0000009200000000000000900000000000000088000000000000008100000000",
            INIT_43 => X"0000006200000000000000650000000000000072000000000000008400000000",
            INIT_44 => X"0000006c000000000000006d0000000000000067000000000000006500000000",
            INIT_45 => X"0000004b00000000000000480000000000000050000000000000006300000000",
            INIT_46 => X"0000003a000000000000003d000000000000004d000000000000005500000000",
            INIT_47 => X"000000270000000000000029000000000000002d000000000000003400000000",
            INIT_48 => X"00000097000000000000009a0000000000000088000000000000007400000000",
            INIT_49 => X"0000007c0000000000000084000000000000008f000000000000009400000000",
            INIT_4A => X"00000057000000000000005b0000000000000067000000000000007600000000",
            INIT_4B => X"000000650000000000000063000000000000005b000000000000005600000000",
            INIT_4C => X"00000052000000000000005e0000000000000063000000000000006500000000",
            INIT_4D => X"00000045000000000000004a0000000000000048000000000000004800000000",
            INIT_4E => X"0000003200000000000000340000000000000044000000000000004e00000000",
            INIT_4F => X"00000030000000000000002f0000000000000030000000000000003300000000",
            INIT_50 => X"00000063000000000000006a0000000000000064000000000000006000000000",
            INIT_51 => X"0000005100000000000000520000000000000056000000000000005c00000000",
            INIT_52 => X"000000540000000000000051000000000000004f000000000000005200000000",
            INIT_53 => X"00000058000000000000005e000000000000005b000000000000005700000000",
            INIT_54 => X"0000004c00000000000000440000000000000044000000000000004d00000000",
            INIT_55 => X"0000003b00000000000000400000000000000048000000000000004a00000000",
            INIT_56 => X"0000003200000000000000310000000000000036000000000000003f00000000",
            INIT_57 => X"0000003000000000000000340000000000000030000000000000003100000000",
            INIT_58 => X"0000003700000000000000360000000000000039000000000000003b00000000",
            INIT_59 => X"00000044000000000000003e000000000000003d000000000000003c00000000",
            INIT_5A => X"0000004d000000000000004f000000000000004f000000000000004e00000000",
            INIT_5B => X"0000004200000000000000450000000000000044000000000000004800000000",
            INIT_5C => X"0000005200000000000000610000000000000047000000000000003d00000000",
            INIT_5D => X"000000390000000000000038000000000000003c000000000000004100000000",
            INIT_5E => X"0000003100000000000000300000000000000031000000000000003500000000",
            INIT_5F => X"0000002300000000000000320000000000000032000000000000003200000000",
            INIT_60 => X"0000002d000000000000002c0000000000000030000000000000003200000000",
            INIT_61 => X"0000003700000000000000350000000000000035000000000000003100000000",
            INIT_62 => X"000000380000000000000038000000000000003b000000000000003a00000000",
            INIT_63 => X"0000004400000000000000470000000000000042000000000000003c00000000",
            INIT_64 => X"0000004b0000000000000068000000000000004b000000000000003b00000000",
            INIT_65 => X"00000033000000000000003a0000000000000038000000000000003500000000",
            INIT_66 => X"0000003300000000000000310000000000000030000000000000003100000000",
            INIT_67 => X"0000001400000000000000250000000000000035000000000000003200000000",
            INIT_68 => X"000000290000000000000028000000000000002c000000000000002d00000000",
            INIT_69 => X"00000030000000000000002e000000000000002e000000000000002c00000000",
            INIT_6A => X"00000041000000000000003f0000000000000039000000000000003300000000",
            INIT_6B => X"0000003d00000000000000440000000000000044000000000000004400000000",
            INIT_6C => X"0000003f000000000000005d0000000000000042000000000000003200000000",
            INIT_6D => X"0000002f00000000000000300000000000000038000000000000003100000000",
            INIT_6E => X"000000330000000000000031000000000000002f000000000000002f00000000",
            INIT_6F => X"00000005000000000000000e000000000000002e000000000000003400000000",
            INIT_70 => X"0000002d0000000000000029000000000000002b000000000000002700000000",
            INIT_71 => X"0000003b00000000000000380000000000000036000000000000003200000000",
            INIT_72 => X"0000004000000000000000420000000000000040000000000000003e00000000",
            INIT_73 => X"00000031000000000000003a000000000000003d000000000000004000000000",
            INIT_74 => X"0000003b00000000000000550000000000000035000000000000002400000000",
            INIT_75 => X"0000002f000000000000002f0000000000000030000000000000003200000000",
            INIT_76 => X"00000032000000000000002d000000000000002e000000000000002e00000000",
            INIT_77 => X"0000000300000000000000030000000000000018000000000000003600000000",
            INIT_78 => X"0000003600000000000000340000000000000032000000000000002f00000000",
            INIT_79 => X"0000003a00000000000000380000000000000038000000000000003800000000",
            INIT_7A => X"0000003200000000000000350000000000000037000000000000003a00000000",
            INIT_7B => X"00000014000000000000001e0000000000000027000000000000002d00000000",
            INIT_7C => X"0000003600000000000000480000000000000021000000000000000b00000000",
            INIT_7D => X"0000002e000000000000002d000000000000002d000000000000002c00000000",
            INIT_7E => X"00000034000000000000002b000000000000002c000000000000002c00000000",
            INIT_7F => X"0000000700000000000000030000000000000008000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "sampleifmap_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000be00000000000000b000000000000000a7000000000000009b00000000",
            INIT_01 => X"000000a600000000000000a800000000000000a600000000000000b100000000",
            INIT_02 => X"000000bb00000000000000bb00000000000000b300000000000000aa00000000",
            INIT_03 => X"000000b800000000000000b800000000000000bb00000000000000bb00000000",
            INIT_04 => X"000000ba00000000000000b800000000000000b400000000000000b600000000",
            INIT_05 => X"000000bd00000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000c000000000000000ca00000000000000c900000000000000c900000000",
            INIT_08 => X"000000bb00000000000000ab00000000000000a3000000000000009900000000",
            INIT_09 => X"0000009f000000000000009a000000000000009b00000000000000b300000000",
            INIT_0A => X"000000af00000000000000ab00000000000000a5000000000000009f00000000",
            INIT_0B => X"000000a500000000000000a200000000000000ab00000000000000a900000000",
            INIT_0C => X"000000a500000000000000a600000000000000a400000000000000aa00000000",
            INIT_0D => X"000000a800000000000000a900000000000000ad00000000000000a700000000",
            INIT_0E => X"000000ca00000000000000be00000000000000ad00000000000000a900000000",
            INIT_0F => X"000000bd00000000000000cb00000000000000ca00000000000000cc00000000",
            INIT_10 => X"000000b800000000000000a800000000000000a0000000000000009b00000000",
            INIT_11 => X"000000bc00000000000000b000000000000000ae00000000000000bb00000000",
            INIT_12 => X"000000be00000000000000b100000000000000b300000000000000b600000000",
            INIT_13 => X"000000b900000000000000bc00000000000000c200000000000000c000000000",
            INIT_14 => X"000000c200000000000000c100000000000000c200000000000000c100000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c500000000000000c300000000",
            INIT_16 => X"000000cf00000000000000ce00000000000000c500000000000000bf00000000",
            INIT_17 => X"000000bd00000000000000cc00000000000000ce00000000000000d000000000",
            INIT_18 => X"000000b100000000000000a6000000000000009d000000000000009700000000",
            INIT_19 => X"000000c500000000000000c700000000000000b900000000000000b400000000",
            INIT_1A => X"000000c600000000000000cd00000000000000cc00000000000000b600000000",
            INIT_1B => X"000000cb00000000000000c400000000000000c500000000000000d200000000",
            INIT_1C => X"000000cb00000000000000d200000000000000cf00000000000000cd00000000",
            INIT_1D => X"000000cc00000000000000c500000000000000d200000000000000cf00000000",
            INIT_1E => X"000000c900000000000000cc00000000000000c600000000000000d000000000",
            INIT_1F => X"000000c000000000000000ce00000000000000cf00000000000000d100000000",
            INIT_20 => X"000000ae00000000000000a8000000000000009e000000000000009700000000",
            INIT_21 => X"000000c400000000000000bf00000000000000b500000000000000b100000000",
            INIT_22 => X"000000b900000000000000bd00000000000000c200000000000000b700000000",
            INIT_23 => X"000000ca00000000000000b900000000000000b900000000000000c400000000",
            INIT_24 => X"000000c000000000000000c800000000000000c700000000000000c700000000",
            INIT_25 => X"000000bc00000000000000be00000000000000c700000000000000c300000000",
            INIT_26 => X"000000c400000000000000c900000000000000c700000000000000c900000000",
            INIT_27 => X"000000c400000000000000cf00000000000000cc00000000000000ce00000000",
            INIT_28 => X"000000ae00000000000000a7000000000000009c000000000000009400000000",
            INIT_29 => X"000000c300000000000000c400000000000000ae00000000000000ab00000000",
            INIT_2A => X"000000b800000000000000bd00000000000000be00000000000000c000000000",
            INIT_2B => X"000000bf00000000000000bd00000000000000bd00000000000000bb00000000",
            INIT_2C => X"000000c600000000000000bb00000000000000c300000000000000be00000000",
            INIT_2D => X"000000c100000000000000c000000000000000bc00000000000000c000000000",
            INIT_2E => X"000000d100000000000000cb00000000000000ce00000000000000cd00000000",
            INIT_2F => X"000000c400000000000000d100000000000000d000000000000000d400000000",
            INIT_30 => X"000000ae00000000000000a50000000000000099000000000000009400000000",
            INIT_31 => X"000000c300000000000000cb00000000000000b000000000000000a800000000",
            INIT_32 => X"000000be00000000000000bb00000000000000bc00000000000000bc00000000",
            INIT_33 => X"000000c300000000000000c500000000000000c200000000000000b600000000",
            INIT_34 => X"000000cd00000000000000c800000000000000c100000000000000c400000000",
            INIT_35 => X"000000c900000000000000c500000000000000c500000000000000c600000000",
            INIT_36 => X"000000c300000000000000c600000000000000c800000000000000c500000000",
            INIT_37 => X"000000c300000000000000cf00000000000000cb00000000000000c500000000",
            INIT_38 => X"000000ac00000000000000a3000000000000009b000000000000009900000000",
            INIT_39 => X"000000d100000000000000c700000000000000bc00000000000000ac00000000",
            INIT_3A => X"000000bf00000000000000bd00000000000000be00000000000000c400000000",
            INIT_3B => X"000000c400000000000000bb00000000000000bc00000000000000c100000000",
            INIT_3C => X"000000ce00000000000000c400000000000000c200000000000000ca00000000",
            INIT_3D => X"000000c800000000000000c400000000000000c900000000000000c200000000",
            INIT_3E => X"000000c900000000000000c800000000000000bb00000000000000b500000000",
            INIT_3F => X"000000bd00000000000000c700000000000000c400000000000000c800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac00000000000000a3000000000000009f00000000000000a000000000",
            INIT_41 => X"000000be00000000000000b000000000000000b000000000000000ae00000000",
            INIT_42 => X"000000b000000000000000b000000000000000af00000000000000b400000000",
            INIT_43 => X"000000b600000000000000ac00000000000000aa00000000000000b500000000",
            INIT_44 => X"000000bb00000000000000b500000000000000b200000000000000bb00000000",
            INIT_45 => X"000000bb00000000000000b400000000000000bc00000000000000b100000000",
            INIT_46 => X"000000bc00000000000000bc00000000000000c400000000000000c700000000",
            INIT_47 => X"000000b800000000000000c200000000000000c000000000000000c500000000",
            INIT_48 => X"000000ac00000000000000a200000000000000a700000000000000ab00000000",
            INIT_49 => X"000000b000000000000000b400000000000000ab00000000000000aa00000000",
            INIT_4A => X"0000009c0000000000000096000000000000009c000000000000009b00000000",
            INIT_4B => X"0000009e00000000000000990000000000000092000000000000009600000000",
            INIT_4C => X"0000009d00000000000000a400000000000000a600000000000000a600000000",
            INIT_4D => X"000000a6000000000000009c00000000000000a2000000000000009d00000000",
            INIT_4E => X"000000bd00000000000000bc00000000000000c700000000000000c800000000",
            INIT_4F => X"000000b600000000000000c200000000000000c100000000000000c500000000",
            INIT_50 => X"000000b000000000000000a800000000000000b400000000000000af00000000",
            INIT_51 => X"000000ae00000000000000b600000000000000b100000000000000ad00000000",
            INIT_52 => X"0000009a000000000000009f00000000000000a0000000000000009c00000000",
            INIT_53 => X"000000ad00000000000000a800000000000000a3000000000000009f00000000",
            INIT_54 => X"000000a200000000000000a000000000000000a400000000000000aa00000000",
            INIT_55 => X"000000ac00000000000000a700000000000000a800000000000000a000000000",
            INIT_56 => X"000000c400000000000000c400000000000000c300000000000000c200000000",
            INIT_57 => X"000000b700000000000000c100000000000000bf00000000000000c500000000",
            INIT_58 => X"000000bb00000000000000b200000000000000bb00000000000000b500000000",
            INIT_59 => X"000000b600000000000000ae00000000000000aa00000000000000b700000000",
            INIT_5A => X"000000b500000000000000b400000000000000b300000000000000b300000000",
            INIT_5B => X"000000c100000000000000c100000000000000bb00000000000000b800000000",
            INIT_5C => X"000000b900000000000000bc00000000000000c000000000000000c100000000",
            INIT_5D => X"000000c000000000000000c000000000000000ba00000000000000b800000000",
            INIT_5E => X"000000bd00000000000000c000000000000000bc00000000000000bb00000000",
            INIT_5F => X"000000ba00000000000000c400000000000000bf00000000000000be00000000",
            INIT_60 => X"000000ab00000000000000ba00000000000000be00000000000000b900000000",
            INIT_61 => X"000000c100000000000000950000000000000084000000000000009900000000",
            INIT_62 => X"000000bc00000000000000ba00000000000000bf00000000000000c600000000",
            INIT_63 => X"000000c400000000000000c300000000000000c100000000000000bf00000000",
            INIT_64 => X"000000bc00000000000000be00000000000000c000000000000000c300000000",
            INIT_65 => X"000000bf00000000000000c000000000000000be00000000000000bc00000000",
            INIT_66 => X"000000c500000000000000c300000000000000c100000000000000bf00000000",
            INIT_67 => X"000000c100000000000000cc00000000000000ca00000000000000ca00000000",
            INIT_68 => X"0000009e00000000000000bc00000000000000c200000000000000ba00000000",
            INIT_69 => X"0000006d000000000000005e0000000000000074000000000000008400000000",
            INIT_6A => X"000000c200000000000000c200000000000000b1000000000000009100000000",
            INIT_6B => X"000000c700000000000000c400000000000000c100000000000000bf00000000",
            INIT_6C => X"000000c600000000000000c800000000000000c700000000000000c700000000",
            INIT_6D => X"000000c600000000000000c700000000000000c400000000000000c400000000",
            INIT_6E => X"000000c400000000000000c400000000000000c400000000000000c500000000",
            INIT_6F => X"000000b900000000000000c600000000000000c500000000000000c600000000",
            INIT_70 => X"000000c600000000000000c400000000000000c500000000000000ba00000000",
            INIT_71 => X"0000005c000000000000008d00000000000000b800000000000000c200000000",
            INIT_72 => X"000000b3000000000000008e0000000000000068000000000000005400000000",
            INIT_73 => X"000000cc00000000000000cc00000000000000c900000000000000c300000000",
            INIT_74 => X"000000c700000000000000cc00000000000000cc00000000000000cc00000000",
            INIT_75 => X"000000bf00000000000000c200000000000000c200000000000000c200000000",
            INIT_76 => X"000000be00000000000000be00000000000000be00000000000000bd00000000",
            INIT_77 => X"000000b500000000000000c000000000000000be00000000000000bf00000000",
            INIT_78 => X"000000c800000000000000c600000000000000c700000000000000b800000000",
            INIT_79 => X"000000b100000000000000c900000000000000c800000000000000c500000000",
            INIT_7A => X"00000080000000000000005d0000000000000054000000000000007500000000",
            INIT_7B => X"000000cd00000000000000d000000000000000ca00000000000000ad00000000",
            INIT_7C => X"000000c700000000000000c700000000000000c800000000000000ca00000000",
            INIT_7D => X"000000c300000000000000c500000000000000c400000000000000c300000000",
            INIT_7E => X"000000bf00000000000000c200000000000000c300000000000000c100000000",
            INIT_7F => X"000000b200000000000000be00000000000000bd00000000000000bf00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "sampleifmap_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d000000000000000cb00000000000000c900000000000000b900000000",
            INIT_01 => X"000000d600000000000000d000000000000000ce00000000000000cd00000000",
            INIT_02 => X"0000005b000000000000004c000000000000005c00000000000000af00000000",
            INIT_03 => X"000000cb00000000000000b5000000000000008c000000000000006900000000",
            INIT_04 => X"000000c200000000000000c500000000000000ca00000000000000ce00000000",
            INIT_05 => X"000000c200000000000000c200000000000000c200000000000000c100000000",
            INIT_06 => X"000000bf00000000000000c100000000000000c300000000000000c200000000",
            INIT_07 => X"000000b400000000000000be00000000000000be00000000000000c100000000",
            INIT_08 => X"000000d600000000000000cf00000000000000cc00000000000000bb00000000",
            INIT_09 => X"000000d000000000000000d300000000000000d400000000000000d400000000",
            INIT_0A => X"000000570000000000000047000000000000007c00000000000000cb00000000",
            INIT_0B => X"0000008400000000000000630000000000000054000000000000005400000000",
            INIT_0C => X"000000cb00000000000000cb00000000000000be00000000000000a700000000",
            INIT_0D => X"000000c400000000000000c500000000000000c000000000000000c300000000",
            INIT_0E => X"000000bf00000000000000c000000000000000c200000000000000c200000000",
            INIT_0F => X"000000b700000000000000c000000000000000bf00000000000000c100000000",
            INIT_10 => X"000000d600000000000000cf00000000000000cf00000000000000be00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000d400000000",
            INIT_12 => X"000000570000000000000048000000000000008900000000000000d300000000",
            INIT_13 => X"0000005300000000000000560000000000000054000000000000005300000000",
            INIT_14 => X"0000009b0000000000000083000000000000006b000000000000005900000000",
            INIT_15 => X"000000cc00000000000000cb00000000000000b600000000000000a300000000",
            INIT_16 => X"000000bf00000000000000c200000000000000c600000000000000ca00000000",
            INIT_17 => X"000000b600000000000000bf00000000000000c000000000000000c100000000",
            INIT_18 => X"000000d700000000000000d100000000000000d200000000000000bf00000000",
            INIT_19 => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1A => X"0000003a000000000000002f000000000000007100000000000000cc00000000",
            INIT_1B => X"0000005d0000000000000057000000000000004c000000000000003f00000000",
            INIT_1C => X"0000003e00000000000000460000000000000050000000000000005a00000000",
            INIT_1D => X"0000009f000000000000007a000000000000004d000000000000003a00000000",
            INIT_1E => X"000000c800000000000000c900000000000000c200000000000000b400000000",
            INIT_1F => X"000000b900000000000000c400000000000000c400000000000000c800000000",
            INIT_20 => X"000000d300000000000000cf00000000000000d000000000000000bf00000000",
            INIT_21 => X"000000d400000000000000d100000000000000d200000000000000d100000000",
            INIT_22 => X"0000002500000000000000410000000000000065000000000000009d00000000",
            INIT_23 => X"00000058000000000000004a0000000000000044000000000000003300000000",
            INIT_24 => X"0000004900000000000000550000000000000056000000000000005b00000000",
            INIT_25 => X"00000048000000000000003e000000000000002e000000000000003700000000",
            INIT_26 => X"0000009e0000000000000085000000000000006b000000000000004e00000000",
            INIT_27 => X"000000ba00000000000000c400000000000000c300000000000000b800000000",
            INIT_28 => X"000000d100000000000000cb00000000000000ca00000000000000ba00000000",
            INIT_29 => X"000000c800000000000000d100000000000000ce00000000000000cf00000000",
            INIT_2A => X"000000640000000000000097000000000000008c000000000000009500000000",
            INIT_2B => X"0000006000000000000000320000000000000035000000000000002d00000000",
            INIT_2C => X"00000048000000000000008000000000000000a0000000000000009c00000000",
            INIT_2D => X"0000004200000000000000590000000000000070000000000000006200000000",
            INIT_2E => X"000000a300000000000000a60000000000000083000000000000004300000000",
            INIT_2F => X"000000b200000000000000bc00000000000000b700000000000000ad00000000",
            INIT_30 => X"000000d200000000000000ca00000000000000c900000000000000b900000000",
            INIT_31 => X"000000d100000000000000d100000000000000d000000000000000d200000000",
            INIT_32 => X"000000bd00000000000000d700000000000000d300000000000000d200000000",
            INIT_33 => X"000000a800000000000000940000000000000092000000000000009000000000",
            INIT_34 => X"0000009a00000000000000c000000000000000ce00000000000000ca00000000",
            INIT_35 => X"0000009f00000000000000b100000000000000b200000000000000a300000000",
            INIT_36 => X"000000c200000000000000bf00000000000000b2000000000000009c00000000",
            INIT_37 => X"000000b000000000000000bc00000000000000c100000000000000c400000000",
            INIT_38 => X"000000c400000000000000c000000000000000bc00000000000000b000000000",
            INIT_39 => X"000000b700000000000000b900000000000000bc00000000000000c000000000",
            INIT_3A => X"000000ad00000000000000b300000000000000b200000000000000b600000000",
            INIT_3B => X"000000ad00000000000000ab00000000000000aa00000000000000aa00000000",
            INIT_3C => X"000000a700000000000000a100000000000000a000000000000000a900000000",
            INIT_3D => X"000000aa00000000000000a500000000000000a100000000000000a500000000",
            INIT_3E => X"00000096000000000000009800000000000000a000000000000000aa00000000",
            INIT_3F => X"0000009c00000000000000a400000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006b000000000000006e0000000000000063000000000000007200000000",
            INIT_41 => X"0000005d000000000000005e0000000000000061000000000000006600000000",
            INIT_42 => X"0000005000000000000000580000000000000055000000000000005800000000",
            INIT_43 => X"000000650000000000000053000000000000004e000000000000004d00000000",
            INIT_44 => X"0000006b000000000000006a000000000000006c000000000000007100000000",
            INIT_45 => X"00000071000000000000006f000000000000006e000000000000006c00000000",
            INIT_46 => X"0000007700000000000000780000000000000077000000000000007500000000",
            INIT_47 => X"0000007c000000000000007a0000000000000079000000000000007800000000",
            INIT_48 => X"000000750000000000000071000000000000006d000000000000007a00000000",
            INIT_49 => X"0000007100000000000000720000000000000070000000000000007300000000",
            INIT_4A => X"0000006d000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006c000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006b00000000000000690000000000000070000000000000007300000000",
            INIT_4D => X"000000680000000000000065000000000000006a000000000000006c00000000",
            INIT_4E => X"0000006d000000000000006d000000000000006b000000000000006a00000000",
            INIT_4F => X"00000065000000000000005e0000000000000066000000000000006700000000",
            INIT_50 => X"00000070000000000000006b0000000000000061000000000000007800000000",
            INIT_51 => X"0000005e00000000000000620000000000000068000000000000006d00000000",
            INIT_52 => X"000000560000000000000058000000000000005d000000000000005e00000000",
            INIT_53 => X"0000004e0000000000000050000000000000004f000000000000005200000000",
            INIT_54 => X"000000450000000000000048000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000042000000000000004300000000",
            INIT_56 => X"0000004000000000000000420000000000000041000000000000004000000000",
            INIT_57 => X"0000004d0000000000000035000000000000003f000000000000004300000000",
            INIT_58 => X"0000004500000000000000410000000000000037000000000000005b00000000",
            INIT_59 => X"0000003d000000000000003f0000000000000042000000000000004200000000",
            INIT_5A => X"00000039000000000000003c0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003a00000000000000400000000000000042000000000000003f00000000",
            INIT_5D => X"0000003c000000000000003b0000000000000039000000000000003800000000",
            INIT_5E => X"0000003900000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000005c000000000000004b0000000000000031000000000000003400000000",
            INIT_60 => X"000000440000000000000042000000000000003c000000000000005d00000000",
            INIT_61 => X"0000004100000000000000400000000000000043000000000000004300000000",
            INIT_62 => X"0000003b000000000000003e0000000000000041000000000000004500000000",
            INIT_63 => X"0000003d000000000000003c000000000000003b000000000000003b00000000",
            INIT_64 => X"00000038000000000000003a000000000000003f000000000000004000000000",
            INIT_65 => X"0000003800000000000000380000000000000037000000000000003700000000",
            INIT_66 => X"000000350000000000000038000000000000003a000000000000003900000000",
            INIT_67 => X"000000510000000000000061000000000000005d000000000000004100000000",
            INIT_68 => X"00000039000000000000003d0000000000000039000000000000005900000000",
            INIT_69 => X"0000003b0000000000000039000000000000003b000000000000003900000000",
            INIT_6A => X"000000360000000000000038000000000000003a000000000000003c00000000",
            INIT_6B => X"0000003d000000000000003b000000000000003d000000000000003c00000000",
            INIT_6C => X"00000039000000000000003a000000000000003d000000000000004100000000",
            INIT_6D => X"0000003d000000000000003d000000000000003c000000000000003c00000000",
            INIT_6E => X"000000460000000000000039000000000000003e000000000000004200000000",
            INIT_6F => X"00000043000000000000003b0000000000000059000000000000006100000000",
            INIT_70 => X"0000003e000000000000003f000000000000003c000000000000005900000000",
            INIT_71 => X"0000003f000000000000003e000000000000003e000000000000003e00000000",
            INIT_72 => X"000000520000000000000041000000000000003d000000000000003e00000000",
            INIT_73 => X"00000051000000000000004e0000000000000051000000000000005400000000",
            INIT_74 => X"0000005300000000000000550000000000000054000000000000005800000000",
            INIT_75 => X"0000004000000000000000420000000000000043000000000000005000000000",
            INIT_76 => X"0000006700000000000000560000000000000038000000000000003400000000",
            INIT_77 => X"0000004b000000000000003d0000000000000039000000000000004c00000000",
            INIT_78 => X"0000003c000000000000003d000000000000003c000000000000005c00000000",
            INIT_79 => X"0000004100000000000000430000000000000042000000000000003f00000000",
            INIT_7A => X"0000004800000000000000410000000000000043000000000000004200000000",
            INIT_7B => X"0000004600000000000000480000000000000049000000000000004900000000",
            INIT_7C => X"0000004b000000000000004b000000000000004a000000000000004900000000",
            INIT_7D => X"0000003e00000000000000400000000000000040000000000000004b00000000",
            INIT_7E => X"0000004000000000000000580000000000000056000000000000004100000000",
            INIT_7F => X"000000490000000000000040000000000000003c000000000000003900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "sampleifmap_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c000000000000000b300000000000000b0000000000000009c00000000",
            INIT_01 => X"000000ad00000000000000ad00000000000000ab00000000000000b900000000",
            INIT_02 => X"000000b800000000000000b600000000000000b300000000000000af00000000",
            INIT_03 => X"000000b500000000000000b600000000000000b800000000000000b900000000",
            INIT_04 => X"000000b900000000000000b700000000000000b300000000000000b300000000",
            INIT_05 => X"000000bd00000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000b700000000000000ca00000000000000c400000000000000c500000000",
            INIT_08 => X"000000c300000000000000b800000000000000b3000000000000009b00000000",
            INIT_09 => X"000000a4000000000000009f00000000000000a200000000000000be00000000",
            INIT_0A => X"000000b000000000000000a900000000000000a500000000000000a300000000",
            INIT_0B => X"000000a700000000000000a400000000000000ae00000000000000ab00000000",
            INIT_0C => X"000000a600000000000000a800000000000000a600000000000000ac00000000",
            INIT_0D => X"000000a900000000000000ab00000000000000af00000000000000a900000000",
            INIT_0E => X"000000cc00000000000000bf00000000000000ae00000000000000aa00000000",
            INIT_0F => X"000000be00000000000000d700000000000000d000000000000000ce00000000",
            INIT_10 => X"000000c400000000000000b900000000000000b2000000000000009a00000000",
            INIT_11 => X"000000a800000000000000b200000000000000c100000000000000cb00000000",
            INIT_12 => X"000000c400000000000000be00000000000000af00000000000000a000000000",
            INIT_13 => X"000000bc00000000000000be00000000000000c500000000000000c300000000",
            INIT_14 => X"000000c300000000000000c200000000000000c300000000000000c400000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c600000000000000c400000000",
            INIT_16 => X"000000cd00000000000000cd00000000000000c400000000000000c000000000",
            INIT_17 => X"000000bf00000000000000d700000000000000d000000000000000ce00000000",
            INIT_18 => X"000000c300000000000000bc00000000000000b2000000000000009a00000000",
            INIT_19 => X"0000008000000000000000bc00000000000000c500000000000000ca00000000",
            INIT_1A => X"0000009b000000000000009a0000000000000098000000000000006c00000000",
            INIT_1B => X"0000009400000000000000950000000000000095000000000000009e00000000",
            INIT_1C => X"000000ad00000000000000a300000000000000a100000000000000a700000000",
            INIT_1D => X"0000009f00000000000000ae00000000000000a300000000000000a800000000",
            INIT_1E => X"000000ce00000000000000cc00000000000000d000000000000000bc00000000",
            INIT_1F => X"000000bc00000000000000d400000000000000cd00000000000000cc00000000",
            INIT_20 => X"000000bf00000000000000bb00000000000000b1000000000000009a00000000",
            INIT_21 => X"0000007e00000000000000bd00000000000000c400000000000000c600000000",
            INIT_22 => X"0000006b000000000000006a000000000000008b000000000000008000000000",
            INIT_23 => X"0000007100000000000000760000000000000078000000000000007300000000",
            INIT_24 => X"0000007e00000000000000720000000000000072000000000000007700000000",
            INIT_25 => X"0000007000000000000000880000000000000070000000000000007600000000",
            INIT_26 => X"000000ce00000000000000c900000000000000cb00000000000000a000000000",
            INIT_27 => X"000000be00000000000000d600000000000000cd00000000000000ce00000000",
            INIT_28 => X"000000bd00000000000000bb00000000000000ae000000000000009700000000",
            INIT_29 => X"0000009300000000000000b700000000000000c800000000000000c500000000",
            INIT_2A => X"000000a5000000000000009100000000000000a800000000000000a900000000",
            INIT_2B => X"0000009d0000000000000095000000000000009200000000000000aa00000000",
            INIT_2C => X"000000bd00000000000000b000000000000000b200000000000000b400000000",
            INIT_2D => X"000000b100000000000000bc00000000000000b300000000000000b000000000",
            INIT_2E => X"000000d000000000000000cf00000000000000d000000000000000c400000000",
            INIT_2F => X"000000be00000000000000d800000000000000d100000000000000d000000000",
            INIT_30 => X"000000bd00000000000000b900000000000000ac000000000000009800000000",
            INIT_31 => X"00000060000000000000009300000000000000c600000000000000c200000000",
            INIT_32 => X"0000009800000000000000900000000000000097000000000000009500000000",
            INIT_33 => X"0000008b00000000000000800000000000000079000000000000009800000000",
            INIT_34 => X"000000a200000000000000aa0000000000000097000000000000009c00000000",
            INIT_35 => X"000000a4000000000000009600000000000000ad000000000000009600000000",
            INIT_36 => X"000000d200000000000000cc00000000000000a6000000000000009c00000000",
            INIT_37 => X"000000bc00000000000000d400000000000000cf00000000000000d300000000",
            INIT_38 => X"000000bb00000000000000b600000000000000ac000000000000009b00000000",
            INIT_39 => X"00000065000000000000007700000000000000b500000000000000c200000000",
            INIT_3A => X"0000007800000000000000830000000000000083000000000000007b00000000",
            INIT_3B => X"0000007f00000000000000870000000000000087000000000000009200000000",
            INIT_3C => X"0000007b0000000000000083000000000000007b000000000000007b00000000",
            INIT_3D => X"0000009f000000000000007b0000000000000084000000000000006d00000000",
            INIT_3E => X"000000c700000000000000bf0000000000000084000000000000007b00000000",
            INIT_3F => X"000000ba00000000000000d000000000000000c900000000000000c900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b900000000000000b400000000000000af00000000000000a100000000",
            INIT_41 => X"000000af00000000000000ab00000000000000ba00000000000000c000000000",
            INIT_42 => X"000000a600000000000000ac00000000000000a500000000000000a200000000",
            INIT_43 => X"000000aa00000000000000ad00000000000000ac00000000000000af00000000",
            INIT_44 => X"000000af00000000000000b200000000000000b200000000000000ac00000000",
            INIT_45 => X"000000be00000000000000b200000000000000ac00000000000000a300000000",
            INIT_46 => X"000000cd00000000000000c800000000000000b000000000000000ac00000000",
            INIT_47 => X"000000b900000000000000d100000000000000c900000000000000c800000000",
            INIT_48 => X"000000ba00000000000000b400000000000000b700000000000000ac00000000",
            INIT_49 => X"000000b700000000000000c200000000000000c000000000000000be00000000",
            INIT_4A => X"000000a300000000000000a200000000000000a500000000000000a000000000",
            INIT_4B => X"000000a200000000000000a4000000000000009e000000000000009f00000000",
            INIT_4C => X"000000a200000000000000ac00000000000000ae00000000000000a700000000",
            INIT_4D => X"000000b600000000000000a500000000000000a300000000000000a000000000",
            INIT_4E => X"000000cd00000000000000ca00000000000000c600000000000000c800000000",
            INIT_4F => X"000000b800000000000000d000000000000000ca00000000000000ca00000000",
            INIT_50 => X"000000be00000000000000ba00000000000000c400000000000000b100000000",
            INIT_51 => X"000000b700000000000000c100000000000000c100000000000000c000000000",
            INIT_52 => X"0000009f00000000000000a500000000000000a700000000000000a300000000",
            INIT_53 => X"000000ac00000000000000aa00000000000000a600000000000000a400000000",
            INIT_54 => X"000000ab00000000000000a600000000000000a600000000000000a800000000",
            INIT_55 => X"000000b200000000000000ab00000000000000ad00000000000000a800000000",
            INIT_56 => X"000000c700000000000000c700000000000000c600000000000000c700000000",
            INIT_57 => X"000000b800000000000000d000000000000000c800000000000000c800000000",
            INIT_58 => X"000000c800000000000000c300000000000000cc00000000000000b700000000",
            INIT_59 => X"000000c600000000000000be00000000000000bb00000000000000c900000000",
            INIT_5A => X"000000c100000000000000c100000000000000c100000000000000c200000000",
            INIT_5B => X"000000c600000000000000c600000000000000c200000000000000c100000000",
            INIT_5C => X"000000c600000000000000c300000000000000c300000000000000c600000000",
            INIT_5D => X"000000c500000000000000c400000000000000c400000000000000c500000000",
            INIT_5E => X"000000c900000000000000c900000000000000cb00000000000000c900000000",
            INIT_5F => X"000000bb00000000000000d100000000000000c800000000000000ca00000000",
            INIT_60 => X"000000b200000000000000c600000000000000cd00000000000000b900000000",
            INIT_61 => X"000000c4000000000000009a000000000000008d00000000000000a600000000",
            INIT_62 => X"000000c500000000000000c700000000000000ca00000000000000ca00000000",
            INIT_63 => X"000000ca00000000000000c900000000000000c700000000000000c500000000",
            INIT_64 => X"000000c400000000000000c600000000000000c700000000000000c900000000",
            INIT_65 => X"000000c600000000000000c700000000000000c600000000000000c400000000",
            INIT_66 => X"000000ce00000000000000cb00000000000000ca00000000000000c700000000",
            INIT_67 => X"000000bd00000000000000d400000000000000ce00000000000000cf00000000",
            INIT_68 => X"000000a500000000000000c800000000000000d000000000000000ba00000000",
            INIT_69 => X"0000006b000000000000005f000000000000007c000000000000009000000000",
            INIT_6A => X"000000c700000000000000c700000000000000b3000000000000008f00000000",
            INIT_6B => X"000000cc00000000000000c900000000000000c600000000000000c500000000",
            INIT_6C => X"000000cc00000000000000ce00000000000000cd00000000000000cc00000000",
            INIT_6D => X"000000cd00000000000000cd00000000000000c900000000000000c900000000",
            INIT_6E => X"000000cb00000000000000cb00000000000000cb00000000000000cc00000000",
            INIT_6F => X"000000b700000000000000cf00000000000000ca00000000000000ca00000000",
            INIT_70 => X"000000cc00000000000000d000000000000000d400000000000000ba00000000",
            INIT_71 => X"0000005b000000000000008f00000000000000c100000000000000ce00000000",
            INIT_72 => X"000000b5000000000000008e0000000000000065000000000000005100000000",
            INIT_73 => X"000000cf00000000000000cf00000000000000cc00000000000000c600000000",
            INIT_74 => X"000000ca00000000000000cf00000000000000cf00000000000000cf00000000",
            INIT_75 => X"000000c500000000000000c600000000000000c500000000000000c500000000",
            INIT_76 => X"000000c500000000000000c500000000000000c500000000000000c500000000",
            INIT_77 => X"000000b500000000000000cc00000000000000c500000000000000c400000000",
            INIT_78 => X"000000ce00000000000000d200000000000000d600000000000000b800000000",
            INIT_79 => X"000000b300000000000000cf00000000000000d400000000000000d100000000",
            INIT_7A => X"00000080000000000000005d0000000000000053000000000000007400000000",
            INIT_7B => X"000000ce00000000000000d200000000000000cb00000000000000ae00000000",
            INIT_7C => X"000000c900000000000000ca00000000000000ca00000000000000cc00000000",
            INIT_7D => X"000000c900000000000000c900000000000000c700000000000000c600000000",
            INIT_7E => X"000000c700000000000000c900000000000000ca00000000000000c800000000",
            INIT_7F => X"000000b400000000000000cb00000000000000c600000000000000c600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "sampleifmap_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d500000000000000d600000000000000d700000000000000ba00000000",
            INIT_01 => X"000000d900000000000000d400000000000000d600000000000000d600000000",
            INIT_02 => X"000000560000000000000049000000000000005b00000000000000af00000000",
            INIT_03 => X"000000cc00000000000000b5000000000000008a000000000000006500000000",
            INIT_04 => X"000000c600000000000000c700000000000000cb00000000000000d000000000",
            INIT_05 => X"000000c800000000000000c900000000000000c900000000000000c700000000",
            INIT_06 => X"000000c900000000000000c900000000000000ca00000000000000c800000000",
            INIT_07 => X"000000b600000000000000cc00000000000000c800000000000000ca00000000",
            INIT_08 => X"000000d900000000000000d800000000000000d800000000000000bb00000000",
            INIT_09 => X"000000d300000000000000d600000000000000d900000000000000db00000000",
            INIT_0A => X"000000520000000000000044000000000000007b00000000000000cc00000000",
            INIT_0B => X"0000008200000000000000610000000000000051000000000000004f00000000",
            INIT_0C => X"000000ca00000000000000c900000000000000bc00000000000000a500000000",
            INIT_0D => X"000000c600000000000000c700000000000000c100000000000000c400000000",
            INIT_0E => X"000000c800000000000000c800000000000000c700000000000000c600000000",
            INIT_0F => X"000000b600000000000000cc00000000000000c700000000000000c900000000",
            INIT_10 => X"000000d600000000000000d500000000000000d900000000000000bc00000000",
            INIT_11 => X"000000d200000000000000d600000000000000d800000000000000d800000000",
            INIT_12 => X"000000530000000000000046000000000000008800000000000000d400000000",
            INIT_13 => X"0000004d00000000000000500000000000000050000000000000004e00000000",
            INIT_14 => X"00000097000000000000007e0000000000000066000000000000005300000000",
            INIT_15 => X"000000cc00000000000000c900000000000000b2000000000000009f00000000",
            INIT_16 => X"000000c600000000000000c800000000000000c900000000000000cb00000000",
            INIT_17 => X"000000b400000000000000c900000000000000c500000000000000c700000000",
            INIT_18 => X"000000d500000000000000d600000000000000da00000000000000bb00000000",
            INIT_19 => X"000000d800000000000000d700000000000000d800000000000000d700000000",
            INIT_1A => X"00000037000000000000002d000000000000007000000000000000cc00000000",
            INIT_1B => X"00000051000000000000004d0000000000000045000000000000003a00000000",
            INIT_1C => X"0000003e0000000000000046000000000000004d000000000000005000000000",
            INIT_1D => X"000000a0000000000000007c000000000000004f000000000000003b00000000",
            INIT_1E => X"000000cd00000000000000cd00000000000000c400000000000000b500000000",
            INIT_1F => X"000000b400000000000000ca00000000000000c800000000000000cb00000000",
            INIT_20 => X"000000d100000000000000d200000000000000d800000000000000bc00000000",
            INIT_21 => X"000000d400000000000000d400000000000000d600000000000000d300000000",
            INIT_22 => X"00000021000000000000003a000000000000005f000000000000009a00000000",
            INIT_23 => X"0000004d0000000000000041000000000000003e000000000000003000000000",
            INIT_24 => X"0000004800000000000000540000000000000054000000000000005200000000",
            INIT_25 => X"00000048000000000000003f000000000000002f000000000000003800000000",
            INIT_26 => X"0000009e0000000000000084000000000000006b000000000000004e00000000",
            INIT_27 => X"000000b600000000000000ca00000000000000c100000000000000b500000000",
            INIT_28 => X"000000cf00000000000000ce00000000000000d200000000000000b800000000",
            INIT_29 => X"000000c800000000000000d400000000000000d300000000000000d100000000",
            INIT_2A => X"00000061000000000000008f0000000000000085000000000000009100000000",
            INIT_2B => X"0000005a000000000000002e0000000000000032000000000000002d00000000",
            INIT_2C => X"00000047000000000000007f000000000000009e000000000000009600000000",
            INIT_2D => X"0000004100000000000000580000000000000070000000000000006100000000",
            INIT_2E => X"000000a200000000000000a50000000000000082000000000000004300000000",
            INIT_2F => X"000000b000000000000000c500000000000000b500000000000000a800000000",
            INIT_30 => X"000000d000000000000000cd00000000000000d200000000000000b700000000",
            INIT_31 => X"000000d200000000000000d500000000000000d400000000000000d300000000",
            INIT_32 => X"000000bf00000000000000d400000000000000d100000000000000d100000000",
            INIT_33 => X"000000a600000000000000930000000000000093000000000000009400000000",
            INIT_34 => X"0000009d00000000000000c300000000000000d000000000000000c800000000",
            INIT_35 => X"000000a200000000000000b400000000000000b500000000000000a600000000",
            INIT_36 => X"000000c500000000000000c100000000000000b4000000000000009f00000000",
            INIT_37 => X"000000b100000000000000c700000000000000c100000000000000c300000000",
            INIT_38 => X"000000c200000000000000c300000000000000c400000000000000ae00000000",
            INIT_39 => X"000000b900000000000000bb00000000000000be00000000000000c200000000",
            INIT_3A => X"000000b500000000000000b700000000000000b500000000000000b800000000",
            INIT_3B => X"000000ad00000000000000ae00000000000000b000000000000000b200000000",
            INIT_3C => X"000000ac00000000000000a600000000000000a400000000000000aa00000000",
            INIT_3D => X"000000b000000000000000aa00000000000000a600000000000000aa00000000",
            INIT_3E => X"0000009b000000000000009d00000000000000a500000000000000af00000000",
            INIT_3F => X"0000009e00000000000000af00000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000070000000000000006c000000000000007000000000",
            INIT_41 => X"0000006000000000000000610000000000000064000000000000006700000000",
            INIT_42 => X"00000057000000000000005e000000000000005a000000000000005c00000000",
            INIT_43 => X"0000006700000000000000570000000000000053000000000000005400000000",
            INIT_44 => X"00000070000000000000006f0000000000000070000000000000007300000000",
            INIT_45 => X"0000007600000000000000740000000000000073000000000000007100000000",
            INIT_46 => X"0000007b000000000000007c000000000000007b000000000000007a00000000",
            INIT_47 => X"0000007c0000000000000084000000000000007a000000000000007900000000",
            INIT_48 => X"0000007000000000000000710000000000000073000000000000007500000000",
            INIT_49 => X"000000710000000000000071000000000000006f000000000000007100000000",
            INIT_4A => X"0000006e000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006b000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006e000000000000006c0000000000000073000000000000007300000000",
            INIT_4D => X"0000006b0000000000000068000000000000006d000000000000006f00000000",
            INIT_4E => X"000000700000000000000070000000000000006e000000000000006d00000000",
            INIT_4F => X"000000650000000000000062000000000000005f000000000000006400000000",
            INIT_50 => X"0000006a00000000000000690000000000000066000000000000007100000000",
            INIT_51 => X"0000005d00000000000000610000000000000066000000000000006a00000000",
            INIT_52 => X"000000550000000000000059000000000000005e000000000000005f00000000",
            INIT_53 => X"0000004e000000000000004f000000000000004e000000000000005200000000",
            INIT_54 => X"000000440000000000000047000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000041000000000000004300000000",
            INIT_56 => X"0000004100000000000000420000000000000042000000000000004100000000",
            INIT_57 => X"0000006400000000000000470000000000000037000000000000003c00000000",
            INIT_58 => X"000000400000000000000041000000000000003c000000000000005400000000",
            INIT_59 => X"0000003c000000000000003e0000000000000040000000000000004000000000",
            INIT_5A => X"00000038000000000000003d0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003b00000000000000410000000000000043000000000000004000000000",
            INIT_5D => X"0000003c000000000000003b000000000000003a000000000000003800000000",
            INIT_5E => X"0000003800000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000008000000000000000750000000000000048000000000000003800000000",
            INIT_60 => X"0000003e000000000000003f000000000000003b000000000000005300000000",
            INIT_61 => X"0000003f000000000000003d0000000000000041000000000000003f00000000",
            INIT_62 => X"00000039000000000000003c000000000000003e000000000000004300000000",
            INIT_63 => X"0000003d000000000000003c000000000000003a000000000000003a00000000",
            INIT_64 => X"0000003e00000000000000400000000000000044000000000000004100000000",
            INIT_65 => X"0000003d000000000000003e000000000000003c000000000000003d00000000",
            INIT_66 => X"00000041000000000000003d000000000000003a000000000000003a00000000",
            INIT_67 => X"0000006300000000000000890000000000000088000000000000005b00000000",
            INIT_68 => X"00000039000000000000003d0000000000000035000000000000004f00000000",
            INIT_69 => X"0000003c000000000000003a000000000000003b000000000000003700000000",
            INIT_6A => X"000000370000000000000039000000000000003c000000000000003d00000000",
            INIT_6B => X"0000003f000000000000003d000000000000003e000000000000003c00000000",
            INIT_6C => X"0000003b000000000000003c000000000000003f000000000000004300000000",
            INIT_6D => X"0000003f0000000000000040000000000000003e000000000000003e00000000",
            INIT_6E => X"0000006e0000000000000047000000000000003c000000000000003e00000000",
            INIT_6F => X"0000004a000000000000004f0000000000000077000000000000008e00000000",
            INIT_70 => X"000000410000000000000042000000000000003a000000000000005200000000",
            INIT_71 => X"0000003e000000000000003e000000000000003e000000000000003f00000000",
            INIT_72 => X"0000004f0000000000000041000000000000003e000000000000003f00000000",
            INIT_73 => X"0000004d000000000000004a000000000000004c000000000000004f00000000",
            INIT_74 => X"0000004e00000000000000500000000000000050000000000000005400000000",
            INIT_75 => X"00000041000000000000003e000000000000003f000000000000004c00000000",
            INIT_76 => X"0000008d000000000000007c0000000000000056000000000000004200000000",
            INIT_77 => X"0000004500000000000000400000000000000042000000000000006600000000",
            INIT_78 => X"0000003a000000000000003a0000000000000034000000000000004e00000000",
            INIT_79 => X"00000039000000000000003b000000000000003a000000000000003a00000000",
            INIT_7A => X"00000045000000000000003a000000000000003b000000000000003a00000000",
            INIT_7B => X"0000004500000000000000460000000000000047000000000000004700000000",
            INIT_7C => X"0000004a00000000000000490000000000000048000000000000004800000000",
            INIT_7D => X"00000044000000000000003f000000000000003f000000000000004900000000",
            INIT_7E => X"0000005800000000000000800000000000000080000000000000005a00000000",
            INIT_7F => X"000000440000000000000041000000000000003f000000000000004200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "sampleifmap_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cd00000000000000c100000000000000bb000000000000009500000000",
            INIT_01 => X"000000b400000000000000b500000000000000b700000000000000ca00000000",
            INIT_02 => X"000000c000000000000000c100000000000000bd00000000000000b600000000",
            INIT_03 => X"000000bd00000000000000bd00000000000000c000000000000000c000000000",
            INIT_04 => X"000000c000000000000000bd00000000000000b900000000000000ba00000000",
            INIT_05 => X"000000be00000000000000c000000000000000c100000000000000c100000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000ab00000000000000d400000000000000d100000000000000ca00000000",
            INIT_08 => X"000000e300000000000000d700000000000000cc000000000000009d00000000",
            INIT_09 => X"000000b300000000000000b300000000000000be00000000000000e000000000",
            INIT_0A => X"000000c300000000000000c300000000000000bb00000000000000b300000000",
            INIT_0B => X"000000b700000000000000b400000000000000be00000000000000bb00000000",
            INIT_0C => X"000000b700000000000000b800000000000000b700000000000000bc00000000",
            INIT_0D => X"000000bc00000000000000bc00000000000000bf00000000000000b900000000",
            INIT_0E => X"000000e000000000000000d300000000000000c200000000000000be00000000",
            INIT_0F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_10 => X"000000db00000000000000d500000000000000c9000000000000009900000000",
            INIT_11 => X"000000b800000000000000c400000000000000d500000000000000df00000000",
            INIT_12 => X"000000d400000000000000d300000000000000c300000000000000b100000000",
            INIT_13 => X"000000ca00000000000000cc00000000000000d200000000000000d000000000",
            INIT_14 => X"000000d100000000000000d000000000000000d100000000000000d100000000",
            INIT_15 => X"000000d000000000000000d000000000000000d400000000000000d200000000",
            INIT_16 => X"000000df00000000000000de00000000000000d500000000000000d000000000",
            INIT_17 => X"000000b800000000000000e000000000000000d700000000000000da00000000",
            INIT_18 => X"000000de00000000000000d300000000000000cf00000000000000a600000000",
            INIT_19 => X"0000008300000000000000c900000000000000dc00000000000000e200000000",
            INIT_1A => X"000000b100000000000000a6000000000000009e000000000000007700000000",
            INIT_1B => X"000000ab00000000000000a600000000000000a700000000000000b200000000",
            INIT_1C => X"000000ba00000000000000b200000000000000b200000000000000b700000000",
            INIT_1D => X"000000a500000000000000b400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000dd00000000000000dc00000000000000e400000000000000cf00000000",
            INIT_1F => X"000000ba00000000000000e600000000000000df00000000000000e000000000",
            INIT_20 => X"000000da00000000000000ca00000000000000cb00000000000000a700000000",
            INIT_21 => X"0000008e00000000000000d600000000000000e100000000000000e000000000",
            INIT_22 => X"0000008100000000000000780000000000000098000000000000009900000000",
            INIT_23 => X"00000083000000000000007c000000000000007e000000000000008100000000",
            INIT_24 => X"0000008a00000000000000820000000000000084000000000000008600000000",
            INIT_25 => X"0000007b000000000000008d0000000000000088000000000000008800000000",
            INIT_26 => X"000000d900000000000000da00000000000000e300000000000000ba00000000",
            INIT_27 => X"000000b900000000000000e300000000000000dc00000000000000de00000000",
            INIT_28 => X"000000d900000000000000cb00000000000000c900000000000000a400000000",
            INIT_29 => X"000000a500000000000000d100000000000000da00000000000000dc00000000",
            INIT_2A => X"000000b4000000000000009c00000000000000b500000000000000c400000000",
            INIT_2B => X"000000ac00000000000000a300000000000000a000000000000000b300000000",
            INIT_2C => X"000000c900000000000000be00000000000000c100000000000000bf00000000",
            INIT_2D => X"000000be00000000000000c600000000000000c000000000000000bf00000000",
            INIT_2E => X"000000e100000000000000e100000000000000e100000000000000d400000000",
            INIT_2F => X"000000bc00000000000000e800000000000000e100000000000000df00000000",
            INIT_30 => X"000000d900000000000000c800000000000000c600000000000000a400000000",
            INIT_31 => X"0000006800000000000000ac00000000000000d600000000000000d900000000",
            INIT_32 => X"000000af00000000000000a600000000000000a5000000000000009e00000000",
            INIT_33 => X"000000a00000000000000097000000000000009000000000000000a500000000",
            INIT_34 => X"000000b600000000000000bd00000000000000ad00000000000000b200000000",
            INIT_35 => X"000000b900000000000000ad00000000000000b700000000000000aa00000000",
            INIT_36 => X"000000e200000000000000dc00000000000000b200000000000000a600000000",
            INIT_37 => X"000000bc00000000000000e700000000000000e000000000000000dd00000000",
            INIT_38 => X"000000d800000000000000c700000000000000c900000000000000a900000000",
            INIT_39 => X"0000006f000000000000009200000000000000cb00000000000000da00000000",
            INIT_3A => X"00000090000000000000009d0000000000000095000000000000008600000000",
            INIT_3B => X"00000090000000000000008f000000000000008f000000000000009b00000000",
            INIT_3C => X"0000008e0000000000000094000000000000008e000000000000009300000000",
            INIT_3D => X"000000b0000000000000008e000000000000008d000000000000007f00000000",
            INIT_3E => X"000000dc00000000000000d10000000000000095000000000000008900000000",
            INIT_3F => X"000000ba00000000000000e400000000000000dc00000000000000d900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d900000000000000c700000000000000ce00000000000000b100000000",
            INIT_41 => X"000000c500000000000000c100000000000000cd00000000000000db00000000",
            INIT_42 => X"000000b800000000000000bb00000000000000b700000000000000b800000000",
            INIT_43 => X"000000bd00000000000000bb00000000000000ba00000000000000c000000000",
            INIT_44 => X"000000bf00000000000000c200000000000000c200000000000000c000000000",
            INIT_45 => X"000000c800000000000000bc00000000000000ba00000000000000b200000000",
            INIT_46 => X"000000db00000000000000d600000000000000c600000000000000c100000000",
            INIT_47 => X"000000b900000000000000e400000000000000dd00000000000000db00000000",
            INIT_48 => X"000000d600000000000000c500000000000000d400000000000000ba00000000",
            INIT_49 => X"000000d200000000000000dc00000000000000d600000000000000d700000000",
            INIT_4A => X"000000ba00000000000000b600000000000000bb00000000000000b900000000",
            INIT_4B => X"000000ba00000000000000b900000000000000b400000000000000b600000000",
            INIT_4C => X"000000b800000000000000c300000000000000c600000000000000c100000000",
            INIT_4D => X"000000c600000000000000b600000000000000b600000000000000b500000000",
            INIT_4E => X"000000df00000000000000dd00000000000000de00000000000000de00000000",
            INIT_4F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_50 => X"000000d800000000000000c800000000000000de00000000000000bc00000000",
            INIT_51 => X"000000cc00000000000000d600000000000000d400000000000000d700000000",
            INIT_52 => X"000000b000000000000000b600000000000000b800000000000000b500000000",
            INIT_53 => X"000000bf00000000000000bc00000000000000b800000000000000b500000000",
            INIT_54 => X"000000b900000000000000b800000000000000ba00000000000000bd00000000",
            INIT_55 => X"000000c900000000000000ba00000000000000b800000000000000b600000000",
            INIT_56 => X"000000db00000000000000dc00000000000000dd00000000000000df00000000",
            INIT_57 => X"000000b800000000000000e300000000000000dc00000000000000db00000000",
            INIT_58 => X"000000e000000000000000cf00000000000000e200000000000000bf00000000",
            INIT_59 => X"000000de00000000000000d700000000000000d100000000000000dc00000000",
            INIT_5A => X"000000d700000000000000d600000000000000d700000000000000d900000000",
            INIT_5B => X"000000df00000000000000df00000000000000db00000000000000d900000000",
            INIT_5C => X"000000da00000000000000db00000000000000dd00000000000000df00000000",
            INIT_5D => X"000000db00000000000000d900000000000000d600000000000000d800000000",
            INIT_5E => X"000000d600000000000000d900000000000000db00000000000000db00000000",
            INIT_5F => X"000000ba00000000000000e300000000000000db00000000000000d700000000",
            INIT_60 => X"000000ce00000000000000d400000000000000dc00000000000000bc00000000",
            INIT_61 => X"000000d900000000000000ac000000000000009900000000000000b500000000",
            INIT_62 => X"000000dc00000000000000dd00000000000000e100000000000000e200000000",
            INIT_63 => X"000000e200000000000000e100000000000000df00000000000000de00000000",
            INIT_64 => X"000000da00000000000000dc00000000000000dd00000000000000e100000000",
            INIT_65 => X"000000da00000000000000dc00000000000000db00000000000000d900000000",
            INIT_66 => X"000000e000000000000000de00000000000000dc00000000000000d900000000",
            INIT_67 => X"000000bb00000000000000e600000000000000e000000000000000e000000000",
            INIT_68 => X"000000c100000000000000d600000000000000df00000000000000bd00000000",
            INIT_69 => X"000000730000000000000063000000000000007e000000000000009d00000000",
            INIT_6A => X"000000dd00000000000000dd00000000000000c6000000000000009d00000000",
            INIT_6B => X"000000e200000000000000df00000000000000dc00000000000000da00000000",
            INIT_6C => X"000000df00000000000000e100000000000000e000000000000000e200000000",
            INIT_6D => X"000000e000000000000000e000000000000000dd00000000000000dc00000000",
            INIT_6E => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_6F => X"000000b700000000000000e200000000000000dd00000000000000dd00000000",
            INIT_70 => X"000000e900000000000000de00000000000000e200000000000000bd00000000",
            INIT_71 => X"0000005a000000000000009200000000000000c400000000000000dc00000000",
            INIT_72 => X"000000ca00000000000000a10000000000000071000000000000005400000000",
            INIT_73 => X"000000e400000000000000e300000000000000e000000000000000da00000000",
            INIT_74 => X"000000dc00000000000000e000000000000000e100000000000000e200000000",
            INIT_75 => X"000000d900000000000000d800000000000000d700000000000000d700000000",
            INIT_76 => X"000000d800000000000000d800000000000000d800000000000000d800000000",
            INIT_77 => X"000000b600000000000000e100000000000000da00000000000000d700000000",
            INIT_78 => X"000000ea00000000000000e000000000000000e500000000000000bb00000000",
            INIT_79 => X"000000b300000000000000da00000000000000e100000000000000e100000000",
            INIT_7A => X"00000091000000000000006a0000000000000058000000000000007300000000",
            INIT_7B => X"000000e100000000000000e400000000000000dd00000000000000c000000000",
            INIT_7C => X"000000d900000000000000da00000000000000db00000000000000df00000000",
            INIT_7D => X"000000db00000000000000d900000000000000d600000000000000d600000000",
            INIT_7E => X"000000da00000000000000dc00000000000000dd00000000000000db00000000",
            INIT_7F => X"000000b700000000000000e200000000000000dc00000000000000d900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "sampleifmap_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e900000000000000de00000000000000e900000000000000be00000000",
            INIT_01 => X"000000e100000000000000e000000000000000e200000000000000e400000000",
            INIT_02 => X"0000005b0000000000000050000000000000006200000000000000b500000000",
            INIT_03 => X"000000d900000000000000c00000000000000092000000000000006a00000000",
            INIT_04 => X"000000da00000000000000dd00000000000000e100000000000000e000000000",
            INIT_05 => X"000000d900000000000000da00000000000000da00000000000000d900000000",
            INIT_06 => X"000000dd00000000000000dd00000000000000dd00000000000000da00000000",
            INIT_07 => X"000000bc00000000000000e300000000000000dc00000000000000dd00000000",
            INIT_08 => X"000000e900000000000000dd00000000000000ea00000000000000bf00000000",
            INIT_09 => X"000000dd00000000000000e200000000000000e300000000000000e700000000",
            INIT_0A => X"0000004f0000000000000049000000000000008200000000000000d500000000",
            INIT_0B => X"0000008800000000000000640000000000000050000000000000004b00000000",
            INIT_0C => X"000000dc00000000000000d700000000000000c800000000000000ad00000000",
            INIT_0D => X"000000de00000000000000df00000000000000d900000000000000d900000000",
            INIT_0E => X"000000db00000000000000db00000000000000dd00000000000000dd00000000",
            INIT_0F => X"000000bd00000000000000e300000000000000db00000000000000da00000000",
            INIT_10 => X"000000e400000000000000d900000000000000e800000000000000bd00000000",
            INIT_11 => X"000000dc00000000000000e200000000000000e100000000000000e300000000",
            INIT_12 => X"00000050000000000000004a000000000000009000000000000000dd00000000",
            INIT_13 => X"0000004c000000000000004e000000000000004c000000000000004a00000000",
            INIT_14 => X"000000a100000000000000810000000000000064000000000000005300000000",
            INIT_15 => X"000000e200000000000000e100000000000000c900000000000000b000000000",
            INIT_16 => X"000000d700000000000000d900000000000000dc00000000000000df00000000",
            INIT_17 => X"000000bb00000000000000e100000000000000d900000000000000d700000000",
            INIT_18 => X"000000e100000000000000d700000000000000e800000000000000bb00000000",
            INIT_19 => X"000000e200000000000000e300000000000000e100000000000000e000000000",
            INIT_1A => X"000000380000000000000032000000000000007700000000000000d500000000",
            INIT_1B => X"00000052000000000000004d0000000000000045000000000000003b00000000",
            INIT_1C => X"0000003f00000000000000420000000000000048000000000000005000000000",
            INIT_1D => X"000000a20000000000000085000000000000005b000000000000004100000000",
            INIT_1E => X"000000df00000000000000da00000000000000cc00000000000000b800000000",
            INIT_1F => X"000000bc00000000000000e300000000000000dd00000000000000dd00000000",
            INIT_20 => X"000000df00000000000000de00000000000000e700000000000000b700000000",
            INIT_21 => X"000000e100000000000000e400000000000000e600000000000000df00000000",
            INIT_22 => X"00000027000000000000003c000000000000006200000000000000a200000000",
            INIT_23 => X"0000004e00000000000000440000000000000043000000000000003500000000",
            INIT_24 => X"0000004800000000000000530000000000000052000000000000005100000000",
            INIT_25 => X"00000043000000000000003f0000000000000031000000000000003900000000",
            INIT_26 => X"000000a8000000000000008b000000000000006d000000000000004b00000000",
            INIT_27 => X"000000c300000000000000df00000000000000d700000000000000c600000000",
            INIT_28 => X"000000de00000000000000e200000000000000e200000000000000b000000000",
            INIT_29 => X"000000d400000000000000e200000000000000e200000000000000de00000000",
            INIT_2A => X"0000006a0000000000000096000000000000008b000000000000009b00000000",
            INIT_2B => X"0000005e00000000000000330000000000000039000000000000003500000000",
            INIT_2C => X"00000049000000000000008200000000000000a1000000000000009a00000000",
            INIT_2D => X"00000043000000000000005a0000000000000072000000000000006300000000",
            INIT_2E => X"000000a900000000000000ab0000000000000086000000000000004500000000",
            INIT_2F => X"000000be00000000000000d000000000000000c500000000000000b700000000",
            INIT_30 => X"000000df00000000000000e100000000000000e100000000000000af00000000",
            INIT_31 => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_32 => X"000000cc00000000000000e400000000000000e000000000000000de00000000",
            INIT_33 => X"000000b300000000000000a0000000000000009f000000000000009f00000000",
            INIT_34 => X"000000a900000000000000cf00000000000000dc00000000000000d600000000",
            INIT_35 => X"000000ad00000000000000c000000000000000c100000000000000b200000000",
            INIT_36 => X"000000d600000000000000d200000000000000c300000000000000ab00000000",
            INIT_37 => X"000000bd00000000000000d200000000000000d100000000000000d800000000",
            INIT_38 => X"000000d100000000000000d700000000000000d400000000000000a600000000",
            INIT_39 => X"000000c700000000000000c900000000000000cc00000000000000ce00000000",
            INIT_3A => X"000000c200000000000000c500000000000000c300000000000000c700000000",
            INIT_3B => X"000000c400000000000000c200000000000000c100000000000000c000000000",
            INIT_3C => X"000000ca00000000000000c400000000000000c200000000000000c400000000",
            INIT_3D => X"000000cd00000000000000c800000000000000c400000000000000c800000000",
            INIT_3E => X"000000bf00000000000000c000000000000000c500000000000000ce00000000",
            INIT_3F => X"000000b500000000000000c900000000000000c500000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007800000000000000820000000000000078000000000000006500000000",
            INIT_41 => X"0000006a000000000000006b0000000000000070000000000000007600000000",
            INIT_42 => X"0000006300000000000000660000000000000062000000000000006500000000",
            INIT_43 => X"00000080000000000000006c0000000000000065000000000000006200000000",
            INIT_44 => X"0000009300000000000000920000000000000092000000000000009000000000",
            INIT_45 => X"0000009e00000000000000980000000000000096000000000000009400000000",
            INIT_46 => X"000000a800000000000000a800000000000000a600000000000000a400000000",
            INIT_47 => X"0000009200000000000000a700000000000000a500000000000000a800000000",
            INIT_48 => X"0000008600000000000000860000000000000082000000000000006f00000000",
            INIT_49 => X"0000008800000000000000890000000000000088000000000000008a00000000",
            INIT_4A => X"0000007e00000000000000830000000000000086000000000000008400000000",
            INIT_4B => X"0000008300000000000000830000000000000080000000000000007f00000000",
            INIT_4C => X"00000081000000000000007f0000000000000086000000000000008a00000000",
            INIT_4D => X"0000007e000000000000007c0000000000000080000000000000008100000000",
            INIT_4E => X"0000008400000000000000840000000000000082000000000000008100000000",
            INIT_4F => X"0000006000000000000000730000000000000073000000000000007700000000",
            INIT_50 => X"0000007800000000000000780000000000000071000000000000006800000000",
            INIT_51 => X"00000064000000000000006c0000000000000076000000000000007a00000000",
            INIT_52 => X"000000590000000000000055000000000000005b000000000000006000000000",
            INIT_53 => X"0000005600000000000000570000000000000055000000000000005800000000",
            INIT_54 => X"000000430000000000000046000000000000004f000000000000005600000000",
            INIT_55 => X"0000003c000000000000003f0000000000000041000000000000004200000000",
            INIT_56 => X"0000003b000000000000003c000000000000003c000000000000003b00000000",
            INIT_57 => X"0000004b000000000000003f0000000000000032000000000000003600000000",
            INIT_58 => X"00000039000000000000003d0000000000000037000000000000003d00000000",
            INIT_59 => X"00000036000000000000003b000000000000003f000000000000003a00000000",
            INIT_5A => X"0000002f000000000000002f0000000000000033000000000000003800000000",
            INIT_5B => X"0000003200000000000000310000000000000032000000000000003000000000",
            INIT_5C => X"0000002f00000000000000350000000000000037000000000000003300000000",
            INIT_5D => X"000000370000000000000032000000000000002e000000000000002d00000000",
            INIT_5E => X"0000003400000000000000340000000000000034000000000000003600000000",
            INIT_5F => X"000000680000000000000068000000000000003a000000000000003000000000",
            INIT_60 => X"0000003c0000000000000041000000000000003d000000000000004400000000",
            INIT_61 => X"000000390000000000000037000000000000003d000000000000003e00000000",
            INIT_62 => X"0000003a00000000000000370000000000000038000000000000003d00000000",
            INIT_63 => X"0000003600000000000000380000000000000038000000000000003b00000000",
            INIT_64 => X"000000340000000000000037000000000000003b000000000000003900000000",
            INIT_65 => X"0000003400000000000000340000000000000033000000000000003300000000",
            INIT_66 => X"0000003900000000000000370000000000000035000000000000003300000000",
            INIT_67 => X"0000004b00000000000000780000000000000071000000000000004b00000000",
            INIT_68 => X"00000035000000000000003b0000000000000034000000000000003e00000000",
            INIT_69 => X"0000003600000000000000340000000000000039000000000000003900000000",
            INIT_6A => X"0000003200000000000000300000000000000032000000000000003600000000",
            INIT_6B => X"0000003500000000000000340000000000000038000000000000003900000000",
            INIT_6C => X"0000003300000000000000340000000000000036000000000000003900000000",
            INIT_6D => X"0000003000000000000000350000000000000037000000000000003600000000",
            INIT_6E => X"0000005f000000000000003d0000000000000034000000000000003200000000",
            INIT_6F => X"00000032000000000000003e0000000000000065000000000000007c00000000",
            INIT_70 => X"00000037000000000000003a0000000000000035000000000000003e00000000",
            INIT_71 => X"0000003c000000000000003c000000000000003d000000000000003b00000000",
            INIT_72 => X"0000004b000000000000003a0000000000000037000000000000003900000000",
            INIT_73 => X"0000004500000000000000440000000000000048000000000000004c00000000",
            INIT_74 => X"00000049000000000000004b000000000000004a000000000000004b00000000",
            INIT_75 => X"000000350000000000000037000000000000003a000000000000004600000000",
            INIT_76 => X"0000007f000000000000006b0000000000000045000000000000003300000000",
            INIT_77 => X"000000330000000000000036000000000000003a000000000000005b00000000",
            INIT_78 => X"0000002e00000000000000330000000000000033000000000000004000000000",
            INIT_79 => X"0000003500000000000000390000000000000038000000000000003300000000",
            INIT_7A => X"0000003e00000000000000320000000000000033000000000000003400000000",
            INIT_7B => X"00000039000000000000003c000000000000003e000000000000004000000000",
            INIT_7C => X"000000400000000000000040000000000000003e000000000000003c00000000",
            INIT_7D => X"0000003700000000000000340000000000000035000000000000004000000000",
            INIT_7E => X"0000004800000000000000690000000000000067000000000000004600000000",
            INIT_7F => X"0000003200000000000000340000000000000032000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "sampleifmap_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e00000000000000300000000000000046000000000000004100000000",
            INIT_01 => X"0000002d000000000000002c0000000000000028000000000000001700000000",
            INIT_02 => X"0000000f000000000000000a0000000000000028000000000000002d00000000",
            INIT_03 => X"0000003000000000000000330000000000000035000000000000002c00000000",
            INIT_04 => X"0000005b000000000000005d000000000000005a000000000000004100000000",
            INIT_05 => X"00000037000000000000003c0000000000000051000000000000005f00000000",
            INIT_06 => X"000000440000000000000029000000000000006f000000000000007000000000",
            INIT_07 => X"0000004300000000000000360000000000000033000000000000004d00000000",
            INIT_08 => X"0000001e000000000000003c000000000000004f000000000000004500000000",
            INIT_09 => X"0000003100000000000000310000000000000041000000000000002900000000",
            INIT_0A => X"0000001900000000000000070000000000000023000000000000003100000000",
            INIT_0B => X"0000003100000000000000370000000000000045000000000000004100000000",
            INIT_0C => X"0000005000000000000000530000000000000055000000000000004d00000000",
            INIT_0D => X"0000003b00000000000000370000000000000051000000000000005700000000",
            INIT_0E => X"0000002f000000000000001f0000000000000079000000000000008300000000",
            INIT_0F => X"0000003d00000000000000410000000000000036000000000000003800000000",
            INIT_10 => X"0000002900000000000000480000000000000054000000000000004900000000",
            INIT_11 => X"000000360000000000000032000000000000004a000000000000004000000000",
            INIT_12 => X"00000024000000000000000b0000000000000020000000000000003600000000",
            INIT_13 => X"00000027000000000000002f0000000000000043000000000000003c00000000",
            INIT_14 => X"0000003e000000000000003b000000000000004d000000000000004b00000000",
            INIT_15 => X"0000003f00000000000000300000000000000055000000000000005300000000",
            INIT_16 => X"0000002900000000000000170000000000000080000000000000008b00000000",
            INIT_17 => X"000000300000000000000049000000000000004e000000000000004600000000",
            INIT_18 => X"000000360000000000000050000000000000004b000000000000005800000000",
            INIT_19 => X"0000003f00000000000000370000000000000044000000000000005000000000",
            INIT_1A => X"000000250000000000000011000000000000001c000000000000003a00000000",
            INIT_1B => X"0000002700000000000000280000000000000033000000000000002b00000000",
            INIT_1C => X"00000046000000000000004b0000000000000062000000000000005500000000",
            INIT_1D => X"0000004400000000000000320000000000000054000000000000005600000000",
            INIT_1E => X"0000004b000000000000002f0000000000000089000000000000008e00000000",
            INIT_1F => X"000000260000000000000041000000000000005d000000000000006400000000",
            INIT_20 => X"00000042000000000000006f0000000000000059000000000000005f00000000",
            INIT_21 => X"00000044000000000000003d000000000000003d000000000000005100000000",
            INIT_22 => X"00000016000000000000000f0000000000000016000000000000003e00000000",
            INIT_23 => X"0000003f00000000000000330000000000000023000000000000001f00000000",
            INIT_24 => X"000000470000000000000048000000000000004b000000000000004800000000",
            INIT_25 => X"0000004e00000000000000330000000000000053000000000000004d00000000",
            INIT_26 => X"000000570000000000000057000000000000009c000000000000009500000000",
            INIT_27 => X"00000058000000000000004b000000000000005f000000000000006300000000",
            INIT_28 => X"0000004d00000000000000520000000000000053000000000000005200000000",
            INIT_29 => X"000000390000000000000040000000000000003a000000000000004700000000",
            INIT_2A => X"0000001c00000000000000110000000000000014000000000000003b00000000",
            INIT_2B => X"000000470000000000000047000000000000003d000000000000003200000000",
            INIT_2C => X"0000003800000000000000440000000000000043000000000000004500000000",
            INIT_2D => X"0000004e00000000000000460000000000000053000000000000002900000000",
            INIT_2E => X"00000059000000000000006200000000000000ac000000000000009c00000000",
            INIT_2F => X"000000630000000000000070000000000000006f000000000000005e00000000",
            INIT_30 => X"0000003b00000000000000200000000000000040000000000000004500000000",
            INIT_31 => X"000000310000000000000049000000000000004a000000000000004800000000",
            INIT_32 => X"0000003e000000000000001d0000000000000012000000000000003100000000",
            INIT_33 => X"0000003f00000000000000560000000000000055000000000000005200000000",
            INIT_34 => X"0000002b000000000000005f0000000000000034000000000000002200000000",
            INIT_35 => X"0000004e0000000000000055000000000000005e000000000000001900000000",
            INIT_36 => X"0000006b000000000000006d00000000000000b400000000000000a600000000",
            INIT_37 => X"0000002f00000000000000560000000000000083000000000000006c00000000",
            INIT_38 => X"0000004600000000000000190000000000000035000000000000003b00000000",
            INIT_39 => X"0000003d0000000000000050000000000000004e000000000000005100000000",
            INIT_3A => X"0000005e0000000000000035000000000000000a000000000000002800000000",
            INIT_3B => X"00000019000000000000004b0000000000000058000000000000005700000000",
            INIT_3C => X"00000039000000000000005c000000000000002d000000000000000d00000000",
            INIT_3D => X"0000006200000000000000590000000000000065000000000000003200000000",
            INIT_3E => X"0000007c000000000000007800000000000000b3000000000000009000000000",
            INIT_3F => X"0000001800000000000000340000000000000080000000000000007c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000660000000000000031000000000000002f000000000000004400000000",
            INIT_41 => X"0000004f000000000000003f0000000000000059000000000000007700000000",
            INIT_42 => X"0000006000000000000000510000000000000022000000000000004200000000",
            INIT_43 => X"0000000e0000000000000029000000000000005a000000000000005900000000",
            INIT_44 => X"000000470000000000000043000000000000005c000000000000003400000000",
            INIT_45 => X"00000073000000000000006e0000000000000071000000000000006f00000000",
            INIT_46 => X"0000007f0000000000000079000000000000009c000000000000008800000000",
            INIT_47 => X"00000016000000000000001f0000000000000073000000000000007c00000000",
            INIT_48 => X"0000007200000000000000370000000000000035000000000000004d00000000",
            INIT_49 => X"000000370000000000000041000000000000007b000000000000008000000000",
            INIT_4A => X"0000006e000000000000006f0000000000000052000000000000004f00000000",
            INIT_4B => X"0000002500000000000000140000000000000045000000000000006a00000000",
            INIT_4C => X"0000006100000000000000530000000000000069000000000000005c00000000",
            INIT_4D => X"0000005c00000000000000730000000000000078000000000000007600000000",
            INIT_4E => X"0000007f000000000000007d0000000000000093000000000000009000000000",
            INIT_4F => X"00000017000000000000000e000000000000005f000000000000007700000000",
            INIT_50 => X"000000700000000000000036000000000000003a000000000000005500000000",
            INIT_51 => X"0000003100000000000000640000000000000084000000000000008100000000",
            INIT_52 => X"0000006d00000000000000680000000000000054000000000000002700000000",
            INIT_53 => X"00000053000000000000003f000000000000005d000000000000007d00000000",
            INIT_54 => X"0000006e0000000000000068000000000000005e000000000000006100000000",
            INIT_55 => X"000000390000000000000055000000000000007f000000000000006d00000000",
            INIT_56 => X"0000007c000000000000007b0000000000000096000000000000009800000000",
            INIT_57 => X"00000015000000000000000c000000000000005d000000000000007200000000",
            INIT_58 => X"0000006b00000000000000320000000000000035000000000000006c00000000",
            INIT_59 => X"0000004b00000000000000800000000000000083000000000000007e00000000",
            INIT_5A => X"0000006b0000000000000055000000000000005b000000000000003300000000",
            INIT_5B => X"000000930000000000000081000000000000006e000000000000008a00000000",
            INIT_5C => X"0000007700000000000000710000000000000078000000000000008400000000",
            INIT_5D => X"0000005d000000000000005a0000000000000073000000000000007500000000",
            INIT_5E => X"0000007d0000000000000071000000000000008d00000000000000a000000000",
            INIT_5F => X"00000009000000000000000e0000000000000065000000000000007900000000",
            INIT_60 => X"0000005c000000000000002b000000000000002a000000000000006000000000",
            INIT_61 => X"0000007700000000000000820000000000000080000000000000006a00000000",
            INIT_62 => X"000000890000000000000072000000000000007b000000000000007800000000",
            INIT_63 => X"000000840000000000000069000000000000006e000000000000009400000000",
            INIT_64 => X"0000008600000000000000800000000000000087000000000000009200000000",
            INIT_65 => X"00000077000000000000007e0000000000000078000000000000008c00000000",
            INIT_66 => X"0000006a00000000000000630000000000000091000000000000009800000000",
            INIT_67 => X"0000002800000000000000120000000000000063000000000000008200000000",
            INIT_68 => X"00000059000000000000003b0000000000000042000000000000006100000000",
            INIT_69 => X"000000880000000000000085000000000000006f000000000000006400000000",
            INIT_6A => X"000000910000000000000096000000000000008c000000000000009300000000",
            INIT_6B => X"0000007f00000000000000830000000000000088000000000000008e00000000",
            INIT_6C => X"000000930000000000000088000000000000007b000000000000007d00000000",
            INIT_6D => X"00000088000000000000009c000000000000008e000000000000009700000000",
            INIT_6E => X"00000070000000000000006d0000000000000090000000000000009200000000",
            INIT_6F => X"000000530000000000000032000000000000005c000000000000008200000000",
            INIT_70 => X"0000005f000000000000004b0000000000000048000000000000006900000000",
            INIT_71 => X"000000850000000000000085000000000000005e000000000000006800000000",
            INIT_72 => X"0000008500000000000000800000000000000087000000000000008f00000000",
            INIT_73 => X"0000009800000000000000a00000000000000096000000000000009300000000",
            INIT_74 => X"0000008700000000000000840000000000000090000000000000009100000000",
            INIT_75 => X"000000a500000000000000a2000000000000008a000000000000008a00000000",
            INIT_76 => X"00000077000000000000007e000000000000007f00000000000000a300000000",
            INIT_77 => X"0000004d000000000000003b000000000000005f000000000000007600000000",
            INIT_78 => X"0000005b00000000000000440000000000000044000000000000005e00000000",
            INIT_79 => X"00000083000000000000007b0000000000000062000000000000006500000000",
            INIT_7A => X"0000004f000000000000008a00000000000000c1000000000000009300000000",
            INIT_7B => X"000000a200000000000000930000000000000093000000000000007c00000000",
            INIT_7C => X"00000090000000000000009800000000000000ab00000000000000b400000000",
            INIT_7D => X"000000b300000000000000940000000000000079000000000000009000000000",
            INIT_7E => X"0000007b000000000000008000000000000000a000000000000000b400000000",
            INIT_7F => X"00000054000000000000001a000000000000003f000000000000007000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "sampleifmap_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000004a000000000000004f000000000000005800000000",
            INIT_01 => X"0000008100000000000000780000000000000078000000000000006e00000000",
            INIT_02 => X"0000005700000000000000c000000000000000b8000000000000007800000000",
            INIT_03 => X"000000a600000000000000a4000000000000009c000000000000007200000000",
            INIT_04 => X"000000b600000000000000b700000000000000a1000000000000009a00000000",
            INIT_05 => X"0000008f000000000000009400000000000000ad00000000000000bb00000000",
            INIT_06 => X"0000007c000000000000008e00000000000000c300000000000000b500000000",
            INIT_07 => X"000000760000000000000029000000000000002c000000000000006b00000000",
            INIT_08 => X"0000006000000000000000670000000000000059000000000000005b00000000",
            INIT_09 => X"0000006a000000000000006f0000000000000064000000000000007400000000",
            INIT_0A => X"000000a800000000000000bb0000000000000080000000000000007200000000",
            INIT_0B => X"000000ac00000000000000ac0000000000000099000000000000008c00000000",
            INIT_0C => X"000000a3000000000000009d00000000000000a400000000000000a700000000",
            INIT_0D => X"0000009c00000000000000ab00000000000000a500000000000000a100000000",
            INIT_0E => X"0000007200000000000000a7000000000000009100000000000000a100000000",
            INIT_0F => X"0000005e000000000000002a000000000000004a000000000000006a00000000",
            INIT_10 => X"0000007a00000000000000780000000000000061000000000000006500000000",
            INIT_11 => X"0000005b000000000000005f000000000000004e000000000000007200000000",
            INIT_12 => X"000000cc0000000000000081000000000000006e000000000000007300000000",
            INIT_13 => X"0000009900000000000000a0000000000000008900000000000000a700000000",
            INIT_14 => X"000000b200000000000000aa00000000000000ba00000000000000b300000000",
            INIT_15 => X"000000a500000000000000a2000000000000009c00000000000000b300000000",
            INIT_16 => X"000000480000000000000068000000000000008c000000000000009c00000000",
            INIT_17 => X"0000007200000000000000460000000000000059000000000000005400000000",
            INIT_18 => X"00000060000000000000007a000000000000006b000000000000006e00000000",
            INIT_19 => X"000000640000000000000048000000000000004c000000000000005a00000000",
            INIT_1A => X"0000008c0000000000000057000000000000007f000000000000006d00000000",
            INIT_1B => X"000000b400000000000000a6000000000000009f00000000000000bd00000000",
            INIT_1C => X"000000bc00000000000000be00000000000000ad00000000000000ae00000000",
            INIT_1D => X"000000a100000000000000a2000000000000009900000000000000a200000000",
            INIT_1E => X"0000004a000000000000004b0000000000000095000000000000009900000000",
            INIT_1F => X"0000008a0000000000000070000000000000003e000000000000004200000000",
            INIT_20 => X"0000004e0000000000000059000000000000006a000000000000007700000000",
            INIT_21 => X"00000067000000000000003c0000000000000047000000000000005900000000",
            INIT_22 => X"000000420000000000000072000000000000005f000000000000004b00000000",
            INIT_23 => X"000000be00000000000000ae00000000000000b5000000000000007f00000000",
            INIT_24 => X"000000c100000000000000b800000000000000ab00000000000000ba00000000",
            INIT_25 => X"000000a500000000000000ab00000000000000a000000000000000a400000000",
            INIT_26 => X"0000005c0000000000000068000000000000008b000000000000009200000000",
            INIT_27 => X"000000730000000000000070000000000000005e000000000000004d00000000",
            INIT_28 => X"00000067000000000000003a000000000000005e000000000000007e00000000",
            INIT_29 => X"0000005f0000000000000048000000000000004c000000000000006a00000000",
            INIT_2A => X"0000006300000000000000780000000000000041000000000000005e00000000",
            INIT_2B => X"000000bc00000000000000c400000000000000a1000000000000005b00000000",
            INIT_2C => X"000000a700000000000000a700000000000000c100000000000000b600000000",
            INIT_2D => X"000000a1000000000000009a00000000000000a000000000000000aa00000000",
            INIT_2E => X"00000051000000000000006e000000000000008a000000000000009100000000",
            INIT_2F => X"00000064000000000000006d0000000000000088000000000000006900000000",
            INIT_30 => X"0000006800000000000000460000000000000052000000000000006f00000000",
            INIT_31 => X"000000540000000000000045000000000000005e000000000000007100000000",
            INIT_32 => X"0000007d0000000000000055000000000000006d000000000000007400000000",
            INIT_33 => X"000000c800000000000000ba000000000000009b000000000000007f00000000",
            INIT_34 => X"0000009d00000000000000b100000000000000bb00000000000000bb00000000",
            INIT_35 => X"000000a600000000000000a400000000000000a2000000000000009400000000",
            INIT_36 => X"000000610000000000000079000000000000009500000000000000a200000000",
            INIT_37 => X"0000006100000000000000610000000000000073000000000000007800000000",
            INIT_38 => X"000000b4000000000000008c000000000000005c000000000000006500000000",
            INIT_39 => X"0000004c0000000000000055000000000000007b000000000000009700000000",
            INIT_3A => X"00000054000000000000005a000000000000007c000000000000006700000000",
            INIT_3B => X"000000c800000000000000ad00000000000000af000000000000009200000000",
            INIT_3C => X"0000009f00000000000000ad00000000000000ad00000000000000bc00000000",
            INIT_3D => X"000000ad00000000000000a300000000000000ac000000000000009f00000000",
            INIT_3E => X"000000830000000000000083000000000000008b00000000000000a400000000",
            INIT_3F => X"000000600000000000000064000000000000005f000000000000007000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000c00000000000000090000000000000007700000000",
            INIT_41 => X"0000006c000000000000007f000000000000009d00000000000000c200000000",
            INIT_42 => X"0000006f000000000000006a000000000000005e000000000000006a00000000",
            INIT_43 => X"000000c500000000000000b000000000000000af000000000000007c00000000",
            INIT_44 => X"000000a500000000000000b000000000000000aa00000000000000b800000000",
            INIT_45 => X"000000a300000000000000af00000000000000c5000000000000009c00000000",
            INIT_46 => X"00000065000000000000007a0000000000000083000000000000009300000000",
            INIT_47 => X"00000066000000000000006b0000000000000060000000000000006400000000",
            INIT_48 => X"000000a9000000000000008a0000000000000074000000000000006e00000000",
            INIT_49 => X"0000008800000000000000a000000000000000c400000000000000c500000000",
            INIT_4A => X"0000008a000000000000005c0000000000000063000000000000008100000000",
            INIT_4B => X"000000a900000000000000b4000000000000009f000000000000009200000000",
            INIT_4C => X"000000b200000000000000af000000000000008d000000000000008e00000000",
            INIT_4D => X"0000009700000000000000b300000000000000bc00000000000000a600000000",
            INIT_4E => X"0000003a0000000000000070000000000000009a000000000000008f00000000",
            INIT_4F => X"0000004900000000000000660000000000000065000000000000005b00000000",
            INIT_50 => X"0000006b000000000000004a0000000000000057000000000000005b00000000",
            INIT_51 => X"000000a300000000000000bf00000000000000b900000000000000a500000000",
            INIT_52 => X"00000066000000000000006a0000000000000080000000000000008600000000",
            INIT_53 => X"0000007400000000000000920000000000000084000000000000007600000000",
            INIT_54 => X"000000b600000000000000a10000000000000063000000000000004d00000000",
            INIT_55 => X"000000a700000000000000ad000000000000009f00000000000000b700000000",
            INIT_56 => X"0000002b000000000000005e0000000000000087000000000000009c00000000",
            INIT_57 => X"0000004d0000000000000044000000000000005c000000000000005b00000000",
            INIT_58 => X"0000002c0000000000000032000000000000005f000000000000005100000000",
            INIT_59 => X"000000bb00000000000000a60000000000000094000000000000005f00000000",
            INIT_5A => X"00000072000000000000007e000000000000009000000000000000ae00000000",
            INIT_5B => X"0000006b00000000000000770000000000000072000000000000006800000000",
            INIT_5C => X"000000b6000000000000009d0000000000000052000000000000005100000000",
            INIT_5D => X"0000009600000000000000a900000000000000b200000000000000a900000000",
            INIT_5E => X"0000003f000000000000002c000000000000006c000000000000009800000000",
            INIT_5F => X"0000005600000000000000500000000000000045000000000000006100000000",
            INIT_60 => X"000000150000000000000034000000000000005f000000000000005a00000000",
            INIT_61 => X"000000b00000000000000092000000000000006d000000000000001c00000000",
            INIT_62 => X"0000007f000000000000008e00000000000000b500000000000000ca00000000",
            INIT_63 => X"0000008200000000000000720000000000000077000000000000007800000000",
            INIT_64 => X"000000a900000000000000900000000000000076000000000000008100000000",
            INIT_65 => X"0000009800000000000000b400000000000000ad000000000000009f00000000",
            INIT_66 => X"00000055000000000000002c0000000000000044000000000000007700000000",
            INIT_67 => X"0000006a00000000000000a70000000000000072000000000000003300000000",
            INIT_68 => X"000000340000000000000039000000000000005b000000000000005f00000000",
            INIT_69 => X"0000009c00000000000000770000000000000031000000000000001800000000",
            INIT_6A => X"0000009b00000000000000ba00000000000000cb00000000000000bb00000000",
            INIT_6B => X"0000007500000000000000740000000000000085000000000000008d00000000",
            INIT_6C => X"00000099000000000000008b0000000000000077000000000000006d00000000",
            INIT_6D => X"0000007d000000000000009c00000000000000a7000000000000009f00000000",
            INIT_6E => X"0000004000000000000000440000000000000041000000000000006500000000",
            INIT_6F => X"0000007a00000000000000aa0000000000000090000000000000003700000000",
            INIT_70 => X"000000490000000000000020000000000000004b000000000000005e00000000",
            INIT_71 => X"0000007300000000000000360000000000000021000000000000002e00000000",
            INIT_72 => X"000000c200000000000000c300000000000000b0000000000000009600000000",
            INIT_73 => X"000000920000000000000088000000000000009b00000000000000b100000000",
            INIT_74 => X"00000077000000000000005e0000000000000065000000000000008b00000000",
            INIT_75 => X"000000690000000000000060000000000000005f000000000000006500000000",
            INIT_76 => X"0000006d000000000000006b0000000000000076000000000000008300000000",
            INIT_77 => X"0000006a000000000000009a000000000000008f000000000000008000000000",
            INIT_78 => X"0000004c00000000000000180000000000000023000000000000004e00000000",
            INIT_79 => X"0000003b000000000000001b0000000000000028000000000000004100000000",
            INIT_7A => X"000000b000000000000000960000000000000088000000000000007800000000",
            INIT_7B => X"000000ba00000000000000a500000000000000b700000000000000c000000000",
            INIT_7C => X"00000056000000000000006b00000000000000aa00000000000000cf00000000",
            INIT_7D => X"0000008c00000000000000700000000000000055000000000000004200000000",
            INIT_7E => X"000000890000000000000089000000000000009500000000000000a900000000",
            INIT_7F => X"00000080000000000000009a000000000000008f000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "sampleifmap_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000000000400000000000000051000000000000004400000000",
            INIT_01 => X"00000050000000000000004b0000000000000039000000000000002100000000",
            INIT_02 => X"0000002200000000000000140000000000000046000000000000005300000000",
            INIT_03 => X"000000420000000000000046000000000000004b000000000000004700000000",
            INIT_04 => X"00000079000000000000007c0000000000000078000000000000005700000000",
            INIT_05 => X"000000520000000000000054000000000000006c000000000000007e00000000",
            INIT_06 => X"0000005b000000000000003b0000000000000081000000000000008800000000",
            INIT_07 => X"00000057000000000000004c0000000000000043000000000000006000000000",
            INIT_08 => X"0000002f000000000000004a0000000000000066000000000000005000000000",
            INIT_09 => X"000000540000000000000054000000000000005c000000000000003800000000",
            INIT_0A => X"000000300000000000000012000000000000003e000000000000005800000000",
            INIT_0B => X"00000049000000000000004d000000000000005c000000000000005d00000000",
            INIT_0C => X"0000006a000000000000006f0000000000000075000000000000006b00000000",
            INIT_0D => X"00000053000000000000004d000000000000006c000000000000007500000000",
            INIT_0E => X"00000041000000000000002d000000000000008b000000000000009700000000",
            INIT_0F => X"00000051000000000000005a0000000000000042000000000000004700000000",
            INIT_10 => X"000000380000000000000058000000000000006d000000000000005f00000000",
            INIT_11 => X"0000005a00000000000000560000000000000069000000000000005400000000",
            INIT_12 => X"0000003c00000000000000140000000000000035000000000000005c00000000",
            INIT_13 => X"0000003c00000000000000420000000000000058000000000000005900000000",
            INIT_14 => X"00000054000000000000004e0000000000000066000000000000006700000000",
            INIT_15 => X"0000005600000000000000420000000000000072000000000000007200000000",
            INIT_16 => X"000000370000000000000023000000000000008f000000000000009e00000000",
            INIT_17 => X"0000003b00000000000000620000000000000062000000000000005400000000",
            INIT_18 => X"0000004900000000000000640000000000000064000000000000007400000000",
            INIT_19 => X"0000006000000000000000580000000000000066000000000000006d00000000",
            INIT_1A => X"00000038000000000000001a000000000000002d000000000000005e00000000",
            INIT_1B => X"0000003700000000000000360000000000000043000000000000004100000000",
            INIT_1C => X"0000006200000000000000610000000000000075000000000000006a00000000",
            INIT_1D => X"0000005b00000000000000450000000000000072000000000000007600000000",
            INIT_1E => X"0000005d0000000000000040000000000000009600000000000000a000000000",
            INIT_1F => X"00000032000000000000005e000000000000007e000000000000007800000000",
            INIT_20 => X"0000005d00000000000000800000000000000068000000000000007800000000",
            INIT_21 => X"0000005e000000000000005a000000000000005e000000000000007200000000",
            INIT_22 => X"00000024000000000000001a0000000000000027000000000000005d00000000",
            INIT_23 => X"0000005600000000000000490000000000000037000000000000002f00000000",
            INIT_24 => X"00000065000000000000006b0000000000000071000000000000006900000000",
            INIT_25 => X"00000067000000000000004a000000000000006d000000000000006700000000",
            INIT_26 => X"00000074000000000000007000000000000000ac00000000000000a200000000",
            INIT_27 => X"0000006c00000000000000670000000000000084000000000000008100000000",
            INIT_28 => X"0000006200000000000000620000000000000066000000000000006900000000",
            INIT_29 => X"0000004e000000000000005b0000000000000059000000000000005f00000000",
            INIT_2A => X"0000002b000000000000001b0000000000000023000000000000005800000000",
            INIT_2B => X"0000006c000000000000006a000000000000005d000000000000004d00000000",
            INIT_2C => X"0000004e00000000000000640000000000000065000000000000006700000000",
            INIT_2D => X"000000660000000000000062000000000000006e000000000000003900000000",
            INIT_2E => X"0000007f000000000000008200000000000000ba00000000000000a700000000",
            INIT_2F => X"0000007800000000000000840000000000000090000000000000008100000000",
            INIT_30 => X"0000004f00000000000000300000000000000060000000000000005e00000000",
            INIT_31 => X"0000003f000000000000005d0000000000000064000000000000005a00000000",
            INIT_32 => X"0000005a0000000000000026000000000000001d000000000000004a00000000",
            INIT_33 => X"0000006300000000000000820000000000000081000000000000007e00000000",
            INIT_34 => X"0000003900000000000000730000000000000047000000000000003a00000000",
            INIT_35 => X"0000006a0000000000000071000000000000007b000000000000002500000000",
            INIT_36 => X"0000008c000000000000008d00000000000000c100000000000000b700000000",
            INIT_37 => X"0000003b000000000000006500000000000000a0000000000000008900000000",
            INIT_38 => X"00000069000000000000002f0000000000000054000000000000005600000000",
            INIT_39 => X"00000047000000000000005e0000000000000061000000000000006700000000",
            INIT_3A => X"0000008b00000000000000490000000000000014000000000000003800000000",
            INIT_3B => X"000000290000000000000072000000000000008c000000000000008a00000000",
            INIT_3C => X"0000004f00000000000000730000000000000041000000000000001a00000000",
            INIT_3D => X"0000008c0000000000000078000000000000007d000000000000003b00000000",
            INIT_3E => X"00000094000000000000009600000000000000c300000000000000b000000000",
            INIT_3F => X"00000018000000000000003f000000000000009b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c000000000000004a000000000000004e000000000000006200000000",
            INIT_41 => X"0000005c00000000000000500000000000000072000000000000009500000000",
            INIT_42 => X"000000900000000000000071000000000000002c000000000000004700000000",
            INIT_43 => X"00000017000000000000003f0000000000000086000000000000008800000000",
            INIT_44 => X"00000056000000000000005e000000000000007c000000000000004500000000",
            INIT_45 => X"000000a5000000000000009b000000000000008b000000000000007000000000",
            INIT_46 => X"00000096000000000000009600000000000000b100000000000000aa00000000",
            INIT_47 => X"000000160000000000000029000000000000008e000000000000009200000000",
            INIT_48 => X"00000094000000000000004e0000000000000051000000000000007400000000",
            INIT_49 => X"000000450000000000000054000000000000009b00000000000000a300000000",
            INIT_4A => X"0000008e0000000000000089000000000000005a000000000000005100000000",
            INIT_4B => X"000000380000000000000021000000000000005d000000000000008a00000000",
            INIT_4C => X"000000800000000000000073000000000000008f000000000000007c00000000",
            INIT_4D => X"00000081000000000000009c000000000000009c000000000000009700000000",
            INIT_4E => X"0000009a000000000000009800000000000000ad00000000000000a700000000",
            INIT_4F => X"0000001800000000000000160000000000000079000000000000009400000000",
            INIT_50 => X"000000910000000000000049000000000000004f000000000000007800000000",
            INIT_51 => X"00000041000000000000007f00000000000000a600000000000000a500000000",
            INIT_52 => X"0000007f000000000000008e0000000000000072000000000000003600000000",
            INIT_53 => X"0000006c0000000000000047000000000000005d000000000000007e00000000",
            INIT_54 => X"000000a100000000000000920000000000000085000000000000008700000000",
            INIT_55 => X"00000057000000000000007500000000000000a5000000000000009c00000000",
            INIT_56 => X"0000009c000000000000009700000000000000af00000000000000a900000000",
            INIT_57 => X"0000001700000000000000130000000000000074000000000000009100000000",
            INIT_58 => X"0000008a00000000000000420000000000000045000000000000007b00000000",
            INIT_59 => X"0000005f00000000000000a500000000000000a800000000000000a100000000",
            INIT_5A => X"00000070000000000000008a000000000000008c000000000000004b00000000",
            INIT_5B => X"000000a200000000000000880000000000000066000000000000006d00000000",
            INIT_5C => X"000000870000000000000097000000000000009a000000000000009900000000",
            INIT_5D => X"0000008800000000000000760000000000000085000000000000007c00000000",
            INIT_5E => X"0000009d000000000000009200000000000000aa00000000000000bd00000000",
            INIT_5F => X"0000000b00000000000000140000000000000077000000000000009400000000",
            INIT_60 => X"00000079000000000000003c0000000000000039000000000000006a00000000",
            INIT_61 => X"0000009800000000000000ad00000000000000a4000000000000008700000000",
            INIT_62 => X"00000076000000000000007f0000000000000093000000000000009000000000",
            INIT_63 => X"0000008b0000000000000066000000000000005c000000000000007300000000",
            INIT_64 => X"000000740000000000000085000000000000008a000000000000008d00000000",
            INIT_65 => X"000000880000000000000077000000000000006b000000000000007800000000",
            INIT_66 => X"00000091000000000000008700000000000000ae00000000000000b000000000",
            INIT_67 => X"0000002b000000000000001a000000000000007200000000000000a100000000",
            INIT_68 => X"00000074000000000000004e0000000000000055000000000000007400000000",
            INIT_69 => X"000000ab00000000000000ac000000000000008c000000000000007f00000000",
            INIT_6A => X"000000780000000000000082000000000000007c000000000000009900000000",
            INIT_6B => X"0000006e00000000000000710000000000000076000000000000007700000000",
            INIT_6C => X"0000007d0000000000000077000000000000006c000000000000006900000000",
            INIT_6D => X"000000750000000000000081000000000000007a000000000000008300000000",
            INIT_6E => X"0000009a000000000000008d00000000000000a2000000000000009000000000",
            INIT_6F => X"0000005f0000000000000041000000000000007000000000000000a600000000",
            INIT_70 => X"0000007800000000000000630000000000000060000000000000008400000000",
            INIT_71 => X"000000a800000000000000a50000000000000072000000000000008200000000",
            INIT_72 => X"000000700000000000000068000000000000006b000000000000008b00000000",
            INIT_73 => X"00000084000000000000008e0000000000000081000000000000007c00000000",
            INIT_74 => X"0000006f000000000000006b0000000000000077000000000000007a00000000",
            INIT_75 => X"00000090000000000000008d0000000000000076000000000000007300000000",
            INIT_76 => X"0000009f0000000000000092000000000000007b000000000000008e00000000",
            INIT_77 => X"0000005e00000000000000480000000000000070000000000000009d00000000",
            INIT_78 => X"00000076000000000000005d000000000000005a000000000000007900000000",
            INIT_79 => X"000000a60000000000000097000000000000007c000000000000007f00000000",
            INIT_7A => X"00000045000000000000007900000000000000ab000000000000009900000000",
            INIT_7B => X"0000008b000000000000007b000000000000007c000000000000006b00000000",
            INIT_7C => X"0000007700000000000000800000000000000090000000000000009b00000000",
            INIT_7D => X"000000a700000000000000830000000000000067000000000000007a00000000",
            INIT_7E => X"000000a00000000000000080000000000000008c000000000000009f00000000",
            INIT_7F => X"000000680000000000000022000000000000004b000000000000009500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "sampleifmap_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007e00000000000000640000000000000064000000000000007000000000",
            INIT_01 => X"000000a300000000000000950000000000000098000000000000008d00000000",
            INIT_02 => X"0000004700000000000000a600000000000000a3000000000000008a00000000",
            INIT_03 => X"0000008d000000000000008b0000000000000085000000000000006400000000",
            INIT_04 => X"0000009e00000000000000a00000000000000088000000000000008100000000",
            INIT_05 => X"0000007e000000000000007d000000000000009700000000000000a300000000",
            INIT_06 => X"0000008f000000000000007a00000000000000b100000000000000a900000000",
            INIT_07 => X"0000008b0000000000000033000000000000003d000000000000008f00000000",
            INIT_08 => X"0000008100000000000000830000000000000070000000000000007000000000",
            INIT_09 => X"000000890000000000000090000000000000007c000000000000009300000000",
            INIT_0A => X"0000009900000000000000a80000000000000079000000000000008f00000000",
            INIT_0B => X"000000930000000000000092000000000000007f000000000000007a00000000",
            INIT_0C => X"0000008a0000000000000084000000000000008b000000000000008d00000000",
            INIT_0D => X"000000860000000000000099000000000000008f000000000000008600000000",
            INIT_0E => X"0000007a00000000000000920000000000000082000000000000009100000000",
            INIT_0F => X"0000006f000000000000003a0000000000000064000000000000008600000000",
            INIT_10 => X"0000008e00000000000000950000000000000076000000000000007900000000",
            INIT_11 => X"00000076000000000000007b0000000000000061000000000000008d00000000",
            INIT_12 => X"000000bb0000000000000079000000000000007e000000000000008f00000000",
            INIT_13 => X"000000820000000000000088000000000000006e000000000000009100000000",
            INIT_14 => X"0000009a000000000000009400000000000000a1000000000000009a00000000",
            INIT_15 => X"0000009100000000000000960000000000000086000000000000009700000000",
            INIT_16 => X"000000570000000000000061000000000000007b000000000000008600000000",
            INIT_17 => X"0000008600000000000000610000000000000077000000000000006700000000",
            INIT_18 => X"0000006f00000000000000970000000000000087000000000000008800000000",
            INIT_19 => X"0000007d000000000000005d0000000000000065000000000000007a00000000",
            INIT_1A => X"0000007d00000000000000600000000000000099000000000000008600000000",
            INIT_1B => X"000000a00000000000000092000000000000008800000000000000a900000000",
            INIT_1C => X"000000a700000000000000a60000000000000094000000000000009600000000",
            INIT_1D => X"0000009100000000000000900000000000000080000000000000008d00000000",
            INIT_1E => X"0000005e000000000000004b0000000000000082000000000000008400000000",
            INIT_1F => X"000000a900000000000000950000000000000057000000000000005300000000",
            INIT_20 => X"0000005e0000000000000070000000000000008c000000000000009400000000",
            INIT_21 => X"0000008200000000000000540000000000000068000000000000007900000000",
            INIT_22 => X"0000004a000000000000008d0000000000000074000000000000006600000000",
            INIT_23 => X"000000aa000000000000009b00000000000000a3000000000000007600000000",
            INIT_24 => X"000000a7000000000000009d000000000000009500000000000000a500000000",
            INIT_25 => X"0000009100000000000000930000000000000089000000000000009200000000",
            INIT_26 => X"00000071000000000000006d000000000000007c000000000000007f00000000",
            INIT_27 => X"000000a1000000000000009c0000000000000077000000000000006000000000",
            INIT_28 => X"0000007d00000000000000480000000000000077000000000000009800000000",
            INIT_29 => X"0000007900000000000000630000000000000065000000000000008100000000",
            INIT_2A => X"0000007d000000000000009a000000000000005b000000000000007800000000",
            INIT_2B => X"000000a900000000000000b50000000000000096000000000000005d00000000",
            INIT_2C => X"0000008f000000000000009100000000000000ad00000000000000a200000000",
            INIT_2D => X"0000008b00000000000000810000000000000087000000000000008f00000000",
            INIT_2E => X"0000006600000000000000750000000000000078000000000000007d00000000",
            INIT_2F => X"00000099000000000000009a00000000000000ab000000000000008100000000",
            INIT_30 => X"0000007b00000000000000520000000000000068000000000000008800000000",
            INIT_31 => X"0000007300000000000000620000000000000076000000000000008800000000",
            INIT_32 => X"000000940000000000000075000000000000008d000000000000009600000000",
            INIT_33 => X"000000b300000000000000ad0000000000000095000000000000008100000000",
            INIT_34 => X"0000008f000000000000009f00000000000000a800000000000000a500000000",
            INIT_35 => X"0000008d000000000000008c000000000000008b000000000000007e00000000",
            INIT_36 => X"0000006d000000000000007a0000000000000085000000000000008800000000",
            INIT_37 => X"00000095000000000000009600000000000000a4000000000000009800000000",
            INIT_38 => X"000000bf0000000000000096000000000000006f000000000000007d00000000",
            INIT_39 => X"0000006f0000000000000079000000000000009e00000000000000ac00000000",
            INIT_3A => X"0000006900000000000000730000000000000099000000000000009100000000",
            INIT_3B => X"000000ac000000000000009a00000000000000a1000000000000009400000000",
            INIT_3C => X"0000008d000000000000009c000000000000009b00000000000000a100000000",
            INIT_3D => X"0000008f00000000000000880000000000000093000000000000008900000000",
            INIT_3E => X"00000086000000000000007b000000000000008c000000000000008900000000",
            INIT_3F => X"00000095000000000000009e0000000000000095000000000000009c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000dc00000000000000c800000000000000a2000000000000009500000000",
            INIT_41 => X"0000009300000000000000aa00000000000000bd00000000000000d100000000",
            INIT_42 => X"00000088000000000000007d000000000000007a000000000000009100000000",
            INIT_43 => X"000000a40000000000000096000000000000009f000000000000008b00000000",
            INIT_44 => X"0000008e000000000000009f000000000000009b000000000000009b00000000",
            INIT_45 => X"00000088000000000000009300000000000000a9000000000000008500000000",
            INIT_46 => X"00000072000000000000006b000000000000007e000000000000007f00000000",
            INIT_47 => X"0000009c00000000000000a0000000000000008f000000000000009a00000000",
            INIT_48 => X"000000be000000000000009d0000000000000089000000000000008b00000000",
            INIT_49 => X"000000b000000000000000bf00000000000000d700000000000000d500000000",
            INIT_4A => X"000000a30000000000000075000000000000008400000000000000a900000000",
            INIT_4B => X"0000008f000000000000009a000000000000009700000000000000ad00000000",
            INIT_4C => X"0000009800000000000000990000000000000081000000000000007c00000000",
            INIT_4D => X"0000007c000000000000009500000000000000a3000000000000009100000000",
            INIT_4E => X"0000004a00000000000000600000000000000083000000000000007700000000",
            INIT_4F => X"0000007800000000000000970000000000000095000000000000009100000000",
            INIT_50 => X"000000860000000000000061000000000000006f000000000000007300000000",
            INIT_51 => X"000000c100000000000000d300000000000000cf00000000000000bf00000000",
            INIT_52 => X"0000007f000000000000009100000000000000ad00000000000000b100000000",
            INIT_53 => X"000000680000000000000086000000000000008f000000000000009000000000",
            INIT_54 => X"0000009b000000000000008b000000000000005c000000000000004900000000",
            INIT_55 => X"0000008e0000000000000094000000000000008a00000000000000a100000000",
            INIT_56 => X"0000003c00000000000000550000000000000075000000000000008300000000",
            INIT_57 => X"0000006d000000000000006f0000000000000091000000000000009200000000",
            INIT_58 => X"0000004000000000000000410000000000000072000000000000006a00000000",
            INIT_59 => X"000000d500000000000000c300000000000000b2000000000000007800000000",
            INIT_5A => X"0000009900000000000000ad00000000000000b900000000000000ca00000000",
            INIT_5B => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_5C => X"0000009a000000000000008e0000000000000060000000000000006c00000000",
            INIT_5D => X"0000007f000000000000009500000000000000a1000000000000009000000000",
            INIT_5E => X"0000006100000000000000310000000000000062000000000000008300000000",
            INIT_5F => X"000000750000000000000076000000000000006c000000000000009300000000",
            INIT_60 => X"00000026000000000000003e0000000000000070000000000000007400000000",
            INIT_61 => X"000000c700000000000000b40000000000000087000000000000002900000000",
            INIT_62 => X"000000b200000000000000b700000000000000cc00000000000000d400000000",
            INIT_63 => X"000000a1000000000000009e00000000000000a400000000000000ab00000000",
            INIT_64 => X"0000008d0000000000000087000000000000008b000000000000009d00000000",
            INIT_65 => X"0000007e000000000000009c0000000000000099000000000000008700000000",
            INIT_66 => X"0000007c000000000000003b0000000000000042000000000000006700000000",
            INIT_67 => X"0000008300000000000000c50000000000000088000000000000005400000000",
            INIT_68 => X"0000004e000000000000004f000000000000007b000000000000007f00000000",
            INIT_69 => X"000000bf00000000000000950000000000000042000000000000002500000000",
            INIT_6A => X"000000c200000000000000d600000000000000db00000000000000d000000000",
            INIT_6B => X"0000009f00000000000000a500000000000000b400000000000000b800000000",
            INIT_6C => X"00000083000000000000007b000000000000007d000000000000008700000000",
            INIT_6D => X"0000007200000000000000870000000000000093000000000000008a00000000",
            INIT_6E => X"0000005b0000000000000055000000000000004f000000000000006c00000000",
            INIT_6F => X"0000008f00000000000000c900000000000000ac000000000000004e00000000",
            INIT_70 => X"0000006b00000000000000340000000000000068000000000000007d00000000",
            INIT_71 => X"00000097000000000000004e0000000000000030000000000000004300000000",
            INIT_72 => X"000000da00000000000000d900000000000000cb00000000000000bd00000000",
            INIT_73 => X"000000b600000000000000b400000000000000c300000000000000cd00000000",
            INIT_74 => X"0000007a000000000000005e000000000000007400000000000000a500000000",
            INIT_75 => X"0000006f00000000000000590000000000000059000000000000006100000000",
            INIT_76 => X"000000860000000000000082000000000000008a000000000000009600000000",
            INIT_77 => X"0000008100000000000000bc00000000000000b5000000000000009f00000000",
            INIT_78 => X"0000007300000000000000280000000000000033000000000000006600000000",
            INIT_79 => X"0000004e0000000000000029000000000000003a000000000000006000000000",
            INIT_7A => X"000000cf00000000000000b900000000000000b500000000000000a000000000",
            INIT_7B => X"000000ce00000000000000c400000000000000d200000000000000da00000000",
            INIT_7C => X"00000071000000000000007c00000000000000b400000000000000d600000000",
            INIT_7D => X"000000a000000000000000840000000000000066000000000000005600000000",
            INIT_7E => X"000000a700000000000000a700000000000000a700000000000000ba00000000",
            INIT_7F => X"0000009c00000000000000b900000000000000b300000000000000b400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "sampleifmap_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000002e0000000000000040000000000000003200000000",
            INIT_01 => X"0000003900000000000000370000000000000024000000000000001600000000",
            INIT_02 => X"00000012000000000000000c0000000000000036000000000000003b00000000",
            INIT_03 => X"000000320000000000000031000000000000002c000000000000002b00000000",
            INIT_04 => X"0000004d0000000000000051000000000000004d000000000000003a00000000",
            INIT_05 => X"000000390000000000000038000000000000004e000000000000005300000000",
            INIT_06 => X"0000003a000000000000001f000000000000005d000000000000006100000000",
            INIT_07 => X"0000004200000000000000350000000000000029000000000000004100000000",
            INIT_08 => X"0000001d00000000000000390000000000000051000000000000003a00000000",
            INIT_09 => X"0000003c000000000000003b000000000000003d000000000000002300000000",
            INIT_0A => X"0000001b0000000000000007000000000000002f000000000000004000000000",
            INIT_0B => X"0000002f000000000000003b000000000000003e000000000000003800000000",
            INIT_0C => X"00000044000000000000004a000000000000004a000000000000004400000000",
            INIT_0D => X"0000003c00000000000000330000000000000051000000000000004e00000000",
            INIT_0E => X"0000002700000000000000150000000000000060000000000000006f00000000",
            INIT_0F => X"000000420000000000000045000000000000002c000000000000002d00000000",
            INIT_10 => X"0000002300000000000000460000000000000057000000000000004800000000",
            INIT_11 => X"00000041000000000000003c0000000000000048000000000000003500000000",
            INIT_12 => X"0000002300000000000000070000000000000026000000000000004500000000",
            INIT_13 => X"0000002100000000000000300000000000000041000000000000003400000000",
            INIT_14 => X"0000003700000000000000320000000000000042000000000000004300000000",
            INIT_15 => X"0000003e000000000000002d0000000000000052000000000000004d00000000",
            INIT_16 => X"0000002600000000000000100000000000000063000000000000007400000000",
            INIT_17 => X"00000033000000000000004d000000000000004b000000000000003f00000000",
            INIT_18 => X"0000002f0000000000000050000000000000004c000000000000005e00000000",
            INIT_19 => X"0000004a00000000000000410000000000000048000000000000004700000000",
            INIT_1A => X"00000022000000000000000c000000000000001e000000000000004800000000",
            INIT_1B => X"0000001e00000000000000230000000000000034000000000000002800000000",
            INIT_1C => X"0000004500000000000000440000000000000057000000000000004b00000000",
            INIT_1D => X"00000043000000000000002e000000000000004d000000000000005100000000",
            INIT_1E => X"00000049000000000000002a000000000000006b000000000000007700000000",
            INIT_1F => X"0000002200000000000000440000000000000060000000000000005f00000000",
            INIT_20 => X"0000003c000000000000006a000000000000004f000000000000006100000000",
            INIT_21 => X"0000004c00000000000000480000000000000044000000000000004b00000000",
            INIT_22 => X"00000011000000000000000c0000000000000018000000000000004900000000",
            INIT_23 => X"0000003b00000000000000330000000000000025000000000000001c00000000",
            INIT_24 => X"00000047000000000000004b000000000000004f000000000000004800000000",
            INIT_25 => X"0000004d000000000000002d0000000000000049000000000000004700000000",
            INIT_26 => X"0000005500000000000000520000000000000081000000000000008000000000",
            INIT_27 => X"0000005000000000000000490000000000000061000000000000005e00000000",
            INIT_28 => X"00000043000000000000004b000000000000004d000000000000005200000000",
            INIT_29 => X"0000003d000000000000004d0000000000000045000000000000003d00000000",
            INIT_2A => X"00000016000000000000000d0000000000000013000000000000004300000000",
            INIT_2B => X"000000490000000000000047000000000000003b000000000000002c00000000",
            INIT_2C => X"0000003500000000000000490000000000000048000000000000004800000000",
            INIT_2D => X"0000004d000000000000003e0000000000000049000000000000002200000000",
            INIT_2E => X"0000005b00000000000000600000000000000093000000000000008800000000",
            INIT_2F => X"0000005c0000000000000068000000000000006e000000000000005c00000000",
            INIT_30 => X"0000003300000000000000190000000000000046000000000000004800000000",
            INIT_31 => X"00000032000000000000004f000000000000004f000000000000003e00000000",
            INIT_32 => X"000000360000000000000018000000000000000f000000000000003800000000",
            INIT_33 => X"0000003e000000000000004d000000000000004b000000000000004900000000",
            INIT_34 => X"0000002a00000000000000600000000000000033000000000000002200000000",
            INIT_35 => X"0000004a00000000000000480000000000000058000000000000001600000000",
            INIT_36 => X"0000006c000000000000006800000000000000a1000000000000009500000000",
            INIT_37 => X"0000002b00000000000000510000000000000083000000000000006b00000000",
            INIT_38 => X"000000460000000000000015000000000000003b000000000000003f00000000",
            INIT_39 => X"0000003a000000000000004b0000000000000048000000000000004d00000000",
            INIT_3A => X"00000051000000000000002f0000000000000008000000000000002900000000",
            INIT_3B => X"00000012000000000000003e000000000000004b000000000000004b00000000",
            INIT_3C => X"0000004000000000000000590000000000000027000000000000000600000000",
            INIT_3D => X"000000530000000000000048000000000000005e000000000000002a00000000",
            INIT_3E => X"00000078000000000000007200000000000000a2000000000000008300000000",
            INIT_3F => X"0000001500000000000000340000000000000085000000000000007600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006800000000000000310000000000000035000000000000004900000000",
            INIT_41 => X"0000004600000000000000390000000000000058000000000000007900000000",
            INIT_42 => X"0000005300000000000000470000000000000017000000000000003300000000",
            INIT_43 => X"000000070000000000000022000000000000004f000000000000004e00000000",
            INIT_44 => X"0000003e000000000000003c0000000000000051000000000000002800000000",
            INIT_45 => X"0000005d000000000000005b0000000000000063000000000000005000000000",
            INIT_46 => X"000000790000000000000078000000000000008d000000000000007300000000",
            INIT_47 => X"000000140000000000000021000000000000007c000000000000007900000000",
            INIT_48 => X"000000760000000000000038000000000000003a000000000000005600000000",
            INIT_49 => X"000000330000000000000040000000000000007f000000000000008300000000",
            INIT_4A => X"0000006300000000000000610000000000000040000000000000003b00000000",
            INIT_4B => X"0000001c000000000000000d000000000000003a000000000000005e00000000",
            INIT_4C => X"000000500000000000000049000000000000005d000000000000005300000000",
            INIT_4D => X"0000004a000000000000005f0000000000000069000000000000006200000000",
            INIT_4E => X"0000007e00000000000000770000000000000084000000000000007400000000",
            INIT_4F => X"00000017000000000000000d0000000000000065000000000000007f00000000",
            INIT_50 => X"000000740000000000000035000000000000003b000000000000005b00000000",
            INIT_51 => X"0000003000000000000000670000000000000087000000000000008400000000",
            INIT_52 => X"000000610000000000000060000000000000004b000000000000002000000000",
            INIT_53 => X"000000490000000000000032000000000000004a000000000000006600000000",
            INIT_54 => X"0000006100000000000000590000000000000052000000000000005a00000000",
            INIT_55 => X"000000310000000000000047000000000000006c000000000000006200000000",
            INIT_56 => X"0000008a0000000000000077000000000000007c000000000000007700000000",
            INIT_57 => X"00000014000000000000000a000000000000005b000000000000007b00000000",
            INIT_58 => X"0000006e000000000000002f0000000000000033000000000000006500000000",
            INIT_59 => X"0000004800000000000000870000000000000087000000000000008100000000",
            INIT_5A => X"0000004f00000000000000520000000000000054000000000000002e00000000",
            INIT_5B => X"0000008700000000000000750000000000000056000000000000005e00000000",
            INIT_5C => X"0000005e000000000000005d0000000000000066000000000000007800000000",
            INIT_5D => X"00000058000000000000004a0000000000000058000000000000005c00000000",
            INIT_5E => X"0000008d00000000000000760000000000000073000000000000008400000000",
            INIT_5F => X"00000007000000000000000b000000000000005b000000000000007700000000",
            INIT_60 => X"0000006000000000000000280000000000000028000000000000005800000000",
            INIT_61 => X"00000077000000000000008b0000000000000083000000000000006b00000000",
            INIT_62 => X"0000005900000000000000570000000000000066000000000000006b00000000",
            INIT_63 => X"0000006c0000000000000051000000000000004a000000000000005f00000000",
            INIT_64 => X"0000005d0000000000000064000000000000006e000000000000007600000000",
            INIT_65 => X"0000005f00000000000000570000000000000055000000000000006600000000",
            INIT_66 => X"0000007100000000000000650000000000000078000000000000007c00000000",
            INIT_67 => X"00000020000000000000000f0000000000000059000000000000007b00000000",
            INIT_68 => X"0000005c0000000000000037000000000000003f000000000000005f00000000",
            INIT_69 => X"00000089000000000000008b000000000000006e000000000000006400000000",
            INIT_6A => X"0000005c00000000000000650000000000000061000000000000007b00000000",
            INIT_6B => X"0000005600000000000000560000000000000058000000000000005a00000000",
            INIT_6C => X"0000006c00000000000000640000000000000058000000000000005500000000",
            INIT_6D => X"0000005f000000000000006e000000000000006c000000000000007200000000",
            INIT_6E => X"00000073000000000000006b0000000000000075000000000000006d00000000",
            INIT_6F => X"0000004c00000000000000310000000000000058000000000000008000000000",
            INIT_70 => X"0000006000000000000000470000000000000045000000000000006a00000000",
            INIT_71 => X"0000008700000000000000860000000000000056000000000000006800000000",
            INIT_72 => X"0000005800000000000000510000000000000057000000000000007400000000",
            INIT_73 => X"0000006a000000000000006e0000000000000060000000000000006000000000",
            INIT_74 => X"0000005c0000000000000057000000000000005f000000000000006200000000",
            INIT_75 => X"00000080000000000000007f000000000000006b000000000000006100000000",
            INIT_76 => X"000000770000000000000074000000000000005e000000000000007a00000000",
            INIT_77 => X"000000460000000000000035000000000000005c000000000000007a00000000",
            INIT_78 => X"0000005c00000000000000400000000000000040000000000000006000000000",
            INIT_79 => X"000000850000000000000079000000000000005f000000000000006700000000",
            INIT_7A => X"0000003300000000000000640000000000000096000000000000008100000000",
            INIT_7B => X"0000007100000000000000620000000000000065000000000000005800000000",
            INIT_7C => X"0000005f00000000000000650000000000000077000000000000008300000000",
            INIT_7D => X"0000009800000000000000710000000000000053000000000000006000000000",
            INIT_7E => X"0000007c00000000000000620000000000000078000000000000009400000000",
            INIT_7F => X"00000048000000000000000d0000000000000039000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "sampleifmap_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005a0000000000000047000000000000004c000000000000005700000000",
            INIT_01 => X"000000820000000000000078000000000000007c000000000000007300000000",
            INIT_02 => X"0000003a0000000000000096000000000000008e000000000000006e00000000",
            INIT_03 => X"0000007800000000000000770000000000000074000000000000005400000000",
            INIT_04 => X"0000008600000000000000850000000000000071000000000000006c00000000",
            INIT_05 => X"0000006e0000000000000067000000000000007e000000000000008900000000",
            INIT_06 => X"00000072000000000000006300000000000000a3000000000000009f00000000",
            INIT_07 => X"0000006b0000000000000021000000000000002a000000000000007500000000",
            INIT_08 => X"0000005d00000000000000640000000000000058000000000000005600000000",
            INIT_09 => X"0000006900000000000000750000000000000063000000000000007500000000",
            INIT_0A => X"0000008b000000000000009b0000000000000066000000000000006e00000000",
            INIT_0B => X"000000810000000000000081000000000000006f000000000000006b00000000",
            INIT_0C => X"00000076000000000000006d0000000000000077000000000000007c00000000",
            INIT_0D => X"00000071000000000000007c0000000000000076000000000000007100000000",
            INIT_0E => X"0000006300000000000000830000000000000075000000000000008300000000",
            INIT_0F => X"0000005700000000000000270000000000000048000000000000006900000000",
            INIT_10 => X"0000007300000000000000780000000000000060000000000000005f00000000",
            INIT_11 => X"0000005600000000000000630000000000000047000000000000006d00000000",
            INIT_12 => X"000000b0000000000000006a0000000000000063000000000000006c00000000",
            INIT_13 => X"00000075000000000000007b000000000000005e000000000000008200000000",
            INIT_14 => X"000000880000000000000081000000000000008d000000000000008900000000",
            INIT_15 => X"000000790000000000000078000000000000006f000000000000008300000000",
            INIT_16 => X"000000430000000000000050000000000000006b000000000000007500000000",
            INIT_17 => X"0000006e00000000000000430000000000000051000000000000004800000000",
            INIT_18 => X"00000057000000000000007d0000000000000070000000000000006d00000000",
            INIT_19 => X"0000005e00000000000000470000000000000048000000000000005800000000",
            INIT_1A => X"0000007300000000000000490000000000000079000000000000006400000000",
            INIT_1B => X"0000009400000000000000870000000000000076000000000000009800000000",
            INIT_1C => X"0000009500000000000000940000000000000082000000000000008500000000",
            INIT_1D => X"0000007a00000000000000790000000000000071000000000000007d00000000",
            INIT_1E => X"0000004e000000000000003a0000000000000071000000000000007200000000",
            INIT_1F => X"0000008a00000000000000730000000000000038000000000000003d00000000",
            INIT_20 => X"0000004300000000000000590000000000000074000000000000007700000000",
            INIT_21 => X"00000066000000000000003c0000000000000048000000000000005800000000",
            INIT_22 => X"00000037000000000000006d0000000000000057000000000000004800000000",
            INIT_23 => X"0000009c000000000000008d0000000000000092000000000000006500000000",
            INIT_24 => X"00000098000000000000008c0000000000000088000000000000009800000000",
            INIT_25 => X"0000007c000000000000007f000000000000007b000000000000008600000000",
            INIT_26 => X"00000062000000000000005d0000000000000069000000000000006d00000000",
            INIT_27 => X"00000077000000000000007a0000000000000062000000000000004d00000000",
            INIT_28 => X"0000005d00000000000000320000000000000061000000000000007e00000000",
            INIT_29 => X"00000060000000000000004b0000000000000046000000000000006000000000",
            INIT_2A => X"000000610000000000000076000000000000003b000000000000005a00000000",
            INIT_2B => X"0000009700000000000000a20000000000000083000000000000004900000000",
            INIT_2C => X"0000007f000000000000008400000000000000a3000000000000009600000000",
            INIT_2D => X"00000075000000000000006e0000000000000076000000000000007d00000000",
            INIT_2E => X"0000004f000000000000005e0000000000000066000000000000006900000000",
            INIT_2F => X"0000006a0000000000000070000000000000008e000000000000006b00000000",
            INIT_30 => X"0000005900000000000000370000000000000051000000000000007000000000",
            INIT_31 => X"000000590000000000000045000000000000004e000000000000005c00000000",
            INIT_32 => X"000000760000000000000053000000000000006b000000000000007700000000",
            INIT_33 => X"0000009c0000000000000097000000000000007d000000000000006b00000000",
            INIT_34 => X"0000007e0000000000000094000000000000009b000000000000009400000000",
            INIT_35 => X"000000750000000000000078000000000000007b000000000000006c00000000",
            INIT_36 => X"0000005600000000000000540000000000000066000000000000007200000000",
            INIT_37 => X"0000006900000000000000630000000000000079000000000000008100000000",
            INIT_38 => X"0000009a00000000000000780000000000000056000000000000006200000000",
            INIT_39 => X"0000004e0000000000000045000000000000005f000000000000007700000000",
            INIT_3A => X"0000004e0000000000000057000000000000007e000000000000007300000000",
            INIT_3B => X"000000960000000000000084000000000000008b000000000000007d00000000",
            INIT_3C => X"0000007e0000000000000092000000000000008e000000000000008d00000000",
            INIT_3D => X"0000007b00000000000000760000000000000084000000000000007900000000",
            INIT_3E => X"0000006f00000000000000520000000000000058000000000000007300000000",
            INIT_3F => X"00000067000000000000006a0000000000000065000000000000007900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a70000000000000088000000000000007400000000",
            INIT_41 => X"0000005c00000000000000600000000000000077000000000000009f00000000",
            INIT_42 => X"0000006f0000000000000066000000000000005a000000000000006600000000",
            INIT_43 => X"0000008f00000000000000830000000000000088000000000000007000000000",
            INIT_44 => X"000000800000000000000096000000000000008e000000000000008600000000",
            INIT_45 => X"000000770000000000000084000000000000009c000000000000007500000000",
            INIT_46 => X"00000053000000000000004e0000000000000059000000000000006600000000",
            INIT_47 => X"0000006c00000000000000710000000000000060000000000000006a00000000",
            INIT_48 => X"000000920000000000000071000000000000006d000000000000006c00000000",
            INIT_49 => X"00000069000000000000007b000000000000009e00000000000000a600000000",
            INIT_4A => X"0000008c00000000000000550000000000000052000000000000006600000000",
            INIT_4B => X"0000007b0000000000000086000000000000007e000000000000009100000000",
            INIT_4C => X"00000089000000000000008a0000000000000073000000000000006800000000",
            INIT_4D => X"0000006a000000000000008a0000000000000096000000000000008300000000",
            INIT_4E => X"0000002d000000000000004a000000000000006f000000000000006100000000",
            INIT_4F => X"0000004b00000000000000690000000000000065000000000000006000000000",
            INIT_50 => X"0000005600000000000000370000000000000055000000000000005800000000",
            INIT_51 => X"0000007e00000000000000970000000000000097000000000000008b00000000",
            INIT_52 => X"0000005700000000000000570000000000000068000000000000006800000000",
            INIT_53 => X"00000052000000000000006e000000000000006e000000000000006f00000000",
            INIT_54 => X"0000008c0000000000000079000000000000004b000000000000003500000000",
            INIT_55 => X"0000007a00000000000000810000000000000078000000000000009100000000",
            INIT_56 => X"00000020000000000000003e0000000000000062000000000000007400000000",
            INIT_57 => X"0000004000000000000000410000000000000062000000000000006100000000",
            INIT_58 => X"000000200000000000000022000000000000005c000000000000005200000000",
            INIT_59 => X"0000009c00000000000000860000000000000075000000000000004b00000000",
            INIT_5A => X"000000570000000000000062000000000000006d000000000000008d00000000",
            INIT_5B => X"0000005f000000000000005b000000000000005a000000000000005200000000",
            INIT_5C => X"0000008b00000000000000790000000000000046000000000000005200000000",
            INIT_5D => X"0000006b0000000000000080000000000000008f000000000000008100000000",
            INIT_5E => X"0000003f000000000000001d000000000000004e000000000000007100000000",
            INIT_5F => X"0000004200000000000000470000000000000047000000000000006300000000",
            INIT_60 => X"0000000d00000000000000230000000000000056000000000000005a00000000",
            INIT_61 => X"000000940000000000000072000000000000004e000000000000000f00000000",
            INIT_62 => X"00000062000000000000006f000000000000008b00000000000000a200000000",
            INIT_63 => X"000000710000000000000056000000000000005b000000000000006100000000",
            INIT_64 => X"0000007e0000000000000073000000000000006a000000000000007800000000",
            INIT_65 => X"0000006a00000000000000870000000000000087000000000000007600000000",
            INIT_66 => X"0000005b0000000000000026000000000000002a000000000000004f00000000",
            INIT_67 => X"0000005300000000000000990000000000000060000000000000002c00000000",
            INIT_68 => X"00000025000000000000002d0000000000000056000000000000005c00000000",
            INIT_69 => X"0000007a0000000000000057000000000000001f000000000000000d00000000",
            INIT_6A => X"0000007a000000000000009e00000000000000ad000000000000009600000000",
            INIT_6B => X"0000005c000000000000005d0000000000000072000000000000007500000000",
            INIT_6C => X"0000007100000000000000670000000000000055000000000000004d00000000",
            INIT_6D => X"0000005b00000000000000730000000000000085000000000000007e00000000",
            INIT_6E => X"0000003c000000000000003b0000000000000032000000000000004e00000000",
            INIT_6F => X"000000620000000000000086000000000000006c000000000000002a00000000",
            INIT_70 => X"0000003800000000000000180000000000000047000000000000005200000000",
            INIT_71 => X"0000005400000000000000230000000000000017000000000000002400000000",
            INIT_72 => X"000000a500000000000000a50000000000000092000000000000007600000000",
            INIT_73 => X"00000079000000000000006f0000000000000082000000000000009600000000",
            INIT_74 => X"00000062000000000000003f0000000000000042000000000000006c00000000",
            INIT_75 => X"0000005600000000000000460000000000000045000000000000004e00000000",
            INIT_76 => X"000000620000000000000060000000000000006c000000000000007500000000",
            INIT_77 => X"00000059000000000000007b0000000000000074000000000000007800000000",
            INIT_78 => X"000000400000000000000011000000000000001b000000000000004100000000",
            INIT_79 => X"00000025000000000000000f000000000000001d000000000000003400000000",
            INIT_7A => X"0000009600000000000000740000000000000064000000000000005900000000",
            INIT_7B => X"0000009c0000000000000088000000000000009800000000000000aa00000000",
            INIT_7C => X"0000004a0000000000000045000000000000007900000000000000a600000000",
            INIT_7D => X"0000007f00000000000000660000000000000047000000000000002f00000000",
            INIT_7E => X"000000820000000000000083000000000000008b000000000000009c00000000",
            INIT_7F => X"0000007500000000000000920000000000000088000000000000009300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "sampleifmap_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000058000000000000004d000000000000008b00000000000000b300000000",
            INIT_01 => X"00000097000000000000009c000000000000009d000000000000008d00000000",
            INIT_02 => X"000000970000000000000090000000000000009e000000000000009c00000000",
            INIT_03 => X"0000007600000000000000790000000000000088000000000000009700000000",
            INIT_04 => X"000000540000000000000054000000000000006c000000000000007e00000000",
            INIT_05 => X"00000053000000000000005e0000000000000062000000000000006200000000",
            INIT_06 => X"0000006000000000000000540000000000000056000000000000005a00000000",
            INIT_07 => X"0000004d000000000000004c0000000000000057000000000000007500000000",
            INIT_08 => X"000000920000000000000080000000000000008500000000000000b800000000",
            INIT_09 => X"000000a7000000000000009e000000000000009f000000000000009f00000000",
            INIT_0A => X"0000009a000000000000009900000000000000a200000000000000a500000000",
            INIT_0B => X"0000007d00000000000000880000000000000096000000000000009600000000",
            INIT_0C => X"00000052000000000000005a000000000000006d000000000000008100000000",
            INIT_0D => X"00000058000000000000005e0000000000000062000000000000005d00000000",
            INIT_0E => X"0000006a000000000000005b000000000000004c000000000000004e00000000",
            INIT_0F => X"0000005a000000000000005b0000000000000062000000000000007600000000",
            INIT_10 => X"000000aa00000000000000b0000000000000009800000000000000b400000000",
            INIT_11 => X"000000a4000000000000009b000000000000009800000000000000a400000000",
            INIT_12 => X"0000009f00000000000000a200000000000000aa00000000000000a200000000",
            INIT_13 => X"0000008c00000000000000920000000000000097000000000000009c00000000",
            INIT_14 => X"000000470000000000000058000000000000007c000000000000009200000000",
            INIT_15 => X"0000006b00000000000000670000000000000062000000000000005500000000",
            INIT_16 => X"0000006f000000000000006f000000000000006d000000000000006500000000",
            INIT_17 => X"0000005f000000000000005d0000000000000065000000000000006f00000000",
            INIT_18 => X"000000b500000000000000b800000000000000ae00000000000000af00000000",
            INIT_19 => X"000000a300000000000000a4000000000000009800000000000000a800000000",
            INIT_1A => X"000000a800000000000000a700000000000000b300000000000000a600000000",
            INIT_1B => X"000000a4000000000000009f00000000000000a200000000000000ae00000000",
            INIT_1C => X"0000003a00000000000000590000000000000089000000000000009700000000",
            INIT_1D => X"0000006b0000000000000063000000000000005a000000000000004800000000",
            INIT_1E => X"00000079000000000000007d0000000000000080000000000000007500000000",
            INIT_1F => X"0000006f000000000000006d0000000000000061000000000000006900000000",
            INIT_20 => X"000000ac00000000000000a700000000000000ae00000000000000af00000000",
            INIT_21 => X"000000af00000000000000b000000000000000a100000000000000a200000000",
            INIT_22 => X"000000b400000000000000b300000000000000b200000000000000b200000000",
            INIT_23 => X"000000a400000000000000a000000000000000a800000000000000b000000000",
            INIT_24 => X"000000450000000000000078000000000000009c00000000000000ad00000000",
            INIT_25 => X"0000005e0000000000000063000000000000005a000000000000004200000000",
            INIT_26 => X"0000007b000000000000007f000000000000007c000000000000006900000000",
            INIT_27 => X"0000007400000000000000710000000000000068000000000000007000000000",
            INIT_28 => X"000000aa000000000000009000000000000000ae00000000000000b500000000",
            INIT_29 => X"000000b300000000000000b000000000000000a600000000000000a900000000",
            INIT_2A => X"000000b500000000000000b400000000000000b400000000000000b400000000",
            INIT_2B => X"00000096000000000000009f00000000000000ae00000000000000b000000000",
            INIT_2C => X"00000074000000000000009b00000000000000af00000000000000b500000000",
            INIT_2D => X"000000700000000000000083000000000000007d000000000000006000000000",
            INIT_2E => X"00000079000000000000007a0000000000000078000000000000007500000000",
            INIT_2F => X"0000007c00000000000000760000000000000078000000000000007900000000",
            INIT_30 => X"000000b2000000000000008a000000000000009c00000000000000c000000000",
            INIT_31 => X"000000af00000000000000b000000000000000ae00000000000000af00000000",
            INIT_32 => X"000000b800000000000000ba00000000000000b400000000000000b800000000",
            INIT_33 => X"0000009900000000000000ad00000000000000bb00000000000000bb00000000",
            INIT_34 => X"000000a700000000000000ad00000000000000ad00000000000000a600000000",
            INIT_35 => X"0000007900000000000000940000000000000095000000000000009600000000",
            INIT_36 => X"0000006f000000000000006d0000000000000075000000000000007300000000",
            INIT_37 => X"00000080000000000000007b000000000000007a000000000000007800000000",
            INIT_38 => X"000000ab000000000000009c000000000000007d00000000000000b900000000",
            INIT_39 => X"000000b800000000000000af00000000000000af00000000000000ad00000000",
            INIT_3A => X"000000c200000000000000c100000000000000b700000000000000bc00000000",
            INIT_3B => X"000000a600000000000000b800000000000000b900000000000000bd00000000",
            INIT_3C => X"000000b000000000000000b100000000000000ac00000000000000a400000000",
            INIT_3D => X"0000007a000000000000008f000000000000008900000000000000aa00000000",
            INIT_3E => X"000000670000000000000060000000000000006e000000000000006b00000000",
            INIT_3F => X"0000007d000000000000007b0000000000000076000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a0000000000000009f0000000000000095000000000000009b00000000",
            INIT_41 => X"000000b400000000000000b200000000000000ad00000000000000ac00000000",
            INIT_42 => X"000000bf00000000000000ba00000000000000ba00000000000000bb00000000",
            INIT_43 => X"000000a000000000000000ac00000000000000af00000000000000bb00000000",
            INIT_44 => X"000000b000000000000000a60000000000000097000000000000009a00000000",
            INIT_45 => X"0000008500000000000000a6000000000000009b00000000000000b700000000",
            INIT_46 => X"0000007700000000000000700000000000000068000000000000006800000000",
            INIT_47 => X"0000007d000000000000007a000000000000007a000000000000007600000000",
            INIT_48 => X"000000a900000000000000930000000000000098000000000000009a00000000",
            INIT_49 => X"000000aa00000000000000b700000000000000b200000000000000b200000000",
            INIT_4A => X"000000c100000000000000c600000000000000bc00000000000000b000000000",
            INIT_4B => X"000000a900000000000000a500000000000000a700000000000000ae00000000",
            INIT_4C => X"000000a90000000000000092000000000000008c000000000000009d00000000",
            INIT_4D => X"0000008d00000000000000ab00000000000000a000000000000000b300000000",
            INIT_4E => X"0000007700000000000000750000000000000068000000000000005f00000000",
            INIT_4F => X"0000007d0000000000000076000000000000007b000000000000007400000000",
            INIT_50 => X"000000b1000000000000009f0000000000000070000000000000008600000000",
            INIT_51 => X"000000ba00000000000000b800000000000000b800000000000000ae00000000",
            INIT_52 => X"000000b000000000000000bf00000000000000c200000000000000ba00000000",
            INIT_53 => X"000000bb00000000000000a7000000000000009e000000000000009b00000000",
            INIT_54 => X"000000970000000000000086000000000000009300000000000000ae00000000",
            INIT_55 => X"0000007c000000000000009b000000000000009c00000000000000a000000000",
            INIT_56 => X"0000006600000000000000690000000000000066000000000000004a00000000",
            INIT_57 => X"0000007f000000000000007b0000000000000075000000000000006b00000000",
            INIT_58 => X"0000009d00000000000000ae000000000000005b000000000000004100000000",
            INIT_59 => X"000000be00000000000000bf00000000000000b1000000000000009300000000",
            INIT_5A => X"000000b000000000000000ac00000000000000b000000000000000bc00000000",
            INIT_5B => X"000000a3000000000000009400000000000000ae00000000000000b800000000",
            INIT_5C => X"000000950000000000000085000000000000009a00000000000000b000000000",
            INIT_5D => X"0000005000000000000000830000000000000095000000000000009800000000",
            INIT_5E => X"0000006600000000000000670000000000000061000000000000004200000000",
            INIT_5F => X"0000007d00000000000000780000000000000071000000000000006700000000",
            INIT_60 => X"000000b100000000000000bf000000000000005c000000000000001500000000",
            INIT_61 => X"000000b600000000000000bd00000000000000ca00000000000000bc00000000",
            INIT_62 => X"000000bc00000000000000a5000000000000009c00000000000000b300000000",
            INIT_63 => X"00000072000000000000009800000000000000ae00000000000000c800000000",
            INIT_64 => X"000000890000000000000078000000000000007f000000000000005f00000000",
            INIT_65 => X"0000004e00000000000000720000000000000088000000000000009700000000",
            INIT_66 => X"0000006200000000000000590000000000000049000000000000004000000000",
            INIT_67 => X"0000007600000000000000750000000000000071000000000000006200000000",
            INIT_68 => X"000000ad00000000000000a80000000000000063000000000000002c00000000",
            INIT_69 => X"000000bb00000000000000bc00000000000000c300000000000000c800000000",
            INIT_6A => X"000000c200000000000000b4000000000000009500000000000000a500000000",
            INIT_6B => X"0000009a00000000000000a800000000000000a800000000000000b900000000",
            INIT_6C => X"0000008a00000000000000910000000000000092000000000000006b00000000",
            INIT_6D => X"000000480000000000000064000000000000007f000000000000009c00000000",
            INIT_6E => X"0000006000000000000000530000000000000040000000000000003900000000",
            INIT_6F => X"0000006f000000000000006c000000000000006a000000000000006200000000",
            INIT_70 => X"0000009f00000000000000750000000000000076000000000000006900000000",
            INIT_71 => X"000000bb00000000000000b400000000000000be00000000000000c400000000",
            INIT_72 => X"000000c100000000000000c600000000000000ad00000000000000ad00000000",
            INIT_73 => X"000000bc00000000000000b400000000000000a500000000000000ab00000000",
            INIT_74 => X"000000b300000000000000ad00000000000000bb00000000000000ae00000000",
            INIT_75 => X"000000480000000000000069000000000000008000000000000000a000000000",
            INIT_76 => X"0000006c00000000000000570000000000000045000000000000004300000000",
            INIT_77 => X"0000006600000000000000610000000000000064000000000000006300000000",
            INIT_78 => X"0000009d00000000000000680000000000000071000000000000008a00000000",
            INIT_79 => X"000000a800000000000000b400000000000000c400000000000000c600000000",
            INIT_7A => X"000000cd00000000000000cb00000000000000bf00000000000000b400000000",
            INIT_7B => X"000000c800000000000000c400000000000000bf00000000000000d200000000",
            INIT_7C => X"000000be00000000000000bc00000000000000bb00000000000000c000000000",
            INIT_7D => X"000000500000000000000071000000000000009900000000000000a800000000",
            INIT_7E => X"0000008700000000000000600000000000000040000000000000004600000000",
            INIT_7F => X"00000062000000000000005a000000000000005a000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "sampleifmap_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000930000000000000073000000000000008a000000000000009600000000",
            INIT_01 => X"0000009600000000000000b000000000000000bb00000000000000be00000000",
            INIT_02 => X"000000c600000000000000d300000000000000c700000000000000ab00000000",
            INIT_03 => X"000000cb00000000000000be00000000000000c200000000000000d300000000",
            INIT_04 => X"000000bd00000000000000b800000000000000ba00000000000000bf00000000",
            INIT_05 => X"00000046000000000000006400000000000000a600000000000000be00000000",
            INIT_06 => X"0000008f000000000000006a0000000000000038000000000000002f00000000",
            INIT_07 => X"0000005e000000000000004a000000000000005c000000000000009500000000",
            INIT_08 => X"000000a50000000000000092000000000000009b000000000000009b00000000",
            INIT_09 => X"0000009100000000000000bf00000000000000c000000000000000bd00000000",
            INIT_0A => X"0000009500000000000000a900000000000000d2000000000000009c00000000",
            INIT_0B => X"000000a800000000000000b200000000000000c200000000000000c000000000",
            INIT_0C => X"000000a700000000000000aa00000000000000b500000000000000a900000000",
            INIT_0D => X"0000002b00000000000000430000000000000075000000000000009a00000000",
            INIT_0E => X"0000008f00000000000000680000000000000031000000000000002200000000",
            INIT_0F => X"00000050000000000000003f000000000000006a000000000000009c00000000",
            INIT_10 => X"000000a6000000000000008a00000000000000a200000000000000a500000000",
            INIT_11 => X"0000008900000000000000ba00000000000000be00000000000000c400000000",
            INIT_12 => X"000000a9000000000000009d00000000000000c9000000000000007400000000",
            INIT_13 => X"0000008f000000000000008000000000000000b600000000000000d200000000",
            INIT_14 => X"00000061000000000000007f0000000000000093000000000000007c00000000",
            INIT_15 => X"00000033000000000000002f0000000000000038000000000000005200000000",
            INIT_16 => X"0000009d00000000000000690000000000000040000000000000002b00000000",
            INIT_17 => X"000000410000000000000039000000000000007b000000000000009d00000000",
            INIT_18 => X"0000009e0000000000000078000000000000009600000000000000a900000000",
            INIT_19 => X"0000009800000000000000be00000000000000be00000000000000be00000000",
            INIT_1A => X"000000b900000000000000bc0000000000000099000000000000003c00000000",
            INIT_1B => X"000000ce000000000000009000000000000000a500000000000000c300000000",
            INIT_1C => X"0000003d0000000000000065000000000000008900000000000000b100000000",
            INIT_1D => X"0000005000000000000000470000000000000033000000000000003700000000",
            INIT_1E => X"000000a0000000000000006e000000000000004a000000000000003700000000",
            INIT_1F => X"000000320000000000000036000000000000008e00000000000000b000000000",
            INIT_20 => X"000000a6000000000000009600000000000000a000000000000000aa00000000",
            INIT_21 => X"0000009a00000000000000ba00000000000000bc00000000000000ba00000000",
            INIT_22 => X"00000092000000000000007e0000000000000031000000000000002000000000",
            INIT_23 => X"000000c0000000000000008c000000000000008c000000000000009b00000000",
            INIT_24 => X"0000003e0000000000000061000000000000009c00000000000000cc00000000",
            INIT_25 => X"0000005700000000000000520000000000000049000000000000004900000000",
            INIT_26 => X"000000a6000000000000006b000000000000003e000000000000003a00000000",
            INIT_27 => X"00000033000000000000004800000000000000a700000000000000bc00000000",
            INIT_28 => X"0000009c000000000000009700000000000000ab00000000000000b200000000",
            INIT_29 => X"0000007c00000000000000a300000000000000b200000000000000b500000000",
            INIT_2A => X"000000370000000000000028000000000000001d000000000000002400000000",
            INIT_2B => X"0000008200000000000000650000000000000063000000000000004e00000000",
            INIT_2C => X"00000037000000000000005f000000000000007b000000000000009000000000",
            INIT_2D => X"00000055000000000000003c0000000000000033000000000000003400000000",
            INIT_2E => X"000000990000000000000066000000000000004d000000000000004e00000000",
            INIT_2F => X"00000037000000000000005900000000000000b100000000000000bb00000000",
            INIT_30 => X"00000098000000000000009200000000000000ab00000000000000b500000000",
            INIT_31 => X"00000069000000000000009500000000000000a700000000000000a900000000",
            INIT_32 => X"0000002e0000000000000042000000000000005e000000000000004f00000000",
            INIT_33 => X"00000078000000000000005c0000000000000047000000000000002f00000000",
            INIT_34 => X"0000002900000000000000380000000000000037000000000000005a00000000",
            INIT_35 => X"00000037000000000000001e0000000000000022000000000000002300000000",
            INIT_36 => X"0000007700000000000000610000000000000056000000000000005200000000",
            INIT_37 => X"0000003c000000000000006a00000000000000ae00000000000000ad00000000",
            INIT_38 => X"000000a3000000000000009e000000000000009c00000000000000b100000000",
            INIT_39 => X"00000089000000000000009400000000000000a0000000000000009c00000000",
            INIT_3A => X"0000006b00000000000000660000000000000076000000000000008f00000000",
            INIT_3B => X"00000067000000000000007d000000000000006d000000000000006e00000000",
            INIT_3C => X"0000001300000000000000100000000000000011000000000000002f00000000",
            INIT_3D => X"00000013000000000000000e000000000000001c000000000000001800000000",
            INIT_3E => X"0000006300000000000000600000000000000041000000000000002b00000000",
            INIT_3F => X"00000043000000000000008500000000000000ad000000000000008c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a7000000000000008b000000000000009e00000000",
            INIT_41 => X"000000c000000000000000ab000000000000008c000000000000009700000000",
            INIT_42 => X"000000880000000000000085000000000000007400000000000000ac00000000",
            INIT_43 => X"00000065000000000000007f000000000000008d000000000000009200000000",
            INIT_44 => X"0000001900000000000000200000000000000025000000000000004100000000",
            INIT_45 => X"0000000f000000000000000a0000000000000011000000000000001800000000",
            INIT_46 => X"0000004e00000000000000610000000000000042000000000000001400000000",
            INIT_47 => X"00000069000000000000009c0000000000000094000000000000006200000000",
            INIT_48 => X"000000ab00000000000000ae00000000000000a400000000000000a000000000",
            INIT_49 => X"000000b100000000000000940000000000000088000000000000009e00000000",
            INIT_4A => X"0000009700000000000000a9000000000000009300000000000000b800000000",
            INIT_4B => X"0000007d000000000000008e000000000000008b000000000000007f00000000",
            INIT_4C => X"0000002b000000000000003f000000000000004d000000000000006700000000",
            INIT_4D => X"0000001a00000000000000110000000000000018000000000000002100000000",
            INIT_4E => X"000000320000000000000048000000000000003e000000000000001f00000000",
            INIT_4F => X"000000880000000000000078000000000000005a000000000000004800000000",
            INIT_50 => X"000000a700000000000000a700000000000000a300000000000000a000000000",
            INIT_51 => X"00000078000000000000008c00000000000000a800000000000000b100000000",
            INIT_52 => X"000000820000000000000076000000000000008f00000000000000ab00000000",
            INIT_53 => X"0000009100000000000000a6000000000000009c000000000000007b00000000",
            INIT_54 => X"0000004e000000000000005b0000000000000069000000000000007c00000000",
            INIT_55 => X"0000004300000000000000380000000000000042000000000000004c00000000",
            INIT_56 => X"0000004900000000000000410000000000000041000000000000004600000000",
            INIT_57 => X"0000006a0000000000000051000000000000007b000000000000006400000000",
            INIT_58 => X"00000093000000000000008c000000000000009f000000000000009c00000000",
            INIT_59 => X"0000007b000000000000009900000000000000aa00000000000000b400000000",
            INIT_5A => X"0000007e0000000000000073000000000000009c000000000000008b00000000",
            INIT_5B => X"000000a200000000000000a8000000000000009e000000000000008300000000",
            INIT_5C => X"00000078000000000000007b0000000000000077000000000000007f00000000",
            INIT_5D => X"0000007700000000000000690000000000000068000000000000007000000000",
            INIT_5E => X"0000006d00000000000000680000000000000069000000000000007400000000",
            INIT_5F => X"00000068000000000000005c0000000000000086000000000000007a00000000",
            INIT_60 => X"0000008b000000000000007b000000000000009e00000000000000a400000000",
            INIT_61 => X"0000008c000000000000008d000000000000009c00000000000000ad00000000",
            INIT_62 => X"000000a100000000000000820000000000000079000000000000008d00000000",
            INIT_63 => X"000000a800000000000000a6000000000000009d000000000000009700000000",
            INIT_64 => X"00000084000000000000008f000000000000008a000000000000009000000000",
            INIT_65 => X"00000094000000000000008a0000000000000085000000000000008100000000",
            INIT_66 => X"0000008400000000000000860000000000000089000000000000008f00000000",
            INIT_67 => X"0000009300000000000000730000000000000064000000000000007800000000",
            INIT_68 => X"000000a800000000000000900000000000000095000000000000008e00000000",
            INIT_69 => X"0000009e000000000000009e00000000000000a100000000000000a700000000",
            INIT_6A => X"000000a90000000000000097000000000000009000000000000000a500000000",
            INIT_6B => X"000000a2000000000000009e00000000000000a000000000000000a100000000",
            INIT_6C => X"0000007f00000000000000890000000000000091000000000000009900000000",
            INIT_6D => X"0000009e00000000000000960000000000000095000000000000008d00000000",
            INIT_6E => X"0000008f00000000000000940000000000000096000000000000009f00000000",
            INIT_6F => X"0000009f000000000000008b0000000000000077000000000000007b00000000",
            INIT_70 => X"000000b900000000000000b300000000000000a6000000000000009800000000",
            INIT_71 => X"000000a800000000000000aa00000000000000a700000000000000a700000000",
            INIT_72 => X"000000b200000000000000ad00000000000000a400000000000000a700000000",
            INIT_73 => X"000000850000000000000089000000000000009d00000000000000a900000000",
            INIT_74 => X"00000088000000000000008c000000000000008f000000000000009200000000",
            INIT_75 => X"0000009d00000000000000980000000000000097000000000000008c00000000",
            INIT_76 => X"000000900000000000000099000000000000009c00000000000000a600000000",
            INIT_77 => X"0000009900000000000000900000000000000083000000000000008500000000",
            INIT_78 => X"000000ab00000000000000b700000000000000b2000000000000009f00000000",
            INIT_79 => X"0000009f0000000000000091000000000000007d000000000000008b00000000",
            INIT_7A => X"0000009c0000000000000095000000000000008b00000000000000a200000000",
            INIT_7B => X"0000007300000000000000830000000000000098000000000000009e00000000",
            INIT_7C => X"0000008f0000000000000094000000000000008e000000000000008400000000",
            INIT_7D => X"000000a1000000000000009c000000000000009d000000000000009000000000",
            INIT_7E => X"0000009c0000000000000094000000000000009f00000000000000a700000000",
            INIT_7F => X"0000009800000000000000990000000000000096000000000000009c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "sampleifmap_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000000000310000000000000060000000000000007600000000",
            INIT_01 => X"000000530000000000000054000000000000005f000000000000006000000000",
            INIT_02 => X"0000005a00000000000000530000000000000061000000000000005f00000000",
            INIT_03 => X"0000004f000000000000004b0000000000000052000000000000005c00000000",
            INIT_04 => X"00000032000000000000003b0000000000000050000000000000005b00000000",
            INIT_05 => X"0000003300000000000000380000000000000038000000000000003700000000",
            INIT_06 => X"0000003a00000000000000330000000000000038000000000000003c00000000",
            INIT_07 => X"0000002f000000000000002f0000000000000035000000000000004c00000000",
            INIT_08 => X"0000006900000000000000590000000000000058000000000000008200000000",
            INIT_09 => X"00000068000000000000005d0000000000000060000000000000006c00000000",
            INIT_0A => X"0000005b000000000000005a0000000000000062000000000000006500000000",
            INIT_0B => X"00000048000000000000004f0000000000000057000000000000005400000000",
            INIT_0C => X"00000032000000000000003d0000000000000048000000000000005200000000",
            INIT_0D => X"0000003300000000000000370000000000000038000000000000003700000000",
            INIT_0E => X"0000004100000000000000350000000000000028000000000000002b00000000",
            INIT_0F => X"00000039000000000000003a000000000000003d000000000000004b00000000",
            INIT_10 => X"0000007a00000000000000810000000000000068000000000000008400000000",
            INIT_11 => X"0000006a000000000000005f0000000000000059000000000000006c00000000",
            INIT_12 => X"0000005e00000000000000620000000000000069000000000000006200000000",
            INIT_13 => X"0000004c000000000000004f0000000000000050000000000000005500000000",
            INIT_14 => X"0000002a0000000000000036000000000000004c000000000000005500000000",
            INIT_15 => X"00000042000000000000003f000000000000003a000000000000003300000000",
            INIT_16 => X"0000004200000000000000430000000000000042000000000000003c00000000",
            INIT_17 => X"000000390000000000000038000000000000003e000000000000004300000000",
            INIT_18 => X"000000840000000000000088000000000000007f000000000000008100000000",
            INIT_19 => X"000000690000000000000068000000000000005a000000000000007000000000",
            INIT_1A => X"0000006600000000000000650000000000000071000000000000006500000000",
            INIT_1B => X"0000005d0000000000000057000000000000005a000000000000006700000000",
            INIT_1C => X"0000001f0000000000000033000000000000004e000000000000004f00000000",
            INIT_1D => X"0000003e00000000000000390000000000000033000000000000002a00000000",
            INIT_1E => X"0000004a000000000000004b000000000000004d000000000000004600000000",
            INIT_1F => X"0000004500000000000000430000000000000037000000000000003c00000000",
            INIT_20 => X"0000007f0000000000000079000000000000007f000000000000008000000000",
            INIT_21 => X"0000007200000000000000720000000000000063000000000000006d00000000",
            INIT_22 => X"000000710000000000000070000000000000006f000000000000006f00000000",
            INIT_23 => X"0000005c00000000000000590000000000000063000000000000006c00000000",
            INIT_24 => X"0000002c000000000000004e0000000000000059000000000000005e00000000",
            INIT_25 => X"0000002e00000000000000380000000000000034000000000000002700000000",
            INIT_26 => X"0000004900000000000000470000000000000043000000000000003500000000",
            INIT_27 => X"000000470000000000000045000000000000003b000000000000004200000000",
            INIT_28 => X"0000007f00000000000000680000000000000083000000000000008900000000",
            INIT_29 => X"000000740000000000000071000000000000006a000000000000007600000000",
            INIT_2A => X"0000007100000000000000740000000000000075000000000000007300000000",
            INIT_2B => X"00000054000000000000005a0000000000000069000000000000006d00000000",
            INIT_2C => X"0000004f00000000000000670000000000000068000000000000006a00000000",
            INIT_2D => X"0000003d0000000000000052000000000000004d000000000000003a00000000",
            INIT_2E => X"000000460000000000000043000000000000003f000000000000003e00000000",
            INIT_2F => X"0000004b00000000000000460000000000000048000000000000004900000000",
            INIT_30 => X"0000008700000000000000660000000000000077000000000000009800000000",
            INIT_31 => X"0000006f00000000000000730000000000000075000000000000007a00000000",
            INIT_32 => X"00000070000000000000007c000000000000007b000000000000007900000000",
            INIT_33 => X"0000005c00000000000000660000000000000071000000000000007300000000",
            INIT_34 => X"0000006e000000000000006d0000000000000065000000000000006400000000",
            INIT_35 => X"00000043000000000000005b0000000000000057000000000000005c00000000",
            INIT_36 => X"0000003b00000000000000380000000000000040000000000000003e00000000",
            INIT_37 => X"0000004e000000000000004a0000000000000048000000000000004500000000",
            INIT_38 => X"0000007e00000000000000780000000000000059000000000000009300000000",
            INIT_39 => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_3A => X"00000073000000000000007c000000000000007a000000000000008000000000",
            INIT_3B => X"00000064000000000000006c000000000000006d000000000000007300000000",
            INIT_3C => X"0000006a000000000000006d0000000000000068000000000000006500000000",
            INIT_3D => X"000000480000000000000057000000000000004b000000000000006600000000",
            INIT_3E => X"00000035000000000000002e000000000000003c000000000000003b00000000",
            INIT_3F => X"0000004b00000000000000490000000000000044000000000000004200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000720000000000000078000000000000006f000000000000007600000000",
            INIT_41 => X"0000007700000000000000750000000000000074000000000000007700000000",
            INIT_42 => X"0000006d000000000000006f000000000000007a000000000000008000000000",
            INIT_43 => X"0000005e00000000000000610000000000000067000000000000007300000000",
            INIT_44 => X"0000006400000000000000610000000000000059000000000000005e00000000",
            INIT_45 => X"000000590000000000000072000000000000005f000000000000006d00000000",
            INIT_46 => X"000000470000000000000040000000000000003a000000000000003e00000000",
            INIT_47 => X"0000004b00000000000000480000000000000048000000000000004600000000",
            INIT_48 => X"0000007800000000000000690000000000000071000000000000007700000000",
            INIT_49 => X"0000006f000000000000007b000000000000007a000000000000007c00000000",
            INIT_4A => X"00000079000000000000007d000000000000007b000000000000007600000000",
            INIT_4B => X"0000006f0000000000000065000000000000006d000000000000007600000000",
            INIT_4C => X"0000006000000000000000520000000000000055000000000000006900000000",
            INIT_4D => X"00000067000000000000007a0000000000000064000000000000006a00000000",
            INIT_4E => X"000000490000000000000047000000000000003e000000000000003d00000000",
            INIT_4F => X"0000004b0000000000000044000000000000004b000000000000004700000000",
            INIT_50 => X"0000007e00000000000000720000000000000048000000000000006400000000",
            INIT_51 => X"0000007e000000000000007c000000000000007f000000000000007800000000",
            INIT_52 => X"0000007b00000000000000800000000000000081000000000000007f00000000",
            INIT_53 => X"0000009000000000000000780000000000000077000000000000007900000000",
            INIT_54 => X"00000058000000000000004f0000000000000063000000000000008300000000",
            INIT_55 => X"0000005b000000000000006c0000000000000061000000000000005f00000000",
            INIT_56 => X"0000003b000000000000003d000000000000003e000000000000002e00000000",
            INIT_57 => X"0000004c00000000000000490000000000000046000000000000004000000000",
            INIT_58 => X"00000069000000000000007f0000000000000034000000000000002200000000",
            INIT_59 => X"000000830000000000000084000000000000007a000000000000005d00000000",
            INIT_5A => X"0000008c00000000000000780000000000000073000000000000008100000000",
            INIT_5B => X"000000850000000000000074000000000000009700000000000000a600000000",
            INIT_5C => X"000000610000000000000056000000000000006e000000000000008d00000000",
            INIT_5D => X"000000310000000000000056000000000000005c000000000000006000000000",
            INIT_5E => X"0000003c000000000000003e000000000000003c000000000000002a00000000",
            INIT_5F => X"0000004a00000000000000450000000000000042000000000000003e00000000",
            INIT_60 => X"0000007d000000000000008e0000000000000040000000000000000400000000",
            INIT_61 => X"00000084000000000000008c000000000000009a000000000000008c00000000",
            INIT_62 => X"0000009c000000000000007b000000000000006b000000000000007f00000000",
            INIT_63 => X"000000530000000000000077000000000000009300000000000000b200000000",
            INIT_64 => X"000000640000000000000053000000000000005b000000000000004000000000",
            INIT_65 => X"00000031000000000000004d000000000000005c000000000000006f00000000",
            INIT_66 => X"000000390000000000000037000000000000002f000000000000002900000000",
            INIT_67 => X"0000004400000000000000420000000000000043000000000000003b00000000",
            INIT_68 => X"0000007b000000000000007a0000000000000048000000000000001800000000",
            INIT_69 => X"0000008d000000000000008f0000000000000096000000000000009c00000000",
            INIT_6A => X"000000a0000000000000008f000000000000006a000000000000007700000000",
            INIT_6B => X"0000007700000000000000800000000000000081000000000000009700000000",
            INIT_6C => X"0000006d00000000000000730000000000000074000000000000004d00000000",
            INIT_6D => X"0000002d0000000000000044000000000000005a000000000000007b00000000",
            INIT_6E => X"000000370000000000000033000000000000002b000000000000002300000000",
            INIT_6F => X"0000003e000000000000003a000000000000003e000000000000003b00000000",
            INIT_70 => X"00000070000000000000004a0000000000000052000000000000004500000000",
            INIT_71 => X"0000008f00000000000000860000000000000091000000000000009600000000",
            INIT_72 => X"0000009c00000000000000a10000000000000084000000000000008300000000",
            INIT_73 => X"0000009700000000000000850000000000000072000000000000007d00000000",
            INIT_74 => X"00000098000000000000009200000000000000a0000000000000009100000000",
            INIT_75 => X"0000002f000000000000004b000000000000005d000000000000008100000000",
            INIT_76 => X"0000004400000000000000380000000000000030000000000000002f00000000",
            INIT_77 => X"000000390000000000000036000000000000003c000000000000003c00000000",
            INIT_78 => X"00000070000000000000003b0000000000000041000000000000005700000000",
            INIT_79 => X"0000007d00000000000000860000000000000096000000000000009800000000",
            INIT_7A => X"000000a500000000000000a7000000000000009b000000000000008f00000000",
            INIT_7B => X"000000a0000000000000008f0000000000000084000000000000009b00000000",
            INIT_7C => X"000000a1000000000000009f000000000000009e00000000000000a200000000",
            INIT_7D => X"0000003900000000000000540000000000000078000000000000008900000000",
            INIT_7E => X"0000005f0000000000000040000000000000002b000000000000003300000000",
            INIT_7F => X"0000003900000000000000360000000000000037000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "sampleifmap_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000660000000000000040000000000000004e000000000000005800000000",
            INIT_01 => X"0000006c0000000000000081000000000000008d000000000000009000000000",
            INIT_02 => X"0000009d00000000000000af00000000000000a5000000000000008b00000000",
            INIT_03 => X"0000009f00000000000000860000000000000086000000000000009e00000000",
            INIT_04 => X"0000009800000000000000930000000000000094000000000000009a00000000",
            INIT_05 => X"0000003100000000000000490000000000000087000000000000009a00000000",
            INIT_06 => X"00000067000000000000004b0000000000000023000000000000001e00000000",
            INIT_07 => X"00000039000000000000002c000000000000003d000000000000006f00000000",
            INIT_08 => X"0000007400000000000000570000000000000057000000000000005600000000",
            INIT_09 => X"0000006900000000000000910000000000000093000000000000008f00000000",
            INIT_0A => X"0000006c000000000000008500000000000000b3000000000000008000000000",
            INIT_0B => X"00000079000000000000007a000000000000008b000000000000009100000000",
            INIT_0C => X"00000079000000000000007c0000000000000087000000000000007d00000000",
            INIT_0D => X"00000018000000000000002a0000000000000058000000000000007200000000",
            INIT_0E => X"000000660000000000000049000000000000001d000000000000001300000000",
            INIT_0F => X"0000002e00000000000000270000000000000050000000000000007500000000",
            INIT_10 => X"00000076000000000000004d000000000000005c000000000000005c00000000",
            INIT_11 => X"0000006200000000000000910000000000000099000000000000009c00000000",
            INIT_12 => X"0000007a000000000000007400000000000000aa000000000000005c00000000",
            INIT_13 => X"00000062000000000000004b000000000000008300000000000000a500000000",
            INIT_14 => X"0000004000000000000000550000000000000061000000000000004c00000000",
            INIT_15 => X"0000001b0000000000000011000000000000001b000000000000003600000000",
            INIT_16 => X"0000007500000000000000450000000000000028000000000000001a00000000",
            INIT_17 => X"0000002800000000000000240000000000000064000000000000007f00000000",
            INIT_18 => X"0000006e000000000000003c0000000000000054000000000000005e00000000",
            INIT_19 => X"00000073000000000000009b00000000000000a3000000000000009c00000000",
            INIT_1A => X"000000890000000000000094000000000000007c000000000000002700000000",
            INIT_1B => X"0000009c00000000000000570000000000000071000000000000009500000000",
            INIT_1C => X"00000027000000000000003d0000000000000050000000000000007800000000",
            INIT_1D => X"0000002e00000000000000220000000000000018000000000000002700000000",
            INIT_1E => X"000000780000000000000045000000000000002d000000000000001f00000000",
            INIT_1F => X"000000200000000000000022000000000000007b000000000000009900000000",
            INIT_20 => X"000000720000000000000059000000000000005d000000000000006100000000",
            INIT_21 => X"00000075000000000000009800000000000000a2000000000000009600000000",
            INIT_22 => X"000000740000000000000064000000000000001d000000000000000d00000000",
            INIT_23 => X"0000007c00000000000000490000000000000056000000000000007300000000",
            INIT_24 => X"0000001b000000000000002f000000000000005b000000000000008600000000",
            INIT_25 => X"0000003200000000000000310000000000000032000000000000003100000000",
            INIT_26 => X"0000007d0000000000000042000000000000001e000000000000001900000000",
            INIT_27 => X"000000200000000000000038000000000000009600000000000000a200000000",
            INIT_28 => X"0000006300000000000000570000000000000068000000000000006a00000000",
            INIT_29 => X"0000005700000000000000810000000000000096000000000000008d00000000",
            INIT_2A => X"000000250000000000000016000000000000000b000000000000000f00000000",
            INIT_2B => X"0000003e00000000000000290000000000000039000000000000003600000000",
            INIT_2C => X"0000001a00000000000000360000000000000048000000000000005300000000",
            INIT_2D => X"0000003300000000000000220000000000000023000000000000002000000000",
            INIT_2E => X"00000070000000000000003e000000000000002b000000000000002800000000",
            INIT_2F => X"0000001f000000000000004a000000000000009e000000000000009b00000000",
            INIT_30 => X"0000005a000000000000004f0000000000000068000000000000007000000000",
            INIT_31 => X"0000004200000000000000730000000000000089000000000000007b00000000",
            INIT_32 => X"0000001700000000000000280000000000000042000000000000002f00000000",
            INIT_33 => X"00000045000000000000002c0000000000000026000000000000001b00000000",
            INIT_34 => X"0000001d0000000000000026000000000000001f000000000000003600000000",
            INIT_35 => X"0000001f000000000000000f0000000000000016000000000000001900000000",
            INIT_36 => X"0000004e000000000000003a0000000000000033000000000000003100000000",
            INIT_37 => X"0000001f00000000000000570000000000000094000000000000008600000000",
            INIT_38 => X"0000006000000000000000590000000000000058000000000000006d00000000",
            INIT_39 => X"0000005e00000000000000730000000000000081000000000000006900000000",
            INIT_3A => X"0000003c00000000000000360000000000000047000000000000006100000000",
            INIT_3B => X"0000003c000000000000004b000000000000003e000000000000004200000000",
            INIT_3C => X"0000000e0000000000000009000000000000000a000000000000001a00000000",
            INIT_3D => X"0000000c000000000000000b0000000000000013000000000000001100000000",
            INIT_3E => X"0000003b000000000000003a000000000000001f000000000000001700000000",
            INIT_3F => X"0000002300000000000000690000000000000088000000000000005e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007000000000000000600000000000000046000000000000005b00000000",
            INIT_41 => X"0000009300000000000000890000000000000068000000000000006000000000",
            INIT_42 => X"000000430000000000000045000000000000003a000000000000007500000000",
            INIT_43 => X"00000035000000000000003f0000000000000045000000000000004a00000000",
            INIT_44 => X"0000000d00000000000000130000000000000019000000000000002900000000",
            INIT_45 => X"00000012000000000000000d0000000000000009000000000000000c00000000",
            INIT_46 => X"00000027000000000000003e0000000000000024000000000000000c00000000",
            INIT_47 => X"0000004700000000000000790000000000000068000000000000003400000000",
            INIT_48 => X"000000620000000000000062000000000000005c000000000000005b00000000",
            INIT_49 => X"0000008600000000000000690000000000000056000000000000006100000000",
            INIT_4A => X"00000061000000000000007c000000000000006b000000000000008e00000000",
            INIT_4B => X"00000049000000000000004e0000000000000049000000000000004400000000",
            INIT_4C => X"0000001c0000000000000026000000000000002b000000000000003e00000000",
            INIT_4D => X"00000014000000000000000b000000000000000e000000000000001600000000",
            INIT_4E => X"000000140000000000000030000000000000002a000000000000001400000000",
            INIT_4F => X"0000006400000000000000580000000000000038000000000000002500000000",
            INIT_50 => X"000000620000000000000061000000000000005e000000000000005b00000000",
            INIT_51 => X"0000004c000000000000005b000000000000006f000000000000007100000000",
            INIT_52 => X"000000510000000000000050000000000000006e000000000000008400000000",
            INIT_53 => X"000000540000000000000063000000000000005f000000000000004700000000",
            INIT_54 => X"000000330000000000000038000000000000003d000000000000004800000000",
            INIT_55 => X"0000002b0000000000000020000000000000002b000000000000003500000000",
            INIT_56 => X"0000002800000000000000250000000000000028000000000000002e00000000",
            INIT_57 => X"000000420000000000000030000000000000005a000000000000004000000000",
            INIT_58 => X"0000005200000000000000500000000000000060000000000000005700000000",
            INIT_59 => X"000000480000000000000062000000000000006d000000000000007100000000",
            INIT_5A => X"0000004600000000000000450000000000000073000000000000005c00000000",
            INIT_5B => X"000000580000000000000060000000000000005e000000000000004a00000000",
            INIT_5C => X"0000004a000000000000004c0000000000000047000000000000004500000000",
            INIT_5D => X"0000004b000000000000003d000000000000003c000000000000004200000000",
            INIT_5E => X"00000041000000000000003f0000000000000040000000000000004900000000",
            INIT_5F => X"0000003a0000000000000036000000000000005e000000000000004c00000000",
            INIT_60 => X"0000004c00000000000000430000000000000061000000000000006000000000",
            INIT_61 => X"00000050000000000000004e000000000000005a000000000000006900000000",
            INIT_62 => X"00000062000000000000004c0000000000000048000000000000005700000000",
            INIT_63 => X"0000005a000000000000005d000000000000005c000000000000005700000000",
            INIT_64 => X"0000004600000000000000550000000000000054000000000000004f00000000",
            INIT_65 => X"00000057000000000000004d0000000000000048000000000000004200000000",
            INIT_66 => X"0000004f00000000000000500000000000000052000000000000005300000000",
            INIT_67 => X"0000005e00000000000000460000000000000035000000000000004300000000",
            INIT_68 => X"0000006500000000000000510000000000000054000000000000004900000000",
            INIT_69 => X"0000005b0000000000000058000000000000005b000000000000006100000000",
            INIT_6A => X"00000063000000000000005b0000000000000059000000000000006900000000",
            INIT_6B => X"0000005a000000000000005d000000000000005d000000000000005900000000",
            INIT_6C => X"0000003c00000000000000490000000000000055000000000000005800000000",
            INIT_6D => X"0000005b00000000000000540000000000000052000000000000004900000000",
            INIT_6E => X"0000005500000000000000570000000000000056000000000000005d00000000",
            INIT_6F => X"0000006400000000000000570000000000000044000000000000004300000000",
            INIT_70 => X"00000071000000000000006a0000000000000060000000000000005300000000",
            INIT_71 => X"0000005f0000000000000060000000000000005f000000000000006000000000",
            INIT_72 => X"00000068000000000000006d0000000000000069000000000000006600000000",
            INIT_73 => X"0000004a0000000000000052000000000000005a000000000000005b00000000",
            INIT_74 => X"0000004a000000000000004d000000000000004e000000000000005200000000",
            INIT_75 => X"0000005c00000000000000570000000000000055000000000000004d00000000",
            INIT_76 => X"00000054000000000000005a0000000000000059000000000000006400000000",
            INIT_77 => X"0000005a0000000000000057000000000000004d000000000000004e00000000",
            INIT_78 => X"000000680000000000000071000000000000006b000000000000005c00000000",
            INIT_79 => X"0000005c000000000000004d0000000000000042000000000000005200000000",
            INIT_7A => X"0000005a000000000000005b0000000000000051000000000000005f00000000",
            INIT_7B => X"0000003d000000000000004d000000000000005b000000000000005800000000",
            INIT_7C => X"000000520000000000000056000000000000004d000000000000004600000000",
            INIT_7D => X"00000060000000000000005b000000000000005c000000000000005300000000",
            INIT_7E => X"0000005b0000000000000057000000000000005c000000000000006500000000",
            INIT_7F => X"00000057000000000000005b000000000000005a000000000000005c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "sampleifmap_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000024000000000000001a000000000000003d000000000000005300000000",
            INIT_01 => X"00000036000000000000003a0000000000000043000000000000004100000000",
            INIT_02 => X"0000003b00000000000000340000000000000041000000000000003f00000000",
            INIT_03 => X"00000034000000000000002e0000000000000035000000000000003e00000000",
            INIT_04 => X"00000027000000000000002b0000000000000041000000000000004700000000",
            INIT_05 => X"00000026000000000000002d000000000000002f000000000000002f00000000",
            INIT_06 => X"00000032000000000000002a000000000000002d000000000000002f00000000",
            INIT_07 => X"000000290000000000000029000000000000002e000000000000004500000000",
            INIT_08 => X"00000046000000000000003a0000000000000035000000000000006100000000",
            INIT_09 => X"0000004d00000000000000440000000000000043000000000000004600000000",
            INIT_0A => X"0000003900000000000000380000000000000041000000000000004400000000",
            INIT_0B => X"0000002e00000000000000320000000000000039000000000000003400000000",
            INIT_0C => X"00000026000000000000002b0000000000000034000000000000003c00000000",
            INIT_0D => X"00000028000000000000002c000000000000002f000000000000002f00000000",
            INIT_0E => X"00000038000000000000002b000000000000001e000000000000002000000000",
            INIT_0F => X"0000003100000000000000330000000000000035000000000000004300000000",
            INIT_10 => X"00000051000000000000005c0000000000000047000000000000006400000000",
            INIT_11 => X"0000004e00000000000000440000000000000039000000000000004400000000",
            INIT_12 => X"0000003b000000000000003f0000000000000047000000000000004000000000",
            INIT_13 => X"0000003000000000000000310000000000000030000000000000003400000000",
            INIT_14 => X"0000001e00000000000000210000000000000032000000000000003b00000000",
            INIT_15 => X"0000003800000000000000350000000000000030000000000000002b00000000",
            INIT_16 => X"0000003800000000000000390000000000000038000000000000003300000000",
            INIT_17 => X"00000031000000000000002f0000000000000035000000000000003900000000",
            INIT_18 => X"000000590000000000000061000000000000005f000000000000006000000000",
            INIT_19 => X"0000004800000000000000490000000000000037000000000000004900000000",
            INIT_1A => X"000000420000000000000042000000000000004e000000000000004100000000",
            INIT_1B => X"0000003f00000000000000360000000000000037000000000000004300000000",
            INIT_1C => X"00000012000000000000001a000000000000002e000000000000002f00000000",
            INIT_1D => X"00000035000000000000002f0000000000000029000000000000002200000000",
            INIT_1E => X"0000003e00000000000000400000000000000044000000000000003d00000000",
            INIT_1F => X"0000003c000000000000003a000000000000002d000000000000003000000000",
            INIT_20 => X"0000005700000000000000540000000000000061000000000000005c00000000",
            INIT_21 => X"0000004b000000000000004c000000000000003f000000000000004900000000",
            INIT_22 => X"0000004b000000000000004b000000000000004a000000000000004a00000000",
            INIT_23 => X"0000003b0000000000000035000000000000003b000000000000004300000000",
            INIT_24 => X"0000001e00000000000000330000000000000034000000000000003b00000000",
            INIT_25 => X"00000027000000000000002e0000000000000029000000000000001f00000000",
            INIT_26 => X"0000003d000000000000003d000000000000003b000000000000002e00000000",
            INIT_27 => X"0000003c000000000000003a0000000000000030000000000000003400000000",
            INIT_28 => X"0000005900000000000000470000000000000066000000000000006500000000",
            INIT_29 => X"0000004c000000000000004c0000000000000046000000000000005100000000",
            INIT_2A => X"00000047000000000000004e0000000000000051000000000000004c00000000",
            INIT_2B => X"0000003100000000000000350000000000000043000000000000004400000000",
            INIT_2C => X"0000003900000000000000480000000000000041000000000000004300000000",
            INIT_2D => X"000000320000000000000042000000000000003e000000000000002b00000000",
            INIT_2E => X"0000003a00000000000000380000000000000036000000000000003800000000",
            INIT_2F => X"00000041000000000000003c000000000000003d000000000000003c00000000",
            INIT_30 => X"0000006300000000000000490000000000000059000000000000007800000000",
            INIT_31 => X"0000004b00000000000000510000000000000050000000000000005300000000",
            INIT_32 => X"0000004200000000000000550000000000000057000000000000005100000000",
            INIT_33 => X"000000350000000000000043000000000000004f000000000000004c00000000",
            INIT_34 => X"0000004d000000000000004a0000000000000040000000000000003c00000000",
            INIT_35 => X"0000002f00000000000000410000000000000040000000000000004100000000",
            INIT_36 => X"00000030000000000000002d0000000000000036000000000000003500000000",
            INIT_37 => X"00000042000000000000003f000000000000003d000000000000003a00000000",
            INIT_38 => X"0000005b000000000000005b000000000000003b000000000000007500000000",
            INIT_39 => X"00000054000000000000004f0000000000000051000000000000005100000000",
            INIT_3A => X"0000004800000000000000560000000000000056000000000000005700000000",
            INIT_3B => X"0000003f000000000000004a000000000000004c000000000000004d00000000",
            INIT_3C => X"00000049000000000000004c0000000000000049000000000000004200000000",
            INIT_3D => X"0000002f0000000000000038000000000000002f000000000000004700000000",
            INIT_3E => X"0000002a00000000000000230000000000000031000000000000002c00000000",
            INIT_3F => X"00000040000000000000003e0000000000000039000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000051000000000000005b0000000000000054000000000000005c00000000",
            INIT_41 => X"000000500000000000000050000000000000004f000000000000005300000000",
            INIT_42 => X"0000004600000000000000490000000000000053000000000000005800000000",
            INIT_43 => X"0000003d00000000000000430000000000000048000000000000005100000000",
            INIT_44 => X"0000004600000000000000460000000000000041000000000000004300000000",
            INIT_45 => X"0000003c000000000000004f0000000000000040000000000000004f00000000",
            INIT_46 => X"0000003b0000000000000034000000000000002d000000000000002c00000000",
            INIT_47 => X"00000040000000000000003d000000000000003d000000000000003a00000000",
            INIT_48 => X"0000005a000000000000004c0000000000000058000000000000006100000000",
            INIT_49 => X"0000004700000000000000530000000000000056000000000000005b00000000",
            INIT_4A => X"0000005300000000000000540000000000000052000000000000004f00000000",
            INIT_4B => X"00000055000000000000004d0000000000000053000000000000005800000000",
            INIT_4C => X"000000460000000000000039000000000000003e000000000000005100000000",
            INIT_4D => X"0000004b00000000000000590000000000000048000000000000005000000000",
            INIT_4E => X"0000003c000000000000003a0000000000000031000000000000002b00000000",
            INIT_4F => X"000000400000000000000039000000000000003f000000000000003a00000000",
            INIT_50 => X"0000006200000000000000560000000000000030000000000000005100000000",
            INIT_51 => X"000000540000000000000052000000000000005b000000000000005900000000",
            INIT_52 => X"0000005000000000000000500000000000000054000000000000005b00000000",
            INIT_53 => X"0000007e00000000000000670000000000000065000000000000005e00000000",
            INIT_54 => X"0000004300000000000000370000000000000049000000000000006b00000000",
            INIT_55 => X"000000440000000000000051000000000000004c000000000000004b00000000",
            INIT_56 => X"0000002d000000000000002f0000000000000031000000000000002000000000",
            INIT_57 => X"00000041000000000000003e000000000000003a000000000000003300000000",
            INIT_58 => X"0000004d0000000000000063000000000000001f000000000000001400000000",
            INIT_59 => X"0000005a000000000000005a0000000000000056000000000000004000000000",
            INIT_5A => X"0000005f00000000000000450000000000000045000000000000005f00000000",
            INIT_5B => X"0000007900000000000000670000000000000088000000000000008f00000000",
            INIT_5C => X"00000050000000000000003f0000000000000052000000000000007600000000",
            INIT_5D => X"000000210000000000000042000000000000004d000000000000005200000000",
            INIT_5E => X"0000002e00000000000000300000000000000030000000000000002100000000",
            INIT_5F => X"0000003f000000000000003b0000000000000036000000000000003000000000",
            INIT_60 => X"0000005c00000000000000700000000000000032000000000000000000000000",
            INIT_61 => X"000000620000000000000069000000000000007a000000000000006e00000000",
            INIT_62 => X"0000007700000000000000540000000000000048000000000000006000000000",
            INIT_63 => X"00000049000000000000005f000000000000007d000000000000009d00000000",
            INIT_64 => X"0000005400000000000000410000000000000047000000000000003400000000",
            INIT_65 => X"0000002a0000000000000041000000000000004f000000000000006000000000",
            INIT_66 => X"0000002900000000000000290000000000000025000000000000002500000000",
            INIT_67 => X"0000003a00000000000000390000000000000038000000000000002d00000000",
            INIT_68 => X"0000005c0000000000000061000000000000003c000000000000001400000000",
            INIT_69 => X"0000006f00000000000000700000000000000078000000000000007d00000000",
            INIT_6A => X"00000080000000000000006e000000000000004c000000000000005900000000",
            INIT_6B => X"0000006c00000000000000620000000000000064000000000000007f00000000",
            INIT_6C => X"0000005b00000000000000620000000000000063000000000000004400000000",
            INIT_6D => X"00000029000000000000003a000000000000004c000000000000006a00000000",
            INIT_6E => X"0000002600000000000000250000000000000023000000000000002100000000",
            INIT_6F => X"0000003500000000000000320000000000000034000000000000002e00000000",
            INIT_70 => X"00000058000000000000003a0000000000000046000000000000003b00000000",
            INIT_71 => X"00000073000000000000006a0000000000000075000000000000007b00000000",
            INIT_72 => X"0000007d00000000000000820000000000000067000000000000006600000000",
            INIT_73 => X"0000008900000000000000660000000000000050000000000000005f00000000",
            INIT_74 => X"00000084000000000000007e000000000000008c000000000000008300000000",
            INIT_75 => X"0000002a0000000000000040000000000000004e000000000000006f00000000",
            INIT_76 => X"00000032000000000000002a0000000000000028000000000000002b00000000",
            INIT_77 => X"00000031000000000000002e0000000000000032000000000000002f00000000",
            INIT_78 => X"0000005e00000000000000320000000000000035000000000000004900000000",
            INIT_79 => X"00000062000000000000006c000000000000007c000000000000007e00000000",
            INIT_7A => X"00000088000000000000008a000000000000007d000000000000007200000000",
            INIT_7B => X"0000008c00000000000000710000000000000062000000000000007b00000000",
            INIT_7C => X"0000008c000000000000008a0000000000000089000000000000008f00000000",
            INIT_7D => X"0000003300000000000000490000000000000069000000000000007500000000",
            INIT_7E => X"0000004d00000000000000320000000000000023000000000000002f00000000",
            INIT_7F => X"00000032000000000000002d000000000000002d000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "sampleifmap_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000056000000000000003a0000000000000041000000000000004800000000",
            INIT_01 => X"0000005300000000000000690000000000000075000000000000007700000000",
            INIT_02 => X"0000008200000000000000930000000000000089000000000000006e00000000",
            INIT_03 => X"00000087000000000000006d000000000000006b000000000000008200000000",
            INIT_04 => X"00000083000000000000007e000000000000007f000000000000008400000000",
            INIT_05 => X"0000002a000000000000003d0000000000000077000000000000008700000000",
            INIT_06 => X"00000055000000000000003c000000000000001b000000000000001a00000000",
            INIT_07 => X"0000003300000000000000240000000000000033000000000000006100000000",
            INIT_08 => X"0000006600000000000000510000000000000048000000000000004700000000",
            INIT_09 => X"00000050000000000000007a000000000000007c000000000000007800000000",
            INIT_0A => X"00000054000000000000006a0000000000000097000000000000006300000000",
            INIT_0B => X"0000005c00000000000000650000000000000079000000000000007c00000000",
            INIT_0C => X"0000006500000000000000680000000000000073000000000000006300000000",
            INIT_0D => X"00000011000000000000001f0000000000000048000000000000005e00000000",
            INIT_0E => X"00000055000000000000003a0000000000000015000000000000000e00000000",
            INIT_0F => X"00000029000000000000001f0000000000000046000000000000006800000000",
            INIT_10 => X"000000640000000000000044000000000000004e000000000000004f00000000",
            INIT_11 => X"0000004b000000000000007d0000000000000088000000000000008600000000",
            INIT_12 => X"00000061000000000000005b0000000000000093000000000000004700000000",
            INIT_13 => X"0000004800000000000000370000000000000071000000000000008e00000000",
            INIT_14 => X"000000320000000000000045000000000000004f000000000000003500000000",
            INIT_15 => X"00000016000000000000000d0000000000000014000000000000002a00000000",
            INIT_16 => X"0000006000000000000000370000000000000023000000000000001400000000",
            INIT_17 => X"00000023000000000000001e000000000000005b000000000000006f00000000",
            INIT_18 => X"0000005800000000000000320000000000000048000000000000005100000000",
            INIT_19 => X"0000005d000000000000008a0000000000000099000000000000008700000000",
            INIT_1A => X"00000071000000000000007f000000000000006f000000000000001f00000000",
            INIT_1B => X"0000008d0000000000000047000000000000005c000000000000007c00000000",
            INIT_1C => X"0000002100000000000000330000000000000041000000000000006700000000",
            INIT_1D => X"0000002c00000000000000240000000000000019000000000000002400000000",
            INIT_1E => X"000000600000000000000036000000000000002b000000000000001a00000000",
            INIT_1F => X"0000001a000000000000001e0000000000000073000000000000008900000000",
            INIT_20 => X"0000005f000000000000004f0000000000000052000000000000005300000000",
            INIT_21 => X"0000006200000000000000860000000000000096000000000000008200000000",
            INIT_22 => X"0000006300000000000000560000000000000017000000000000000a00000000",
            INIT_23 => X"000000740000000000000042000000000000004c000000000000006500000000",
            INIT_24 => X"000000170000000000000027000000000000004e000000000000007a00000000",
            INIT_25 => X"0000002e000000000000002f000000000000002f000000000000002e00000000",
            INIT_26 => X"000000670000000000000034000000000000001b000000000000001400000000",
            INIT_27 => X"00000019000000000000002f0000000000000089000000000000009200000000",
            INIT_28 => X"00000053000000000000004e000000000000005c000000000000005c00000000",
            INIT_29 => X"00000046000000000000006e0000000000000087000000000000007b00000000",
            INIT_2A => X"0000001d00000000000000100000000000000008000000000000000c00000000",
            INIT_2B => X"0000003800000000000000250000000000000034000000000000002f00000000",
            INIT_2C => X"00000012000000000000002b0000000000000039000000000000004600000000",
            INIT_2D => X"0000002c000000000000001d000000000000001c000000000000001900000000",
            INIT_2E => X"0000005e00000000000000310000000000000026000000000000002100000000",
            INIT_2F => X"00000018000000000000003d000000000000008d000000000000008c00000000",
            INIT_30 => X"0000004e0000000000000046000000000000005d000000000000006100000000",
            INIT_31 => X"0000003000000000000000600000000000000076000000000000006b00000000",
            INIT_32 => X"000000130000000000000022000000000000003a000000000000002500000000",
            INIT_33 => X"0000003b0000000000000026000000000000001f000000000000001300000000",
            INIT_34 => X"00000012000000000000001b0000000000000013000000000000002700000000",
            INIT_35 => X"00000018000000000000000a0000000000000011000000000000001100000000",
            INIT_36 => X"000000400000000000000030000000000000002c000000000000002a00000000",
            INIT_37 => X"0000001800000000000000460000000000000080000000000000007800000000",
            INIT_38 => X"000000580000000000000052000000000000004d000000000000005e00000000",
            INIT_39 => X"0000004b000000000000005f000000000000006b000000000000005b00000000",
            INIT_3A => X"0000003900000000000000300000000000000037000000000000004a00000000",
            INIT_3B => X"0000003300000000000000430000000000000035000000000000003a00000000",
            INIT_3C => X"0000000800000000000000030000000000000004000000000000001000000000",
            INIT_3D => X"0000000600000000000000070000000000000013000000000000000e00000000",
            INIT_3E => X"0000002f00000000000000300000000000000017000000000000001100000000",
            INIT_3F => X"0000001b00000000000000570000000000000073000000000000005100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000057000000000000003b000000000000004b00000000",
            INIT_41 => X"0000007e00000000000000750000000000000052000000000000005300000000",
            INIT_42 => X"0000003e00000000000000390000000000000022000000000000005500000000",
            INIT_43 => X"0000002e0000000000000039000000000000003d000000000000004200000000",
            INIT_44 => X"0000000d00000000000000120000000000000017000000000000002400000000",
            INIT_45 => X"0000000e000000000000000c000000000000000e000000000000000f00000000",
            INIT_46 => X"0000001e0000000000000036000000000000001c000000000000000700000000",
            INIT_47 => X"0000003e00000000000000680000000000000055000000000000002800000000",
            INIT_48 => X"000000560000000000000051000000000000004d000000000000004d00000000",
            INIT_49 => X"0000007000000000000000570000000000000045000000000000005500000000",
            INIT_4A => X"0000004f0000000000000064000000000000004f000000000000006f00000000",
            INIT_4B => X"0000003a00000000000000450000000000000043000000000000003b00000000",
            INIT_4C => X"0000001500000000000000200000000000000026000000000000003300000000",
            INIT_4D => X"0000000e0000000000000006000000000000000c000000000000001100000000",
            INIT_4E => X"0000000f00000000000000290000000000000022000000000000000f00000000",
            INIT_4F => X"0000005a000000000000004c000000000000002e000000000000001f00000000",
            INIT_50 => X"0000005500000000000000520000000000000051000000000000004f00000000",
            INIT_51 => X"00000039000000000000004a0000000000000060000000000000006500000000",
            INIT_52 => X"0000003e000000000000003a0000000000000057000000000000006d00000000",
            INIT_53 => X"00000044000000000000005a0000000000000058000000000000003d00000000",
            INIT_54 => X"0000002a000000000000002f0000000000000035000000000000003b00000000",
            INIT_55 => X"0000002300000000000000180000000000000023000000000000002c00000000",
            INIT_56 => X"0000001f000000000000001b000000000000001d000000000000002600000000",
            INIT_57 => X"0000003800000000000000270000000000000052000000000000003900000000",
            INIT_58 => X"0000004a000000000000004a0000000000000057000000000000004c00000000",
            INIT_59 => X"000000390000000000000053000000000000005f000000000000006600000000",
            INIT_5A => X"0000003a00000000000000370000000000000063000000000000004d00000000",
            INIT_5B => X"0000004d00000000000000570000000000000054000000000000003f00000000",
            INIT_5C => X"000000440000000000000043000000000000003c000000000000003900000000",
            INIT_5D => X"0000003f00000000000000310000000000000031000000000000003b00000000",
            INIT_5E => X"0000003300000000000000300000000000000031000000000000003c00000000",
            INIT_5F => X"0000002f000000000000002d0000000000000054000000000000003f00000000",
            INIT_60 => X"000000450000000000000040000000000000005a000000000000005500000000",
            INIT_61 => X"000000440000000000000041000000000000004e000000000000005e00000000",
            INIT_62 => X"0000005a0000000000000042000000000000003c000000000000004c00000000",
            INIT_63 => X"000000510000000000000053000000000000004e000000000000004a00000000",
            INIT_64 => X"00000040000000000000004c0000000000000047000000000000004300000000",
            INIT_65 => X"00000048000000000000003e0000000000000039000000000000003b00000000",
            INIT_66 => X"0000003e00000000000000400000000000000042000000000000004400000000",
            INIT_67 => X"00000053000000000000003d0000000000000029000000000000003200000000",
            INIT_68 => X"0000005c0000000000000049000000000000004b000000000000003d00000000",
            INIT_69 => X"00000050000000000000004e0000000000000051000000000000005700000000",
            INIT_6A => X"000000590000000000000050000000000000004c000000000000005d00000000",
            INIT_6B => X"00000050000000000000004e000000000000004c000000000000004a00000000",
            INIT_6C => X"00000035000000000000003e0000000000000045000000000000004a00000000",
            INIT_6D => X"0000004b00000000000000440000000000000042000000000000004000000000",
            INIT_6E => X"0000004400000000000000480000000000000048000000000000004d00000000",
            INIT_6F => X"00000059000000000000004e0000000000000038000000000000003200000000",
            INIT_70 => X"00000064000000000000005a0000000000000051000000000000004600000000",
            INIT_71 => X"0000005500000000000000570000000000000055000000000000005600000000",
            INIT_72 => X"0000005a000000000000005d0000000000000057000000000000005600000000",
            INIT_73 => X"0000003c000000000000003f0000000000000046000000000000004a00000000",
            INIT_74 => X"0000003e000000000000003e000000000000003c000000000000004200000000",
            INIT_75 => X"0000004c00000000000000470000000000000046000000000000004100000000",
            INIT_76 => X"00000047000000000000004e000000000000004d000000000000005500000000",
            INIT_77 => X"0000004f000000000000004d0000000000000041000000000000003e00000000",
            INIT_78 => X"00000059000000000000005f000000000000005d000000000000004f00000000",
            INIT_79 => X"0000005100000000000000460000000000000039000000000000004600000000",
            INIT_7A => X"0000004700000000000000470000000000000040000000000000005300000000",
            INIT_7B => X"0000002f000000000000003d000000000000004c000000000000004a00000000",
            INIT_7C => X"000000460000000000000048000000000000003f000000000000003800000000",
            INIT_7D => X"00000050000000000000004b000000000000004c000000000000004500000000",
            INIT_7E => X"0000004e0000000000000049000000000000004f000000000000005600000000",
            INIT_7F => X"00000049000000000000004f000000000000004c000000000000004f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "sampleifmap_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d900000000000000d100000000000000b900000000000000a000000000",
            INIT_01 => X"000000f600000000000000f900000000000000f600000000000000e600000000",
            INIT_02 => X"000000dd00000000000000e600000000000000f300000000000000f800000000",
            INIT_03 => X"000000c700000000000000d800000000000000dd00000000000000da00000000",
            INIT_04 => X"000000b400000000000000b800000000000000bb00000000000000bc00000000",
            INIT_05 => X"0000008b0000000000000079000000000000009000000000000000a600000000",
            INIT_06 => X"0000004f00000000000000660000000000000066000000000000006a00000000",
            INIT_07 => X"0000005e000000000000005b0000000000000065000000000000005e00000000",
            INIT_08 => X"000000e600000000000000f200000000000000ef00000000000000e100000000",
            INIT_09 => X"000000eb00000000000000f300000000000000f500000000000000e800000000",
            INIT_0A => X"000000cd00000000000000d800000000000000e600000000000000ed00000000",
            INIT_0B => X"000000ba00000000000000c800000000000000cb00000000000000c900000000",
            INIT_0C => X"0000007f00000000000000a100000000000000ab00000000000000af00000000",
            INIT_0D => X"00000087000000000000007a000000000000008d000000000000008e00000000",
            INIT_0E => X"0000003400000000000000250000000000000052000000000000007600000000",
            INIT_0F => X"000000640000000000000061000000000000006b000000000000005f00000000",
            INIT_10 => X"000000dc00000000000000f100000000000000f900000000000000fc00000000",
            INIT_11 => X"000000d600000000000000df00000000000000e200000000000000d900000000",
            INIT_12 => X"000000b800000000000000c300000000000000cf00000000000000d500000000",
            INIT_13 => X"000000a700000000000000b300000000000000b600000000000000b300000000",
            INIT_14 => X"0000008100000000000000940000000000000098000000000000009f00000000",
            INIT_15 => X"000000720000000000000080000000000000008c000000000000008000000000",
            INIT_16 => X"0000002600000000000000040000000000000028000000000000005700000000",
            INIT_17 => X"0000006900000000000000690000000000000073000000000000006300000000",
            INIT_18 => X"000000d300000000000000de00000000000000e100000000000000e900000000",
            INIT_19 => X"000000c000000000000000c800000000000000cb00000000000000d300000000",
            INIT_1A => X"000000a400000000000000ae00000000000000b700000000000000bb00000000",
            INIT_1B => X"0000009900000000000000a000000000000000a500000000000000a000000000",
            INIT_1C => X"0000008a000000000000008c000000000000008d000000000000009100000000",
            INIT_1D => X"00000069000000000000007f000000000000007d000000000000007d00000000",
            INIT_1E => X"00000037000000000000001a0000000000000025000000000000003b00000000",
            INIT_1F => X"0000006d00000000000000700000000000000078000000000000007000000000",
            INIT_20 => X"000000c900000000000000cf00000000000000c300000000000000cf00000000",
            INIT_21 => X"000000ab00000000000000b300000000000000b400000000000000be00000000",
            INIT_22 => X"000000920000000000000099000000000000009f00000000000000a300000000",
            INIT_23 => X"0000008d00000000000000930000000000000097000000000000009100000000",
            INIT_24 => X"0000008700000000000000830000000000000088000000000000008700000000",
            INIT_25 => X"0000005a0000000000000084000000000000007a000000000000008100000000",
            INIT_26 => X"000000560000000000000030000000000000003d000000000000003a00000000",
            INIT_27 => X"0000006d00000000000000720000000000000078000000000000007500000000",
            INIT_28 => X"000000a200000000000000aa00000000000000ab00000000000000b600000000",
            INIT_29 => X"00000097000000000000009f000000000000009c000000000000009900000000",
            INIT_2A => X"0000008a000000000000008c000000000000008d000000000000009000000000",
            INIT_2B => X"0000008a000000000000008a000000000000008d000000000000008b00000000",
            INIT_2C => X"0000008a0000000000000086000000000000008c000000000000008700000000",
            INIT_2D => X"0000004500000000000000660000000000000089000000000000008c00000000",
            INIT_2E => X"000000740000000000000043000000000000003e000000000000004b00000000",
            INIT_2F => X"0000006e00000000000000700000000000000080000000000000008100000000",
            INIT_30 => X"0000008600000000000000880000000000000088000000000000008d00000000",
            INIT_31 => X"00000085000000000000008c0000000000000086000000000000008800000000",
            INIT_32 => X"0000008d000000000000008b0000000000000089000000000000008700000000",
            INIT_33 => X"00000091000000000000008e0000000000000092000000000000008f00000000",
            INIT_34 => X"0000008f000000000000008a0000000000000091000000000000009100000000",
            INIT_35 => X"00000021000000000000002f000000000000006b000000000000008e00000000",
            INIT_36 => X"0000007f000000000000006c000000000000004b000000000000004800000000",
            INIT_37 => X"00000070000000000000006f0000000000000084000000000000008400000000",
            INIT_38 => X"000000810000000000000080000000000000007d000000000000007600000000",
            INIT_39 => X"00000084000000000000008a0000000000000083000000000000008800000000",
            INIT_3A => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_3B => X"00000099000000000000009a000000000000009e000000000000009600000000",
            INIT_3C => X"0000009400000000000000930000000000000095000000000000009200000000",
            INIT_3D => X"00000011000000000000000d0000000000000042000000000000008000000000",
            INIT_3E => X"0000007a00000000000000800000000000000075000000000000005000000000",
            INIT_3F => X"0000007000000000000000720000000000000080000000000000007b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000850000000000000084000000000000007e000000000000007300000000",
            INIT_41 => X"00000089000000000000008f0000000000000087000000000000008b00000000",
            INIT_42 => X"0000009800000000000000950000000000000091000000000000008b00000000",
            INIT_43 => X"000000aa00000000000000a3000000000000009a000000000000009400000000",
            INIT_44 => X"00000094000000000000009d00000000000000a2000000000000009e00000000",
            INIT_45 => X"0000001e000000000000000e000000000000002c000000000000007300000000",
            INIT_46 => X"0000007e0000000000000088000000000000008b000000000000006900000000",
            INIT_47 => X"0000006f0000000000000074000000000000007a000000000000007700000000",
            INIT_48 => X"0000008800000000000000880000000000000080000000000000007600000000",
            INIT_49 => X"0000008d00000000000000910000000000000088000000000000008d00000000",
            INIT_4A => X"000000a5000000000000009a0000000000000093000000000000008d00000000",
            INIT_4B => X"000000a700000000000000a2000000000000009a000000000000009d00000000",
            INIT_4C => X"0000008a00000000000000910000000000000093000000000000009b00000000",
            INIT_4D => X"00000037000000000000002e0000000000000038000000000000006300000000",
            INIT_4E => X"0000007e000000000000007a000000000000007c000000000000006d00000000",
            INIT_4F => X"0000006e00000000000000750000000000000074000000000000007300000000",
            INIT_50 => X"00000089000000000000008b0000000000000084000000000000007d00000000",
            INIT_51 => X"0000008c00000000000000900000000000000088000000000000008e00000000",
            INIT_52 => X"0000009900000000000000960000000000000090000000000000008b00000000",
            INIT_53 => X"000000980000000000000090000000000000008b000000000000008300000000",
            INIT_54 => X"000000d600000000000000d300000000000000ba00000000000000a600000000",
            INIT_55 => X"0000002a0000000000000045000000000000005c000000000000008000000000",
            INIT_56 => X"000000730000000000000063000000000000005f000000000000005500000000",
            INIT_57 => X"0000006b0000000000000071000000000000006f000000000000007000000000",
            INIT_58 => X"0000008a000000000000008e0000000000000089000000000000008500000000",
            INIT_59 => X"0000008a000000000000008e0000000000000088000000000000008d00000000",
            INIT_5A => X"000000840000000000000088000000000000008f000000000000008900000000",
            INIT_5B => X"000000cb00000000000000c900000000000000b6000000000000008e00000000",
            INIT_5C => X"000000c000000000000000cf00000000000000ce00000000000000d200000000",
            INIT_5D => X"0000002a000000000000009200000000000000bd00000000000000a200000000",
            INIT_5E => X"0000007200000000000000670000000000000028000000000000001b00000000",
            INIT_5F => X"00000068000000000000006c000000000000006a000000000000006d00000000",
            INIT_60 => X"0000008b000000000000008f000000000000008b000000000000008c00000000",
            INIT_61 => X"00000089000000000000008a000000000000008c000000000000008f00000000",
            INIT_62 => X"000000a400000000000000900000000000000085000000000000008700000000",
            INIT_63 => X"00000073000000000000008900000000000000a000000000000000ab00000000",
            INIT_64 => X"0000003b000000000000004b000000000000005d000000000000006a00000000",
            INIT_65 => X"0000005f00000000000000c900000000000000dc000000000000006f00000000",
            INIT_66 => X"00000074000000000000003e0000000000000007000000000000000d00000000",
            INIT_67 => X"0000006400000000000000690000000000000065000000000000006300000000",
            INIT_68 => X"0000008c000000000000008f000000000000008a000000000000009000000000",
            INIT_69 => X"0000008700000000000000820000000000000092000000000000009200000000",
            INIT_6A => X"0000006e000000000000008c0000000000000091000000000000008200000000",
            INIT_6B => X"000000130000000000000031000000000000005c000000000000005e00000000",
            INIT_6C => X"0000001200000000000000190000000000000032000000000000001d00000000",
            INIT_6D => X"0000009d00000000000000d200000000000000d1000000000000007800000000",
            INIT_6E => X"0000004400000000000000130000000000000006000000000000002600000000",
            INIT_6F => X"0000005f00000000000000630000000000000052000000000000004500000000",
            INIT_70 => X"0000008e0000000000000092000000000000008b000000000000009100000000",
            INIT_71 => X"000000800000000000000079000000000000008e000000000000009000000000",
            INIT_72 => X"000000440000000000000054000000000000007f000000000000008500000000",
            INIT_73 => X"00000016000000000000002e0000000000000052000000000000005600000000",
            INIT_74 => X"00000041000000000000001e0000000000000032000000000000001300000000",
            INIT_75 => X"000000cb00000000000000cd00000000000000c900000000000000af00000000",
            INIT_76 => X"0000001600000000000000120000000000000010000000000000006600000000",
            INIT_77 => X"00000058000000000000004f0000000000000038000000000000002300000000",
            INIT_78 => X"000000900000000000000094000000000000008b000000000000008f00000000",
            INIT_79 => X"00000083000000000000008b0000000000000084000000000000008a00000000",
            INIT_7A => X"0000005600000000000000480000000000000042000000000000007500000000",
            INIT_7B => X"000000220000000000000028000000000000004e000000000000006a00000000",
            INIT_7C => X"000000b600000000000000730000000000000046000000000000002400000000",
            INIT_7D => X"000000c300000000000000cd00000000000000c500000000000000cb00000000",
            INIT_7E => X"000000120000000000000025000000000000003d000000000000006c00000000",
            INIT_7F => X"000000530000000000000064000000000000004f000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "sampleifmap_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000900000000000000093000000000000008b000000000000008e00000000",
            INIT_01 => X"0000007900000000000000840000000000000072000000000000008500000000",
            INIT_02 => X"00000045000000000000003c0000000000000059000000000000005100000000",
            INIT_03 => X"0000009b00000000000000530000000000000044000000000000005500000000",
            INIT_04 => X"000000eb00000000000000ed00000000000000db00000000000000c000000000",
            INIT_05 => X"0000007200000000000000d300000000000000d700000000000000d700000000",
            INIT_06 => X"000000140000000000000035000000000000005d000000000000003000000000",
            INIT_07 => X"00000054000000000000008f000000000000008b000000000000004100000000",
            INIT_08 => X"00000089000000000000008e000000000000008d000000000000008f00000000",
            INIT_09 => X"00000043000000000000003a0000000000000045000000000000007400000000",
            INIT_0A => X"0000001c000000000000001d000000000000004b000000000000005100000000",
            INIT_0B => X"000000f2000000000000008c0000000000000019000000000000002400000000",
            INIT_0C => X"000000dc00000000000000e300000000000000eb00000000000000ec00000000",
            INIT_0D => X"0000003a000000000000009500000000000000df00000000000000db00000000",
            INIT_0E => X"0000004e000000000000004e0000000000000054000000000000003900000000",
            INIT_0F => X"0000005b00000000000000a700000000000000a1000000000000008500000000",
            INIT_10 => X"000000860000000000000088000000000000008c000000000000008f00000000",
            INIT_11 => X"00000034000000000000002d0000000000000047000000000000008d00000000",
            INIT_12 => X"0000001600000000000000170000000000000021000000000000004300000000",
            INIT_13 => X"000000d9000000000000009b0000000000000029000000000000002f00000000",
            INIT_14 => X"000000d000000000000000bf00000000000000be00000000000000c700000000",
            INIT_15 => X"0000006700000000000000ad00000000000000df00000000000000dc00000000",
            INIT_16 => X"0000009500000000000000870000000000000073000000000000005d00000000",
            INIT_17 => X"0000005900000000000000a50000000000000094000000000000009800000000",
            INIT_18 => X"000000b5000000000000007e000000000000008c000000000000008f00000000",
            INIT_19 => X"0000002b0000000000000021000000000000004c00000000000000bd00000000",
            INIT_1A => X"0000001700000000000000100000000000000015000000000000003900000000",
            INIT_1B => X"000000c2000000000000009e0000000000000042000000000000003900000000",
            INIT_1C => X"000000c900000000000000c400000000000000b300000000000000b600000000",
            INIT_1D => X"000000b300000000000000de00000000000000ce00000000000000c200000000",
            INIT_1E => X"000000970000000000000095000000000000009c000000000000009700000000",
            INIT_1F => X"0000004200000000000000880000000000000092000000000000009600000000",
            INIT_20 => X"000000ea000000000000009a0000000000000085000000000000008c00000000",
            INIT_21 => X"0000002a0000000000000026000000000000005a00000000000000b500000000",
            INIT_22 => X"0000000b000000000000000b000000000000000b000000000000003400000000",
            INIT_23 => X"000000ba00000000000000a00000000000000031000000000000001400000000",
            INIT_24 => X"0000007300000000000000b900000000000000b900000000000000b000000000",
            INIT_25 => X"000000c400000000000000a1000000000000005a000000000000004500000000",
            INIT_26 => X"0000009900000000000000a000000000000000aa00000000000000b700000000",
            INIT_27 => X"00000026000000000000004d0000000000000088000000000000009300000000",
            INIT_28 => X"000000a300000000000000a30000000000000080000000000000008200000000",
            INIT_29 => X"0000002e000000000000002d000000000000006a000000000000008b00000000",
            INIT_2A => X"0000000f00000000000000090000000000000003000000000000001c00000000",
            INIT_2B => X"000000b400000000000000a20000000000000036000000000000001e00000000",
            INIT_2C => X"00000015000000000000007100000000000000be00000000000000ac00000000",
            INIT_2D => X"0000009500000000000000300000000000000015000000000000001400000000",
            INIT_2E => X"00000085000000000000008e00000000000000ab00000000000000bb00000000",
            INIT_2F => X"0000002700000000000000150000000000000043000000000000008000000000",
            INIT_30 => X"0000001a00000000000000670000000000000084000000000000007c00000000",
            INIT_31 => X"000000300000000000000034000000000000006c000000000000004800000000",
            INIT_32 => X"0000003b000000000000000b0000000000000007000000000000001200000000",
            INIT_33 => X"000000b000000000000000a50000000000000063000000000000005a00000000",
            INIT_34 => X"0000001d000000000000002a00000000000000a900000000000000b100000000",
            INIT_35 => X"00000046000000000000000e0000000000000026000000000000002f00000000",
            INIT_36 => X"0000007500000000000000750000000000000088000000000000009500000000",
            INIT_37 => X"000000300000000000000015000000000000000e000000000000003c00000000",
            INIT_38 => X"0000001e0000000000000049000000000000007c000000000000007900000000",
            INIT_39 => X"0000001f00000000000000440000000000000072000000000000003b00000000",
            INIT_3A => X"000000480000000000000018000000000000000e000000000000000d00000000",
            INIT_3B => X"000000bb00000000000000bb000000000000006c000000000000004f00000000",
            INIT_3C => X"0000002b000000000000001b000000000000008b00000000000000bf00000000",
            INIT_3D => X"0000001b000000000000001c000000000000001b000000000000001e00000000",
            INIT_3E => X"00000059000000000000007b0000000000000084000000000000006c00000000",
            INIT_3F => X"0000003b000000000000002a0000000000000015000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003f00000000000000470000000000000066000000000000006d00000000",
            INIT_41 => X"0000001c000000000000004d0000000000000071000000000000003c00000000",
            INIT_42 => X"000000470000000000000030000000000000001f000000000000001000000000",
            INIT_43 => X"000000b300000000000000bd0000000000000088000000000000004600000000",
            INIT_44 => X"00000036000000000000001f000000000000007400000000000000b400000000",
            INIT_45 => X"0000000e000000000000001b0000000000000029000000000000003500000000",
            INIT_46 => X"0000003c000000000000007c0000000000000085000000000000004800000000",
            INIT_47 => X"0000003b00000000000000320000000000000022000000000000001200000000",
            INIT_48 => X"0000003c000000000000003d0000000000000051000000000000005700000000",
            INIT_49 => X"00000015000000000000004b0000000000000069000000000000003a00000000",
            INIT_4A => X"00000060000000000000004c000000000000002e000000000000001400000000",
            INIT_4B => X"000000a300000000000000a40000000000000091000000000000006100000000",
            INIT_4C => X"000000390000000000000020000000000000007100000000000000aa00000000",
            INIT_4D => X"0000001100000000000000250000000000000031000000000000004700000000",
            INIT_4E => X"000000210000000000000060000000000000006c000000000000002900000000",
            INIT_4F => X"000000320000000000000028000000000000001d000000000000000c00000000",
            INIT_50 => X"0000003c00000000000000400000000000000049000000000000004900000000",
            INIT_51 => X"0000002f0000000000000057000000000000005f000000000000003900000000",
            INIT_52 => X"000000a500000000000000890000000000000062000000000000003d00000000",
            INIT_53 => X"000000b600000000000000b700000000000000b000000000000000a900000000",
            INIT_54 => X"000000360000000000000022000000000000007c00000000000000b600000000",
            INIT_55 => X"0000001b0000000000000033000000000000005c000000000000006000000000",
            INIT_56 => X"0000000c000000000000003b0000000000000046000000000000001100000000",
            INIT_57 => X"00000028000000000000001d0000000000000012000000000000000600000000",
            INIT_58 => X"0000004e00000000000000450000000000000049000000000000004900000000",
            INIT_59 => X"0000002f00000000000000450000000000000059000000000000004100000000",
            INIT_5A => X"00000056000000000000004a000000000000003c000000000000003400000000",
            INIT_5B => X"0000006000000000000000620000000000000060000000000000005b00000000",
            INIT_5C => X"0000003c00000000000000200000000000000053000000000000006200000000",
            INIT_5D => X"00000014000000000000001d000000000000003e000000000000003b00000000",
            INIT_5E => X"00000003000000000000000a0000000000000011000000000000000400000000",
            INIT_5F => X"000000210000000000000011000000000000000a000000000000000700000000",
            INIT_60 => X"0000003600000000000000480000000000000053000000000000004b00000000",
            INIT_61 => X"00000004000000000000000f0000000000000027000000000000002d00000000",
            INIT_62 => X"0000000700000000000000050000000000000002000000000000000300000000",
            INIT_63 => X"0000000b000000000000000a0000000000000008000000000000000700000000",
            INIT_64 => X"000000420000000000000008000000000000000d000000000000000b00000000",
            INIT_65 => X"0000000f0000000000000038000000000000002f000000000000004300000000",
            INIT_66 => X"0000000300000000000000010000000000000002000000000000000200000000",
            INIT_67 => X"00000020000000000000000f000000000000000a000000000000000600000000",
            INIT_68 => X"0000002f00000000000000510000000000000059000000000000005000000000",
            INIT_69 => X"000000190000000000000010000000000000000a000000000000001500000000",
            INIT_6A => X"0000000e000000000000000e000000000000000a000000000000000e00000000",
            INIT_6B => X"0000000c000000000000000e000000000000000e000000000000000e00000000",
            INIT_6C => X"0000001700000000000000060000000000000009000000000000000a00000000",
            INIT_6D => X"00000007000000000000002a0000000000000048000000000000003e00000000",
            INIT_6E => X"0000000500000000000000050000000000000004000000000000000300000000",
            INIT_6F => X"000000210000000000000015000000000000000b000000000000000700000000",
            INIT_70 => X"000000370000000000000049000000000000004f000000000000004900000000",
            INIT_71 => X"0000003a000000000000003b000000000000002f000000000000002e00000000",
            INIT_72 => X"0000001c00000000000000190000000000000011000000000000001a00000000",
            INIT_73 => X"0000001c000000000000001d0000000000000020000000000000001f00000000",
            INIT_74 => X"0000000c00000000000000100000000000000015000000000000001800000000",
            INIT_75 => X"0000000600000000000000080000000000000016000000000000001400000000",
            INIT_76 => X"0000000800000000000000080000000000000007000000000000000800000000",
            INIT_77 => X"0000001f000000000000001b000000000000000f000000000000000b00000000",
            INIT_78 => X"0000004e000000000000004c0000000000000048000000000000004500000000",
            INIT_79 => X"0000003800000000000000480000000000000053000000000000005800000000",
            INIT_7A => X"0000002a000000000000002b0000000000000026000000000000002000000000",
            INIT_7B => X"0000003100000000000000320000000000000033000000000000002f00000000",
            INIT_7C => X"0000001c000000000000001e0000000000000026000000000000002c00000000",
            INIT_7D => X"0000000c00000000000000130000000000000022000000000000002200000000",
            INIT_7E => X"0000000d000000000000000f0000000000000010000000000000000e00000000",
            INIT_7F => X"0000001d000000000000001e000000000000001a000000000000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "sampleifmap_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003a00000000000000390000000000000031000000000000002500000000",
            INIT_01 => X"000000510000000000000050000000000000004e000000000000004200000000",
            INIT_02 => X"0000004200000000000000490000000000000052000000000000005600000000",
            INIT_03 => X"0000003800000000000000430000000000000043000000000000004100000000",
            INIT_04 => X"0000007300000000000000400000000000000032000000000000003200000000",
            INIT_05 => X"0000002700000000000000320000000000000038000000000000003400000000",
            INIT_06 => X"00000024000000000000002e0000000000000022000000000000001600000000",
            INIT_07 => X"0000001300000000000000150000000000000012000000000000001d00000000",
            INIT_08 => X"00000044000000000000004d0000000000000048000000000000004300000000",
            INIT_09 => X"000000420000000000000048000000000000004a000000000000004300000000",
            INIT_0A => X"0000003400000000000000390000000000000040000000000000004400000000",
            INIT_0B => X"0000002e00000000000000370000000000000036000000000000003200000000",
            INIT_0C => X"000000290000000000000027000000000000002a000000000000002900000000",
            INIT_0D => X"00000021000000000000001e0000000000000023000000000000002800000000",
            INIT_0E => X"0000001b000000000000001e000000000000002e000000000000002200000000",
            INIT_0F => X"0000001200000000000000160000000000000015000000000000001c00000000",
            INIT_10 => X"0000003e00000000000000480000000000000044000000000000004800000000",
            INIT_11 => X"000000310000000000000038000000000000003d000000000000003a00000000",
            INIT_12 => X"00000028000000000000002b000000000000002d000000000000003000000000",
            INIT_13 => X"00000026000000000000002b000000000000002a000000000000002600000000",
            INIT_14 => X"0000001c000000000000001e0000000000000023000000000000002200000000",
            INIT_15 => X"00000022000000000000001f0000000000000021000000000000002300000000",
            INIT_16 => X"0000000e000000000000000d0000000000000022000000000000003000000000",
            INIT_17 => X"0000001100000000000000130000000000000014000000000000001500000000",
            INIT_18 => X"0000003c000000000000003d0000000000000036000000000000003800000000",
            INIT_19 => X"00000024000000000000002b0000000000000030000000000000003e00000000",
            INIT_1A => X"0000002000000000000000220000000000000023000000000000002300000000",
            INIT_1B => X"0000002000000000000000220000000000000021000000000000001f00000000",
            INIT_1C => X"0000001d000000000000001b000000000000001e000000000000001d00000000",
            INIT_1D => X"00000025000000000000001d000000000000001c000000000000002000000000",
            INIT_1E => X"0000000f000000000000000b0000000000000012000000000000002a00000000",
            INIT_1F => X"0000001100000000000000100000000000000013000000000000001600000000",
            INIT_20 => X"0000003b00000000000000420000000000000039000000000000003900000000",
            INIT_21 => X"0000001b00000000000000200000000000000024000000000000003400000000",
            INIT_22 => X"0000001a000000000000001c000000000000001d000000000000001c00000000",
            INIT_23 => X"0000001e000000000000001c000000000000001a000000000000001a00000000",
            INIT_24 => X"0000001c000000000000001c000000000000001c000000000000001c00000000",
            INIT_25 => X"0000002a00000000000000430000000000000030000000000000001c00000000",
            INIT_26 => X"00000019000000000000000d0000000000000012000000000000001900000000",
            INIT_27 => X"000000110000000000000013000000000000001f000000000000001b00000000",
            INIT_28 => X"00000021000000000000002f000000000000003a000000000000003b00000000",
            INIT_29 => X"000000160000000000000019000000000000001a000000000000001a00000000",
            INIT_2A => X"00000019000000000000001a0000000000000019000000000000001700000000",
            INIT_2B => X"0000001f000000000000001b0000000000000018000000000000001800000000",
            INIT_2C => X"0000001e0000000000000021000000000000001e000000000000001d00000000",
            INIT_2D => X"0000003c000000000000005e000000000000005d000000000000002100000000",
            INIT_2E => X"0000002c000000000000001e000000000000001b000000000000002900000000",
            INIT_2F => X"000000130000000000000018000000000000002d000000000000002b00000000",
            INIT_30 => X"000000140000000000000017000000000000001c000000000000002200000000",
            INIT_31 => X"0000001500000000000000160000000000000017000000000000001600000000",
            INIT_32 => X"0000001a00000000000000190000000000000016000000000000001600000000",
            INIT_33 => X"00000023000000000000001d0000000000000019000000000000001800000000",
            INIT_34 => X"0000001e0000000000000023000000000000001f000000000000002000000000",
            INIT_35 => X"0000002500000000000000370000000000000059000000000000003300000000",
            INIT_36 => X"0000002d000000000000002b0000000000000028000000000000003800000000",
            INIT_37 => X"000000150000000000000017000000000000001e000000000000002400000000",
            INIT_38 => X"0000001200000000000000100000000000000011000000000000001100000000",
            INIT_39 => X"0000001600000000000000160000000000000017000000000000001600000000",
            INIT_3A => X"0000001b000000000000001a0000000000000017000000000000001800000000",
            INIT_3B => X"00000027000000000000001d000000000000001b000000000000001900000000",
            INIT_3C => X"000000300000000000000033000000000000002d000000000000002800000000",
            INIT_3D => X"0000000b00000000000000120000000000000040000000000000004100000000",
            INIT_3E => X"00000020000000000000001f0000000000000025000000000000002200000000",
            INIT_3F => X"0000001500000000000000160000000000000016000000000000001900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000000000120000000000000012000000000000001100000000",
            INIT_41 => X"0000001700000000000000170000000000000016000000000000001500000000",
            INIT_42 => X"0000001e000000000000001c0000000000000018000000000000001900000000",
            INIT_43 => X"0000003b00000000000000330000000000000038000000000000002500000000",
            INIT_44 => X"000000360000000000000037000000000000003a000000000000003b00000000",
            INIT_45 => X"0000001000000000000000110000000000000028000000000000003d00000000",
            INIT_46 => X"0000001b00000000000000180000000000000019000000000000001a00000000",
            INIT_47 => X"0000001400000000000000150000000000000017000000000000001a00000000",
            INIT_48 => X"0000001200000000000000120000000000000012000000000000001300000000",
            INIT_49 => X"0000001800000000000000160000000000000014000000000000001500000000",
            INIT_4A => X"0000003100000000000000200000000000000019000000000000001800000000",
            INIT_4B => X"000000340000000000000039000000000000004c000000000000003e00000000",
            INIT_4C => X"0000003a0000000000000032000000000000002e000000000000003100000000",
            INIT_4D => X"0000002c00000000000000300000000000000031000000000000003800000000",
            INIT_4E => X"0000001900000000000000190000000000000023000000000000002900000000",
            INIT_4F => X"0000001400000000000000140000000000000018000000000000001900000000",
            INIT_50 => X"0000001200000000000000130000000000000012000000000000001400000000",
            INIT_51 => X"0000001700000000000000150000000000000015000000000000001500000000",
            INIT_52 => X"0000003500000000000000240000000000000019000000000000001900000000",
            INIT_53 => X"0000004a000000000000003e0000000000000042000000000000003100000000",
            INIT_54 => X"000000b800000000000000a60000000000000089000000000000006800000000",
            INIT_55 => X"00000021000000000000004b0000000000000068000000000000007c00000000",
            INIT_56 => X"000000190000000000000026000000000000003d000000000000003800000000",
            INIT_57 => X"0000001300000000000000120000000000000019000000000000001800000000",
            INIT_58 => X"0000001300000000000000140000000000000012000000000000001500000000",
            INIT_59 => X"0000001800000000000000160000000000000018000000000000001800000000",
            INIT_5A => X"00000030000000000000001f000000000000001d000000000000001900000000",
            INIT_5B => X"000000be00000000000000b20000000000000097000000000000005500000000",
            INIT_5C => X"000000c500000000000000ca00000000000000cd00000000000000cd00000000",
            INIT_5D => X"00000016000000000000009800000000000000d000000000000000b200000000",
            INIT_5E => X"0000002800000000000000460000000000000025000000000000001800000000",
            INIT_5F => X"0000001100000000000000110000000000000016000000000000001500000000",
            INIT_60 => X"0000001500000000000000160000000000000014000000000000001400000000",
            INIT_61 => X"0000001a00000000000000190000000000000018000000000000001800000000",
            INIT_62 => X"0000007000000000000000420000000000000020000000000000001900000000",
            INIT_63 => X"00000075000000000000008c000000000000009b000000000000009000000000",
            INIT_64 => X"0000003d00000000000000470000000000000058000000000000006400000000",
            INIT_65 => X"0000004e00000000000000d500000000000000e8000000000000007500000000",
            INIT_66 => X"000000460000000000000032000000000000000a000000000000000f00000000",
            INIT_67 => X"0000001000000000000000110000000000000015000000000000001a00000000",
            INIT_68 => X"0000001600000000000000190000000000000016000000000000001400000000",
            INIT_69 => X"0000001a00000000000000190000000000000017000000000000001700000000",
            INIT_6A => X"0000005b00000000000000670000000000000048000000000000001a00000000",
            INIT_6B => X"0000001200000000000000340000000000000056000000000000005000000000",
            INIT_6C => X"00000010000000000000000f0000000000000022000000000000001100000000",
            INIT_6D => X"0000009b00000000000000e000000000000000dd000000000000007c00000000",
            INIT_6E => X"0000003b00000000000000160000000000000007000000000000002400000000",
            INIT_6F => X"0000001000000000000000120000000000000013000000000000002100000000",
            INIT_70 => X"00000016000000000000001b0000000000000017000000000000001800000000",
            INIT_71 => X"0000001500000000000000130000000000000019000000000000001800000000",
            INIT_72 => X"00000029000000000000003a0000000000000055000000000000003700000000",
            INIT_73 => X"000000180000000000000032000000000000004e000000000000003d00000000",
            INIT_74 => X"00000049000000000000001e000000000000002b000000000000000b00000000",
            INIT_75 => X"000000cd00000000000000d100000000000000d800000000000000bf00000000",
            INIT_76 => X"000000170000000000000010000000000000000e000000000000006700000000",
            INIT_77 => X"0000001200000000000000140000000000000016000000000000001b00000000",
            INIT_78 => X"00000017000000000000001a0000000000000016000000000000001a00000000",
            INIT_79 => X"00000034000000000000003c0000000000000025000000000000001900000000",
            INIT_7A => X"0000003b00000000000000380000000000000034000000000000004c00000000",
            INIT_7B => X"00000026000000000000002e000000000000004d000000000000005000000000",
            INIT_7C => X"000000c4000000000000007c0000000000000049000000000000002300000000",
            INIT_7D => X"000000d200000000000000d900000000000000d800000000000000df00000000",
            INIT_7E => X"0000000e00000000000000150000000000000039000000000000007600000000",
            INIT_7F => X"00000011000000000000003e0000000000000047000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "sampleifmap_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001700000000000000190000000000000014000000000000001900000000",
            INIT_01 => X"0000005c00000000000000600000000000000035000000000000002100000000",
            INIT_02 => X"00000042000000000000003e000000000000005d000000000000004900000000",
            INIT_03 => X"000000a2000000000000005a0000000000000047000000000000005100000000",
            INIT_04 => X"000000f500000000000000f500000000000000df00000000000000c400000000",
            INIT_05 => X"0000007900000000000000de00000000000000e400000000000000e300000000",
            INIT_06 => X"000000090000000000000011000000000000003b000000000000002500000000",
            INIT_07 => X"000000130000000000000075000000000000008c000000000000004800000000",
            INIT_08 => X"0000001a00000000000000180000000000000015000000000000001900000000",
            INIT_09 => X"000000450000000000000035000000000000002c000000000000002800000000",
            INIT_0A => X"0000002900000000000000250000000000000052000000000000005800000000",
            INIT_0B => X"000000fb00000000000000940000000000000020000000000000003100000000",
            INIT_0C => X"000000e200000000000000e900000000000000f200000000000000f600000000",
            INIT_0D => X"0000001f000000000000008b00000000000000e200000000000000e100000000",
            INIT_0E => X"0000004300000000000000280000000000000019000000000000000b00000000",
            INIT_0F => X"00000022000000000000009700000000000000a2000000000000008500000000",
            INIT_10 => X"0000002600000000000000160000000000000013000000000000001600000000",
            INIT_11 => X"00000036000000000000002e0000000000000046000000000000005d00000000",
            INIT_12 => X"0000001b00000000000000180000000000000026000000000000004b00000000",
            INIT_13 => X"000000e300000000000000a30000000000000031000000000000003800000000",
            INIT_14 => X"000000da00000000000000cb00000000000000cd00000000000000d600000000",
            INIT_15 => X"0000004a00000000000000a300000000000000e400000000000000e500000000",
            INIT_16 => X"000000950000000000000080000000000000005a000000000000003900000000",
            INIT_17 => X"0000003300000000000000a00000000000000096000000000000009700000000",
            INIT_18 => X"0000007c0000000000000026000000000000000f000000000000001300000000",
            INIT_19 => X"0000002a0000000000000024000000000000005a00000000000000af00000000",
            INIT_1A => X"00000015000000000000000b0000000000000017000000000000003f00000000",
            INIT_1B => X"000000d000000000000000aa000000000000004f000000000000004000000000",
            INIT_1C => X"000000d600000000000000d300000000000000c500000000000000c700000000",
            INIT_1D => X"000000b100000000000000e300000000000000d900000000000000ce00000000",
            INIT_1E => X"000000a200000000000000a700000000000000a8000000000000009800000000",
            INIT_1F => X"0000002a00000000000000880000000000000097000000000000009a00000000",
            INIT_20 => X"000000dc0000000000000065000000000000000a000000000000001200000000",
            INIT_21 => X"0000002e000000000000002f000000000000006f00000000000000be00000000",
            INIT_22 => X"0000000e0000000000000009000000000000000a000000000000003900000000",
            INIT_23 => X"000000cc00000000000000b10000000000000042000000000000001f00000000",
            INIT_24 => X"0000007c00000000000000c600000000000000ca00000000000000c200000000",
            INIT_25 => X"000000d300000000000000ac0000000000000066000000000000004f00000000",
            INIT_26 => X"000000a900000000000000b100000000000000b800000000000000c800000000",
            INIT_27 => X"00000011000000000000004a000000000000008c000000000000009c00000000",
            INIT_28 => X"000000a500000000000000840000000000000014000000000000000e00000000",
            INIT_29 => X"0000003400000000000000370000000000000080000000000000009600000000",
            INIT_2A => X"00000016000000000000000a0000000000000003000000000000001e00000000",
            INIT_2B => X"000000c600000000000000b40000000000000048000000000000002d00000000",
            INIT_2C => X"00000019000000000000007b00000000000000cd00000000000000be00000000",
            INIT_2D => X"000000a30000000000000038000000000000001e000000000000001a00000000",
            INIT_2E => X"00000093000000000000009e00000000000000b800000000000000ca00000000",
            INIT_2F => X"00000011000000000000000d0000000000000044000000000000008800000000",
            INIT_30 => X"0000002100000000000000530000000000000023000000000000000a00000000",
            INIT_31 => X"00000035000000000000003e0000000000000082000000000000005300000000",
            INIT_32 => X"0000004800000000000000100000000000000007000000000000001300000000",
            INIT_33 => X"000000c200000000000000b70000000000000075000000000000006c00000000",
            INIT_34 => X"0000001e000000000000002f00000000000000b700000000000000c300000000",
            INIT_35 => X"0000004f0000000000000014000000000000002b000000000000003100000000",
            INIT_36 => X"000000810000000000000084000000000000009400000000000000a100000000",
            INIT_37 => X"000000180000000000000009000000000000000a000000000000004000000000",
            INIT_38 => X"0000002300000000000000370000000000000021000000000000000a00000000",
            INIT_39 => X"00000024000000000000004e0000000000000088000000000000004600000000",
            INIT_3A => X"0000005800000000000000220000000000000011000000000000000f00000000",
            INIT_3B => X"000000cd00000000000000cd000000000000007e000000000000006100000000",
            INIT_3C => X"0000002b0000000000000020000000000000009800000000000000d000000000",
            INIT_3D => X"0000001f0000000000000020000000000000001f000000000000002000000000",
            INIT_3E => X"00000063000000000000008a0000000000000091000000000000007500000000",
            INIT_3F => X"000000210000000000000019000000000000000c000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004100000000000000360000000000000015000000000000000a00000000",
            INIT_41 => X"0000002100000000000000570000000000000088000000000000004700000000",
            INIT_42 => X"00000057000000000000003f0000000000000027000000000000001500000000",
            INIT_43 => X"000000c500000000000000cf000000000000009a000000000000005600000000",
            INIT_44 => X"000000380000000000000025000000000000008100000000000000c600000000",
            INIT_45 => X"0000000f000000000000001c000000000000002c000000000000003700000000",
            INIT_46 => X"00000043000000000000008b0000000000000093000000000000004d00000000",
            INIT_47 => X"0000001f000000000000001c0000000000000014000000000000000e00000000",
            INIT_48 => X"0000003e000000000000002f000000000000000e000000000000000700000000",
            INIT_49 => X"0000001c00000000000000560000000000000080000000000000004500000000",
            INIT_4A => X"0000006f000000000000005e000000000000003c000000000000001e00000000",
            INIT_4B => X"000000b400000000000000b600000000000000a2000000000000006f00000000",
            INIT_4C => X"0000003c0000000000000029000000000000007f00000000000000bc00000000",
            INIT_4D => X"0000000f00000000000000230000000000000035000000000000004b00000000",
            INIT_4E => X"00000026000000000000006f000000000000007a000000000000002c00000000",
            INIT_4F => X"000000160000000000000010000000000000000d000000000000000700000000",
            INIT_50 => X"0000003b00000000000000270000000000000011000000000000000b00000000",
            INIT_51 => X"0000003d00000000000000680000000000000075000000000000004600000000",
            INIT_52 => X"000000b7000000000000009f0000000000000079000000000000005100000000",
            INIT_53 => X"000000c700000000000000c900000000000000c300000000000000b900000000",
            INIT_54 => X"0000003c000000000000002a000000000000008800000000000000c600000000",
            INIT_55 => X"0000001c00000000000000340000000000000062000000000000006600000000",
            INIT_56 => X"000000100000000000000045000000000000004f000000000000001500000000",
            INIT_57 => X"00000016000000000000000c0000000000000007000000000000000300000000",
            INIT_58 => X"00000043000000000000001d0000000000000014000000000000001300000000",
            INIT_59 => X"0000003c00000000000000550000000000000067000000000000004900000000",
            INIT_5A => X"00000064000000000000005b0000000000000050000000000000004500000000",
            INIT_5B => X"0000006d00000000000000710000000000000071000000000000006800000000",
            INIT_5C => X"0000004100000000000000250000000000000059000000000000006d00000000",
            INIT_5D => X"00000017000000000000001f0000000000000042000000000000004000000000",
            INIT_5E => X"00000005000000000000000e0000000000000014000000000000000800000000",
            INIT_5F => X"00000018000000000000000b0000000000000006000000000000000600000000",
            INIT_60 => X"00000025000000000000001d000000000000001c000000000000001700000000",
            INIT_61 => X"000000070000000000000016000000000000002c000000000000002c00000000",
            INIT_62 => X"0000000c000000000000000c000000000000000a000000000000000a00000000",
            INIT_63 => X"0000001000000000000000110000000000000010000000000000000d00000000",
            INIT_64 => X"000000430000000000000009000000000000000f000000000000000f00000000",
            INIT_65 => X"0000001000000000000000380000000000000030000000000000004400000000",
            INIT_66 => X"0000000400000000000000030000000000000003000000000000000400000000",
            INIT_67 => X"00000019000000000000000e0000000000000009000000000000000600000000",
            INIT_68 => X"0000002000000000000000270000000000000025000000000000002100000000",
            INIT_69 => X"0000002000000000000000190000000000000012000000000000001700000000",
            INIT_6A => X"0000001700000000000000170000000000000015000000000000001700000000",
            INIT_6B => X"0000000f00000000000000130000000000000015000000000000001700000000",
            INIT_6C => X"000000180000000000000007000000000000000a000000000000000b00000000",
            INIT_6D => X"0000000800000000000000290000000000000047000000000000003e00000000",
            INIT_6E => X"0000000600000000000000050000000000000005000000000000000400000000",
            INIT_6F => X"0000001d0000000000000018000000000000000e000000000000000900000000",
            INIT_70 => X"0000003200000000000000290000000000000025000000000000002300000000",
            INIT_71 => X"0000004d00000000000000510000000000000043000000000000003c00000000",
            INIT_72 => X"00000030000000000000002d0000000000000024000000000000002c00000000",
            INIT_73 => X"000000230000000000000027000000000000002c000000000000003100000000",
            INIT_74 => X"000000100000000000000015000000000000001b000000000000001d00000000",
            INIT_75 => X"00000009000000000000000a0000000000000019000000000000001700000000",
            INIT_76 => X"0000000b000000000000000a0000000000000009000000000000000b00000000",
            INIT_77 => X"0000001e000000000000001f0000000000000014000000000000000e00000000",
            INIT_78 => X"00000057000000000000003b000000000000002a000000000000002a00000000",
            INIT_79 => X"000000520000000000000066000000000000006f000000000000006d00000000",
            INIT_7A => X"000000470000000000000045000000000000003e000000000000003700000000",
            INIT_7B => X"0000004300000000000000460000000000000048000000000000004a00000000",
            INIT_7C => X"00000029000000000000002b0000000000000033000000000000003b00000000",
            INIT_7D => X"000000120000000000000018000000000000002c000000000000002f00000000",
            INIT_7E => X"0000001300000000000000150000000000000016000000000000001400000000",
            INIT_7F => X"0000001e0000000000000020000000000000001c000000000000001600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "sampleifmap_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000a000000000000000e000000000000000b000000000000000d00000000",
            INIT_01 => X"000000020000000000000005000000000000000a000000000000000900000000",
            INIT_02 => X"0000000200000000000000010000000000000003000000000000000300000000",
            INIT_03 => X"0000000000000000000000050000000000000006000000000000000400000000",
            INIT_04 => X"0000005600000000000000230000000000000000000000000000000100000000",
            INIT_05 => X"00000008000000000000001d0000000000000017000000000000001600000000",
            INIT_06 => X"0000001d0000000000000027000000000000001b000000000000000d00000000",
            INIT_07 => X"0000000500000000000000060000000000000008000000000000001300000000",
            INIT_08 => X"00000004000000000000000a000000000000000c000000000000000d00000000",
            INIT_09 => X"0000000000000000000000030000000000000008000000000000000700000000",
            INIT_0A => X"0000000100000000000000010000000000000002000000000000000400000000",
            INIT_0B => X"0000000100000000000000040000000000000004000000000000000200000000",
            INIT_0C => X"0000001300000000000000100000000000000001000000000000000100000000",
            INIT_0D => X"0000000700000000000000060000000000000006000000000000000700000000",
            INIT_0E => X"000000160000000000000017000000000000002e000000000000002100000000",
            INIT_0F => X"0000000600000000000000040000000000000008000000000000001300000000",
            INIT_10 => X"0000000000000000000000030000000000000004000000000000000700000000",
            INIT_11 => X"0000000000000000000000010000000000000004000000000000000400000000",
            INIT_12 => X"0000000400000000000000040000000000000004000000000000000400000000",
            INIT_13 => X"0000000300000000000000050000000000000006000000000000000400000000",
            INIT_14 => X"00000009000000000000000c0000000000000003000000000000000400000000",
            INIT_15 => X"0000000a00000000000000060000000000000007000000000000000400000000",
            INIT_16 => X"0000000c000000000000000d0000000000000023000000000000002800000000",
            INIT_17 => X"0000000600000000000000030000000000000006000000000000000f00000000",
            INIT_18 => X"0000000b00000000000000080000000000000003000000000000000100000000",
            INIT_19 => X"0000000300000000000000030000000000000004000000000000001200000000",
            INIT_1A => X"0000000700000000000000080000000000000006000000000000000500000000",
            INIT_1B => X"0000000600000000000000060000000000000009000000000000000800000000",
            INIT_1C => X"00000009000000000000000a0000000000000005000000000000000700000000",
            INIT_1D => X"000000170000000000000010000000000000000a000000000000000400000000",
            INIT_1E => X"0000000e00000000000000110000000000000016000000000000001e00000000",
            INIT_1F => X"0000000800000000000000050000000000000006000000000000000f00000000",
            INIT_20 => X"0000001a000000000000001d0000000000000013000000000000000c00000000",
            INIT_21 => X"0000000800000000000000070000000000000006000000000000001700000000",
            INIT_22 => X"0000000800000000000000090000000000000008000000000000000700000000",
            INIT_23 => X"000000080000000000000007000000000000000a000000000000000900000000",
            INIT_24 => X"0000000700000000000000080000000000000007000000000000000900000000",
            INIT_25 => X"0000002700000000000000400000000000000025000000000000000800000000",
            INIT_26 => X"00000015000000000000000e0000000000000010000000000000001000000000",
            INIT_27 => X"00000009000000000000000d000000000000000f000000000000000e00000000",
            INIT_28 => X"0000000c0000000000000016000000000000001e000000000000001800000000",
            INIT_29 => X"0000000800000000000000090000000000000006000000000000000900000000",
            INIT_2A => X"0000000a00000000000000090000000000000005000000000000000500000000",
            INIT_2B => X"000000090000000000000007000000000000000a000000000000000b00000000",
            INIT_2C => X"00000007000000000000000b000000000000000b000000000000000a00000000",
            INIT_2D => X"0000003b000000000000005d0000000000000055000000000000001400000000",
            INIT_2E => X"000000200000000000000013000000000000000e000000000000002200000000",
            INIT_2F => X"000000090000000000000010000000000000001b000000000000001700000000",
            INIT_30 => X"00000007000000000000000a000000000000000b000000000000000c00000000",
            INIT_31 => X"00000007000000000000000a0000000000000008000000000000000800000000",
            INIT_32 => X"0000000e000000000000000a0000000000000005000000000000000600000000",
            INIT_33 => X"0000000c000000000000000a000000000000000c000000000000000d00000000",
            INIT_34 => X"00000007000000000000000e000000000000000e000000000000000900000000",
            INIT_35 => X"00000028000000000000003c0000000000000056000000000000002500000000",
            INIT_36 => X"0000001c000000000000001c000000000000001c000000000000003500000000",
            INIT_37 => X"0000000700000000000000060000000000000010000000000000001400000000",
            INIT_38 => X"0000000700000000000000060000000000000006000000000000000300000000",
            INIT_39 => X"00000009000000000000000c000000000000000a000000000000000b00000000",
            INIT_3A => X"0000000e000000000000000c0000000000000008000000000000000900000000",
            INIT_3B => X"0000001300000000000000100000000000000012000000000000000e00000000",
            INIT_3C => X"00000016000000000000001a0000000000000015000000000000001000000000",
            INIT_3D => X"0000000a0000000000000014000000000000003e000000000000003100000000",
            INIT_3E => X"0000000d0000000000000010000000000000001a000000000000001e00000000",
            INIT_3F => X"0000000700000000000000040000000000000008000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000080000000000000009000000000000000a000000000000000700000000",
            INIT_41 => X"0000000b000000000000000e000000000000000a000000000000000b00000000",
            INIT_42 => X"0000000f000000000000000e000000000000000c000000000000000d00000000",
            INIT_43 => X"0000002800000000000000220000000000000024000000000000001300000000",
            INIT_44 => X"0000002200000000000000220000000000000020000000000000002400000000",
            INIT_45 => X"00000009000000000000000f000000000000002b000000000000003300000000",
            INIT_46 => X"0000000a0000000000000009000000000000000c000000000000001400000000",
            INIT_47 => X"0000000800000000000000080000000000000008000000000000000800000000",
            INIT_48 => X"00000008000000000000000b000000000000000c000000000000000c00000000",
            INIT_49 => X"0000000d000000000000000e000000000000000a000000000000000c00000000",
            INIT_4A => X"000000220000000000000014000000000000000e000000000000000e00000000",
            INIT_4B => X"0000002600000000000000280000000000000031000000000000002700000000",
            INIT_4C => X"000000320000000000000027000000000000001b000000000000002000000000",
            INIT_4D => X"000000260000000000000034000000000000003b000000000000003600000000",
            INIT_4E => X"0000000c000000000000000b0000000000000015000000000000002300000000",
            INIT_4F => X"0000000a000000000000000b0000000000000009000000000000000600000000",
            INIT_50 => X"00000009000000000000000b000000000000000b000000000000000c00000000",
            INIT_51 => X"0000000d000000000000000d000000000000000a000000000000000c00000000",
            INIT_52 => X"00000028000000000000001b0000000000000010000000000000000d00000000",
            INIT_53 => X"0000003f00000000000000320000000000000032000000000000002000000000",
            INIT_54 => X"000000b400000000000000a10000000000000077000000000000005800000000",
            INIT_55 => X"0000002200000000000000540000000000000071000000000000007900000000",
            INIT_56 => X"00000011000000000000001d0000000000000031000000000000003200000000",
            INIT_57 => X"0000000a000000000000000c000000000000000a000000000000000900000000",
            INIT_58 => X"0000000b000000000000000e000000000000000a000000000000000900000000",
            INIT_59 => X"0000000c000000000000000d000000000000000c000000000000000e00000000",
            INIT_5A => X"0000002700000000000000180000000000000012000000000000000c00000000",
            INIT_5B => X"000000ba00000000000000af0000000000000093000000000000004d00000000",
            INIT_5C => X"000000ca00000000000000d200000000000000c800000000000000c800000000",
            INIT_5D => X"0000001c000000000000009e00000000000000d500000000000000b100000000",
            INIT_5E => X"0000002500000000000000460000000000000022000000000000001300000000",
            INIT_5F => X"00000009000000000000000b0000000000000009000000000000000a00000000",
            INIT_60 => X"0000000d000000000000000f000000000000000a000000000000000800000000",
            INIT_61 => X"0000000e000000000000000d000000000000000e000000000000001000000000",
            INIT_62 => X"0000006c000000000000003e0000000000000018000000000000000c00000000",
            INIT_63 => X"0000007d000000000000009300000000000000a2000000000000008e00000000",
            INIT_64 => X"0000004a0000000000000054000000000000005e000000000000006e00000000",
            INIT_65 => X"0000005400000000000000d700000000000000f1000000000000007e00000000",
            INIT_66 => X"0000004900000000000000340000000000000009000000000000000c00000000",
            INIT_67 => X"000000080000000000000009000000000000000d000000000000001900000000",
            INIT_68 => X"0000000e000000000000000f000000000000000b000000000000000b00000000",
            INIT_69 => X"0000000e000000000000000c0000000000000010000000000000001100000000",
            INIT_6A => X"0000005d00000000000000670000000000000044000000000000001400000000",
            INIT_6B => X"00000019000000000000003d000000000000005f000000000000005600000000",
            INIT_6C => X"0000001700000000000000110000000000000023000000000000001600000000",
            INIT_6D => X"000000a700000000000000eb00000000000000eb000000000000008900000000",
            INIT_6E => X"0000004200000000000000170000000000000007000000000000002a00000000",
            INIT_6F => X"0000000700000000000000090000000000000011000000000000002800000000",
            INIT_70 => X"0000000e0000000000000012000000000000000d000000000000000f00000000",
            INIT_71 => X"00000012000000000000000b0000000000000012000000000000001000000000",
            INIT_72 => X"0000002e000000000000003b0000000000000053000000000000003600000000",
            INIT_73 => X"0000001b00000000000000370000000000000053000000000000004400000000",
            INIT_74 => X"0000004c000000000000001c0000000000000027000000000000000c00000000",
            INIT_75 => X"000000e000000000000000e700000000000000e800000000000000c800000000",
            INIT_76 => X"0000001a00000000000000130000000000000016000000000000007300000000",
            INIT_77 => X"00000008000000000000000d0000000000000016000000000000001f00000000",
            INIT_78 => X"0000000e0000000000000013000000000000000d000000000000001000000000",
            INIT_79 => X"000000370000000000000039000000000000001e000000000000000e00000000",
            INIT_7A => X"0000003c00000000000000390000000000000035000000000000004f00000000",
            INIT_7B => X"000000290000000000000032000000000000004e000000000000005200000000",
            INIT_7C => X"000000c8000000000000007c0000000000000047000000000000002300000000",
            INIT_7D => X"000000dd00000000000000ec00000000000000e600000000000000e700000000",
            INIT_7E => X"0000000e000000000000001a0000000000000044000000000000007e00000000",
            INIT_7F => X"00000009000000000000003f0000000000000049000000000000002000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "sampleifmap_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000110000000000000013000000000000000e000000000000001100000000",
            INIT_01 => X"0000005c000000000000005d000000000000002f000000000000001800000000",
            INIT_02 => X"0000003d000000000000003c0000000000000062000000000000004f00000000",
            INIT_03 => X"000000a6000000000000005e0000000000000047000000000000004c00000000",
            INIT_04 => X"000000fc00000000000000fa00000000000000e200000000000000c600000000",
            INIT_05 => X"0000007c00000000000000e700000000000000f000000000000000ed00000000",
            INIT_06 => X"0000000c000000000000001c000000000000004a000000000000002a00000000",
            INIT_07 => X"00000011000000000000007e0000000000000095000000000000004c00000000",
            INIT_08 => X"0000001500000000000000120000000000000010000000000000001200000000",
            INIT_09 => X"000000480000000000000038000000000000002a000000000000002400000000",
            INIT_0A => X"0000002400000000000000240000000000000058000000000000006000000000",
            INIT_0B => X"00000100000000000000009a0000000000000022000000000000002d00000000",
            INIT_0C => X"000000ed00000000000000f400000000000000f900000000000000fa00000000",
            INIT_0D => X"00000027000000000000009600000000000000ee00000000000000ed00000000",
            INIT_0E => X"0000004d000000000000003b000000000000002e000000000000001500000000",
            INIT_0F => X"0000002600000000000000a300000000000000ae000000000000008e00000000",
            INIT_10 => X"0000002200000000000000100000000000000010000000000000001100000000",
            INIT_11 => X"00000042000000000000003c0000000000000049000000000000005c00000000",
            INIT_12 => X"00000021000000000000001c000000000000002c000000000000005400000000",
            INIT_13 => X"000000f000000000000000ae0000000000000037000000000000003e00000000",
            INIT_14 => X"000000e700000000000000d900000000000000d900000000000000e100000000",
            INIT_15 => X"0000005600000000000000b100000000000000ee00000000000000ef00000000",
            INIT_16 => X"000000a40000000000000092000000000000006a000000000000004500000000",
            INIT_17 => X"0000003700000000000000a900000000000000a100000000000000a400000000",
            INIT_18 => X"0000007d0000000000000020000000000000000a000000000000000d00000000",
            INIT_19 => X"000000380000000000000035000000000000006200000000000000b400000000",
            INIT_1A => X"0000001b000000000000000e000000000000001c000000000000004800000000",
            INIT_1B => X"000000e000000000000000b90000000000000059000000000000004900000000",
            INIT_1C => X"000000e300000000000000e400000000000000d500000000000000d500000000",
            INIT_1D => X"000000c000000000000000f200000000000000e100000000000000d700000000",
            INIT_1E => X"000000b000000000000000b500000000000000b400000000000000a500000000",
            INIT_1F => X"0000002a000000000000008d000000000000009f00000000000000a600000000",
            INIT_20 => X"000000e500000000000000650000000000000007000000000000000c00000000",
            INIT_21 => X"00000039000000000000003e000000000000007b00000000000000c900000000",
            INIT_22 => X"0000000f0000000000000009000000000000000f000000000000004100000000",
            INIT_23 => X"000000da00000000000000bf000000000000004f000000000000002600000000",
            INIT_24 => X"0000008a00000000000000d800000000000000db00000000000000d000000000",
            INIT_25 => X"000000e400000000000000b8000000000000006d000000000000005800000000",
            INIT_26 => X"000000b500000000000000bf00000000000000c900000000000000da00000000",
            INIT_27 => X"0000000e000000000000004d000000000000009300000000000000a600000000",
            INIT_28 => X"000000b3000000000000008b0000000000000018000000000000000d00000000",
            INIT_29 => X"0000003d0000000000000045000000000000008d00000000000000a200000000",
            INIT_2A => X"0000001b000000000000000b0000000000000004000000000000002300000000",
            INIT_2B => X"000000d400000000000000c20000000000000056000000000000003600000000",
            INIT_2C => X"00000024000000000000008800000000000000db00000000000000cc00000000",
            INIT_2D => X"000000b100000000000000400000000000000022000000000000002000000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000cc00000000000000dd00000000",
            INIT_2F => X"0000000d000000000000000f0000000000000049000000000000009000000000",
            INIT_30 => X"00000031000000000000005b0000000000000027000000000000000900000000",
            INIT_31 => X"0000003e000000000000004c000000000000008f000000000000006000000000",
            INIT_32 => X"0000005100000000000000150000000000000007000000000000001500000000",
            INIT_33 => X"000000d000000000000000c50000000000000083000000000000007900000000",
            INIT_34 => X"00000026000000000000003800000000000000c100000000000000d100000000",
            INIT_35 => X"000000590000000000000019000000000000002e000000000000003700000000",
            INIT_36 => X"0000008d000000000000009500000000000000a900000000000000b200000000",
            INIT_37 => X"000000140000000000000008000000000000000e000000000000004800000000",
            INIT_38 => X"00000030000000000000003b0000000000000022000000000000000500000000",
            INIT_39 => X"0000002d000000000000005c0000000000000095000000000000005300000000",
            INIT_3A => X"00000064000000000000002a0000000000000013000000000000000f00000000",
            INIT_3B => X"000000db00000000000000db000000000000008c000000000000006f00000000",
            INIT_3C => X"00000033000000000000002600000000000000a000000000000000de00000000",
            INIT_3D => X"0000002700000000000000240000000000000023000000000000002500000000",
            INIT_3E => X"0000006e000000000000009b00000000000000a4000000000000008200000000",
            INIT_3F => X"0000001e0000000000000016000000000000000c000000000000001d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d000000000000003a0000000000000017000000000000000700000000",
            INIT_41 => X"0000002a00000000000000650000000000000094000000000000005400000000",
            INIT_42 => X"00000065000000000000004a000000000000002b000000000000001600000000",
            INIT_43 => X"000000d300000000000000dd00000000000000a8000000000000006400000000",
            INIT_44 => X"00000040000000000000002b000000000000008900000000000000d400000000",
            INIT_45 => X"0000001500000000000000230000000000000034000000000000003f00000000",
            INIT_46 => X"0000004e000000000000009a00000000000000a2000000000000005600000000",
            INIT_47 => X"0000001c00000000000000180000000000000012000000000000001300000000",
            INIT_48 => X"0000004c00000000000000370000000000000015000000000000000900000000",
            INIT_49 => X"000000250000000000000065000000000000008c000000000000005200000000",
            INIT_4A => X"0000007f000000000000006c0000000000000043000000000000002100000000",
            INIT_4B => X"000000c200000000000000c300000000000000b0000000000000007e00000000",
            INIT_4C => X"000000460000000000000030000000000000008700000000000000c900000000",
            INIT_4D => X"00000015000000000000002e0000000000000041000000000000005600000000",
            INIT_4E => X"00000031000000000000007b0000000000000083000000000000003200000000",
            INIT_4F => X"00000014000000000000000b000000000000000a000000000000000b00000000",
            INIT_50 => X"0000004900000000000000310000000000000017000000000000000b00000000",
            INIT_51 => X"0000004b00000000000000780000000000000084000000000000005700000000",
            INIT_52 => X"000000c800000000000000b10000000000000086000000000000005d00000000",
            INIT_53 => X"000000d500000000000000d400000000000000cf00000000000000c800000000",
            INIT_54 => X"000000480000000000000035000000000000009400000000000000d600000000",
            INIT_55 => X"000000220000000000000040000000000000006e000000000000007100000000",
            INIT_56 => X"00000016000000000000004c0000000000000055000000000000001800000000",
            INIT_57 => X"00000016000000000000000d0000000000000009000000000000000700000000",
            INIT_58 => X"0000004e00000000000000250000000000000016000000000000000f00000000",
            INIT_59 => X"0000004800000000000000600000000000000073000000000000005700000000",
            INIT_5A => X"000000720000000000000069000000000000005d000000000000005200000000",
            INIT_5B => X"0000007b000000000000007e000000000000007d000000000000007700000000",
            INIT_5C => X"0000004c00000000000000300000000000000066000000000000007c00000000",
            INIT_5D => X"0000001b0000000000000029000000000000004e000000000000004b00000000",
            INIT_5E => X"0000000600000000000000100000000000000018000000000000000900000000",
            INIT_5F => X"00000019000000000000000f000000000000000a000000000000000800000000",
            INIT_60 => X"0000002b0000000000000023000000000000001f000000000000001500000000",
            INIT_61 => X"0000000c00000000000000190000000000000030000000000000003200000000",
            INIT_62 => X"000000110000000000000011000000000000000e000000000000000e00000000",
            INIT_63 => X"00000019000000000000001a0000000000000018000000000000001400000000",
            INIT_64 => X"0000004a000000000000000d0000000000000014000000000000001800000000",
            INIT_65 => X"000000120000000000000041000000000000003b000000000000004e00000000",
            INIT_66 => X"0000000300000000000000040000000000000005000000000000000300000000",
            INIT_67 => X"0000001a000000000000000d0000000000000009000000000000000500000000",
            INIT_68 => X"00000025000000000000002c0000000000000028000000000000002100000000",
            INIT_69 => X"00000025000000000000001e0000000000000017000000000000001e00000000",
            INIT_6A => X"0000001c000000000000001c0000000000000019000000000000001c00000000",
            INIT_6B => X"0000001300000000000000170000000000000018000000000000001b00000000",
            INIT_6C => X"0000001c00000000000000060000000000000009000000000000000f00000000",
            INIT_6D => X"00000008000000000000002f0000000000000053000000000000004700000000",
            INIT_6E => X"0000000400000000000000050000000000000005000000000000000200000000",
            INIT_6F => X"0000001c0000000000000015000000000000000b000000000000000600000000",
            INIT_70 => X"0000003b00000000000000300000000000000029000000000000002500000000",
            INIT_71 => X"00000059000000000000005c000000000000004f000000000000004900000000",
            INIT_72 => X"0000003b0000000000000038000000000000002f000000000000003800000000",
            INIT_73 => X"00000028000000000000002b0000000000000030000000000000003900000000",
            INIT_74 => X"000000150000000000000015000000000000001b000000000000002300000000",
            INIT_75 => X"0000000800000000000000100000000000000025000000000000002100000000",
            INIT_76 => X"0000000a000000000000000a0000000000000009000000000000000800000000",
            INIT_77 => X"0000001c000000000000001d0000000000000012000000000000000d00000000",
            INIT_78 => X"0000006500000000000000460000000000000031000000000000002c00000000",
            INIT_79 => X"0000006300000000000000760000000000000080000000000000008000000000",
            INIT_7A => X"000000550000000000000054000000000000004e000000000000004700000000",
            INIT_7B => X"0000004f00000000000000510000000000000053000000000000005700000000",
            INIT_7C => X"000000310000000000000031000000000000003c000000000000004700000000",
            INIT_7D => X"0000001300000000000000200000000000000038000000000000003a00000000",
            INIT_7E => X"0000001500000000000000180000000000000018000000000000001300000000",
            INIT_7F => X"0000001c0000000000000022000000000000001f000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "sampleifmap_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004d00000000000000510000000000000052000000000000005300000000",
            INIT_01 => X"0000005c000000000000005b0000000000000055000000000000005100000000",
            INIT_02 => X"0000005c0000000000000065000000000000005f000000000000005c00000000",
            INIT_03 => X"0000004c00000000000000500000000000000052000000000000005700000000",
            INIT_04 => X"0000003e000000000000003f0000000000000041000000000000004400000000",
            INIT_05 => X"0000002f00000000000000340000000000000038000000000000003c00000000",
            INIT_06 => X"0000002200000000000000230000000000000025000000000000002a00000000",
            INIT_07 => X"000000150000000000000019000000000000001d000000000000002400000000",
            INIT_08 => X"0000004d00000000000000530000000000000053000000000000005400000000",
            INIT_09 => X"0000005d000000000000005a0000000000000054000000000000005000000000",
            INIT_0A => X"00000061000000000000005f0000000000000058000000000000005a00000000",
            INIT_0B => X"0000004c000000000000004e0000000000000052000000000000005800000000",
            INIT_0C => X"0000004200000000000000400000000000000044000000000000004700000000",
            INIT_0D => X"0000002e00000000000000340000000000000036000000000000003d00000000",
            INIT_0E => X"0000002300000000000000240000000000000026000000000000002a00000000",
            INIT_0F => X"0000001f000000000000001d000000000000001e000000000000002400000000",
            INIT_10 => X"0000004b00000000000000500000000000000051000000000000005200000000",
            INIT_11 => X"0000004c00000000000000580000000000000054000000000000004b00000000",
            INIT_12 => X"0000006300000000000000570000000000000056000000000000005200000000",
            INIT_13 => X"0000004c000000000000004d0000000000000058000000000000006500000000",
            INIT_14 => X"0000004000000000000000400000000000000044000000000000004900000000",
            INIT_15 => X"0000002d00000000000000340000000000000037000000000000003a00000000",
            INIT_16 => X"0000002c00000000000000290000000000000028000000000000002b00000000",
            INIT_17 => X"0000003500000000000000310000000000000030000000000000003100000000",
            INIT_18 => X"0000004e00000000000000500000000000000051000000000000005300000000",
            INIT_19 => X"0000003200000000000000500000000000000057000000000000004a00000000",
            INIT_1A => X"0000005b00000000000000570000000000000061000000000000005500000000",
            INIT_1B => X"0000005000000000000000580000000000000066000000000000006800000000",
            INIT_1C => X"0000003f000000000000003f0000000000000040000000000000004900000000",
            INIT_1D => X"0000003a00000000000000390000000000000038000000000000003b00000000",
            INIT_1E => X"000000470000000000000044000000000000003f000000000000003d00000000",
            INIT_1F => X"0000004500000000000000450000000000000047000000000000004900000000",
            INIT_20 => X"0000004f000000000000004f000000000000004f000000000000004f00000000",
            INIT_21 => X"00000037000000000000004c0000000000000053000000000000004a00000000",
            INIT_22 => X"0000004b000000000000004b0000000000000054000000000000005300000000",
            INIT_23 => X"00000057000000000000005a0000000000000059000000000000004e00000000",
            INIT_24 => X"0000004600000000000000430000000000000042000000000000005300000000",
            INIT_25 => X"0000005700000000000000540000000000000050000000000000004e00000000",
            INIT_26 => X"0000005900000000000000590000000000000056000000000000005700000000",
            INIT_27 => X"00000049000000000000004f0000000000000054000000000000005800000000",
            INIT_28 => X"0000004d000000000000004b000000000000004a000000000000004c00000000",
            INIT_29 => X"0000004600000000000000460000000000000049000000000000004900000000",
            INIT_2A => X"0000004900000000000000470000000000000045000000000000004600000000",
            INIT_2B => X"00000051000000000000004e000000000000004e000000000000004b00000000",
            INIT_2C => X"0000006200000000000000600000000000000059000000000000005a00000000",
            INIT_2D => X"0000006800000000000000660000000000000068000000000000006400000000",
            INIT_2E => X"0000005e0000000000000061000000000000005f000000000000006300000000",
            INIT_2F => X"0000004200000000000000490000000000000050000000000000005700000000",
            INIT_30 => X"0000004900000000000000470000000000000048000000000000004a00000000",
            INIT_31 => X"00000033000000000000002b000000000000003e000000000000004a00000000",
            INIT_32 => X"0000004700000000000000440000000000000040000000000000004400000000",
            INIT_33 => X"0000005e0000000000000051000000000000004a000000000000004b00000000",
            INIT_34 => X"00000072000000000000006e0000000000000062000000000000006000000000",
            INIT_35 => X"0000006d00000000000000680000000000000064000000000000006600000000",
            INIT_36 => X"000000500000000000000055000000000000005b000000000000006300000000",
            INIT_37 => X"0000004300000000000000460000000000000049000000000000004c00000000",
            INIT_38 => X"0000004800000000000000470000000000000048000000000000004700000000",
            INIT_39 => X"00000029000000000000002a000000000000003a000000000000004700000000",
            INIT_3A => X"0000003f000000000000003a0000000000000036000000000000003900000000",
            INIT_3B => X"0000006000000000000000520000000000000047000000000000004100000000",
            INIT_3C => X"00000067000000000000005d000000000000005e000000000000006900000000",
            INIT_3D => X"00000061000000000000006c000000000000006a000000000000006700000000",
            INIT_3E => X"000000500000000000000054000000000000005b000000000000005d00000000",
            INIT_3F => X"0000004d000000000000004f0000000000000050000000000000005000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000052000000000000004b0000000000000049000000000000004900000000",
            INIT_41 => X"0000002e00000000000000570000000000000067000000000000005800000000",
            INIT_42 => X"0000005200000000000000450000000000000038000000000000003800000000",
            INIT_43 => X"00000057000000000000005a0000000000000057000000000000005100000000",
            INIT_44 => X"0000005b000000000000005e0000000000000063000000000000006200000000",
            INIT_45 => X"00000066000000000000006a0000000000000066000000000000006100000000",
            INIT_46 => X"0000005c00000000000000610000000000000063000000000000005e00000000",
            INIT_47 => X"0000005f000000000000005b0000000000000059000000000000005900000000",
            INIT_48 => X"0000007b000000000000006d000000000000005f000000000000005600000000",
            INIT_49 => X"0000003300000000000000680000000000000099000000000000008800000000",
            INIT_4A => X"000000610000000000000049000000000000003b000000000000003c00000000",
            INIT_4B => X"0000005a0000000000000066000000000000006c000000000000006500000000",
            INIT_4C => X"0000005d00000000000000610000000000000061000000000000005f00000000",
            INIT_4D => X"0000006e00000000000000690000000000000063000000000000005d00000000",
            INIT_4E => X"0000006c000000000000006c0000000000000069000000000000006700000000",
            INIT_4F => X"0000006e000000000000006e000000000000006e000000000000006d00000000",
            INIT_50 => X"0000009d0000000000000096000000000000008b000000000000007f00000000",
            INIT_51 => X"00000032000000000000005700000000000000a200000000000000a000000000",
            INIT_52 => X"0000005800000000000000350000000000000038000000000000004300000000",
            INIT_53 => X"0000005a000000000000006b0000000000000070000000000000006500000000",
            INIT_54 => X"00000060000000000000005e0000000000000060000000000000005e00000000",
            INIT_55 => X"000000650000000000000060000000000000005f000000000000006000000000",
            INIT_56 => X"0000007e000000000000007d0000000000000071000000000000006800000000",
            INIT_57 => X"0000007000000000000000740000000000000077000000000000007b00000000",
            INIT_58 => X"000000a2000000000000009f000000000000009d000000000000009800000000",
            INIT_59 => X"0000002c000000000000005a000000000000009f00000000000000a000000000",
            INIT_5A => X"00000056000000000000003a0000000000000045000000000000004800000000",
            INIT_5B => X"0000005c0000000000000061000000000000005a000000000000006700000000",
            INIT_5C => X"0000005e000000000000005f0000000000000060000000000000005a00000000",
            INIT_5D => X"0000005c00000000000000570000000000000062000000000000006300000000",
            INIT_5E => X"0000008300000000000000830000000000000070000000000000006100000000",
            INIT_5F => X"0000006c00000000000000740000000000000079000000000000007f00000000",
            INIT_60 => X"0000009d00000000000000a0000000000000009e000000000000009b00000000",
            INIT_61 => X"0000003000000000000000720000000000000094000000000000009800000000",
            INIT_62 => X"00000067000000000000005e0000000000000058000000000000004400000000",
            INIT_63 => X"0000005d00000000000000580000000000000060000000000000007300000000",
            INIT_64 => X"0000005e00000000000000620000000000000065000000000000005900000000",
            INIT_65 => X"0000005500000000000000540000000000000065000000000000006300000000",
            INIT_66 => X"00000084000000000000007d000000000000006e000000000000006900000000",
            INIT_67 => X"0000005f000000000000006b0000000000000076000000000000007f00000000",
            INIT_68 => X"0000009200000000000000950000000000000094000000000000009400000000",
            INIT_69 => X"000000500000000000000088000000000000008e000000000000009000000000",
            INIT_6A => X"00000068000000000000005e0000000000000048000000000000002f00000000",
            INIT_6B => X"0000005e000000000000005c0000000000000071000000000000007200000000",
            INIT_6C => X"0000005d00000000000000610000000000000067000000000000005d00000000",
            INIT_6D => X"0000005200000000000000550000000000000061000000000000006000000000",
            INIT_6E => X"00000079000000000000006f000000000000006b000000000000006b00000000",
            INIT_6F => X"0000004d00000000000000570000000000000064000000000000007000000000",
            INIT_70 => X"0000008c000000000000008a0000000000000087000000000000008600000000",
            INIT_71 => X"0000008900000000000000970000000000000093000000000000008e00000000",
            INIT_72 => X"0000003e00000000000000320000000000000049000000000000005d00000000",
            INIT_73 => X"00000062000000000000005a000000000000005e000000000000005900000000",
            INIT_74 => X"0000006100000000000000670000000000000069000000000000006600000000",
            INIT_75 => X"000000530000000000000056000000000000005e000000000000005e00000000",
            INIT_76 => X"00000066000000000000005c0000000000000065000000000000005f00000000",
            INIT_77 => X"0000004b000000000000004a0000000000000052000000000000005f00000000",
            INIT_78 => X"00000090000000000000008b0000000000000086000000000000008300000000",
            INIT_79 => X"00000098000000000000009a000000000000009f000000000000009800000000",
            INIT_7A => X"0000003900000000000000350000000000000076000000000000009e00000000",
            INIT_7B => X"00000066000000000000005f0000000000000064000000000000006700000000",
            INIT_7C => X"0000006a000000000000006f0000000000000074000000000000006e00000000",
            INIT_7D => X"000000550000000000000057000000000000005b000000000000006100000000",
            INIT_7E => X"0000005300000000000000550000000000000062000000000000005400000000",
            INIT_7F => X"0000005f000000000000005a0000000000000055000000000000005300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "sampleifmap_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a000000000000000980000000000000090000000000000008700000000",
            INIT_01 => X"00000073000000000000008900000000000000a100000000000000a400000000",
            INIT_02 => X"0000006e00000000000000800000000000000091000000000000009d00000000",
            INIT_03 => X"000000670000000000000068000000000000007a000000000000007b00000000",
            INIT_04 => X"00000068000000000000006c000000000000006d000000000000006900000000",
            INIT_05 => X"000000570000000000000058000000000000005a000000000000006100000000",
            INIT_06 => X"000000550000000000000057000000000000005c000000000000004f00000000",
            INIT_07 => X"0000005e00000000000000690000000000000069000000000000006500000000",
            INIT_08 => X"000000a4000000000000009f000000000000009a000000000000009400000000",
            INIT_09 => X"0000007f00000000000000b000000000000000b300000000000000aa00000000",
            INIT_0A => X"00000098000000000000009d00000000000000c500000000000000b000000000",
            INIT_0B => X"0000006700000000000000800000000000000091000000000000007100000000",
            INIT_0C => X"0000006600000000000000680000000000000065000000000000006700000000",
            INIT_0D => X"00000059000000000000005b000000000000005f000000000000006100000000",
            INIT_0E => X"0000005b000000000000005b0000000000000056000000000000004f00000000",
            INIT_0F => X"0000004600000000000000560000000000000068000000000000006d00000000",
            INIT_10 => X"000000c500000000000000b200000000000000a4000000000000009b00000000",
            INIT_11 => X"000000c400000000000000f800000000000000ee00000000000000dd00000000",
            INIT_12 => X"000000b800000000000000b000000000000000c8000000000000009c00000000",
            INIT_13 => X"0000006a0000000000000089000000000000008e000000000000006c00000000",
            INIT_14 => X"0000006500000000000000640000000000000063000000000000006400000000",
            INIT_15 => X"00000059000000000000005f0000000000000063000000000000006500000000",
            INIT_16 => X"00000053000000000000005c0000000000000051000000000000005000000000",
            INIT_17 => X"0000004700000000000000490000000000000052000000000000005800000000",
            INIT_18 => X"000000f900000000000000eb00000000000000d600000000000000bf00000000",
            INIT_19 => X"000000f400000000000000fb00000000000000f600000000000000fd00000000",
            INIT_1A => X"000000c300000000000000ac000000000000009e00000000000000a000000000",
            INIT_1B => X"0000006e000000000000008b0000000000000072000000000000007100000000",
            INIT_1C => X"0000006300000000000000610000000000000062000000000000006200000000",
            INIT_1D => X"0000005c00000000000000660000000000000068000000000000006700000000",
            INIT_1E => X"000000490000000000000055000000000000004e000000000000005300000000",
            INIT_1F => X"00000048000000000000004a0000000000000050000000000000004b00000000",
            INIT_20 => X"000000fe00000000000000fd00000000000000fc00000000000000f500000000",
            INIT_21 => X"000000c900000000000000ba00000000000000bb00000000000000f300000000",
            INIT_22 => X"0000009c00000000000000970000000000000080000000000000009100000000",
            INIT_23 => X"000000720000000000000080000000000000006a000000000000007400000000",
            INIT_24 => X"0000006700000000000000650000000000000067000000000000006800000000",
            INIT_25 => X"0000005c0000000000000069000000000000006e000000000000006c00000000",
            INIT_26 => X"000000550000000000000054000000000000004c000000000000005200000000",
            INIT_27 => X"00000049000000000000004d0000000000000053000000000000004e00000000",
            INIT_28 => X"0000010000000000000000fc00000000000000fc00000000000000fb00000000",
            INIT_29 => X"00000072000000000000006b000000000000007e00000000000000e900000000",
            INIT_2A => X"0000006e00000000000000780000000000000073000000000000006900000000",
            INIT_2B => X"0000006700000000000000680000000000000063000000000000006300000000",
            INIT_2C => X"0000006b000000000000006b000000000000006e000000000000006d00000000",
            INIT_2D => X"000000560000000000000060000000000000006e000000000000007000000000",
            INIT_2E => X"00000068000000000000005a000000000000004c000000000000004e00000000",
            INIT_2F => X"0000004f00000000000000520000000000000052000000000000005b00000000",
            INIT_30 => X"000000eb00000000000000f600000000000000f800000000000000f800000000",
            INIT_31 => X"000000760000000000000072000000000000007c00000000000000c800000000",
            INIT_32 => X"0000004f00000000000000530000000000000057000000000000005d00000000",
            INIT_33 => X"00000044000000000000004b0000000000000056000000000000005000000000",
            INIT_34 => X"0000006100000000000000620000000000000064000000000000005f00000000",
            INIT_35 => X"0000006100000000000000610000000000000061000000000000006200000000",
            INIT_36 => X"0000006f000000000000005b0000000000000057000000000000005b00000000",
            INIT_37 => X"0000005200000000000000520000000000000055000000000000006e00000000",
            INIT_38 => X"0000009600000000000000b500000000000000d600000000000000eb00000000",
            INIT_39 => X"0000008400000000000000850000000000000088000000000000008a00000000",
            INIT_3A => X"0000003c0000000000000039000000000000003d000000000000006400000000",
            INIT_3B => X"0000003a00000000000000600000000000000059000000000000004300000000",
            INIT_3C => X"0000005000000000000000470000000000000045000000000000003300000000",
            INIT_3D => X"0000006500000000000000680000000000000065000000000000005e00000000",
            INIT_3E => X"0000006d000000000000005e0000000000000057000000000000005d00000000",
            INIT_3F => X"0000005100000000000000510000000000000062000000000000007700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009900000000",
            INIT_41 => X"00000067000000000000006f000000000000007a000000000000007c00000000",
            INIT_42 => X"000000340000000000000039000000000000005a000000000000006a00000000",
            INIT_43 => X"00000053000000000000006a0000000000000066000000000000004500000000",
            INIT_44 => X"00000055000000000000004d0000000000000047000000000000004000000000",
            INIT_45 => X"0000006d00000000000000660000000000000067000000000000006400000000",
            INIT_46 => X"00000063000000000000005d0000000000000057000000000000006a00000000",
            INIT_47 => X"00000050000000000000005c0000000000000073000000000000007100000000",
            INIT_48 => X"0000006d0000000000000072000000000000006f000000000000006d00000000",
            INIT_49 => X"0000006d00000000000000660000000000000061000000000000006500000000",
            INIT_4A => X"0000005500000000000000670000000000000078000000000000007500000000",
            INIT_4B => X"00000059000000000000005f0000000000000065000000000000005d00000000",
            INIT_4C => X"0000005a0000000000000052000000000000004b000000000000004a00000000",
            INIT_4D => X"0000006600000000000000690000000000000077000000000000007200000000",
            INIT_4E => X"00000062000000000000005e000000000000006b000000000000006f00000000",
            INIT_4F => X"0000004f000000000000006b0000000000000075000000000000006500000000",
            INIT_50 => X"0000005b000000000000005d0000000000000062000000000000006900000000",
            INIT_51 => X"00000071000000000000006f000000000000006a000000000000006300000000",
            INIT_52 => X"0000005f00000000000000610000000000000068000000000000007000000000",
            INIT_53 => X"0000005c0000000000000054000000000000004c000000000000005000000000",
            INIT_54 => X"00000059000000000000004f0000000000000048000000000000005100000000",
            INIT_55 => X"0000005e0000000000000069000000000000007b000000000000007500000000",
            INIT_56 => X"0000006500000000000000670000000000000067000000000000006000000000",
            INIT_57 => X"0000005a000000000000006f0000000000000069000000000000006000000000",
            INIT_58 => X"00000065000000000000005e0000000000000057000000000000005700000000",
            INIT_59 => X"00000064000000000000006b000000000000006e000000000000006c00000000",
            INIT_5A => X"0000006800000000000000560000000000000051000000000000005b00000000",
            INIT_5B => X"0000005c000000000000004c0000000000000049000000000000005d00000000",
            INIT_5C => X"0000004f000000000000004f000000000000004d000000000000005800000000",
            INIT_5D => X"00000056000000000000005d0000000000000064000000000000005b00000000",
            INIT_5E => X"000000600000000000000061000000000000005c000000000000005700000000",
            INIT_5F => X"0000006500000000000000660000000000000060000000000000006000000000",
            INIT_60 => X"0000006900000000000000670000000000000060000000000000005a00000000",
            INIT_61 => X"000000500000000000000056000000000000005f000000000000006500000000",
            INIT_62 => X"0000006a00000000000000600000000000000055000000000000005100000000",
            INIT_63 => X"0000005d00000000000000600000000000000055000000000000006200000000",
            INIT_64 => X"0000004c000000000000004f0000000000000051000000000000005800000000",
            INIT_65 => X"0000005b0000000000000054000000000000004c000000000000004700000000",
            INIT_66 => X"0000005a00000000000000530000000000000056000000000000005c00000000",
            INIT_67 => X"00000060000000000000005b0000000000000060000000000000006200000000",
            INIT_68 => X"00000056000000000000005f0000000000000063000000000000006400000000",
            INIT_69 => X"0000004f000000000000004f000000000000004f000000000000005000000000",
            INIT_6A => X"0000006c00000000000000620000000000000053000000000000005200000000",
            INIT_6B => X"0000005900000000000000610000000000000060000000000000006300000000",
            INIT_6C => X"00000051000000000000004f0000000000000054000000000000005c00000000",
            INIT_6D => X"000000590000000000000052000000000000004a000000000000004c00000000",
            INIT_6E => X"0000005600000000000000520000000000000055000000000000005a00000000",
            INIT_6F => X"000000530000000000000053000000000000005c000000000000005d00000000",
            INIT_70 => X"000000470000000000000049000000000000004e000000000000005700000000",
            INIT_71 => X"0000005300000000000000590000000000000057000000000000004d00000000",
            INIT_72 => X"0000006a0000000000000061000000000000004f000000000000005100000000",
            INIT_73 => X"0000005c00000000000000590000000000000067000000000000006400000000",
            INIT_74 => X"0000005900000000000000580000000000000057000000000000006000000000",
            INIT_75 => X"000000530000000000000054000000000000004f000000000000005200000000",
            INIT_76 => X"000000530000000000000056000000000000005a000000000000005600000000",
            INIT_77 => X"00000049000000000000004f0000000000000056000000000000005600000000",
            INIT_78 => X"000000490000000000000046000000000000003f000000000000003e00000000",
            INIT_79 => X"0000005100000000000000530000000000000056000000000000005400000000",
            INIT_7A => X"0000006b000000000000005e000000000000004a000000000000004e00000000",
            INIT_7B => X"00000058000000000000005b0000000000000068000000000000005f00000000",
            INIT_7C => X"0000005900000000000000580000000000000058000000000000005b00000000",
            INIT_7D => X"0000005300000000000000550000000000000050000000000000005500000000",
            INIT_7E => X"0000005000000000000000560000000000000059000000000000005400000000",
            INIT_7F => X"00000048000000000000004c000000000000004d000000000000004c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "sampleifmap_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000005d000000000000005e000000000000005e00000000",
            INIT_01 => X"000000600000000000000060000000000000005a000000000000005a00000000",
            INIT_02 => X"00000065000000000000006e0000000000000066000000000000006100000000",
            INIT_03 => X"0000005200000000000000550000000000000058000000000000005e00000000",
            INIT_04 => X"000000480000000000000049000000000000004b000000000000004e00000000",
            INIT_05 => X"00000038000000000000003d0000000000000041000000000000004500000000",
            INIT_06 => X"000000270000000000000029000000000000002e000000000000003300000000",
            INIT_07 => X"00000019000000000000001d0000000000000022000000000000002800000000",
            INIT_08 => X"00000059000000000000005f000000000000005f000000000000006000000000",
            INIT_09 => X"00000062000000000000005f0000000000000059000000000000005900000000",
            INIT_0A => X"0000006b000000000000006a0000000000000060000000000000006100000000",
            INIT_0B => X"0000005200000000000000550000000000000059000000000000006000000000",
            INIT_0C => X"000000490000000000000047000000000000004b000000000000004f00000000",
            INIT_0D => X"00000035000000000000003b000000000000003d000000000000004400000000",
            INIT_0E => X"000000250000000000000027000000000000002c000000000000003100000000",
            INIT_0F => X"0000001f000000000000001f0000000000000020000000000000002600000000",
            INIT_10 => X"00000057000000000000005c000000000000005c000000000000005e00000000",
            INIT_11 => X"00000051000000000000005d000000000000005a000000000000005400000000",
            INIT_12 => X"0000006e00000000000000630000000000000060000000000000005900000000",
            INIT_13 => X"0000005400000000000000560000000000000062000000000000007000000000",
            INIT_14 => X"0000004600000000000000440000000000000049000000000000004f00000000",
            INIT_15 => X"000000300000000000000036000000000000003a000000000000003f00000000",
            INIT_16 => X"0000002b0000000000000029000000000000002b000000000000002e00000000",
            INIT_17 => X"000000310000000000000030000000000000002e000000000000002f00000000",
            INIT_18 => X"0000005a000000000000005c000000000000005d000000000000005f00000000",
            INIT_19 => X"000000390000000000000056000000000000005d000000000000005300000000",
            INIT_1A => X"000000680000000000000063000000000000006b000000000000005d00000000",
            INIT_1B => X"0000005a00000000000000650000000000000072000000000000007400000000",
            INIT_1C => X"0000004200000000000000420000000000000043000000000000004e00000000",
            INIT_1D => X"0000003900000000000000380000000000000038000000000000003e00000000",
            INIT_1E => X"000000420000000000000041000000000000003e000000000000003c00000000",
            INIT_1F => X"0000003d000000000000003f0000000000000041000000000000004300000000",
            INIT_20 => X"0000005b000000000000005b000000000000005b000000000000005c00000000",
            INIT_21 => X"0000003e00000000000000520000000000000059000000000000005300000000",
            INIT_22 => X"000000580000000000000058000000000000005f000000000000005c00000000",
            INIT_23 => X"0000006400000000000000690000000000000068000000000000005c00000000",
            INIT_24 => X"0000004800000000000000450000000000000046000000000000005b00000000",
            INIT_25 => X"000000530000000000000050000000000000004d000000000000005000000000",
            INIT_26 => X"0000005000000000000000510000000000000051000000000000005300000000",
            INIT_27 => X"0000003f0000000000000046000000000000004b000000000000004f00000000",
            INIT_28 => X"0000005900000000000000570000000000000056000000000000005800000000",
            INIT_29 => X"0000004d000000000000004c000000000000004f000000000000005200000000",
            INIT_2A => X"0000005700000000000000550000000000000052000000000000005000000000",
            INIT_2B => X"0000005f000000000000005e000000000000005e000000000000005a00000000",
            INIT_2C => X"000000630000000000000062000000000000005e000000000000006300000000",
            INIT_2D => X"0000006200000000000000600000000000000064000000000000006400000000",
            INIT_2E => X"0000005300000000000000580000000000000058000000000000005d00000000",
            INIT_2F => X"00000037000000000000003e0000000000000045000000000000004c00000000",
            INIT_30 => X"0000005400000000000000520000000000000054000000000000005500000000",
            INIT_31 => X"00000037000000000000002a000000000000003d000000000000005100000000",
            INIT_32 => X"0000005900000000000000580000000000000057000000000000005300000000",
            INIT_33 => X"00000065000000000000005d0000000000000057000000000000005b00000000",
            INIT_34 => X"0000007300000000000000700000000000000064000000000000006200000000",
            INIT_35 => X"0000006700000000000000670000000000000067000000000000006900000000",
            INIT_36 => X"0000004a000000000000004e0000000000000050000000000000005b00000000",
            INIT_37 => X"000000360000000000000039000000000000003f000000000000004400000000",
            INIT_38 => X"0000005400000000000000520000000000000053000000000000005200000000",
            INIT_39 => X"0000002c00000000000000260000000000000037000000000000004c00000000",
            INIT_3A => X"0000005100000000000000520000000000000055000000000000004c00000000",
            INIT_3B => X"00000063000000000000005b0000000000000053000000000000005000000000",
            INIT_3C => X"0000006c00000000000000610000000000000060000000000000006700000000",
            INIT_3D => X"0000005e00000000000000710000000000000072000000000000006d00000000",
            INIT_3E => X"0000004b000000000000004d000000000000004d000000000000005200000000",
            INIT_3F => X"0000003b00000000000000400000000000000044000000000000004700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005b00000000000000540000000000000052000000000000005100000000",
            INIT_41 => X"0000003100000000000000550000000000000068000000000000005e00000000",
            INIT_42 => X"00000063000000000000005b0000000000000054000000000000004900000000",
            INIT_43 => X"0000005e00000000000000650000000000000064000000000000006100000000",
            INIT_44 => X"0000006200000000000000650000000000000068000000000000006500000000",
            INIT_45 => X"000000670000000000000072000000000000006f000000000000006a00000000",
            INIT_46 => X"0000004e00000000000000520000000000000055000000000000005700000000",
            INIT_47 => X"0000004800000000000000470000000000000046000000000000004a00000000",
            INIT_48 => X"0000008000000000000000730000000000000065000000000000005c00000000",
            INIT_49 => X"000000360000000000000068000000000000009d000000000000008e00000000",
            INIT_4A => X"00000071000000000000005d0000000000000054000000000000004b00000000",
            INIT_4B => X"000000650000000000000075000000000000007c000000000000007500000000",
            INIT_4C => X"00000067000000000000006b000000000000006a000000000000006700000000",
            INIT_4D => X"000000760000000000000074000000000000006e000000000000006800000000",
            INIT_4E => X"000000540000000000000055000000000000005a000000000000006400000000",
            INIT_4F => X"0000005200000000000000550000000000000055000000000000005500000000",
            INIT_50 => X"000000a00000000000000099000000000000008e000000000000008200000000",
            INIT_51 => X"00000035000000000000005900000000000000aa00000000000000a600000000",
            INIT_52 => X"000000680000000000000046000000000000004d000000000000005000000000",
            INIT_53 => X"0000006b000000000000007f0000000000000082000000000000007700000000",
            INIT_54 => X"0000006a0000000000000069000000000000006c000000000000006a00000000",
            INIT_55 => X"00000072000000000000006e0000000000000069000000000000006a00000000",
            INIT_56 => X"0000006000000000000000620000000000000062000000000000006900000000",
            INIT_57 => X"000000550000000000000059000000000000005b000000000000005e00000000",
            INIT_58 => X"000000a400000000000000a2000000000000009f000000000000009a00000000",
            INIT_59 => X"0000002e000000000000005d00000000000000a900000000000000a700000000",
            INIT_5A => X"00000067000000000000004a0000000000000056000000000000005100000000",
            INIT_5B => X"00000072000000000000007a0000000000000070000000000000007b00000000",
            INIT_5C => X"00000067000000000000006a000000000000006d000000000000006a00000000",
            INIT_5D => X"0000006e00000000000000670000000000000069000000000000006b00000000",
            INIT_5E => X"0000006300000000000000650000000000000061000000000000006600000000",
            INIT_5F => X"00000055000000000000005a000000000000005e000000000000006000000000",
            INIT_60 => X"0000009e00000000000000a1000000000000009f000000000000009d00000000",
            INIT_61 => X"000000300000000000000075000000000000009f000000000000009e00000000",
            INIT_62 => X"00000078000000000000006c0000000000000065000000000000004900000000",
            INIT_63 => X"0000007500000000000000740000000000000078000000000000008700000000",
            INIT_64 => X"00000066000000000000006c0000000000000073000000000000006b00000000",
            INIT_65 => X"000000690000000000000064000000000000006a000000000000006900000000",
            INIT_66 => X"0000006500000000000000600000000000000060000000000000007000000000",
            INIT_67 => X"0000004c0000000000000055000000000000005d000000000000006200000000",
            INIT_68 => X"0000009300000000000000970000000000000098000000000000009900000000",
            INIT_69 => X"0000004c00000000000000870000000000000093000000000000009300000000",
            INIT_6A => X"0000007500000000000000670000000000000049000000000000002c00000000",
            INIT_6B => X"0000007100000000000000730000000000000085000000000000008300000000",
            INIT_6C => X"0000006b00000000000000710000000000000077000000000000006c00000000",
            INIT_6D => X"000000640000000000000065000000000000006a000000000000006a00000000",
            INIT_6E => X"00000062000000000000005d0000000000000069000000000000007500000000",
            INIT_6F => X"00000040000000000000004a0000000000000055000000000000005d00000000",
            INIT_70 => X"0000008e000000000000008e000000000000008e000000000000008f00000000",
            INIT_71 => X"0000008300000000000000950000000000000094000000000000008f00000000",
            INIT_72 => X"0000004600000000000000350000000000000041000000000000005400000000",
            INIT_73 => X"0000006d0000000000000068000000000000006b000000000000006300000000",
            INIT_74 => X"00000075000000000000007d000000000000007c000000000000007200000000",
            INIT_75 => X"000000620000000000000065000000000000006c000000000000006e00000000",
            INIT_76 => X"0000005a0000000000000058000000000000006f000000000000006c00000000",
            INIT_77 => X"0000003f00000000000000410000000000000048000000000000005500000000",
            INIT_78 => X"00000091000000000000008e000000000000008d000000000000008c00000000",
            INIT_79 => X"00000093000000000000009900000000000000a0000000000000009900000000",
            INIT_7A => X"0000003a0000000000000034000000000000006f000000000000009700000000",
            INIT_7B => X"0000006e00000000000000650000000000000068000000000000006a00000000",
            INIT_7C => X"0000008000000000000000870000000000000089000000000000007b00000000",
            INIT_7D => X"000000650000000000000068000000000000006c000000000000007300000000",
            INIT_7E => X"0000004e0000000000000059000000000000006f000000000000006300000000",
            INIT_7F => X"0000004d000000000000004a0000000000000048000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "sampleifmap_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000000000009b0000000000000095000000000000008f00000000",
            INIT_01 => X"00000072000000000000008800000000000000a000000000000000a400000000",
            INIT_02 => X"00000068000000000000007a000000000000008f000000000000009b00000000",
            INIT_03 => X"0000006c00000000000000660000000000000077000000000000007600000000",
            INIT_04 => X"0000008000000000000000850000000000000084000000000000007800000000",
            INIT_05 => X"0000006a000000000000006b000000000000006d000000000000007500000000",
            INIT_06 => X"000000560000000000000062000000000000006c000000000000006100000000",
            INIT_07 => X"00000044000000000000004f0000000000000054000000000000005a00000000",
            INIT_08 => X"000000a1000000000000009f000000000000009d000000000000009a00000000",
            INIT_09 => X"0000008100000000000000b000000000000000b100000000000000a700000000",
            INIT_0A => X"0000008e000000000000009700000000000000c700000000000000b300000000",
            INIT_0B => X"0000006c000000000000007b0000000000000089000000000000006800000000",
            INIT_0C => X"000000800000000000000083000000000000007e000000000000007900000000",
            INIT_0D => X"0000006e00000000000000700000000000000073000000000000007700000000",
            INIT_0E => X"0000005e000000000000006a0000000000000069000000000000006300000000",
            INIT_0F => X"000000270000000000000034000000000000004a000000000000005c00000000",
            INIT_10 => X"000000c100000000000000b000000000000000a4000000000000009d00000000",
            INIT_11 => X"000000c700000000000000f700000000000000ec00000000000000da00000000",
            INIT_12 => X"000000b100000000000000ad00000000000000ce00000000000000a300000000",
            INIT_13 => X"0000007100000000000000860000000000000088000000000000006500000000",
            INIT_14 => X"000000810000000000000082000000000000007e000000000000007700000000",
            INIT_15 => X"000000710000000000000076000000000000007a000000000000007d00000000",
            INIT_16 => X"00000050000000000000006a0000000000000067000000000000006800000000",
            INIT_17 => X"000000270000000000000025000000000000002c000000000000003e00000000",
            INIT_18 => X"000000f600000000000000e800000000000000d400000000000000c000000000",
            INIT_19 => X"000000f700000000000000fa00000000000000f200000000000000fa00000000",
            INIT_1A => X"000000c100000000000000ae00000000000000aa00000000000000a900000000",
            INIT_1B => X"00000078000000000000008b0000000000000070000000000000006e00000000",
            INIT_1C => X"000000800000000000000080000000000000007e000000000000007600000000",
            INIT_1D => X"00000074000000000000007e000000000000007f000000000000008000000000",
            INIT_1E => X"0000003e00000000000000600000000000000066000000000000006c00000000",
            INIT_1F => X"0000002b00000000000000270000000000000025000000000000002a00000000",
            INIT_20 => X"000000fb00000000000000fa00000000000000fb00000000000000f500000000",
            INIT_21 => X"000000d200000000000000be00000000000000ba00000000000000f100000000",
            INIT_22 => X"000000a0000000000000009c000000000000009200000000000000a100000000",
            INIT_23 => X"0000007a00000000000000870000000000000073000000000000007d00000000",
            INIT_24 => X"000000800000000000000081000000000000007f000000000000007800000000",
            INIT_25 => X"00000074000000000000007d000000000000007f000000000000007f00000000",
            INIT_26 => X"0000004200000000000000570000000000000062000000000000006a00000000",
            INIT_27 => X"000000290000000000000029000000000000002a000000000000002d00000000",
            INIT_28 => X"000000fe00000000000000fb00000000000000fb00000000000000fb00000000",
            INIT_29 => X"000000820000000000000074000000000000008300000000000000ea00000000",
            INIT_2A => X"0000007c0000000000000082000000000000008a000000000000007f00000000",
            INIT_2B => X"0000006b00000000000000720000000000000077000000000000007a00000000",
            INIT_2C => X"0000007f00000000000000820000000000000080000000000000007600000000",
            INIT_2D => X"0000006c000000000000006f0000000000000077000000000000007d00000000",
            INIT_2E => X"000000500000000000000052000000000000005a000000000000006300000000",
            INIT_2F => X"00000029000000000000002c000000000000002f000000000000003d00000000",
            INIT_30 => X"000000ef00000000000000f900000000000000fc00000000000000fc00000000",
            INIT_31 => X"00000083000000000000007b000000000000008000000000000000cb00000000",
            INIT_32 => X"000000670000000000000066000000000000006c000000000000006f00000000",
            INIT_33 => X"0000004400000000000000510000000000000069000000000000006a00000000",
            INIT_34 => X"0000007400000000000000780000000000000075000000000000006600000000",
            INIT_35 => X"000000730000000000000070000000000000006b000000000000006e00000000",
            INIT_36 => X"00000054000000000000004b0000000000000059000000000000006800000000",
            INIT_37 => X"0000002d000000000000002d0000000000000034000000000000005100000000",
            INIT_38 => X"000000a000000000000000bf00000000000000df00000000000000f500000000",
            INIT_39 => X"0000008a00000000000000890000000000000089000000000000009000000000",
            INIT_3A => X"000000570000000000000051000000000000004b000000000000006d00000000",
            INIT_3B => X"0000003a00000000000000630000000000000066000000000000005a00000000",
            INIT_3C => X"00000065000000000000005f0000000000000056000000000000003a00000000",
            INIT_3D => X"00000074000000000000007a0000000000000074000000000000006d00000000",
            INIT_3E => X"000000500000000000000046000000000000004d000000000000006100000000",
            INIT_3F => X"0000002f000000000000002f0000000000000042000000000000005900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000840000000000000086000000000000008d00000000000000a500000000",
            INIT_41 => X"000000690000000000000070000000000000007b000000000000008200000000",
            INIT_42 => X"00000047000000000000004a000000000000005e000000000000006b00000000",
            INIT_43 => X"00000056000000000000006f000000000000006e000000000000005300000000",
            INIT_44 => X"0000006c0000000000000066000000000000005a000000000000004800000000",
            INIT_45 => X"0000007c000000000000007b000000000000007b000000000000007600000000",
            INIT_46 => X"0000004400000000000000420000000000000049000000000000006c00000000",
            INIT_47 => X"00000030000000000000003d0000000000000054000000000000005200000000",
            INIT_48 => X"00000075000000000000007a0000000000000078000000000000007500000000",
            INIT_49 => X"0000006a00000000000000650000000000000061000000000000006a00000000",
            INIT_4A => X"00000057000000000000006a0000000000000073000000000000007000000000",
            INIT_4B => X"0000006100000000000000680000000000000068000000000000005c00000000",
            INIT_4C => X"00000072000000000000006c000000000000005f000000000000005400000000",
            INIT_4D => X"0000007a0000000000000082000000000000008e000000000000008600000000",
            INIT_4E => X"0000004000000000000000450000000000000064000000000000007700000000",
            INIT_4F => X"00000032000000000000004f0000000000000057000000000000004500000000",
            INIT_50 => X"0000005e00000000000000600000000000000066000000000000006c00000000",
            INIT_51 => X"0000006b000000000000006e000000000000006b000000000000006500000000",
            INIT_52 => X"000000510000000000000056000000000000005d000000000000006700000000",
            INIT_53 => X"00000068000000000000005d0000000000000048000000000000004200000000",
            INIT_54 => X"00000071000000000000006b000000000000005f000000000000005e00000000",
            INIT_55 => X"0000007a00000000000000850000000000000094000000000000008900000000",
            INIT_56 => X"000000420000000000000051000000000000006b000000000000007200000000",
            INIT_57 => X"0000003f0000000000000055000000000000004b000000000000004000000000",
            INIT_58 => X"00000063000000000000005d0000000000000057000000000000005800000000",
            INIT_59 => X"000000570000000000000065000000000000006c000000000000006b00000000",
            INIT_5A => X"000000530000000000000041000000000000003c000000000000004900000000",
            INIT_5B => X"0000005e000000000000004e000000000000003f000000000000004a00000000",
            INIT_5C => X"0000005d000000000000005f0000000000000057000000000000005900000000",
            INIT_5D => X"00000072000000000000007a000000000000007b000000000000006900000000",
            INIT_5E => X"0000003b000000000000004e0000000000000068000000000000006d00000000",
            INIT_5F => X"0000004b000000000000004a000000000000003f000000000000003c00000000",
            INIT_60 => X"0000005f0000000000000061000000000000005f000000000000005d00000000",
            INIT_61 => X"0000003800000000000000450000000000000054000000000000005b00000000",
            INIT_62 => X"0000005500000000000000420000000000000031000000000000003200000000",
            INIT_63 => X"0000004800000000000000550000000000000049000000000000005300000000",
            INIT_64 => X"000000440000000000000043000000000000003e000000000000003e00000000",
            INIT_65 => X"0000006800000000000000640000000000000058000000000000004500000000",
            INIT_66 => X"000000330000000000000040000000000000005a000000000000006500000000",
            INIT_67 => X"00000045000000000000003a0000000000000036000000000000003500000000",
            INIT_68 => X"000000440000000000000051000000000000005b000000000000006000000000",
            INIT_69 => X"0000003000000000000000340000000000000037000000000000003b00000000",
            INIT_6A => X"000000520000000000000040000000000000002e000000000000002f00000000",
            INIT_6B => X"00000039000000000000004d000000000000004f000000000000005200000000",
            INIT_6C => X"0000003a00000000000000340000000000000032000000000000003500000000",
            INIT_6D => X"0000004a0000000000000047000000000000003f000000000000003a00000000",
            INIT_6E => X"0000002e00000000000000340000000000000041000000000000004800000000",
            INIT_6F => X"0000003600000000000000300000000000000031000000000000003000000000",
            INIT_70 => X"0000002b0000000000000031000000000000003c000000000000004900000000",
            INIT_71 => X"0000003000000000000000340000000000000030000000000000002c00000000",
            INIT_72 => X"00000049000000000000003a000000000000002c000000000000003000000000",
            INIT_73 => X"00000035000000000000003e000000000000004f000000000000004b00000000",
            INIT_74 => X"000000390000000000000034000000000000002e000000000000003200000000",
            INIT_75 => X"0000002f0000000000000033000000000000002f000000000000003400000000",
            INIT_76 => X"0000002a000000000000002e0000000000000031000000000000002f00000000",
            INIT_77 => X"0000002a000000000000002b000000000000002d000000000000002b00000000",
            INIT_78 => X"0000002500000000000000270000000000000025000000000000002900000000",
            INIT_79 => X"0000002d00000000000000290000000000000029000000000000002a00000000",
            INIT_7A => X"000000470000000000000036000000000000002b000000000000002f00000000",
            INIT_7B => X"0000002e000000000000003b000000000000004c000000000000004300000000",
            INIT_7C => X"00000030000000000000002d000000000000002a000000000000002b00000000",
            INIT_7D => X"0000002d0000000000000031000000000000002d000000000000002f00000000",
            INIT_7E => X"00000027000000000000002a000000000000002d000000000000002b00000000",
            INIT_7F => X"0000002600000000000000280000000000000028000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "sampleifmap_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004f00000000000000530000000000000054000000000000005500000000",
            INIT_01 => X"0000005f000000000000005d0000000000000052000000000000005000000000",
            INIT_02 => X"00000048000000000000004f0000000000000055000000000000005a00000000",
            INIT_03 => X"0000004f0000000000000054000000000000004e000000000000004b00000000",
            INIT_04 => X"0000003d000000000000003c000000000000003e000000000000004400000000",
            INIT_05 => X"000000330000000000000038000000000000003b000000000000003c00000000",
            INIT_06 => X"0000002300000000000000250000000000000029000000000000002e00000000",
            INIT_07 => X"000000150000000000000019000000000000001e000000000000002400000000",
            INIT_08 => X"0000004f00000000000000550000000000000055000000000000005600000000",
            INIT_09 => X"0000005d000000000000005a0000000000000050000000000000004e00000000",
            INIT_0A => X"0000004700000000000000460000000000000049000000000000005400000000",
            INIT_0B => X"0000004800000000000000470000000000000045000000000000004400000000",
            INIT_0C => X"0000003e000000000000003e0000000000000043000000000000004600000000",
            INIT_0D => X"0000002e00000000000000340000000000000035000000000000003800000000",
            INIT_0E => X"0000002000000000000000220000000000000025000000000000002900000000",
            INIT_0F => X"0000001b000000000000001a000000000000001b000000000000002100000000",
            INIT_10 => X"0000004e00000000000000520000000000000053000000000000005400000000",
            INIT_11 => X"0000004800000000000000560000000000000050000000000000004900000000",
            INIT_12 => X"0000004300000000000000380000000000000041000000000000004600000000",
            INIT_13 => X"0000003c0000000000000036000000000000003f000000000000004800000000",
            INIT_14 => X"0000003a000000000000003d0000000000000041000000000000004200000000",
            INIT_15 => X"00000026000000000000002d000000000000002f000000000000003000000000",
            INIT_16 => X"0000002500000000000000220000000000000021000000000000002400000000",
            INIT_17 => X"0000002c000000000000002a0000000000000029000000000000002a00000000",
            INIT_18 => X"0000005000000000000000520000000000000053000000000000005500000000",
            INIT_19 => X"0000002b000000000000004d0000000000000052000000000000004800000000",
            INIT_1A => X"0000003400000000000000320000000000000045000000000000004300000000",
            INIT_1B => X"0000002f0000000000000032000000000000003f000000000000004100000000",
            INIT_1C => X"0000003600000000000000390000000000000034000000000000003200000000",
            INIT_1D => X"0000002c000000000000002b000000000000002b000000000000002d00000000",
            INIT_1E => X"0000003b00000000000000380000000000000032000000000000002f00000000",
            INIT_1F => X"000000370000000000000038000000000000003b000000000000003c00000000",
            INIT_20 => X"0000005100000000000000510000000000000051000000000000005200000000",
            INIT_21 => X"0000002c0000000000000046000000000000004c000000000000004800000000",
            INIT_22 => X"0000001d00000000000000220000000000000033000000000000003d00000000",
            INIT_23 => X"0000002300000000000000260000000000000027000000000000001f00000000",
            INIT_24 => X"0000003b0000000000000039000000000000002b000000000000002900000000",
            INIT_25 => X"000000440000000000000041000000000000003d000000000000003d00000000",
            INIT_26 => X"0000004800000000000000470000000000000042000000000000004400000000",
            INIT_27 => X"00000038000000000000003e0000000000000043000000000000004700000000",
            INIT_28 => X"0000004f000000000000004c000000000000004c000000000000004d00000000",
            INIT_29 => X"00000038000000000000003e0000000000000042000000000000004700000000",
            INIT_2A => X"00000017000000000000001a0000000000000021000000000000002c00000000",
            INIT_2B => X"0000000e000000000000000f0000000000000014000000000000001600000000",
            INIT_2C => X"00000054000000000000004f0000000000000035000000000000001f00000000",
            INIT_2D => X"00000050000000000000004e0000000000000052000000000000005300000000",
            INIT_2E => X"0000004b000000000000004d0000000000000048000000000000004c00000000",
            INIT_2F => X"0000002e0000000000000035000000000000003c000000000000004400000000",
            INIT_30 => X"0000004800000000000000460000000000000047000000000000004900000000",
            INIT_31 => X"0000002000000000000000200000000000000037000000000000004700000000",
            INIT_32 => X"0000001300000000000000140000000000000018000000000000002600000000",
            INIT_33 => X"00000015000000000000000e000000000000000b000000000000001200000000",
            INIT_34 => X"0000005900000000000000460000000000000029000000000000001800000000",
            INIT_35 => X"00000052000000000000004f0000000000000050000000000000005600000000",
            INIT_36 => X"0000004300000000000000480000000000000048000000000000004b00000000",
            INIT_37 => X"0000002a000000000000002d0000000000000034000000000000003b00000000",
            INIT_38 => X"0000004500000000000000440000000000000045000000000000004400000000",
            INIT_39 => X"00000011000000000000001c0000000000000033000000000000004300000000",
            INIT_3A => X"0000000b000000000000000a000000000000000c000000000000001700000000",
            INIT_3B => X"000000180000000000000011000000000000000b000000000000000900000000",
            INIT_3C => X"0000003f00000000000000210000000000000016000000000000001c00000000",
            INIT_3D => X"00000040000000000000004d000000000000004f000000000000004d00000000",
            INIT_3E => X"0000004200000000000000480000000000000049000000000000004100000000",
            INIT_3F => X"0000002b000000000000002f0000000000000036000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004e00000000000000470000000000000045000000000000004400000000",
            INIT_41 => X"000000130000000000000046000000000000005d000000000000005200000000",
            INIT_42 => X"000000250000000000000019000000000000000c000000000000001200000000",
            INIT_43 => X"0000001400000000000000210000000000000021000000000000002000000000",
            INIT_44 => X"0000002100000000000000190000000000000018000000000000001600000000",
            INIT_45 => X"0000003b000000000000003c0000000000000038000000000000003100000000",
            INIT_46 => X"0000003f0000000000000049000000000000004b000000000000003b00000000",
            INIT_47 => X"0000003500000000000000340000000000000034000000000000003900000000",
            INIT_48 => X"0000007500000000000000670000000000000059000000000000005000000000",
            INIT_49 => X"000000160000000000000055000000000000008d000000000000008000000000",
            INIT_4A => X"000000380000000000000021000000000000000f000000000000001500000000",
            INIT_4B => X"0000001c0000000000000035000000000000003d000000000000003900000000",
            INIT_4C => X"0000001400000000000000160000000000000016000000000000001500000000",
            INIT_4D => X"0000003a000000000000002d0000000000000023000000000000001800000000",
            INIT_4E => X"0000004100000000000000460000000000000048000000000000003d00000000",
            INIT_4F => X"0000003d000000000000003f0000000000000040000000000000004100000000",
            INIT_50 => X"00000095000000000000008e0000000000000083000000000000007700000000",
            INIT_51 => X"0000001800000000000000470000000000000098000000000000009800000000",
            INIT_52 => X"0000003100000000000000150000000000000011000000000000001e00000000",
            INIT_53 => X"00000021000000000000003f0000000000000044000000000000003c00000000",
            INIT_54 => X"000000110000000000000015000000000000001b000000000000001900000000",
            INIT_55 => X"0000002b000000000000001c0000000000000014000000000000000f00000000",
            INIT_56 => X"0000004a000000000000004d0000000000000046000000000000003700000000",
            INIT_57 => X"0000004100000000000000440000000000000047000000000000004900000000",
            INIT_58 => X"0000009900000000000000960000000000000094000000000000008f00000000",
            INIT_59 => X"00000017000000000000004f0000000000000099000000000000009900000000",
            INIT_5A => X"0000002e00000000000000190000000000000022000000000000002800000000",
            INIT_5B => X"0000002700000000000000370000000000000030000000000000003d00000000",
            INIT_5C => X"00000015000000000000001f0000000000000024000000000000001d00000000",
            INIT_5D => X"0000001f00000000000000120000000000000015000000000000001300000000",
            INIT_5E => X"0000004d000000000000004c000000000000003b000000000000002a00000000",
            INIT_5F => X"00000045000000000000004a000000000000004c000000000000004d00000000",
            INIT_60 => X"0000009400000000000000970000000000000095000000000000009200000000",
            INIT_61 => X"00000020000000000000006b0000000000000092000000000000009200000000",
            INIT_62 => X"0000003b00000000000000340000000000000037000000000000002b00000000",
            INIT_63 => X"00000029000000000000002c0000000000000034000000000000004700000000",
            INIT_64 => X"0000001e000000000000002c0000000000000032000000000000002200000000",
            INIT_65 => X"000000190000000000000012000000000000001c000000000000001a00000000",
            INIT_66 => X"0000005100000000000000450000000000000032000000000000002e00000000",
            INIT_67 => X"000000420000000000000049000000000000004f000000000000005100000000",
            INIT_68 => X"0000008b000000000000008f000000000000008f000000000000009000000000",
            INIT_69 => X"00000040000000000000007e0000000000000089000000000000008a00000000",
            INIT_6A => X"00000041000000000000003d000000000000002e000000000000001a00000000",
            INIT_6B => X"0000002400000000000000280000000000000040000000000000004600000000",
            INIT_6C => X"0000002800000000000000330000000000000036000000000000002400000000",
            INIT_6D => X"000000130000000000000012000000000000001d000000000000002100000000",
            INIT_6E => X"0000004e000000000000003c0000000000000033000000000000002f00000000",
            INIT_6F => X"000000370000000000000040000000000000004a000000000000004f00000000",
            INIT_70 => X"0000008600000000000000860000000000000084000000000000008500000000",
            INIT_71 => X"0000007700000000000000890000000000000088000000000000008600000000",
            INIT_72 => X"00000021000000000000001b0000000000000031000000000000004700000000",
            INIT_73 => X"000000220000000000000020000000000000002a000000000000002e00000000",
            INIT_74 => X"00000032000000000000003d0000000000000039000000000000002800000000",
            INIT_75 => X"000000110000000000000011000000000000001c000000000000002700000000",
            INIT_76 => X"0000004100000000000000300000000000000033000000000000002400000000",
            INIT_77 => X"000000320000000000000036000000000000003e000000000000004600000000",
            INIT_78 => X"000000850000000000000081000000000000007f000000000000007d00000000",
            INIT_79 => X"0000008100000000000000880000000000000091000000000000008c00000000",
            INIT_7A => X"0000001e000000000000001e000000000000005a000000000000008400000000",
            INIT_7B => X"0000002700000000000000270000000000000033000000000000004000000000",
            INIT_7C => X"0000003d00000000000000450000000000000045000000000000003100000000",
            INIT_7D => X"000000130000000000000014000000000000001c000000000000002c00000000",
            INIT_7E => X"0000002d00000000000000290000000000000030000000000000001900000000",
            INIT_7F => X"0000003d000000000000003c0000000000000039000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "sampleifmap_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000091000000000000008b0000000000000084000000000000007d00000000",
            INIT_01 => X"0000005a00000000000000750000000000000091000000000000009500000000",
            INIT_02 => X"0000005000000000000000620000000000000072000000000000008000000000",
            INIT_03 => X"000000280000000000000031000000000000004d000000000000005700000000",
            INIT_04 => X"0000003c0000000000000044000000000000003f000000000000002e00000000",
            INIT_05 => X"000000170000000000000019000000000000001f000000000000002d00000000",
            INIT_06 => X"0000002d000000000000002b000000000000002a000000000000001500000000",
            INIT_07 => X"00000032000000000000003e0000000000000042000000000000004000000000",
            INIT_08 => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_09 => X"00000068000000000000009e00000000000000a4000000000000009a00000000",
            INIT_0A => X"00000077000000000000007a00000000000000a6000000000000009500000000",
            INIT_0B => X"00000029000000000000004b0000000000000067000000000000005000000000",
            INIT_0C => X"0000003c00000000000000410000000000000038000000000000002d00000000",
            INIT_0D => X"0000001b000000000000001f0000000000000028000000000000003000000000",
            INIT_0E => X"00000032000000000000002f0000000000000023000000000000001500000000",
            INIT_0F => X"0000001400000000000000230000000000000039000000000000004100000000",
            INIT_10 => X"000000b600000000000000a40000000000000097000000000000009000000000",
            INIT_11 => X"000000b200000000000000eb00000000000000e600000000000000d200000000",
            INIT_12 => X"00000095000000000000008a00000000000000ab000000000000008500000000",
            INIT_13 => X"0000002d00000000000000550000000000000067000000000000004d00000000",
            INIT_14 => X"0000003c000000000000003f0000000000000038000000000000002b00000000",
            INIT_15 => X"0000001d00000000000000270000000000000030000000000000003500000000",
            INIT_16 => X"00000027000000000000002f000000000000001d000000000000001700000000",
            INIT_17 => X"000000150000000000000016000000000000001f000000000000002700000000",
            INIT_18 => X"000000f000000000000000e100000000000000cd00000000000000b700000000",
            INIT_19 => X"000000e600000000000000f200000000000000f200000000000000f800000000",
            INIT_1A => X"0000009f00000000000000840000000000000084000000000000008d00000000",
            INIT_1B => X"000000310000000000000056000000000000004d000000000000005300000000",
            INIT_1C => X"0000003a000000000000003c0000000000000037000000000000002a00000000",
            INIT_1D => X"00000021000000000000002f0000000000000037000000000000003900000000",
            INIT_1E => X"0000001c0000000000000027000000000000001a000000000000001900000000",
            INIT_1F => X"0000001b000000000000001c000000000000001d000000000000001900000000",
            INIT_20 => X"000000f900000000000000f700000000000000f800000000000000f100000000",
            INIT_21 => X"000000b500000000000000ab00000000000000b000000000000000ec00000000",
            INIT_22 => X"0000007600000000000000720000000000000062000000000000007800000000",
            INIT_23 => X"000000340000000000000047000000000000003c000000000000004d00000000",
            INIT_24 => X"0000003a00000000000000390000000000000036000000000000002e00000000",
            INIT_25 => X"0000002000000000000000300000000000000039000000000000003b00000000",
            INIT_26 => X"0000002500000000000000250000000000000017000000000000001800000000",
            INIT_27 => X"0000001a000000000000001f0000000000000020000000000000001c00000000",
            INIT_28 => X"000000fd00000000000000f900000000000000f900000000000000f800000000",
            INIT_29 => X"000000550000000000000053000000000000006a00000000000000e000000000",
            INIT_2A => X"000000410000000000000051000000000000004e000000000000004700000000",
            INIT_2B => X"000000310000000000000034000000000000002e000000000000003000000000",
            INIT_2C => X"0000003900000000000000360000000000000037000000000000003300000000",
            INIT_2D => X"0000001b00000000000000240000000000000033000000000000003d00000000",
            INIT_2E => X"0000003600000000000000270000000000000016000000000000001500000000",
            INIT_2F => X"0000001c000000000000001f000000000000001f000000000000002800000000",
            INIT_30 => X"000000eb00000000000000f500000000000000f800000000000000f700000000",
            INIT_31 => X"0000005e0000000000000060000000000000006d00000000000000c200000000",
            INIT_32 => X"0000001900000000000000230000000000000035000000000000004100000000",
            INIT_33 => X"00000020000000000000002d000000000000002b000000000000001c00000000",
            INIT_34 => X"0000002f000000000000002f0000000000000033000000000000002e00000000",
            INIT_35 => X"00000029000000000000002b000000000000002d000000000000003000000000",
            INIT_36 => X"0000003a0000000000000024000000000000001e000000000000002200000000",
            INIT_37 => X"0000001e000000000000001d0000000000000021000000000000003900000000",
            INIT_38 => X"0000009800000000000000b600000000000000d700000000000000ec00000000",
            INIT_39 => X"00000074000000000000007a0000000000000081000000000000008800000000",
            INIT_3A => X"00000009000000000000000d0000000000000023000000000000005100000000",
            INIT_3B => X"0000002200000000000000490000000000000034000000000000001400000000",
            INIT_3C => X"00000020000000000000001a000000000000001c000000000000001100000000",
            INIT_3D => X"00000031000000000000003b000000000000003b000000000000002f00000000",
            INIT_3E => X"000000340000000000000022000000000000001a000000000000002300000000",
            INIT_3F => X"0000001d000000000000001c000000000000002c000000000000003f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009a00000000",
            INIT_41 => X"0000005c00000000000000680000000000000076000000000000007b00000000",
            INIT_42 => X"00000012000000000000001f0000000000000046000000000000005a00000000",
            INIT_43 => X"000000340000000000000045000000000000003d000000000000001d00000000",
            INIT_44 => X"0000002800000000000000240000000000000024000000000000002200000000",
            INIT_45 => X"0000003d00000000000000410000000000000047000000000000003a00000000",
            INIT_46 => X"00000028000000000000001f0000000000000017000000000000003000000000",
            INIT_47 => X"0000001c0000000000000027000000000000003c000000000000003800000000",
            INIT_48 => X"00000068000000000000006d000000000000006b000000000000006900000000",
            INIT_49 => X"0000005d000000000000005b0000000000000058000000000000005f00000000",
            INIT_4A => X"0000003e00000000000000560000000000000062000000000000006000000000",
            INIT_4B => X"00000031000000000000002f0000000000000038000000000000003800000000",
            INIT_4C => X"00000030000000000000002a0000000000000025000000000000002800000000",
            INIT_4D => X"000000390000000000000048000000000000005b000000000000004c00000000",
            INIT_4E => X"00000023000000000000001d000000000000002c000000000000003600000000",
            INIT_4F => X"0000001d0000000000000037000000000000003d000000000000002a00000000",
            INIT_50 => X"0000005100000000000000530000000000000059000000000000005f00000000",
            INIT_51 => X"00000058000000000000005b0000000000000058000000000000005600000000",
            INIT_52 => X"0000003e00000000000000440000000000000049000000000000005300000000",
            INIT_53 => X"00000034000000000000002c0000000000000023000000000000002800000000",
            INIT_54 => X"000000310000000000000027000000000000001e000000000000002800000000",
            INIT_55 => X"000000320000000000000047000000000000005f000000000000005100000000",
            INIT_56 => X"000000230000000000000025000000000000002a000000000000002900000000",
            INIT_57 => X"00000028000000000000003a0000000000000030000000000000002200000000",
            INIT_58 => X"00000055000000000000004f0000000000000049000000000000004b00000000",
            INIT_59 => X"00000040000000000000004c0000000000000053000000000000005700000000",
            INIT_5A => X"0000003b000000000000002a0000000000000027000000000000003300000000",
            INIT_5B => X"0000003100000000000000290000000000000022000000000000003200000000",
            INIT_5C => X"000000270000000000000024000000000000001e000000000000002600000000",
            INIT_5D => X"0000002d000000000000003c0000000000000045000000000000003700000000",
            INIT_5E => X"0000001d00000000000000220000000000000026000000000000002600000000",
            INIT_5F => X"0000003300000000000000300000000000000024000000000000002000000000",
            INIT_60 => X"0000004d000000000000004f000000000000004e000000000000004c00000000",
            INIT_61 => X"00000021000000000000002c0000000000000039000000000000004400000000",
            INIT_62 => X"0000003d000000000000002e000000000000001e000000000000001d00000000",
            INIT_63 => X"0000002600000000000000320000000000000029000000000000003700000000",
            INIT_64 => X"0000001e000000000000001d000000000000001a000000000000001d00000000",
            INIT_65 => X"00000030000000000000002e0000000000000025000000000000001d00000000",
            INIT_66 => X"0000001800000000000000190000000000000025000000000000002e00000000",
            INIT_67 => X"0000002f00000000000000240000000000000020000000000000001e00000000",
            INIT_68 => X"000000320000000000000040000000000000004a000000000000005000000000",
            INIT_69 => X"0000001b000000000000001e0000000000000020000000000000002600000000",
            INIT_6A => X"0000003c000000000000002d000000000000001b000000000000001b00000000",
            INIT_6B => X"0000001d000000000000002c000000000000002f000000000000003500000000",
            INIT_6C => X"0000001c00000000000000170000000000000017000000000000001c00000000",
            INIT_6D => X"0000002500000000000000200000000000000018000000000000001900000000",
            INIT_6E => X"000000150000000000000015000000000000001d000000000000002300000000",
            INIT_6F => X"00000022000000000000001c000000000000001e000000000000001a00000000",
            INIT_70 => X"0000001a0000000000000021000000000000002d000000000000003a00000000",
            INIT_71 => X"0000001c0000000000000021000000000000001d000000000000001a00000000",
            INIT_72 => X"0000003300000000000000270000000000000018000000000000001b00000000",
            INIT_73 => X"0000001c00000000000000210000000000000032000000000000003100000000",
            INIT_74 => X"0000001d00000000000000190000000000000015000000000000001b00000000",
            INIT_75 => X"0000001700000000000000190000000000000015000000000000001800000000",
            INIT_76 => X"000000120000000000000016000000000000001a000000000000001700000000",
            INIT_77 => X"000000170000000000000019000000000000001a000000000000001500000000",
            INIT_78 => X"0000001500000000000000180000000000000017000000000000001b00000000",
            INIT_79 => X"0000001900000000000000180000000000000019000000000000001a00000000",
            INIT_7A => X"0000003000000000000000210000000000000016000000000000001a00000000",
            INIT_7B => X"0000001800000000000000230000000000000033000000000000002a00000000",
            INIT_7C => X"0000001800000000000000150000000000000014000000000000001500000000",
            INIT_7D => X"00000019000000000000001d0000000000000017000000000000001700000000",
            INIT_7E => X"000000120000000000000016000000000000001b000000000000001800000000",
            INIT_7F => X"0000001600000000000000180000000000000016000000000000001100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "sampleifmap_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004100000000000000150000000000000013000000000000001700000000",
            INIT_01 => X"000000b200000000000000b700000000000000bc00000000000000a400000000",
            INIT_02 => X"000000ba00000000000000ba00000000000000ac00000000000000aa00000000",
            INIT_03 => X"000000b700000000000000b600000000000000b700000000000000b800000000",
            INIT_04 => X"0000005c000000000000007f00000000000000a400000000000000b400000000",
            INIT_05 => X"000000c20000000000000099000000000000006e000000000000006b00000000",
            INIT_06 => X"000000c600000000000000c500000000000000c900000000000000c300000000",
            INIT_07 => X"000000c500000000000000c700000000000000c800000000000000c900000000",
            INIT_08 => X"0000002e00000000000000150000000000000013000000000000001700000000",
            INIT_09 => X"000000b200000000000000bf00000000000000ca000000000000009900000000",
            INIT_0A => X"000000b700000000000000a9000000000000009e00000000000000a400000000",
            INIT_0B => X"000000b200000000000000b400000000000000b800000000000000ba00000000",
            INIT_0C => X"00000056000000000000008a00000000000000ad00000000000000b400000000",
            INIT_0D => X"000000ce00000000000000b4000000000000006a000000000000004a00000000",
            INIT_0E => X"000000ce00000000000000d000000000000000d500000000000000cf00000000",
            INIT_0F => X"000000ca00000000000000cc00000000000000cd00000000000000cf00000000",
            INIT_10 => X"0000001f00000000000000170000000000000014000000000000001700000000",
            INIT_11 => X"000000a800000000000000b900000000000000c8000000000000007f00000000",
            INIT_12 => X"000000a2000000000000009a000000000000009e000000000000009f00000000",
            INIT_13 => X"000000b200000000000000b300000000000000b200000000000000b200000000",
            INIT_14 => X"0000007d00000000000000b600000000000000be00000000000000b500000000",
            INIT_15 => X"000000d100000000000000c50000000000000072000000000000004700000000",
            INIT_16 => X"000000d300000000000000d500000000000000d800000000000000d500000000",
            INIT_17 => X"000000ce00000000000000d000000000000000d300000000000000d400000000",
            INIT_18 => X"0000001700000000000000180000000000000015000000000000001700000000",
            INIT_19 => X"000000a000000000000000af00000000000000bd000000000000006300000000",
            INIT_1A => X"0000009500000000000000a600000000000000a800000000000000a800000000",
            INIT_1B => X"000000c300000000000000bf00000000000000ba00000000000000aa00000000",
            INIT_1C => X"0000008d00000000000000bc00000000000000c800000000000000c300000000",
            INIT_1D => X"000000d600000000000000d20000000000000092000000000000006300000000",
            INIT_1E => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1F => X"000000d600000000000000d700000000000000d900000000000000d900000000",
            INIT_20 => X"0000001500000000000000170000000000000017000000000000001900000000",
            INIT_21 => X"0000009700000000000000a500000000000000aa000000000000004800000000",
            INIT_22 => X"0000009b00000000000000b900000000000000b700000000000000af00000000",
            INIT_23 => X"000000bc00000000000000a9000000000000009d000000000000009200000000",
            INIT_24 => X"0000008d00000000000000b200000000000000c400000000000000c500000000",
            INIT_25 => X"000000db00000000000000d300000000000000ac000000000000007900000000",
            INIT_26 => X"000000d900000000000000d900000000000000d900000000000000dd00000000",
            INIT_27 => X"000000ce00000000000000d100000000000000d400000000000000d600000000",
            INIT_28 => X"00000017000000000000001a000000000000001b000000000000001a00000000",
            INIT_29 => X"0000009a00000000000000a4000000000000008f000000000000003100000000",
            INIT_2A => X"000000a600000000000000c800000000000000c200000000000000a900000000",
            INIT_2B => X"000000970000000000000080000000000000007d000000000000008200000000",
            INIT_2C => X"0000008f000000000000009400000000000000a500000000000000a500000000",
            INIT_2D => X"000000c900000000000000bc00000000000000b6000000000000009300000000",
            INIT_2E => X"000000db00000000000000d500000000000000d900000000000000d400000000",
            INIT_2F => X"000000d300000000000000d700000000000000d700000000000000dc00000000",
            INIT_30 => X"00000019000000000000001b000000000000001a000000000000001e00000000",
            INIT_31 => X"000000ab00000000000000b4000000000000007d000000000000002500000000",
            INIT_32 => X"000000b300000000000000ca00000000000000c500000000000000a900000000",
            INIT_33 => X"00000082000000000000007a0000000000000071000000000000008b00000000",
            INIT_34 => X"0000008c000000000000007a0000000000000085000000000000007700000000",
            INIT_35 => X"000000c900000000000000bf00000000000000cb00000000000000b900000000",
            INIT_36 => X"000000db00000000000000d700000000000000da00000000000000d700000000",
            INIT_37 => X"000000e000000000000000dc00000000000000da00000000000000dc00000000",
            INIT_38 => X"00000024000000000000001f0000000000000030000000000000005e00000000",
            INIT_39 => X"000000a800000000000000c100000000000000af000000000000006400000000",
            INIT_3A => X"000000c300000000000000c600000000000000c000000000000000a300000000",
            INIT_3B => X"00000084000000000000008e000000000000009100000000000000ae00000000",
            INIT_3C => X"0000008b000000000000007a0000000000000079000000000000006a00000000",
            INIT_3D => X"000000d500000000000000bd00000000000000d100000000000000c000000000",
            INIT_3E => X"000000e800000000000000ef00000000000000ed00000000000000f200000000",
            INIT_3F => X"000000e500000000000000de00000000000000d500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007a0000000000000072000000000000009e00000000000000b400000000",
            INIT_41 => X"000000a000000000000000be00000000000000be00000000000000b100000000",
            INIT_42 => X"000000c800000000000000c500000000000000ad000000000000008500000000",
            INIT_43 => X"0000009200000000000000a700000000000000b900000000000000c200000000",
            INIT_44 => X"0000008d00000000000000850000000000000081000000000000008100000000",
            INIT_45 => X"000000dc00000000000000bd00000000000000c900000000000000b100000000",
            INIT_46 => X"000000d500000000000000e800000000000000eb00000000000000f100000000",
            INIT_47 => X"000000ea00000000000000e100000000000000c700000000000000bd00000000",
            INIT_48 => X"000000ba00000000000000b200000000000000c000000000000000c500000000",
            INIT_49 => X"0000009d00000000000000c500000000000000c300000000000000c100000000",
            INIT_4A => X"000000bf00000000000000b900000000000000a3000000000000008000000000",
            INIT_4B => X"0000009700000000000000b200000000000000c300000000000000c100000000",
            INIT_4C => X"0000008600000000000000830000000000000081000000000000007200000000",
            INIT_4D => X"000000ea00000000000000d000000000000000c200000000000000aa00000000",
            INIT_4E => X"000000c900000000000000eb00000000000000f000000000000000ec00000000",
            INIT_4F => X"000000eb00000000000000d000000000000000bb00000000000000b900000000",
            INIT_50 => X"000000c000000000000000bb00000000000000c400000000000000ca00000000",
            INIT_51 => X"0000009700000000000000c500000000000000cd00000000000000c800000000",
            INIT_52 => X"000000bd00000000000000b800000000000000af000000000000009500000000",
            INIT_53 => X"0000008800000000000000a800000000000000bb00000000000000c100000000",
            INIT_54 => X"0000008100000000000000800000000000000080000000000000007500000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b500000000000000a700000000",
            INIT_56 => X"000000ce00000000000000ee00000000000000f300000000000000f300000000",
            INIT_57 => X"000000dd00000000000000c100000000000000bb00000000000000ba00000000",
            INIT_58 => X"000000c000000000000000c500000000000000cd00000000000000cd00000000",
            INIT_59 => X"000000a000000000000000c200000000000000d000000000000000cb00000000",
            INIT_5A => X"000000bf00000000000000c100000000000000bf00000000000000a800000000",
            INIT_5B => X"00000077000000000000009200000000000000ac00000000000000c100000000",
            INIT_5C => X"000000870000000000000085000000000000008e000000000000007c00000000",
            INIT_5D => X"000000ea00000000000000bf00000000000000b000000000000000a700000000",
            INIT_5E => X"000000d700000000000000ec00000000000000f100000000000000f300000000",
            INIT_5F => X"000000c400000000000000b900000000000000b800000000000000ba00000000",
            INIT_60 => X"000000c100000000000000c800000000000000cc00000000000000ce00000000",
            INIT_61 => X"000000b400000000000000bf00000000000000c700000000000000c500000000",
            INIT_62 => X"000000ad00000000000000b700000000000000b300000000000000ac00000000",
            INIT_63 => X"00000083000000000000009800000000000000ae00000000000000ae00000000",
            INIT_64 => X"0000009a000000000000008e00000000000000a6000000000000008d00000000",
            INIT_65 => X"000000e600000000000000bf00000000000000ac00000000000000a900000000",
            INIT_66 => X"000000e400000000000000ef00000000000000f100000000000000f000000000",
            INIT_67 => X"000000c000000000000000b800000000000000ba00000000000000c800000000",
            INIT_68 => X"000000bf00000000000000c600000000000000ca00000000000000d200000000",
            INIT_69 => X"000000ca00000000000000b100000000000000b400000000000000c900000000",
            INIT_6A => X"0000008e000000000000008e000000000000009a00000000000000ab00000000",
            INIT_6B => X"0000009c000000000000009300000000000000a800000000000000a800000000",
            INIT_6C => X"000000a4000000000000009600000000000000a900000000000000af00000000",
            INIT_6D => X"000000e600000000000000c500000000000000a0000000000000009e00000000",
            INIT_6E => X"000000f200000000000000f400000000000000f100000000000000f100000000",
            INIT_6F => X"000000d700000000000000c300000000000000bf00000000000000e200000000",
            INIT_70 => X"000000c000000000000000c700000000000000c900000000000000d300000000",
            INIT_71 => X"000000d700000000000000a100000000000000aa00000000000000cf00000000",
            INIT_72 => X"000000ac00000000000000ad00000000000000ba00000000000000bd00000000",
            INIT_73 => X"0000007f000000000000008900000000000000b100000000000000be00000000",
            INIT_74 => X"000000a0000000000000009600000000000000ae00000000000000b400000000",
            INIT_75 => X"000000ec00000000000000c100000000000000b000000000000000af00000000",
            INIT_76 => X"000000fb00000000000000f300000000000000f200000000000000f500000000",
            INIT_77 => X"000000e100000000000000d400000000000000c900000000000000ef00000000",
            INIT_78 => X"000000c100000000000000c500000000000000c400000000000000d300000000",
            INIT_79 => X"000000d9000000000000009a00000000000000b500000000000000d100000000",
            INIT_7A => X"000000b900000000000000c300000000000000c500000000000000ce00000000",
            INIT_7B => X"0000009800000000000000a600000000000000ad00000000000000aa00000000",
            INIT_7C => X"0000009800000000000000a600000000000000b800000000000000a300000000",
            INIT_7D => X"000000cc00000000000000af00000000000000b500000000000000c000000000",
            INIT_7E => X"000000f700000000000000f400000000000000f300000000000000ee00000000",
            INIT_7F => X"000000e200000000000000e200000000000000d500000000000000df00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "sampleifmap_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b500000000000000b400000000000000c200000000000000d600000000",
            INIT_01 => X"000000c6000000000000009b00000000000000c400000000000000c500000000",
            INIT_02 => X"000000b700000000000000ae00000000000000c000000000000000d600000000",
            INIT_03 => X"000000b200000000000000ae00000000000000a100000000000000ad00000000",
            INIT_04 => X"0000009300000000000000bd00000000000000a4000000000000008000000000",
            INIT_05 => X"00000076000000000000009c00000000000000b400000000000000a700000000",
            INIT_06 => X"000000eb00000000000000ef00000000000000d7000000000000009d00000000",
            INIT_07 => X"000000e400000000000000ea00000000000000d600000000000000ce00000000",
            INIT_08 => X"000000a300000000000000a600000000000000c600000000000000d700000000",
            INIT_09 => X"000000b900000000000000be00000000000000ca00000000000000b400000000",
            INIT_0A => X"000000d600000000000000cd00000000000000d200000000000000cf00000000",
            INIT_0B => X"000000ad00000000000000b000000000000000ae00000000000000c100000000",
            INIT_0C => X"0000009900000000000000bf0000000000000089000000000000008100000000",
            INIT_0D => X"0000008700000000000000ab00000000000000c800000000000000a300000000",
            INIT_0E => X"000000c100000000000000b80000000000000090000000000000007400000000",
            INIT_0F => X"000000eb00000000000000ef00000000000000d200000000000000bb00000000",
            INIT_10 => X"000000a400000000000000ae00000000000000cd00000000000000d800000000",
            INIT_11 => X"000000c200000000000000d200000000000000cb00000000000000b900000000",
            INIT_12 => X"000000e200000000000000da00000000000000d300000000000000bf00000000",
            INIT_13 => X"000000b300000000000000be00000000000000cb00000000000000e100000000",
            INIT_14 => X"0000009e00000000000000a80000000000000079000000000000009700000000",
            INIT_15 => X"000000ac00000000000000aa00000000000000c200000000000000a700000000",
            INIT_16 => X"000000a900000000000000990000000000000083000000000000009a00000000",
            INIT_17 => X"000000ec00000000000000de00000000000000b800000000000000a200000000",
            INIT_18 => X"000000b400000000000000c000000000000000d000000000000000d800000000",
            INIT_19 => X"000000d200000000000000d100000000000000ca00000000000000c500000000",
            INIT_1A => X"000000cc00000000000000c500000000000000bd00000000000000ba00000000",
            INIT_1B => X"000000b500000000000000cf00000000000000d500000000000000d100000000",
            INIT_1C => X"000000af0000000000000092000000000000009500000000000000b200000000",
            INIT_1D => X"000000ab000000000000009c00000000000000ae00000000000000b700000000",
            INIT_1E => X"000000b400000000000000a9000000000000009400000000000000a300000000",
            INIT_1F => X"000000cc00000000000000ac00000000000000a000000000000000a600000000",
            INIT_20 => X"000000b600000000000000ca00000000000000d500000000000000da00000000",
            INIT_21 => X"000000ca00000000000000c900000000000000cb00000000000000bf00000000",
            INIT_22 => X"000000c000000000000000c100000000000000c300000000000000ca00000000",
            INIT_23 => X"000000c700000000000000cf00000000000000c600000000000000b200000000",
            INIT_24 => X"000000bb00000000000000a600000000000000cb00000000000000d300000000",
            INIT_25 => X"000000a60000000000000093000000000000009b00000000000000b100000000",
            INIT_26 => X"000000af00000000000000b600000000000000ab00000000000000a700000000",
            INIT_27 => X"000000a7000000000000009f000000000000009c000000000000009c00000000",
            INIT_28 => X"000000ba00000000000000d100000000000000d700000000000000d900000000",
            INIT_29 => X"000000c800000000000000d000000000000000c800000000000000b300000000",
            INIT_2A => X"000000ba00000000000000d200000000000000d700000000000000d100000000",
            INIT_2B => X"000000c200000000000000c400000000000000b600000000000000a100000000",
            INIT_2C => X"000000b900000000000000be00000000000000cf00000000000000cb00000000",
            INIT_2D => X"000000a6000000000000009b000000000000008e000000000000009b00000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000b300000000000000ac00000000",
            INIT_2F => X"0000008f000000000000009e000000000000009e000000000000009600000000",
            INIT_30 => X"000000c000000000000000d600000000000000d500000000000000d600000000",
            INIT_31 => X"000000d900000000000000da00000000000000c500000000000000a900000000",
            INIT_32 => X"000000c300000000000000d400000000000000d900000000000000d700000000",
            INIT_33 => X"000000bf00000000000000c300000000000000b300000000000000aa00000000",
            INIT_34 => X"000000aa00000000000000c000000000000000c000000000000000be00000000",
            INIT_35 => X"000000aa00000000000000a7000000000000008e000000000000008400000000",
            INIT_36 => X"0000009d00000000000000ad00000000000000b300000000000000aa00000000",
            INIT_37 => X"0000007d00000000000000860000000000000093000000000000009d00000000",
            INIT_38 => X"000000ca00000000000000d300000000000000d100000000000000d500000000",
            INIT_39 => X"000000de00000000000000d800000000000000c100000000000000a800000000",
            INIT_3A => X"000000cd00000000000000d300000000000000de00000000000000df00000000",
            INIT_3B => X"000000c600000000000000c900000000000000c200000000000000c200000000",
            INIT_3C => X"0000009900000000000000bc00000000000000c400000000000000c600000000",
            INIT_3D => X"000000a700000000000000ab000000000000009b000000000000008600000000",
            INIT_3E => X"000000a500000000000000b200000000000000bd00000000000000a600000000",
            INIT_3F => X"000000890000000000000085000000000000008e00000000000000a300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ca00000000000000ce00000000000000ce00000000000000d300000000",
            INIT_41 => X"000000d500000000000000d300000000000000bf00000000000000af00000000",
            INIT_42 => X"000000ab00000000000000c600000000000000d800000000000000d600000000",
            INIT_43 => X"000000c900000000000000c900000000000000ce00000000000000c200000000",
            INIT_44 => X"0000009600000000000000b100000000000000c500000000000000c800000000",
            INIT_45 => X"0000009d00000000000000a7000000000000009e000000000000009000000000",
            INIT_46 => X"000000a800000000000000b000000000000000b5000000000000009f00000000",
            INIT_47 => X"0000009000000000000000950000000000000096000000000000009800000000",
            INIT_48 => X"000000c100000000000000c900000000000000cc00000000000000d200000000",
            INIT_49 => X"000000d200000000000000d000000000000000bc00000000000000b500000000",
            INIT_4A => X"0000007a00000000000000a000000000000000ce00000000000000cd00000000",
            INIT_4B => X"000000c200000000000000c600000000000000d000000000000000b100000000",
            INIT_4C => X"0000009600000000000000a600000000000000b800000000000000c100000000",
            INIT_4D => X"0000009900000000000000a0000000000000009c000000000000008b00000000",
            INIT_4E => X"0000009b000000000000009f00000000000000a0000000000000009b00000000",
            INIT_4F => X"00000083000000000000008c0000000000000098000000000000009800000000",
            INIT_50 => X"000000bb00000000000000c600000000000000ca00000000000000d200000000",
            INIT_51 => X"000000d600000000000000cd00000000000000b200000000000000ae00000000",
            INIT_52 => X"0000008300000000000000a400000000000000cb00000000000000d100000000",
            INIT_53 => X"000000b600000000000000bb00000000000000ca00000000000000b400000000",
            INIT_54 => X"0000008b000000000000009d00000000000000a900000000000000b600000000",
            INIT_55 => X"00000090000000000000009a0000000000000099000000000000008600000000",
            INIT_56 => X"0000008d0000000000000083000000000000008d000000000000009700000000",
            INIT_57 => X"000000930000000000000096000000000000009b000000000000009d00000000",
            INIT_58 => X"000000b500000000000000c200000000000000c800000000000000d200000000",
            INIT_59 => X"000000d700000000000000c400000000000000a800000000000000a800000000",
            INIT_5A => X"000000b800000000000000bd00000000000000c700000000000000d400000000",
            INIT_5B => X"000000ac00000000000000ad00000000000000b900000000000000cb00000000",
            INIT_5C => X"000000760000000000000093000000000000009b00000000000000a300000000",
            INIT_5D => X"0000008d00000000000000910000000000000094000000000000008300000000",
            INIT_5E => X"00000085000000000000007f0000000000000084000000000000009000000000",
            INIT_5F => X"0000009c00000000000000a200000000000000a3000000000000009500000000",
            INIT_60 => X"000000b400000000000000bd00000000000000c200000000000000d000000000",
            INIT_61 => X"000000d300000000000000bd000000000000009e00000000000000a200000000",
            INIT_62 => X"000000c700000000000000c200000000000000c500000000000000d300000000",
            INIT_63 => X"000000a400000000000000a300000000000000ac00000000000000bf00000000",
            INIT_64 => X"0000006d00000000000000820000000000000093000000000000009e00000000",
            INIT_65 => X"0000009100000000000000900000000000000090000000000000008900000000",
            INIT_66 => X"00000086000000000000007c0000000000000084000000000000009000000000",
            INIT_67 => X"00000093000000000000009f00000000000000a2000000000000009700000000",
            INIT_68 => X"000000b500000000000000b000000000000000b100000000000000c200000000",
            INIT_69 => X"000000cd00000000000000b3000000000000008f000000000000009f00000000",
            INIT_6A => X"000000be00000000000000c200000000000000c700000000000000d000000000",
            INIT_6B => X"000000a1000000000000009c00000000000000a500000000000000b500000000",
            INIT_6C => X"0000007200000000000000700000000000000088000000000000009500000000",
            INIT_6D => X"00000092000000000000008a0000000000000085000000000000008900000000",
            INIT_6E => X"0000009000000000000000830000000000000083000000000000009200000000",
            INIT_6F => X"0000008d00000000000000940000000000000095000000000000009600000000",
            INIT_70 => X"000000b200000000000000a5000000000000009d00000000000000ac00000000",
            INIT_71 => X"000000c7000000000000009c000000000000008500000000000000a700000000",
            INIT_72 => X"000000c200000000000000c700000000000000c700000000000000ce00000000",
            INIT_73 => X"0000008b0000000000000084000000000000008500000000000000a000000000",
            INIT_74 => X"0000007e000000000000006b000000000000007e000000000000008c00000000",
            INIT_75 => X"00000095000000000000008a0000000000000081000000000000008200000000",
            INIT_76 => X"0000008e0000000000000091000000000000008c000000000000008d00000000",
            INIT_77 => X"000000980000000000000095000000000000008c000000000000008800000000",
            INIT_78 => X"0000009b00000000000000900000000000000086000000000000009700000000",
            INIT_79 => X"000000b70000000000000082000000000000007d000000000000009e00000000",
            INIT_7A => X"000000a500000000000000b700000000000000bf00000000000000c500000000",
            INIT_7B => X"00000069000000000000005e0000000000000067000000000000008000000000",
            INIT_7C => X"0000007c00000000000000750000000000000070000000000000007700000000",
            INIT_7D => X"0000008f000000000000008b000000000000007d000000000000007900000000",
            INIT_7E => X"0000007d0000000000000081000000000000008c000000000000008b00000000",
            INIT_7F => X"00000096000000000000009b0000000000000095000000000000008400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "sampleifmap_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002f00000000000000100000000000000015000000000000001300000000",
            INIT_01 => X"0000008e00000000000000930000000000000093000000000000008300000000",
            INIT_02 => X"0000008e00000000000000900000000000000089000000000000008700000000",
            INIT_03 => X"0000008f000000000000008c000000000000008c000000000000008d00000000",
            INIT_04 => X"000000490000000000000060000000000000007e000000000000008c00000000",
            INIT_05 => X"000000a40000000000000082000000000000005d000000000000005f00000000",
            INIT_06 => X"0000009d000000000000009b000000000000009c000000000000009b00000000",
            INIT_07 => X"000000970000000000000098000000000000009b000000000000009e00000000",
            INIT_08 => X"0000001f00000000000000110000000000000014000000000000001400000000",
            INIT_09 => X"00000092000000000000009b00000000000000a1000000000000007a00000000",
            INIT_0A => X"00000095000000000000008b0000000000000088000000000000008a00000000",
            INIT_0B => X"0000009700000000000000920000000000000096000000000000009800000000",
            INIT_0C => X"0000004900000000000000750000000000000096000000000000009f00000000",
            INIT_0D => X"000000af000000000000009c0000000000000058000000000000004100000000",
            INIT_0E => X"000000ad00000000000000ab00000000000000a900000000000000a800000000",
            INIT_0F => X"000000a300000000000000a400000000000000a800000000000000ac00000000",
            INIT_10 => X"0000001500000000000000140000000000000014000000000000001400000000",
            INIT_11 => X"0000008c000000000000009700000000000000a2000000000000006600000000",
            INIT_12 => X"0000008b00000000000000880000000000000095000000000000008d00000000",
            INIT_13 => X"0000009f00000000000000980000000000000099000000000000009a00000000",
            INIT_14 => X"0000006d00000000000000a100000000000000ab00000000000000a600000000",
            INIT_15 => X"000000b700000000000000b10000000000000061000000000000003a00000000",
            INIT_16 => X"000000b200000000000000b100000000000000b200000000000000b300000000",
            INIT_17 => X"000000a600000000000000a900000000000000ad00000000000000b100000000",
            INIT_18 => X"0000001100000000000000150000000000000014000000000000001400000000",
            INIT_19 => X"00000082000000000000008c0000000000000099000000000000004f00000000",
            INIT_1A => X"00000087000000000000009d00000000000000a4000000000000009700000000",
            INIT_1B => X"000000b000000000000000a900000000000000a6000000000000009900000000",
            INIT_1C => X"0000007600000000000000a100000000000000af00000000000000b000000000",
            INIT_1D => X"000000c300000000000000c40000000000000085000000000000005200000000",
            INIT_1E => X"000000b300000000000000b400000000000000b700000000000000bd00000000",
            INIT_1F => X"000000ab00000000000000ad00000000000000b100000000000000b300000000",
            INIT_20 => X"0000001300000000000000150000000000000014000000000000001500000000",
            INIT_21 => X"0000007700000000000000820000000000000089000000000000003800000000",
            INIT_22 => X"0000009200000000000000b300000000000000b2000000000000009c00000000",
            INIT_23 => X"000000a70000000000000094000000000000008b000000000000008400000000",
            INIT_24 => X"00000078000000000000009800000000000000a900000000000000af00000000",
            INIT_25 => X"000000d200000000000000ce00000000000000a7000000000000006d00000000",
            INIT_26 => X"000000bf00000000000000c300000000000000c900000000000000d100000000",
            INIT_27 => X"000000ac00000000000000b100000000000000b600000000000000ba00000000",
            INIT_28 => X"0000001600000000000000170000000000000016000000000000001600000000",
            INIT_29 => X"0000007800000000000000820000000000000073000000000000002600000000",
            INIT_2A => X"0000009e00000000000000c300000000000000b9000000000000009200000000",
            INIT_2B => X"00000084000000000000006b000000000000006c000000000000007600000000",
            INIT_2C => X"000000840000000000000081000000000000008f000000000000009200000000",
            INIT_2D => X"000000c700000000000000be00000000000000b7000000000000008f00000000",
            INIT_2E => X"000000d100000000000000cc00000000000000d100000000000000cf00000000",
            INIT_2F => X"000000c200000000000000c700000000000000ca00000000000000d100000000",
            INIT_30 => X"0000001400000000000000150000000000000013000000000000001800000000",
            INIT_31 => X"0000009400000000000000a10000000000000071000000000000001e00000000",
            INIT_32 => X"000000aa00000000000000c200000000000000ba000000000000009700000000",
            INIT_33 => X"0000007100000000000000690000000000000062000000000000008000000000",
            INIT_34 => X"00000080000000000000006b0000000000000074000000000000006800000000",
            INIT_35 => X"000000c500000000000000c000000000000000ca00000000000000b200000000",
            INIT_36 => X"000000d700000000000000d100000000000000cf00000000000000ce00000000",
            INIT_37 => X"000000da00000000000000d700000000000000d600000000000000d800000000",
            INIT_38 => X"0000001d00000000000000180000000000000029000000000000005800000000",
            INIT_39 => X"0000009c00000000000000ba00000000000000ae000000000000006000000000",
            INIT_3A => X"000000ba00000000000000bd00000000000000b5000000000000009500000000",
            INIT_3B => X"000000760000000000000081000000000000008400000000000000a400000000",
            INIT_3C => X"0000007c000000000000006c000000000000006b000000000000005c00000000",
            INIT_3D => X"000000ce00000000000000bb00000000000000cc00000000000000b400000000",
            INIT_3E => X"000000e400000000000000e700000000000000e000000000000000e600000000",
            INIT_3F => X"000000e200000000000000dc00000000000000d300000000000000cd00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000075000000000000006d000000000000009900000000000000b100000000",
            INIT_41 => X"0000009300000000000000b700000000000000bd00000000000000af00000000",
            INIT_42 => X"000000c000000000000000bc00000000000000a1000000000000007800000000",
            INIT_43 => X"00000083000000000000009a00000000000000ad00000000000000b800000000",
            INIT_44 => X"0000007f00000000000000770000000000000073000000000000007300000000",
            INIT_45 => X"000000d800000000000000bc00000000000000c500000000000000a600000000",
            INIT_46 => X"000000d300000000000000e300000000000000e200000000000000e900000000",
            INIT_47 => X"000000e800000000000000e000000000000000c600000000000000bc00000000",
            INIT_48 => X"000000b600000000000000af00000000000000bc00000000000000c200000000",
            INIT_49 => X"0000009000000000000000be00000000000000c200000000000000bf00000000",
            INIT_4A => X"000000b600000000000000b10000000000000098000000000000007300000000",
            INIT_4B => X"0000008a00000000000000a400000000000000b600000000000000b700000000",
            INIT_4C => X"0000007b00000000000000770000000000000076000000000000006600000000",
            INIT_4D => X"000000e900000000000000d000000000000000bd00000000000000a000000000",
            INIT_4E => X"000000cb00000000000000ea00000000000000eb00000000000000e800000000",
            INIT_4F => X"000000eb00000000000000d100000000000000bd00000000000000bb00000000",
            INIT_50 => X"000000bb00000000000000b700000000000000c000000000000000c700000000",
            INIT_51 => X"0000008a00000000000000bf00000000000000cd00000000000000c600000000",
            INIT_52 => X"000000b500000000000000b000000000000000a5000000000000008800000000",
            INIT_53 => X"0000007c000000000000009a00000000000000af00000000000000b800000000",
            INIT_54 => X"0000007800000000000000770000000000000076000000000000006b00000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b0000000000000009e00000000",
            INIT_56 => X"000000d400000000000000f200000000000000f400000000000000f300000000",
            INIT_57 => X"000000e000000000000000c600000000000000c000000000000000c000000000",
            INIT_58 => X"000000bb00000000000000c100000000000000c900000000000000c900000000",
            INIT_59 => X"0000009200000000000000bc00000000000000d100000000000000c900000000",
            INIT_5A => X"000000b700000000000000b900000000000000b6000000000000009b00000000",
            INIT_5B => X"0000006b0000000000000084000000000000009f00000000000000b700000000",
            INIT_5C => X"0000007e000000000000007c0000000000000085000000000000007300000000",
            INIT_5D => X"000000eb00000000000000bd00000000000000aa000000000000009e00000000",
            INIT_5E => X"000000de00000000000000f200000000000000f600000000000000f600000000",
            INIT_5F => X"000000ca00000000000000c000000000000000c000000000000000c200000000",
            INIT_60 => X"000000bd00000000000000c500000000000000c900000000000000cb00000000",
            INIT_61 => X"000000a500000000000000b700000000000000c600000000000000c400000000",
            INIT_62 => X"000000a500000000000000b000000000000000aa000000000000009f00000000",
            INIT_63 => X"00000078000000000000008a00000000000000a200000000000000a400000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008500000000",
            INIT_65 => X"000000e700000000000000bd00000000000000a500000000000000a100000000",
            INIT_66 => X"000000ea00000000000000f700000000000000f800000000000000f400000000",
            INIT_67 => X"000000c700000000000000c100000000000000c300000000000000d000000000",
            INIT_68 => X"000000b900000000000000c400000000000000ca00000000000000d000000000",
            INIT_69 => X"000000b9000000000000009c00000000000000a700000000000000c100000000",
            INIT_6A => X"000000870000000000000087000000000000009100000000000000a100000000",
            INIT_6B => X"0000008f0000000000000089000000000000009e00000000000000a100000000",
            INIT_6C => X"000000a2000000000000009500000000000000a400000000000000a400000000",
            INIT_6D => X"000000e400000000000000c3000000000000009d000000000000009900000000",
            INIT_6E => X"000000f500000000000000f900000000000000f700000000000000f200000000",
            INIT_6F => X"000000de00000000000000cc00000000000000c700000000000000e800000000",
            INIT_70 => X"000000b600000000000000c500000000000000cc00000000000000d200000000",
            INIT_71 => X"000000c1000000000000007d000000000000008e00000000000000bf00000000",
            INIT_72 => X"000000a700000000000000a600000000000000b100000000000000b500000000",
            INIT_73 => X"00000072000000000000008200000000000000aa00000000000000b800000000",
            INIT_74 => X"0000009e000000000000009800000000000000aa00000000000000a500000000",
            INIT_75 => X"000000e700000000000000bd00000000000000ae00000000000000ab00000000",
            INIT_76 => X"000000fb00000000000000f500000000000000f400000000000000f200000000",
            INIT_77 => X"000000e900000000000000dd00000000000000cf00000000000000f200000000",
            INIT_78 => X"000000b900000000000000c500000000000000c800000000000000d400000000",
            INIT_79 => X"000000c00000000000000070000000000000009100000000000000bd00000000",
            INIT_7A => X"000000b400000000000000bd00000000000000be00000000000000c700000000",
            INIT_7B => X"0000008900000000000000a000000000000000a700000000000000a400000000",
            INIT_7C => X"0000009100000000000000a200000000000000b0000000000000009200000000",
            INIT_7D => X"000000c300000000000000a800000000000000b100000000000000b800000000",
            INIT_7E => X"000000f900000000000000f500000000000000f100000000000000e800000000",
            INIT_7F => X"000000eb00000000000000ec00000000000000dd00000000000000e400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "sampleifmap_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ae00000000000000b600000000000000c700000000000000d800000000",
            INIT_01 => X"000000ad000000000000006e000000000000009b00000000000000b000000000",
            INIT_02 => X"000000b200000000000000a800000000000000ba00000000000000d000000000",
            INIT_03 => X"000000a400000000000000a7000000000000009b00000000000000a800000000",
            INIT_04 => X"0000008600000000000000b10000000000000096000000000000006e00000000",
            INIT_05 => X"00000068000000000000009000000000000000ab000000000000009a00000000",
            INIT_06 => X"000000ed00000000000000ee00000000000000d1000000000000009100000000",
            INIT_07 => X"000000ed00000000000000f300000000000000dd00000000000000d200000000",
            INIT_08 => X"0000009e00000000000000a900000000000000ce00000000000000db00000000",
            INIT_09 => X"000000a2000000000000009500000000000000a700000000000000a300000000",
            INIT_0A => X"000000d100000000000000c800000000000000cd00000000000000ca00000000",
            INIT_0B => X"000000a100000000000000aa00000000000000a800000000000000bc00000000",
            INIT_0C => X"0000008700000000000000ad0000000000000078000000000000007000000000",
            INIT_0D => X"00000073000000000000009b00000000000000ba000000000000009300000000",
            INIT_0E => X"000000bc00000000000000b20000000000000084000000000000006200000000",
            INIT_0F => X"000000ef00000000000000f300000000000000d400000000000000b900000000",
            INIT_10 => X"000000a100000000000000b300000000000000d600000000000000dd00000000",
            INIT_11 => X"000000b100000000000000b300000000000000b500000000000000af00000000",
            INIT_12 => X"000000dd00000000000000d400000000000000cf00000000000000bd00000000",
            INIT_13 => X"000000ab00000000000000b800000000000000c500000000000000dc00000000",
            INIT_14 => X"0000008c00000000000000950000000000000067000000000000008b00000000",
            INIT_15 => X"00000093000000000000009400000000000000b1000000000000009700000000",
            INIT_16 => X"0000009c000000000000008a0000000000000070000000000000008300000000",
            INIT_17 => X"000000ea00000000000000d900000000000000b1000000000000009700000000",
            INIT_18 => X"000000b200000000000000c600000000000000da00000000000000df00000000",
            INIT_19 => X"000000c800000000000000be00000000000000c200000000000000c200000000",
            INIT_1A => X"000000c700000000000000bf00000000000000b800000000000000ba00000000",
            INIT_1B => X"000000b100000000000000c800000000000000d000000000000000cb00000000",
            INIT_1C => X"0000009e000000000000007f000000000000008700000000000000ab00000000",
            INIT_1D => X"0000008f0000000000000083000000000000009b00000000000000a800000000",
            INIT_1E => X"0000009f0000000000000094000000000000007e000000000000008900000000",
            INIT_1F => X"000000c5000000000000009e0000000000000090000000000000009300000000",
            INIT_20 => X"000000b700000000000000d000000000000000dd00000000000000e100000000",
            INIT_21 => X"000000c200000000000000be00000000000000c700000000000000bf00000000",
            INIT_22 => X"000000ba00000000000000be00000000000000bc00000000000000c600000000",
            INIT_23 => X"000000bf00000000000000c600000000000000c100000000000000ab00000000",
            INIT_24 => X"000000a9000000000000009400000000000000bf00000000000000cf00000000",
            INIT_25 => X"0000008d000000000000007b000000000000008700000000000000a000000000",
            INIT_26 => X"00000098000000000000009f0000000000000095000000000000008e00000000",
            INIT_27 => X"0000009a000000000000008c0000000000000088000000000000008700000000",
            INIT_28 => X"000000be00000000000000d600000000000000dd00000000000000de00000000",
            INIT_29 => X"000000be00000000000000c800000000000000c300000000000000b300000000",
            INIT_2A => X"000000b200000000000000d100000000000000cd00000000000000c600000000",
            INIT_2B => X"000000b500000000000000b600000000000000b3000000000000009700000000",
            INIT_2C => X"000000a500000000000000ae00000000000000c400000000000000c500000000",
            INIT_2D => X"000000930000000000000089000000000000007c000000000000008600000000",
            INIT_2E => X"0000008b000000000000009900000000000000a1000000000000009900000000",
            INIT_2F => X"0000007d000000000000008b000000000000008b000000000000008300000000",
            INIT_30 => X"000000c600000000000000db00000000000000da00000000000000db00000000",
            INIT_31 => X"000000cf00000000000000d200000000000000bf00000000000000aa00000000",
            INIT_32 => X"000000b400000000000000cf00000000000000ce00000000000000cb00000000",
            INIT_33 => X"000000b000000000000000b400000000000000ae000000000000009c00000000",
            INIT_34 => X"0000009600000000000000b000000000000000b500000000000000b600000000",
            INIT_35 => X"000000980000000000000096000000000000007d000000000000006f00000000",
            INIT_36 => X"0000008a000000000000009a00000000000000a1000000000000009800000000",
            INIT_37 => X"0000006a00000000000000730000000000000080000000000000008a00000000",
            INIT_38 => X"000000cf00000000000000d900000000000000d600000000000000da00000000",
            INIT_39 => X"000000d500000000000000d200000000000000bc00000000000000aa00000000",
            INIT_3A => X"000000b600000000000000c700000000000000d300000000000000d400000000",
            INIT_3B => X"000000b500000000000000ba00000000000000ba00000000000000ae00000000",
            INIT_3C => X"0000008500000000000000ab00000000000000b600000000000000ba00000000",
            INIT_3D => X"00000095000000000000009a0000000000000089000000000000007200000000",
            INIT_3E => X"00000092000000000000009f00000000000000ab000000000000009400000000",
            INIT_3F => X"000000760000000000000073000000000000007b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000d400000000000000d400000000000000d800000000",
            INIT_41 => X"000000cd00000000000000cf00000000000000bd00000000000000b300000000",
            INIT_42 => X"0000008a00000000000000b100000000000000cd00000000000000cd00000000",
            INIT_43 => X"000000b600000000000000bb00000000000000c300000000000000a700000000",
            INIT_44 => X"00000082000000000000009e00000000000000b500000000000000b900000000",
            INIT_45 => X"0000008c0000000000000096000000000000008d000000000000007d00000000",
            INIT_46 => X"00000095000000000000009d00000000000000a3000000000000008d00000000",
            INIT_47 => X"0000007c00000000000000820000000000000083000000000000008500000000",
            INIT_48 => X"000000c800000000000000d000000000000000d200000000000000d700000000",
            INIT_49 => X"000000cc00000000000000ce00000000000000be00000000000000bb00000000",
            INIT_4A => X"00000050000000000000008300000000000000c400000000000000c600000000",
            INIT_4B => X"000000ae00000000000000b800000000000000c2000000000000009100000000",
            INIT_4C => X"00000083000000000000009300000000000000a500000000000000ae00000000",
            INIT_4D => X"00000088000000000000008f000000000000008b000000000000007800000000",
            INIT_4E => X"00000088000000000000008c000000000000008e000000000000008900000000",
            INIT_4F => X"0000007000000000000000790000000000000085000000000000008500000000",
            INIT_50 => X"000000c200000000000000cd00000000000000d000000000000000d700000000",
            INIT_51 => X"000000d100000000000000cd00000000000000b700000000000000b500000000",
            INIT_52 => X"00000051000000000000008100000000000000c200000000000000cc00000000",
            INIT_53 => X"000000a100000000000000ab00000000000000ba000000000000008e00000000",
            INIT_54 => X"000000780000000000000089000000000000009500000000000000a100000000",
            INIT_55 => X"0000007e00000000000000890000000000000087000000000000007300000000",
            INIT_56 => X"0000007a0000000000000070000000000000007b000000000000008500000000",
            INIT_57 => X"0000008000000000000000830000000000000088000000000000008a00000000",
            INIT_58 => X"000000bc00000000000000c800000000000000cd00000000000000d600000000",
            INIT_59 => X"000000d400000000000000c600000000000000af00000000000000b000000000",
            INIT_5A => X"0000008e00000000000000a000000000000000c000000000000000d000000000",
            INIT_5B => X"00000095000000000000009b00000000000000a800000000000000aa00000000",
            INIT_5C => X"00000064000000000000007f0000000000000085000000000000008d00000000",
            INIT_5D => X"0000007b00000000000000800000000000000083000000000000007100000000",
            INIT_5E => X"00000072000000000000006c0000000000000072000000000000007e00000000",
            INIT_5F => X"0000008900000000000000900000000000000090000000000000008200000000",
            INIT_60 => X"000000b700000000000000c000000000000000c400000000000000d200000000",
            INIT_61 => X"000000d200000000000000c000000000000000a600000000000000a900000000",
            INIT_62 => X"000000b400000000000000b600000000000000c000000000000000d100000000",
            INIT_63 => X"0000008c000000000000008d000000000000009900000000000000ab00000000",
            INIT_64 => X"0000005c000000000000006f000000000000007d000000000000008600000000",
            INIT_65 => X"0000007f000000000000007e000000000000007e000000000000007800000000",
            INIT_66 => X"0000007400000000000000690000000000000072000000000000007e00000000",
            INIT_67 => X"00000081000000000000008d0000000000000090000000000000008500000000",
            INIT_68 => X"000000b900000000000000b300000000000000b300000000000000c400000000",
            INIT_69 => X"000000cc00000000000000b5000000000000009700000000000000a600000000",
            INIT_6A => X"000000b300000000000000ba00000000000000c200000000000000cd00000000",
            INIT_6B => X"000000880000000000000085000000000000009200000000000000a600000000",
            INIT_6C => X"00000061000000000000005d0000000000000072000000000000007e00000000",
            INIT_6D => X"0000008000000000000000780000000000000073000000000000007800000000",
            INIT_6E => X"0000007e00000000000000710000000000000071000000000000008000000000",
            INIT_6F => X"0000007b00000000000000820000000000000083000000000000008400000000",
            INIT_70 => X"000000b800000000000000aa00000000000000a100000000000000b100000000",
            INIT_71 => X"000000c3000000000000009c000000000000008c00000000000000ae00000000",
            INIT_72 => X"000000b600000000000000bf00000000000000c100000000000000c900000000",
            INIT_73 => X"00000073000000000000006c0000000000000071000000000000009100000000",
            INIT_74 => X"0000006e0000000000000059000000000000006a000000000000007600000000",
            INIT_75 => X"0000008300000000000000780000000000000070000000000000007200000000",
            INIT_76 => X"0000007c000000000000007f000000000000007a000000000000007b00000000",
            INIT_77 => X"000000860000000000000082000000000000007a000000000000007500000000",
            INIT_78 => X"000000a10000000000000097000000000000008c000000000000009d00000000",
            INIT_79 => X"000000b10000000000000080000000000000008200000000000000a600000000",
            INIT_7A => X"0000009a00000000000000af00000000000000b700000000000000bf00000000",
            INIT_7B => X"0000005300000000000000470000000000000053000000000000007000000000",
            INIT_7C => X"0000006e0000000000000065000000000000005e000000000000006300000000",
            INIT_7D => X"0000007e0000000000000079000000000000006c000000000000006c00000000",
            INIT_7E => X"0000006b000000000000006f000000000000007a000000000000007900000000",
            INIT_7F => X"0000008400000000000000890000000000000084000000000000007300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "sampleifmap_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000280000000000000013000000000000001c000000000000001700000000",
            INIT_01 => X"00000074000000000000006d0000000000000073000000000000007100000000",
            INIT_02 => X"00000069000000000000006a0000000000000067000000000000007100000000",
            INIT_03 => X"0000006b00000000000000690000000000000069000000000000006900000000",
            INIT_04 => X"0000003a000000000000004c0000000000000063000000000000006a00000000",
            INIT_05 => X"0000008900000000000000720000000000000056000000000000005400000000",
            INIT_06 => X"0000007d000000000000007c000000000000007d000000000000007c00000000",
            INIT_07 => X"00000078000000000000007a000000000000007d000000000000007f00000000",
            INIT_08 => X"0000001a0000000000000014000000000000001b000000000000001800000000",
            INIT_09 => X"0000007c00000000000000760000000000000082000000000000006a00000000",
            INIT_0A => X"00000075000000000000006d0000000000000072000000000000007d00000000",
            INIT_0B => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_0C => X"00000044000000000000006a0000000000000083000000000000008500000000",
            INIT_0D => X"00000096000000000000008c0000000000000051000000000000003e00000000",
            INIT_0E => X"000000880000000000000089000000000000008c000000000000008a00000000",
            INIT_0F => X"0000008000000000000000810000000000000085000000000000008800000000",
            INIT_10 => X"000000120000000000000017000000000000001a000000000000001800000000",
            INIT_11 => X"0000007b00000000000000740000000000000083000000000000005800000000",
            INIT_12 => X"000000740000000000000074000000000000008d000000000000008b00000000",
            INIT_13 => X"00000084000000000000007d000000000000007f000000000000008100000000",
            INIT_14 => X"000000690000000000000098000000000000009a000000000000008e00000000",
            INIT_15 => X"0000009e000000000000009f0000000000000059000000000000003700000000",
            INIT_16 => X"0000008e00000000000000920000000000000097000000000000009700000000",
            INIT_17 => X"000000840000000000000088000000000000008b000000000000008e00000000",
            INIT_18 => X"0000001200000000000000190000000000000019000000000000001800000000",
            INIT_19 => X"00000073000000000000006a000000000000007c000000000000004500000000",
            INIT_1A => X"00000078000000000000009200000000000000a6000000000000009c00000000",
            INIT_1B => X"0000009700000000000000950000000000000094000000000000008900000000",
            INIT_1C => X"0000006d0000000000000094000000000000009c000000000000009600000000",
            INIT_1D => X"000000a900000000000000b1000000000000007a000000000000004a00000000",
            INIT_1E => X"000000950000000000000098000000000000009d00000000000000a100000000",
            INIT_1F => X"0000008e00000000000000910000000000000094000000000000009600000000",
            INIT_20 => X"0000001700000000000000190000000000000018000000000000001900000000",
            INIT_21 => X"000000680000000000000060000000000000006d000000000000003300000000",
            INIT_22 => X"0000008d00000000000000b200000000000000b800000000000000a100000000",
            INIT_23 => X"0000009300000000000000860000000000000080000000000000007c00000000",
            INIT_24 => X"0000006c00000000000000890000000000000096000000000000009700000000",
            INIT_25 => X"000000b500000000000000b70000000000000098000000000000006000000000",
            INIT_26 => X"000000a400000000000000a800000000000000ae00000000000000b300000000",
            INIT_27 => X"000000930000000000000098000000000000009c00000000000000a000000000",
            INIT_28 => X"0000001c000000000000001b000000000000001a000000000000001a00000000",
            INIT_29 => X"00000066000000000000005f0000000000000059000000000000002300000000",
            INIT_2A => X"0000009f00000000000000c700000000000000c1000000000000009600000000",
            INIT_2B => X"0000007600000000000000620000000000000066000000000000007400000000",
            INIT_2C => X"0000007a00000000000000770000000000000083000000000000008200000000",
            INIT_2D => X"000000aa00000000000000a600000000000000a7000000000000008400000000",
            INIT_2E => X"000000b700000000000000b300000000000000b700000000000000b200000000",
            INIT_2F => X"000000a900000000000000af00000000000000b100000000000000b700000000",
            INIT_30 => X"0000001a00000000000000190000000000000016000000000000001a00000000",
            INIT_31 => X"0000007b0000000000000080000000000000005c000000000000001d00000000",
            INIT_32 => X"000000ab00000000000000c700000000000000c3000000000000009300000000",
            INIT_33 => X"0000006a0000000000000063000000000000005e000000000000007e00000000",
            INIT_34 => X"0000007a0000000000000065000000000000006d000000000000006000000000",
            INIT_35 => X"000000b000000000000000aa00000000000000c000000000000000ac00000000",
            INIT_36 => X"000000ca00000000000000c500000000000000c400000000000000c300000000",
            INIT_37 => X"000000c200000000000000bf00000000000000bf00000000000000c500000000",
            INIT_38 => X"0000001900000000000000110000000000000021000000000000004d00000000",
            INIT_39 => X"0000007e000000000000009b000000000000009a000000000000005800000000",
            INIT_3A => X"000000b900000000000000c100000000000000be000000000000008c00000000",
            INIT_3B => X"00000071000000000000007b000000000000008100000000000000a300000000",
            INIT_3C => X"0000007900000000000000680000000000000067000000000000005800000000",
            INIT_3D => X"000000bd00000000000000a500000000000000c600000000000000b100000000",
            INIT_3E => X"000000da00000000000000e000000000000000db00000000000000e400000000",
            INIT_3F => X"000000cd00000000000000c400000000000000bb00000000000000ba00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006000000000000000560000000000000080000000000000009500000000",
            INIT_41 => X"00000077000000000000009900000000000000a7000000000000009b00000000",
            INIT_42 => X"000000bf00000000000000bf00000000000000a8000000000000006f00000000",
            INIT_43 => X"0000007f000000000000009400000000000000aa00000000000000b700000000",
            INIT_44 => X"0000007c00000000000000740000000000000070000000000000007000000000",
            INIT_45 => X"000000c100000000000000a200000000000000bb00000000000000a300000000",
            INIT_46 => X"000000bb00000000000000cf00000000000000d500000000000000df00000000",
            INIT_47 => X"000000d200000000000000c400000000000000a6000000000000009d00000000",
            INIT_48 => X"0000009b0000000000000092000000000000009e00000000000000a100000000",
            INIT_49 => X"00000075000000000000009f00000000000000a900000000000000a700000000",
            INIT_4A => X"000000b500000000000000b3000000000000009b000000000000006800000000",
            INIT_4B => X"00000087000000000000009f00000000000000b400000000000000b600000000",
            INIT_4C => X"0000007900000000000000750000000000000074000000000000006400000000",
            INIT_4D => X"000000cc00000000000000b200000000000000b2000000000000009e00000000",
            INIT_4E => X"000000a700000000000000cb00000000000000d600000000000000d800000000",
            INIT_4F => X"000000cf00000000000000b00000000000000096000000000000009300000000",
            INIT_50 => X"000000a5000000000000009e00000000000000a500000000000000aa00000000",
            INIT_51 => X"0000007000000000000000a000000000000000b000000000000000af00000000",
            INIT_52 => X"000000b400000000000000b100000000000000a4000000000000007b00000000",
            INIT_53 => X"00000079000000000000009500000000000000ac00000000000000b600000000",
            INIT_54 => X"0000007600000000000000750000000000000074000000000000006a00000000",
            INIT_55 => X"000000d100000000000000af00000000000000a6000000000000009c00000000",
            INIT_56 => X"000000a900000000000000cd00000000000000d800000000000000de00000000",
            INIT_57 => X"000000ba000000000000009f0000000000000093000000000000009100000000",
            INIT_58 => X"000000a600000000000000a900000000000000ae00000000000000ac00000000",
            INIT_59 => X"0000007a000000000000009d00000000000000b000000000000000b000000000",
            INIT_5A => X"000000b600000000000000b900000000000000b1000000000000008d00000000",
            INIT_5B => X"00000068000000000000007f000000000000009d00000000000000b600000000",
            INIT_5C => X"0000007d000000000000007b0000000000000084000000000000007300000000",
            INIT_5D => X"000000ce00000000000000a300000000000000a4000000000000009f00000000",
            INIT_5E => X"000000b500000000000000cd00000000000000d900000000000000e000000000",
            INIT_5F => X"0000009c0000000000000093000000000000008e000000000000009200000000",
            INIT_60 => X"000000a000000000000000a500000000000000a700000000000000a700000000",
            INIT_61 => X"0000008f000000000000009900000000000000a400000000000000a500000000",
            INIT_62 => X"000000a400000000000000ae00000000000000a3000000000000009100000000",
            INIT_63 => X"000000760000000000000085000000000000009f00000000000000a300000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008600000000",
            INIT_65 => X"000000cd00000000000000a800000000000000a300000000000000a300000000",
            INIT_66 => X"000000c700000000000000d600000000000000dc00000000000000df00000000",
            INIT_67 => X"000000980000000000000090000000000000009000000000000000a300000000",
            INIT_68 => X"0000009b00000000000000a000000000000000a200000000000000a900000000",
            INIT_69 => X"000000a40000000000000083000000000000008800000000000000a300000000",
            INIT_6A => X"0000008500000000000000840000000000000088000000000000009200000000",
            INIT_6B => X"000000920000000000000087000000000000009e000000000000009f00000000",
            INIT_6C => X"0000009e000000000000009000000000000000a200000000000000a700000000",
            INIT_6D => X"000000cb00000000000000b00000000000000098000000000000009800000000",
            INIT_6E => X"000000da00000000000000dd00000000000000d800000000000000d700000000",
            INIT_6F => X"000000b600000000000000a2000000000000009f00000000000000c500000000",
            INIT_70 => X"0000009d00000000000000a200000000000000a400000000000000ae00000000",
            INIT_71 => X"000000b2000000000000006d000000000000007800000000000000a800000000",
            INIT_72 => X"000000a300000000000000a100000000000000a700000000000000a600000000",
            INIT_73 => X"00000078000000000000008400000000000000ab00000000000000b600000000",
            INIT_74 => X"00000095000000000000008c00000000000000a300000000000000a900000000",
            INIT_75 => X"000000cc00000000000000aa00000000000000a400000000000000a600000000",
            INIT_76 => X"000000e400000000000000da00000000000000d500000000000000d300000000",
            INIT_77 => X"000000c700000000000000bb00000000000000b000000000000000d600000000",
            INIT_78 => X"0000009f00000000000000a100000000000000a000000000000000af00000000",
            INIT_79 => X"000000b70000000000000068000000000000008400000000000000aa00000000",
            INIT_7A => X"000000b000000000000000b800000000000000b600000000000000bc00000000",
            INIT_7B => X"0000008d00000000000000a300000000000000a800000000000000a200000000",
            INIT_7C => X"00000085000000000000009200000000000000a5000000000000009100000000",
            INIT_7D => X"000000a9000000000000009600000000000000a500000000000000af00000000",
            INIT_7E => X"000000dd00000000000000d900000000000000d400000000000000ca00000000",
            INIT_7F => X"000000c700000000000000c700000000000000ba00000000000000c400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "sampleifmap_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000940000000000000092000000000000009f00000000000000b300000000",
            INIT_01 => X"000000a8000000000000006d000000000000009700000000000000a100000000",
            INIT_02 => X"000000ae00000000000000a400000000000000b500000000000000c700000000",
            INIT_03 => X"000000a600000000000000aa000000000000009c00000000000000a500000000",
            INIT_04 => X"00000077000000000000009f0000000000000088000000000000006900000000",
            INIT_05 => X"00000050000000000000007e000000000000009e000000000000008f00000000",
            INIT_06 => X"000000cd00000000000000d100000000000000b7000000000000007600000000",
            INIT_07 => X"000000c500000000000000c900000000000000b700000000000000af00000000",
            INIT_08 => X"00000083000000000000008500000000000000a400000000000000b500000000",
            INIT_09 => X"0000009f000000000000009700000000000000a5000000000000009500000000",
            INIT_0A => X"000000cd00000000000000c400000000000000c700000000000000c200000000",
            INIT_0B => X"000000a200000000000000ac00000000000000a800000000000000b900000000",
            INIT_0C => X"00000077000000000000009b0000000000000069000000000000006800000000",
            INIT_0D => X"0000005c000000000000008800000000000000ad000000000000008600000000",
            INIT_0E => X"0000009e0000000000000098000000000000006f000000000000004b00000000",
            INIT_0F => X"000000c800000000000000cb00000000000000b0000000000000009800000000",
            INIT_10 => X"00000085000000000000008e00000000000000ac00000000000000b700000000",
            INIT_11 => X"000000aa00000000000000b100000000000000b0000000000000009f00000000",
            INIT_12 => X"000000d900000000000000cf00000000000000c500000000000000b100000000",
            INIT_13 => X"000000aa00000000000000bb00000000000000c600000000000000d900000000",
            INIT_14 => X"0000007e0000000000000085000000000000005a000000000000008300000000",
            INIT_15 => X"0000007e000000000000008200000000000000a2000000000000008b00000000",
            INIT_16 => X"0000008400000000000000760000000000000060000000000000006f00000000",
            INIT_17 => X"000000c700000000000000b80000000000000092000000000000007c00000000",
            INIT_18 => X"0000009500000000000000a100000000000000b000000000000000b900000000",
            INIT_19 => X"000000bc00000000000000b600000000000000b700000000000000af00000000",
            INIT_1A => X"000000c200000000000000b900000000000000aa00000000000000aa00000000",
            INIT_1B => X"000000af00000000000000ca00000000000000d000000000000000c900000000",
            INIT_1C => X"000000910000000000000071000000000000007b00000000000000a400000000",
            INIT_1D => X"0000007b0000000000000071000000000000008c000000000000009d00000000",
            INIT_1E => X"0000008e00000000000000860000000000000070000000000000007700000000",
            INIT_1F => X"000000a600000000000000840000000000000079000000000000007f00000000",
            INIT_20 => X"0000009b00000000000000ad00000000000000b700000000000000bd00000000",
            INIT_21 => X"000000b200000000000000b100000000000000ba00000000000000ab00000000",
            INIT_22 => X"000000b100000000000000b200000000000000ac00000000000000b400000000",
            INIT_23 => X"000000bd00000000000000c300000000000000bc00000000000000a400000000",
            INIT_24 => X"0000009d000000000000008800000000000000b600000000000000c900000000",
            INIT_25 => X"0000007c000000000000006a0000000000000078000000000000009300000000",
            INIT_26 => X"0000008a0000000000000094000000000000008a000000000000008000000000",
            INIT_27 => X"00000082000000000000007a0000000000000077000000000000007800000000",
            INIT_28 => X"000000a100000000000000b700000000000000bc00000000000000bd00000000",
            INIT_29 => X"000000b000000000000000bb00000000000000b7000000000000009e00000000",
            INIT_2A => X"000000a400000000000000c000000000000000bf00000000000000b800000000",
            INIT_2B => X"000000b100000000000000ad00000000000000a6000000000000008b00000000",
            INIT_2C => X"0000009600000000000000a200000000000000bc00000000000000c000000000",
            INIT_2D => X"000000850000000000000079000000000000006b000000000000007600000000",
            INIT_2E => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_2F => X"0000006c000000000000007d000000000000007c000000000000007500000000",
            INIT_30 => X"000000a600000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_31 => X"000000c500000000000000c700000000000000b4000000000000009400000000",
            INIT_32 => X"000000a800000000000000c000000000000000c300000000000000c100000000",
            INIT_33 => X"000000aa00000000000000a9000000000000009f000000000000009100000000",
            INIT_34 => X"0000008600000000000000a300000000000000ac00000000000000af00000000",
            INIT_35 => X"0000008b0000000000000086000000000000006c000000000000005d00000000",
            INIT_36 => X"0000007c000000000000008e0000000000000097000000000000008d00000000",
            INIT_37 => X"0000005b00000000000000650000000000000072000000000000007c00000000",
            INIT_38 => X"000000ac00000000000000b700000000000000b500000000000000ba00000000",
            INIT_39 => X"000000cf00000000000000c900000000000000b0000000000000008f00000000",
            INIT_3A => X"000000af00000000000000bd00000000000000cb00000000000000ce00000000",
            INIT_3B => X"000000ac00000000000000ae00000000000000ab00000000000000a500000000",
            INIT_3C => X"00000075000000000000009e00000000000000ab00000000000000b200000000",
            INIT_3D => X"00000088000000000000008a0000000000000078000000000000006100000000",
            INIT_3E => X"00000084000000000000009200000000000000a1000000000000008a00000000",
            INIT_3F => X"000000680000000000000064000000000000006d000000000000008200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a900000000000000af00000000000000b200000000000000b800000000",
            INIT_41 => X"000000ca00000000000000c600000000000000aa000000000000009200000000",
            INIT_42 => X"0000008800000000000000ab00000000000000c500000000000000c800000000",
            INIT_43 => X"000000aa00000000000000ab00000000000000b400000000000000a100000000",
            INIT_44 => X"00000073000000000000009000000000000000a800000000000000ad00000000",
            INIT_45 => X"0000007e0000000000000086000000000000007c000000000000006c00000000",
            INIT_46 => X"0000008700000000000000910000000000000099000000000000008200000000",
            INIT_47 => X"0000006f00000000000000740000000000000075000000000000007700000000",
            INIT_48 => X"0000009d00000000000000a800000000000000b000000000000000b800000000",
            INIT_49 => X"000000c800000000000000c000000000000000a2000000000000009300000000",
            INIT_4A => X"00000052000000000000008100000000000000b900000000000000bf00000000",
            INIT_4B => X"0000009f00000000000000a600000000000000b3000000000000008d00000000",
            INIT_4C => X"0000007400000000000000840000000000000096000000000000009f00000000",
            INIT_4D => X"0000007a000000000000007f000000000000007a000000000000006900000000",
            INIT_4E => X"0000007a00000000000000800000000000000084000000000000007f00000000",
            INIT_4F => X"00000062000000000000006b0000000000000077000000000000007700000000",
            INIT_50 => X"0000009400000000000000a300000000000000ac00000000000000b800000000",
            INIT_51 => X"000000ca00000000000000ba0000000000000092000000000000008600000000",
            INIT_52 => X"00000058000000000000008200000000000000b200000000000000c000000000",
            INIT_53 => X"00000090000000000000009800000000000000ac000000000000008c00000000",
            INIT_54 => X"00000069000000000000007a0000000000000084000000000000009100000000",
            INIT_55 => X"0000007000000000000000790000000000000077000000000000006400000000",
            INIT_56 => X"0000006c00000000000000640000000000000071000000000000007a00000000",
            INIT_57 => X"000000720000000000000075000000000000007a000000000000007c00000000",
            INIT_58 => X"0000008e000000000000009e00000000000000a900000000000000b700000000",
            INIT_59 => X"000000cc00000000000000b20000000000000084000000000000007e00000000",
            INIT_5A => X"00000090000000000000009d00000000000000af00000000000000c300000000",
            INIT_5B => X"000000830000000000000087000000000000009800000000000000a400000000",
            INIT_5C => X"00000054000000000000006f0000000000000074000000000000007c00000000",
            INIT_5D => X"0000006d00000000000000710000000000000073000000000000006100000000",
            INIT_5E => X"00000064000000000000005f0000000000000066000000000000007200000000",
            INIT_5F => X"0000007b00000000000000820000000000000082000000000000007400000000",
            INIT_60 => X"0000008e000000000000009900000000000000a100000000000000b100000000",
            INIT_61 => X"000000cc00000000000000b2000000000000007a000000000000007700000000",
            INIT_62 => X"000000a800000000000000aa00000000000000b400000000000000c500000000",
            INIT_63 => X"0000007b000000000000007a0000000000000087000000000000009d00000000",
            INIT_64 => X"0000004b000000000000005e000000000000006d000000000000007700000000",
            INIT_65 => X"000000710000000000000070000000000000006f000000000000006800000000",
            INIT_66 => X"00000066000000000000005c0000000000000064000000000000007000000000",
            INIT_67 => X"00000073000000000000007e0000000000000082000000000000007700000000",
            INIT_68 => X"00000091000000000000008d000000000000009000000000000000a300000000",
            INIT_69 => X"000000c800000000000000a9000000000000006b000000000000007400000000",
            INIT_6A => X"000000a300000000000000ac00000000000000b700000000000000c200000000",
            INIT_6B => X"0000007900000000000000730000000000000081000000000000009600000000",
            INIT_6C => X"00000051000000000000004e0000000000000064000000000000007000000000",
            INIT_6D => X"00000072000000000000006a0000000000000065000000000000006800000000",
            INIT_6E => X"0000007000000000000000630000000000000063000000000000007200000000",
            INIT_6F => X"0000006e00000000000000740000000000000075000000000000007600000000",
            INIT_70 => X"0000008f0000000000000083000000000000007e000000000000008e00000000",
            INIT_71 => X"000000c00000000000000091000000000000005f000000000000007c00000000",
            INIT_72 => X"000000a800000000000000b200000000000000b700000000000000be00000000",
            INIT_73 => X"00000065000000000000005c0000000000000062000000000000008200000000",
            INIT_74 => X"0000005f000000000000004b000000000000005c000000000000006800000000",
            INIT_75 => X"00000074000000000000006a0000000000000061000000000000006300000000",
            INIT_76 => X"0000006e0000000000000071000000000000006c000000000000006d00000000",
            INIT_77 => X"000000770000000000000074000000000000006c000000000000006700000000",
            INIT_78 => X"0000007800000000000000700000000000000068000000000000007b00000000",
            INIT_79 => X"000000ae00000000000000760000000000000057000000000000007400000000",
            INIT_7A => X"0000008d00000000000000a400000000000000ae00000000000000b500000000",
            INIT_7B => X"0000004600000000000000390000000000000045000000000000006300000000",
            INIT_7C => X"0000006000000000000000580000000000000051000000000000005700000000",
            INIT_7D => X"00000070000000000000006b000000000000005e000000000000005d00000000",
            INIT_7E => X"0000005d0000000000000061000000000000006c000000000000006b00000000",
            INIT_7F => X"00000076000000000000007b0000000000000076000000000000006500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "sampleifmap_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c700000000000000cd00000000000000d200000000000000d900000000",
            INIT_01 => X"000000bd00000000000000cf00000000000000d600000000000000da00000000",
            INIT_02 => X"000000a900000000000000a600000000000000ae00000000000000bb00000000",
            INIT_03 => X"0000008f000000000000008c000000000000009a000000000000009600000000",
            INIT_04 => X"000000df00000000000000db00000000000000bf00000000000000a700000000",
            INIT_05 => X"000000e100000000000000e200000000000000d700000000000000db00000000",
            INIT_06 => X"000000bb00000000000000af00000000000000be00000000000000db00000000",
            INIT_07 => X"000000a200000000000000a100000000000000aa00000000000000c800000000",
            INIT_08 => X"000000d700000000000000dc00000000000000dd00000000000000de00000000",
            INIT_09 => X"000000b300000000000000d300000000000000e100000000000000d800000000",
            INIT_0A => X"000000bc00000000000000be00000000000000c000000000000000b400000000",
            INIT_0B => X"000000db00000000000000d100000000000000ce00000000000000c700000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000eb00000000000000e500000000",
            INIT_0D => X"000000e500000000000000e100000000000000e200000000000000e900000000",
            INIT_0E => X"000000cd00000000000000d000000000000000d400000000000000e700000000",
            INIT_0F => X"000000c800000000000000ba00000000000000b700000000000000d800000000",
            INIT_10 => X"000000e800000000000000e700000000000000e900000000000000ea00000000",
            INIT_11 => X"000000ad00000000000000d900000000000000ef00000000000000e900000000",
            INIT_12 => X"000000b700000000000000ad00000000000000b400000000000000a400000000",
            INIT_13 => X"000000e000000000000000d400000000000000bc00000000000000be00000000",
            INIT_14 => X"000000e100000000000000e300000000000000eb00000000000000da00000000",
            INIT_15 => X"000000e100000000000000d600000000000000df00000000000000e500000000",
            INIT_16 => X"000000d800000000000000e600000000000000e800000000000000ea00000000",
            INIT_17 => X"000000d300000000000000d000000000000000ca00000000000000d100000000",
            INIT_18 => X"000000f200000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009e00000000000000e400000000000000f300000000000000f400000000",
            INIT_1A => X"0000009f0000000000000083000000000000009d000000000000009200000000",
            INIT_1B => X"0000009f00000000000000a20000000000000088000000000000009100000000",
            INIT_1C => X"000000d300000000000000c300000000000000cb00000000000000a900000000",
            INIT_1D => X"000000e200000000000000d000000000000000cb00000000000000d100000000",
            INIT_1E => X"000000d500000000000000e400000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e000000000000000db00000000000000c700000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000007500000000000000cf00000000000000f100000000000000f500000000",
            INIT_22 => X"0000006b0000000000000059000000000000006c000000000000006300000000",
            INIT_23 => X"0000005c0000000000000064000000000000005b000000000000006400000000",
            INIT_24 => X"00000095000000000000007c000000000000007c000000000000006600000000",
            INIT_25 => X"000000e900000000000000ca00000000000000b900000000000000b600000000",
            INIT_26 => X"000000cd00000000000000e300000000000000e200000000000000e100000000",
            INIT_27 => X"000000de00000000000000e200000000000000d500000000000000c200000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007e00000000000000d800000000000000ed00000000000000f500000000",
            INIT_2A => X"00000066000000000000005b000000000000005a000000000000004800000000",
            INIT_2B => X"00000063000000000000006b0000000000000067000000000000006500000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005900000000",
            INIT_2D => X"000000eb00000000000000d800000000000000be000000000000007e00000000",
            INIT_2E => X"000000c400000000000000d800000000000000df00000000000000e700000000",
            INIT_2F => X"000000ec00000000000000d900000000000000bd00000000000000ae00000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009e00000000000000d900000000000000db00000000000000f100000000",
            INIT_32 => X"0000009700000000000000840000000000000072000000000000005000000000",
            INIT_33 => X"0000008a000000000000008f0000000000000084000000000000008c00000000",
            INIT_34 => X"000000780000000000000072000000000000007a000000000000008200000000",
            INIT_35 => X"000000e900000000000000dd000000000000009b000000000000006e00000000",
            INIT_36 => X"000000c000000000000000c600000000000000e000000000000000eb00000000",
            INIT_37 => X"000000eb00000000000000cc00000000000000ab00000000000000a700000000",
            INIT_38 => X"000000f600000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009900000000000000d700000000000000c700000000000000e300000000",
            INIT_3A => X"000000ca00000000000000bb0000000000000092000000000000005100000000",
            INIT_3B => X"000000830000000000000083000000000000009e00000000000000cf00000000",
            INIT_3C => X"000000840000000000000083000000000000008d000000000000008100000000",
            INIT_3D => X"000000d7000000000000009f0000000000000084000000000000009f00000000",
            INIT_3E => X"000000d100000000000000d400000000000000d700000000000000e500000000",
            INIT_3F => X"000000dd00000000000000b200000000000000ab00000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000008200000000000000da00000000000000ce00000000000000e300000000",
            INIT_42 => X"0000008100000000000000800000000000000082000000000000005100000000",
            INIT_43 => X"0000007d0000000000000074000000000000009100000000000000b800000000",
            INIT_44 => X"0000007d000000000000008e0000000000000089000000000000007c00000000",
            INIT_45 => X"000000c600000000000000900000000000000093000000000000009900000000",
            INIT_46 => X"000000dc00000000000000e900000000000000db00000000000000d600000000",
            INIT_47 => X"000000c900000000000000a900000000000000a400000000000000b800000000",
            INIT_48 => X"000000f200000000000000f400000000000000f300000000000000f300000000",
            INIT_49 => X"0000006e00000000000000a800000000000000be00000000000000e400000000",
            INIT_4A => X"0000006e00000000000000770000000000000086000000000000005300000000",
            INIT_4B => X"0000007800000000000000730000000000000080000000000000008f00000000",
            INIT_4C => X"0000007d00000000000000920000000000000083000000000000007d00000000",
            INIT_4D => X"000000c4000000000000008c000000000000009b000000000000009500000000",
            INIT_4E => X"000000e900000000000000f000000000000000f000000000000000e900000000",
            INIT_4F => X"000000dc00000000000000d700000000000000c800000000000000c800000000",
            INIT_50 => X"000000f500000000000000f400000000000000f100000000000000ef00000000",
            INIT_51 => X"0000005f0000000000000082000000000000008500000000000000dc00000000",
            INIT_52 => X"0000006c00000000000000740000000000000074000000000000004e00000000",
            INIT_53 => X"0000006c000000000000006d000000000000006b000000000000006d00000000",
            INIT_54 => X"0000007300000000000000780000000000000078000000000000007300000000",
            INIT_55 => X"000000a7000000000000008f0000000000000096000000000000008800000000",
            INIT_56 => X"000000f300000000000000f500000000000000e400000000000000d000000000",
            INIT_57 => X"000000f400000000000000f500000000000000f500000000000000f400000000",
            INIT_58 => X"000000f400000000000000f200000000000000e900000000000000de00000000",
            INIT_59 => X"0000005900000000000000a500000000000000a900000000000000d800000000",
            INIT_5A => X"00000064000000000000005b0000000000000043000000000000003d00000000",
            INIT_5B => X"000000600000000000000062000000000000005f000000000000005f00000000",
            INIT_5C => X"00000061000000000000005a000000000000005f000000000000006000000000",
            INIT_5D => X"0000007e00000000000000810000000000000079000000000000006900000000",
            INIT_5E => X"000000f300000000000000f800000000000000d8000000000000009b00000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e300000000000000ec00000000000000df00000000000000d000000000",
            INIT_61 => X"0000006400000000000000b500000000000000b700000000000000bf00000000",
            INIT_62 => X"0000006500000000000000580000000000000038000000000000003700000000",
            INIT_63 => X"0000005400000000000000560000000000000063000000000000006f00000000",
            INIT_64 => X"00000071000000000000005d0000000000000054000000000000005200000000",
            INIT_65 => X"0000008100000000000000700000000000000062000000000000006d00000000",
            INIT_66 => X"000000f400000000000000f500000000000000e200000000000000ae00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c300000000000000db00000000000000cc00000000000000c800000000",
            INIT_69 => X"00000066000000000000009c000000000000009a00000000000000aa00000000",
            INIT_6A => X"00000066000000000000006c0000000000000063000000000000006800000000",
            INIT_6B => X"00000055000000000000005e0000000000000075000000000000007300000000",
            INIT_6C => X"0000008c000000000000007a000000000000006a000000000000005a00000000",
            INIT_6D => X"0000007c000000000000006c0000000000000068000000000000008000000000",
            INIT_6E => X"000000d400000000000000c300000000000000b3000000000000009600000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a900000000000000cf00000000000000d200000000000000c800000000",
            INIT_71 => X"0000008a0000000000000093000000000000009400000000000000a400000000",
            INIT_72 => X"0000005d000000000000006a000000000000005c000000000000008100000000",
            INIT_73 => X"0000004d0000000000000054000000000000005d000000000000005900000000",
            INIT_74 => X"0000005100000000000000510000000000000051000000000000004c00000000",
            INIT_75 => X"00000052000000000000004b000000000000004a000000000000004f00000000",
            INIT_76 => X"0000008f000000000000008c000000000000007b000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bf00000000",
            INIT_78 => X"0000007700000000000000c400000000000000e200000000000000d200000000",
            INIT_79 => X"000000c000000000000000ba0000000000000096000000000000007000000000",
            INIT_7A => X"00000037000000000000004d000000000000004d000000000000006c00000000",
            INIT_7B => X"0000003f000000000000003c000000000000002f000000000000002d00000000",
            INIT_7C => X"00000036000000000000003b000000000000003f000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000032000000000000003100000000",
            INIT_7E => X"00000067000000000000005b000000000000004b000000000000004700000000",
            INIT_7F => X"000000f400000000000000f600000000000000e1000000000000008700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "sampleifmap_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006000000000000000b400000000000000c100000000000000c700000000",
            INIT_01 => X"000000a100000000000000c00000000000000091000000000000005d00000000",
            INIT_02 => X"00000062000000000000005c0000000000000049000000000000005600000000",
            INIT_03 => X"00000047000000000000004f000000000000004f000000000000006800000000",
            INIT_04 => X"0000001b000000000000001e000000000000001c000000000000002500000000",
            INIT_05 => X"0000001c00000000000000160000000000000032000000000000003400000000",
            INIT_06 => X"00000068000000000000005b0000000000000035000000000000001800000000",
            INIT_07 => X"000000f300000000000000f700000000000000ce000000000000008000000000",
            INIT_08 => X"0000007100000000000000c200000000000000c700000000000000d300000000",
            INIT_09 => X"00000047000000000000009f000000000000009d000000000000007800000000",
            INIT_0A => X"0000007c0000000000000074000000000000005a000000000000004400000000",
            INIT_0B => X"0000006600000000000000800000000000000079000000000000009500000000",
            INIT_0C => X"0000006400000000000000700000000000000062000000000000004e00000000",
            INIT_0D => X"00000063000000000000005c0000000000000093000000000000009400000000",
            INIT_0E => X"0000008e0000000000000087000000000000006c000000000000005e00000000",
            INIT_0F => X"000000f500000000000000f200000000000000b7000000000000009c00000000",
            INIT_10 => X"0000006600000000000000b700000000000000ca00000000000000dc00000000",
            INIT_11 => X"0000001e000000000000008400000000000000a5000000000000006e00000000",
            INIT_12 => X"00000053000000000000006b0000000000000062000000000000003900000000",
            INIT_13 => X"0000006400000000000000810000000000000065000000000000005200000000",
            INIT_14 => X"0000009f000000000000009e00000000000000ae000000000000009900000000",
            INIT_15 => X"000000a300000000000000a200000000000000a800000000000000ac00000000",
            INIT_16 => X"00000077000000000000009c00000000000000af00000000000000a000000000",
            INIT_17 => X"000000f700000000000000e40000000000000087000000000000007200000000",
            INIT_18 => X"0000006200000000000000bc00000000000000cf00000000000000db00000000",
            INIT_19 => X"0000002a000000000000006f000000000000008d000000000000005300000000",
            INIT_1A => X"0000003e000000000000004c0000000000000048000000000000003a00000000",
            INIT_1B => X"0000005d00000000000000400000000000000038000000000000003500000000",
            INIT_1C => X"00000065000000000000005b000000000000007c00000000000000a000000000",
            INIT_1D => X"000000670000000000000067000000000000006b000000000000007400000000",
            INIT_1E => X"00000043000000000000007e000000000000009b000000000000006300000000",
            INIT_1F => X"000000f800000000000000d90000000000000076000000000000005100000000",
            INIT_20 => X"0000006500000000000000c700000000000000d200000000000000d900000000",
            INIT_21 => X"0000003c000000000000005d0000000000000058000000000000003800000000",
            INIT_22 => X"00000046000000000000003f000000000000002e000000000000003800000000",
            INIT_23 => X"0000004100000000000000400000000000000036000000000000003c00000000",
            INIT_24 => X"0000006700000000000000690000000000000072000000000000006300000000",
            INIT_25 => X"00000061000000000000005d0000000000000060000000000000006400000000",
            INIT_26 => X"000000490000000000000064000000000000006f000000000000006600000000",
            INIT_27 => X"000000f900000000000000d40000000000000072000000000000005200000000",
            INIT_28 => X"0000007500000000000000ca00000000000000cd00000000000000d100000000",
            INIT_29 => X"0000004400000000000000510000000000000046000000000000005300000000",
            INIT_2A => X"00000033000000000000002b0000000000000023000000000000003200000000",
            INIT_2B => X"0000003f0000000000000057000000000000004d000000000000004400000000",
            INIT_2C => X"0000004800000000000000520000000000000047000000000000003400000000",
            INIT_2D => X"0000005d000000000000003e0000000000000043000000000000004000000000",
            INIT_2E => X"0000006c0000000000000053000000000000003c000000000000005800000000",
            INIT_2F => X"000000fa00000000000000cc000000000000006c000000000000007000000000",
            INIT_30 => X"0000006800000000000000c500000000000000ca00000000000000cd00000000",
            INIT_31 => X"000000490000000000000047000000000000006f000000000000005d00000000",
            INIT_32 => X"0000002200000000000000260000000000000029000000000000003f00000000",
            INIT_33 => X"0000004f000000000000008e0000000000000063000000000000004b00000000",
            INIT_34 => X"0000007600000000000000930000000000000056000000000000001e00000000",
            INIT_35 => X"0000009900000000000000660000000000000072000000000000006300000000",
            INIT_36 => X"0000008d000000000000004a000000000000003f00000000000000b200000000",
            INIT_37 => X"000000f600000000000000c3000000000000005a000000000000007700000000",
            INIT_38 => X"0000005700000000000000b900000000000000c200000000000000c600000000",
            INIT_39 => X"000000630000000000000061000000000000006c000000000000003100000000",
            INIT_3A => X"0000002400000000000000270000000000000033000000000000005f00000000",
            INIT_3B => X"0000003700000000000000570000000000000032000000000000002800000000",
            INIT_3C => X"0000007f0000000000000097000000000000004f000000000000002000000000",
            INIT_3D => X"0000009c00000000000000740000000000000088000000000000007a00000000",
            INIT_3E => X"0000004a00000000000000350000000000000037000000000000009f00000000",
            INIT_3F => X"000000f000000000000000c2000000000000004e000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d00000000000000a900000000000000b400000000000000b600000000",
            INIT_41 => X"00000090000000000000006c000000000000003b000000000000002500000000",
            INIT_42 => X"00000020000000000000002b000000000000003c000000000000006a00000000",
            INIT_43 => X"00000021000000000000001e000000000000001c000000000000001d00000000",
            INIT_44 => X"00000058000000000000003a000000000000002a000000000000002700000000",
            INIT_45 => X"00000075000000000000007a0000000000000079000000000000006a00000000",
            INIT_46 => X"000000320000000000000033000000000000002f000000000000004300000000",
            INIT_47 => X"000000e100000000000000ba0000000000000050000000000000003300000000",
            INIT_48 => X"0000007d00000000000000a400000000000000a500000000000000a800000000",
            INIT_49 => X"0000008d000000000000006f0000000000000060000000000000005b00000000",
            INIT_4A => X"000000240000000000000037000000000000004a000000000000006000000000",
            INIT_4B => X"0000001f000000000000001d000000000000001e000000000000001e00000000",
            INIT_4C => X"000000ae00000000000000400000000000000018000000000000002300000000",
            INIT_4D => X"000000b500000000000000b300000000000000cb00000000000000cd00000000",
            INIT_4E => X"00000030000000000000002b0000000000000026000000000000005700000000",
            INIT_4F => X"000000d300000000000000ae000000000000005b000000000000004200000000",
            INIT_50 => X"000000b400000000000000af00000000000000a300000000000000a200000000",
            INIT_51 => X"0000008d000000000000006c0000000000000076000000000000009800000000",
            INIT_52 => X"00000030000000000000004e0000000000000053000000000000005b00000000",
            INIT_53 => X"0000001d00000000000000190000000000000018000000000000001900000000",
            INIT_54 => X"000000a400000000000000470000000000000026000000000000002700000000",
            INIT_55 => X"000000a600000000000000a900000000000000b100000000000000b800000000",
            INIT_56 => X"00000031000000000000001e000000000000001e000000000000005100000000",
            INIT_57 => X"000000ce00000000000000a9000000000000005f000000000000004e00000000",
            INIT_58 => X"000000a600000000000000b300000000000000ac000000000000009a00000000",
            INIT_59 => X"0000009200000000000000670000000000000075000000000000009200000000",
            INIT_5A => X"0000003600000000000000520000000000000055000000000000005700000000",
            INIT_5B => X"000000250000000000000021000000000000001e000000000000002000000000",
            INIT_5C => X"000000650000000000000056000000000000004d000000000000003600000000",
            INIT_5D => X"00000089000000000000008e0000000000000079000000000000006b00000000",
            INIT_5E => X"000000360000000000000021000000000000001e000000000000003c00000000",
            INIT_5F => X"000000c700000000000000a5000000000000005b000000000000004e00000000",
            INIT_60 => X"00000094000000000000009e00000000000000a900000000000000a600000000",
            INIT_61 => X"0000007100000000000000670000000000000085000000000000008f00000000",
            INIT_62 => X"0000003c000000000000004b0000000000000051000000000000004f00000000",
            INIT_63 => X"0000002c000000000000002a0000000000000027000000000000002a00000000",
            INIT_64 => X"0000004d00000000000000410000000000000036000000000000003000000000",
            INIT_65 => X"0000008b0000000000000083000000000000006e000000000000005a00000000",
            INIT_66 => X"000000360000000000000026000000000000001d000000000000003500000000",
            INIT_67 => X"000000c400000000000000a9000000000000005b000000000000004600000000",
            INIT_68 => X"0000008d0000000000000093000000000000009700000000000000a200000000",
            INIT_69 => X"0000004e000000000000006b0000000000000085000000000000008900000000",
            INIT_6A => X"0000003c0000000000000046000000000000004e000000000000004800000000",
            INIT_6B => X"00000030000000000000002e000000000000002a000000000000003200000000",
            INIT_6C => X"00000042000000000000003b0000000000000033000000000000003100000000",
            INIT_6D => X"0000007100000000000000650000000000000059000000000000004c00000000",
            INIT_6E => X"000000340000000000000023000000000000001d000000000000004500000000",
            INIT_6F => X"000000ba00000000000000ae0000000000000062000000000000003f00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009400000000",
            INIT_71 => X"0000003c000000000000006a000000000000008c000000000000008f00000000",
            INIT_72 => X"000000370000000000000042000000000000004a000000000000004200000000",
            INIT_73 => X"0000003a00000000000000360000000000000034000000000000003900000000",
            INIT_74 => X"000000460000000000000041000000000000003a000000000000003a00000000",
            INIT_75 => X"0000005d00000000000000570000000000000050000000000000004900000000",
            INIT_76 => X"0000003700000000000000260000000000000025000000000000004d00000000",
            INIT_77 => X"000000b400000000000000b30000000000000083000000000000004a00000000",
            INIT_78 => X"000000a200000000000000a00000000000000095000000000000009000000000",
            INIT_79 => X"0000003d000000000000007e0000000000000092000000000000009e00000000",
            INIT_7A => X"00000043000000000000003a0000000000000039000000000000003900000000",
            INIT_7B => X"0000004800000000000000490000000000000045000000000000004600000000",
            INIT_7C => X"0000006200000000000000590000000000000049000000000000004400000000",
            INIT_7D => X"0000006100000000000000630000000000000061000000000000005e00000000",
            INIT_7E => X"0000004700000000000000400000000000000045000000000000005200000000",
            INIT_7F => X"000000ba00000000000000b600000000000000a4000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "sampleifmap_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ca00000000000000d000000000000000d000000000000000d700000000",
            INIT_01 => X"000000b900000000000000ca00000000000000d100000000000000d700000000",
            INIT_02 => X"000000a0000000000000009800000000000000a800000000000000b800000000",
            INIT_03 => X"0000009d000000000000009a00000000000000a7000000000000009d00000000",
            INIT_04 => X"000000e100000000000000e100000000000000cb00000000000000b500000000",
            INIT_05 => X"000000e400000000000000e500000000000000db00000000000000de00000000",
            INIT_06 => X"000000c400000000000000b800000000000000c500000000000000dd00000000",
            INIT_07 => X"000000a500000000000000b000000000000000b800000000000000d000000000",
            INIT_08 => X"000000d900000000000000e100000000000000e000000000000000e200000000",
            INIT_09 => X"000000ab00000000000000cc00000000000000dd00000000000000d500000000",
            INIT_0A => X"000000b100000000000000b200000000000000bd00000000000000b400000000",
            INIT_0B => X"000000e000000000000000d000000000000000cd00000000000000c400000000",
            INIT_0C => X"000000f300000000000000f200000000000000f000000000000000ec00000000",
            INIT_0D => X"000000e700000000000000e400000000000000e500000000000000ee00000000",
            INIT_0E => X"000000d200000000000000d400000000000000d600000000000000e700000000",
            INIT_0F => X"000000c500000000000000bf00000000000000be00000000000000de00000000",
            INIT_10 => X"000000eb00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_11 => X"000000a600000000000000d600000000000000ef00000000000000ea00000000",
            INIT_12 => X"000000b100000000000000a800000000000000b100000000000000a600000000",
            INIT_13 => X"000000df00000000000000ce00000000000000b700000000000000b800000000",
            INIT_14 => X"000000e800000000000000e300000000000000ec00000000000000dc00000000",
            INIT_15 => X"000000e000000000000000d900000000000000e400000000000000eb00000000",
            INIT_16 => X"000000dd00000000000000e600000000000000e900000000000000e900000000",
            INIT_17 => X"000000d200000000000000d100000000000000ce00000000000000d900000000",
            INIT_18 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009900000000000000e300000000000000f400000000000000f400000000",
            INIT_1A => X"0000009f0000000000000082000000000000009b000000000000009200000000",
            INIT_1B => X"000000a000000000000000a2000000000000008a000000000000009000000000",
            INIT_1C => X"000000dc00000000000000c200000000000000cd00000000000000ac00000000",
            INIT_1D => X"000000e000000000000000d300000000000000d300000000000000de00000000",
            INIT_1E => X"000000db00000000000000e500000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e200000000000000df00000000000000cf00000000",
            INIT_20 => X"000000f400000000000000f400000000000000f400000000000000f500000000",
            INIT_21 => X"0000007000000000000000cd00000000000000f000000000000000f500000000",
            INIT_22 => X"0000006d000000000000005b000000000000006d000000000000006200000000",
            INIT_23 => X"0000005c0000000000000064000000000000005c000000000000006500000000",
            INIT_24 => X"0000009a000000000000007c000000000000007d000000000000006800000000",
            INIT_25 => X"000000e300000000000000c900000000000000c200000000000000c200000000",
            INIT_26 => X"000000d300000000000000e300000000000000de00000000000000dc00000000",
            INIT_27 => X"000000e100000000000000e800000000000000dc00000000000000cb00000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007b00000000000000d400000000000000eb00000000000000f600000000",
            INIT_2A => X"00000069000000000000005f000000000000005d000000000000004700000000",
            INIT_2B => X"00000066000000000000006e000000000000006a000000000000006700000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005b00000000",
            INIT_2D => X"000000e600000000000000d900000000000000c5000000000000008100000000",
            INIT_2E => X"000000c600000000000000d600000000000000da00000000000000dd00000000",
            INIT_2F => X"000000ed00000000000000e200000000000000c500000000000000b400000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009c00000000000000d500000000000000d600000000000000f000000000",
            INIT_32 => X"0000009a00000000000000890000000000000077000000000000004f00000000",
            INIT_33 => X"00000096000000000000009b000000000000008b000000000000009000000000",
            INIT_34 => X"0000007e00000000000000790000000000000080000000000000008e00000000",
            INIT_35 => X"000000e900000000000000e100000000000000a0000000000000007200000000",
            INIT_36 => X"000000ba00000000000000c000000000000000da00000000000000e900000000",
            INIT_37 => X"000000ec00000000000000d400000000000000b000000000000000a500000000",
            INIT_38 => X"000000f700000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009600000000000000d300000000000000c100000000000000e200000000",
            INIT_3A => X"000000c800000000000000bc0000000000000098000000000000005100000000",
            INIT_3B => X"00000090000000000000008d00000000000000a500000000000000cd00000000",
            INIT_3C => X"0000008f000000000000008d0000000000000096000000000000008e00000000",
            INIT_3D => X"000000d600000000000000a3000000000000008c00000000000000a700000000",
            INIT_3E => X"000000d200000000000000d300000000000000d100000000000000e000000000",
            INIT_3F => X"000000dc00000000000000af00000000000000ae00000000000000c700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000007f00000000000000d800000000000000ca00000000000000e100000000",
            INIT_42 => X"0000008700000000000000840000000000000086000000000000005100000000",
            INIT_43 => X"00000087000000000000007c000000000000009700000000000000b900000000",
            INIT_44 => X"0000008800000000000000960000000000000091000000000000008600000000",
            INIT_45 => X"000000c0000000000000008e000000000000009e00000000000000a400000000",
            INIT_46 => X"000000d700000000000000e700000000000000d800000000000000cf00000000",
            INIT_47 => X"000000c4000000000000009c000000000000009e00000000000000b100000000",
            INIT_48 => X"000000f200000000000000f400000000000000f200000000000000f200000000",
            INIT_49 => X"0000006e00000000000000a800000000000000bd00000000000000e300000000",
            INIT_4A => X"000000760000000000000080000000000000008c000000000000005300000000",
            INIT_4B => X"00000081000000000000007c0000000000000087000000000000009300000000",
            INIT_4C => X"000000860000000000000097000000000000008b000000000000008500000000",
            INIT_4D => X"000000c1000000000000009100000000000000a4000000000000009e00000000",
            INIT_4E => X"000000e600000000000000ef00000000000000ef00000000000000e500000000",
            INIT_4F => X"000000d700000000000000cc00000000000000be00000000000000c100000000",
            INIT_50 => X"000000f400000000000000f300000000000000ef00000000000000e800000000",
            INIT_51 => X"0000005e0000000000000080000000000000008100000000000000da00000000",
            INIT_52 => X"00000070000000000000007a000000000000007a000000000000004f00000000",
            INIT_53 => X"0000007300000000000000730000000000000070000000000000007100000000",
            INIT_54 => X"0000007e000000000000007f0000000000000080000000000000007c00000000",
            INIT_55 => X"000000aa0000000000000099000000000000009e000000000000009000000000",
            INIT_56 => X"000000f400000000000000f600000000000000e300000000000000ce00000000",
            INIT_57 => X"000000f400000000000000f500000000000000f300000000000000f300000000",
            INIT_58 => X"000000f200000000000000f200000000000000e300000000000000cd00000000",
            INIT_59 => X"00000058000000000000009f00000000000000a100000000000000d300000000",
            INIT_5A => X"00000066000000000000005e0000000000000045000000000000003c00000000",
            INIT_5B => X"0000006600000000000000670000000000000061000000000000006200000000",
            INIT_5C => X"00000067000000000000005f0000000000000064000000000000006800000000",
            INIT_5D => X"000000800000000000000089000000000000007f000000000000007100000000",
            INIT_5E => X"000000f300000000000000f800000000000000d7000000000000009900000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000dc00000000000000e400000000000000d500000000000000bc00000000",
            INIT_61 => X"0000006300000000000000ad00000000000000aa00000000000000b400000000",
            INIT_62 => X"00000066000000000000005a0000000000000039000000000000003700000000",
            INIT_63 => X"0000005500000000000000580000000000000067000000000000007200000000",
            INIT_64 => X"00000073000000000000005d0000000000000055000000000000005500000000",
            INIT_65 => X"0000008600000000000000760000000000000065000000000000007000000000",
            INIT_66 => X"000000f400000000000000f500000000000000e100000000000000b000000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000b500000000000000ca00000000000000bc00000000000000b800000000",
            INIT_69 => X"00000063000000000000008d0000000000000086000000000000009800000000",
            INIT_6A => X"00000067000000000000006f0000000000000066000000000000006700000000",
            INIT_6B => X"0000005600000000000000600000000000000078000000000000007600000000",
            INIT_6C => X"00000092000000000000007d000000000000006b000000000000005c00000000",
            INIT_6D => X"0000007f000000000000006e000000000000006a000000000000008400000000",
            INIT_6E => X"000000d200000000000000c300000000000000b3000000000000009800000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ee00000000",
            INIT_70 => X"0000009800000000000000bd00000000000000c200000000000000b600000000",
            INIT_71 => X"0000007e000000000000007f000000000000007b000000000000009200000000",
            INIT_72 => X"0000005e0000000000000069000000000000005d000000000000007c00000000",
            INIT_73 => X"0000004f0000000000000055000000000000005d000000000000005a00000000",
            INIT_74 => X"0000005500000000000000540000000000000053000000000000004e00000000",
            INIT_75 => X"00000053000000000000004c000000000000004b000000000000005100000000",
            INIT_76 => X"0000008a000000000000008a000000000000007a000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bc00000000",
            INIT_78 => X"0000006500000000000000a700000000000000cc00000000000000bd00000000",
            INIT_79 => X"000000ae00000000000000a9000000000000007d000000000000006500000000",
            INIT_7A => X"00000036000000000000004f000000000000004d000000000000006700000000",
            INIT_7B => X"0000003e000000000000003b000000000000002f000000000000002b00000000",
            INIT_7C => X"000000340000000000000039000000000000003e000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000030000000000000002f00000000",
            INIT_7E => X"00000061000000000000005a000000000000004a000000000000004600000000",
            INIT_7F => X"000000f400000000000000f600000000000000df000000000000008000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "sampleifmap_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000054000000000000009700000000000000a400000000000000ae00000000",
            INIT_01 => X"0000009200000000000000ac000000000000007c000000000000005200000000",
            INIT_02 => X"0000005a00000000000000570000000000000049000000000000005300000000",
            INIT_03 => X"00000044000000000000004c000000000000004b000000000000006400000000",
            INIT_04 => X"00000017000000000000001a0000000000000017000000000000002100000000",
            INIT_05 => X"000000190000000000000014000000000000002f000000000000003000000000",
            INIT_06 => X"0000006400000000000000560000000000000032000000000000001500000000",
            INIT_07 => X"000000f300000000000000f700000000000000ca000000000000007800000000",
            INIT_08 => X"0000006800000000000000b300000000000000b400000000000000c000000000",
            INIT_09 => X"00000040000000000000008e0000000000000087000000000000006800000000",
            INIT_0A => X"00000078000000000000006c0000000000000057000000000000004100000000",
            INIT_0B => X"00000062000000000000007d0000000000000076000000000000009500000000",
            INIT_0C => X"00000060000000000000006a0000000000000059000000000000004600000000",
            INIT_0D => X"0000006000000000000000590000000000000090000000000000009000000000",
            INIT_0E => X"0000008b00000000000000820000000000000067000000000000005a00000000",
            INIT_0F => X"000000f400000000000000f100000000000000b2000000000000009700000000",
            INIT_10 => X"0000005e00000000000000ab00000000000000bd00000000000000d100000000",
            INIT_11 => X"0000001c00000000000000760000000000000092000000000000006200000000",
            INIT_12 => X"0000004f0000000000000067000000000000005f000000000000003600000000",
            INIT_13 => X"0000005f00000000000000800000000000000064000000000000005300000000",
            INIT_14 => X"0000009e000000000000009b00000000000000aa000000000000009200000000",
            INIT_15 => X"000000a100000000000000a000000000000000a800000000000000ab00000000",
            INIT_16 => X"00000077000000000000009b00000000000000ac000000000000009e00000000",
            INIT_17 => X"000000f700000000000000e20000000000000080000000000000006f00000000",
            INIT_18 => X"0000005b00000000000000b000000000000000c100000000000000d000000000",
            INIT_19 => X"000000280000000000000064000000000000007f000000000000004c00000000",
            INIT_1A => X"0000003900000000000000490000000000000044000000000000003500000000",
            INIT_1B => X"00000059000000000000003d0000000000000035000000000000003200000000",
            INIT_1C => X"0000006200000000000000570000000000000077000000000000009c00000000",
            INIT_1D => X"0000006400000000000000630000000000000068000000000000007100000000",
            INIT_1E => X"0000003f000000000000007a0000000000000098000000000000006000000000",
            INIT_1F => X"000000f800000000000000d60000000000000070000000000000004d00000000",
            INIT_20 => X"0000005f00000000000000be00000000000000c300000000000000ca00000000",
            INIT_21 => X"000000380000000000000053000000000000004e000000000000003300000000",
            INIT_22 => X"00000044000000000000003c0000000000000027000000000000003300000000",
            INIT_23 => X"0000003d000000000000003b0000000000000033000000000000003900000000",
            INIT_24 => X"000000650000000000000066000000000000006e000000000000005f00000000",
            INIT_25 => X"00000060000000000000005c000000000000005f000000000000006300000000",
            INIT_26 => X"000000460000000000000060000000000000006c000000000000006400000000",
            INIT_27 => X"000000f900000000000000d0000000000000006c000000000000004f00000000",
            INIT_28 => X"0000006e00000000000000c000000000000000c000000000000000c200000000",
            INIT_29 => X"0000003f0000000000000049000000000000003e000000000000004c00000000",
            INIT_2A => X"000000300000000000000028000000000000001d000000000000002e00000000",
            INIT_2B => X"0000003b00000000000000530000000000000048000000000000004100000000",
            INIT_2C => X"00000043000000000000004d0000000000000043000000000000003000000000",
            INIT_2D => X"00000058000000000000003b0000000000000040000000000000003c00000000",
            INIT_2E => X"00000069000000000000004e0000000000000036000000000000005200000000",
            INIT_2F => X"000000f900000000000000c90000000000000065000000000000006b00000000",
            INIT_30 => X"0000006100000000000000bb00000000000000be00000000000000c300000000",
            INIT_31 => X"0000004300000000000000410000000000000063000000000000005500000000",
            INIT_32 => X"0000002000000000000000230000000000000026000000000000003a00000000",
            INIT_33 => X"0000004c000000000000008d0000000000000060000000000000004800000000",
            INIT_34 => X"00000071000000000000008c000000000000004f000000000000001900000000",
            INIT_35 => X"000000920000000000000061000000000000006d000000000000005e00000000",
            INIT_36 => X"0000008a0000000000000045000000000000003a00000000000000ab00000000",
            INIT_37 => X"000000f400000000000000c00000000000000053000000000000007400000000",
            INIT_38 => X"0000005200000000000000b000000000000000b700000000000000bd00000000",
            INIT_39 => X"0000005e00000000000000590000000000000063000000000000002c00000000",
            INIT_3A => X"0000002100000000000000240000000000000030000000000000005a00000000",
            INIT_3B => X"000000340000000000000055000000000000002f000000000000002600000000",
            INIT_3C => X"0000007b0000000000000091000000000000004a000000000000001c00000000",
            INIT_3D => X"0000009700000000000000710000000000000086000000000000007700000000",
            INIT_3E => X"0000004700000000000000320000000000000033000000000000009c00000000",
            INIT_3F => X"000000ee00000000000000c00000000000000047000000000000003b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004800000000000000a300000000000000ad00000000000000ae00000000",
            INIT_41 => X"0000008b00000000000000650000000000000036000000000000002200000000",
            INIT_42 => X"0000001e0000000000000028000000000000003a000000000000006600000000",
            INIT_43 => X"0000001e000000000000001a0000000000000019000000000000001a00000000",
            INIT_44 => X"0000005600000000000000350000000000000026000000000000002500000000",
            INIT_45 => X"0000007200000000000000760000000000000075000000000000006800000000",
            INIT_46 => X"0000002e0000000000000030000000000000002b000000000000003e00000000",
            INIT_47 => X"000000df00000000000000b8000000000000004b000000000000002f00000000",
            INIT_48 => X"00000078000000000000009e00000000000000a000000000000000a200000000",
            INIT_49 => X"0000008800000000000000670000000000000059000000000000005700000000",
            INIT_4A => X"0000002200000000000000340000000000000048000000000000005c00000000",
            INIT_4B => X"0000001d000000000000001b000000000000001b000000000000001c00000000",
            INIT_4C => X"000000af000000000000003d0000000000000015000000000000002000000000",
            INIT_4D => X"000000b400000000000000b100000000000000ca00000000000000cf00000000",
            INIT_4E => X"0000002c00000000000000280000000000000022000000000000005400000000",
            INIT_4F => X"000000d100000000000000ab0000000000000057000000000000003e00000000",
            INIT_50 => X"000000b000000000000000a8000000000000009c000000000000009c00000000",
            INIT_51 => X"0000008800000000000000660000000000000070000000000000009300000000",
            INIT_52 => X"0000002d000000000000004b0000000000000051000000000000005600000000",
            INIT_53 => X"0000001a00000000000000170000000000000016000000000000001600000000",
            INIT_54 => X"000000a400000000000000450000000000000022000000000000002300000000",
            INIT_55 => X"000000a500000000000000a900000000000000b100000000000000b900000000",
            INIT_56 => X"0000002d000000000000001a0000000000000019000000000000004e00000000",
            INIT_57 => X"000000cc00000000000000a7000000000000005c000000000000004b00000000",
            INIT_58 => X"000000a100000000000000ad00000000000000a7000000000000009500000000",
            INIT_59 => X"0000008e00000000000000630000000000000071000000000000008d00000000",
            INIT_5A => X"00000033000000000000004f0000000000000053000000000000005300000000",
            INIT_5B => X"00000022000000000000001f000000000000001c000000000000001d00000000",
            INIT_5C => X"0000006100000000000000510000000000000048000000000000003200000000",
            INIT_5D => X"00000085000000000000008a0000000000000074000000000000006600000000",
            INIT_5E => X"00000032000000000000001d000000000000001b000000000000003700000000",
            INIT_5F => X"000000c600000000000000a40000000000000059000000000000004c00000000",
            INIT_60 => X"00000090000000000000009b00000000000000a600000000000000a400000000",
            INIT_61 => X"0000006c00000000000000630000000000000082000000000000008b00000000",
            INIT_62 => X"0000003800000000000000480000000000000050000000000000004c00000000",
            INIT_63 => X"0000002900000000000000270000000000000024000000000000002600000000",
            INIT_64 => X"00000048000000000000003d0000000000000033000000000000002d00000000",
            INIT_65 => X"00000083000000000000007c0000000000000067000000000000005400000000",
            INIT_66 => X"000000320000000000000021000000000000001a000000000000003100000000",
            INIT_67 => X"000000c300000000000000a90000000000000059000000000000004500000000",
            INIT_68 => X"0000008d0000000000000092000000000000009400000000000000a000000000",
            INIT_69 => X"0000004900000000000000660000000000000082000000000000008700000000",
            INIT_6A => X"000000380000000000000042000000000000004d000000000000004500000000",
            INIT_6B => X"0000002d000000000000002b0000000000000028000000000000002f00000000",
            INIT_6C => X"0000003d00000000000000360000000000000030000000000000002e00000000",
            INIT_6D => X"0000006a000000000000005e0000000000000054000000000000004600000000",
            INIT_6E => X"00000030000000000000001f000000000000001a000000000000004000000000",
            INIT_6F => X"000000ba00000000000000af0000000000000062000000000000003d00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009300000000",
            INIT_71 => X"000000390000000000000068000000000000008b000000000000008f00000000",
            INIT_72 => X"00000034000000000000003f000000000000004a000000000000004000000000",
            INIT_73 => X"0000003600000000000000330000000000000031000000000000003700000000",
            INIT_74 => X"00000042000000000000003d0000000000000036000000000000003600000000",
            INIT_75 => X"000000570000000000000051000000000000004a000000000000004400000000",
            INIT_76 => X"0000003400000000000000230000000000000021000000000000004800000000",
            INIT_77 => X"000000b500000000000000b60000000000000084000000000000004800000000",
            INIT_78 => X"000000a300000000000000a10000000000000096000000000000009200000000",
            INIT_79 => X"0000003a000000000000007c0000000000000091000000000000009d00000000",
            INIT_7A => X"0000004100000000000000390000000000000038000000000000003700000000",
            INIT_7B => X"0000004500000000000000460000000000000042000000000000004300000000",
            INIT_7C => X"0000005f00000000000000570000000000000048000000000000004300000000",
            INIT_7D => X"0000005e0000000000000060000000000000005f000000000000005c00000000",
            INIT_7E => X"00000046000000000000003e0000000000000044000000000000005100000000",
            INIT_7F => X"000000b900000000000000b600000000000000a3000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "sampleifmap_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000bf00000000000000ca00000000000000d100000000",
            INIT_01 => X"000000af00000000000000c600000000000000d100000000000000d100000000",
            INIT_02 => X"000000a0000000000000009d00000000000000a500000000000000ab00000000",
            INIT_03 => X"0000008f000000000000008d000000000000009a000000000000009500000000",
            INIT_04 => X"000000db00000000000000d600000000000000bc00000000000000a400000000",
            INIT_05 => X"000000d600000000000000d900000000000000ca00000000000000d100000000",
            INIT_06 => X"000000ad00000000000000a100000000000000b100000000000000d000000000",
            INIT_07 => X"000000950000000000000095000000000000009d00000000000000b700000000",
            INIT_08 => X"000000cd00000000000000d200000000000000d400000000000000d400000000",
            INIT_09 => X"000000a300000000000000c800000000000000db00000000000000cf00000000",
            INIT_0A => X"000000b600000000000000b800000000000000b600000000000000a500000000",
            INIT_0B => X"000000d700000000000000cd00000000000000c900000000000000c200000000",
            INIT_0C => X"000000e400000000000000e300000000000000e300000000000000df00000000",
            INIT_0D => X"000000d700000000000000d300000000000000d400000000000000dd00000000",
            INIT_0E => X"000000bb00000000000000c300000000000000cd00000000000000df00000000",
            INIT_0F => X"000000ba00000000000000ad00000000000000aa00000000000000c600000000",
            INIT_10 => X"000000e200000000000000e300000000000000e500000000000000e600000000",
            INIT_11 => X"000000a400000000000000d300000000000000ec00000000000000e300000000",
            INIT_12 => X"000000b800000000000000b700000000000000ad000000000000009f00000000",
            INIT_13 => X"000000e000000000000000cf00000000000000bf00000000000000bc00000000",
            INIT_14 => X"000000d600000000000000e000000000000000e500000000000000db00000000",
            INIT_15 => X"000000d300000000000000c800000000000000d000000000000000d600000000",
            INIT_16 => X"000000c500000000000000db00000000000000e000000000000000de00000000",
            INIT_17 => X"000000c600000000000000c500000000000000bc00000000000000b900000000",
            INIT_18 => X"000000f100000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"000000af00000000000000e300000000000000f100000000000000f200000000",
            INIT_1A => X"000000bb00000000000000a100000000000000b000000000000000a800000000",
            INIT_1B => X"000000b600000000000000b800000000000000a000000000000000ae00000000",
            INIT_1C => X"000000ca00000000000000d000000000000000d500000000000000b900000000",
            INIT_1D => X"000000d400000000000000c400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000bb00000000000000d500000000000000dc00000000000000d700000000",
            INIT_1F => X"000000c800000000000000d400000000000000c500000000000000a900000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000008400000000000000cd00000000000000f100000000000000f500000000",
            INIT_22 => X"000000a7000000000000008a00000000000000a1000000000000008b00000000",
            INIT_23 => X"0000008d000000000000009b000000000000008b000000000000009f00000000",
            INIT_24 => X"000000a4000000000000009900000000000000a6000000000000008e00000000",
            INIT_25 => X"000000e000000000000000c400000000000000a900000000000000a900000000",
            INIT_26 => X"000000b100000000000000d400000000000000d100000000000000d100000000",
            INIT_27 => X"000000d200000000000000cc00000000000000b800000000000000a000000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000008100000000000000d700000000000000ee00000000000000f600000000",
            INIT_2A => X"000000aa00000000000000a0000000000000009c000000000000007100000000",
            INIT_2B => X"000000a700000000000000b100000000000000aa00000000000000aa00000000",
            INIT_2C => X"0000008f0000000000000098000000000000009d000000000000009d00000000",
            INIT_2D => X"000000e400000000000000cd00000000000000b3000000000000009400000000",
            INIT_2E => X"000000aa00000000000000c100000000000000ce00000000000000da00000000",
            INIT_2F => X"000000df00000000000000c000000000000000a0000000000000009300000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"000000b400000000000000dd00000000000000dd00000000000000f100000000",
            INIT_32 => X"000000cf00000000000000c400000000000000b4000000000000008300000000",
            INIT_33 => X"000000d300000000000000d900000000000000cb00000000000000c800000000",
            INIT_34 => X"000000bf00000000000000c000000000000000c300000000000000cc00000000",
            INIT_35 => X"000000e100000000000000cd00000000000000a600000000000000a300000000",
            INIT_36 => X"000000a900000000000000b100000000000000d500000000000000e300000000",
            INIT_37 => X"000000da00000000000000b20000000000000092000000000000009100000000",
            INIT_38 => X"000000f700000000000000f200000000000000f200000000000000f400000000",
            INIT_39 => X"000000c000000000000000d900000000000000ca00000000000000e600000000",
            INIT_3A => X"000000e800000000000000e000000000000000c2000000000000008600000000",
            INIT_3B => X"000000d100000000000000ce00000000000000d700000000000000ea00000000",
            INIT_3C => X"000000cf00000000000000ca00000000000000d000000000000000cf00000000",
            INIT_3D => X"000000cc000000000000009a00000000000000b400000000000000e000000000",
            INIT_3E => X"000000bc00000000000000c400000000000000c900000000000000dc00000000",
            INIT_3F => X"000000c7000000000000009a000000000000009200000000000000ab00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f300000000000000f300000000000000f500000000",
            INIT_41 => X"000000ae00000000000000df00000000000000d100000000000000e300000000",
            INIT_42 => X"000000c100000000000000c100000000000000ba000000000000008700000000",
            INIT_43 => X"000000c900000000000000c100000000000000cc00000000000000dd00000000",
            INIT_44 => X"000000c600000000000000cd00000000000000cd00000000000000ca00000000",
            INIT_45 => X"000000bc00000000000000a300000000000000d000000000000000dc00000000",
            INIT_46 => X"000000cb00000000000000df00000000000000d100000000000000cb00000000",
            INIT_47 => X"000000b20000000000000094000000000000008b00000000000000a100000000",
            INIT_48 => X"000000f200000000000000f300000000000000f100000000000000f200000000",
            INIT_49 => X"000000a400000000000000c200000000000000cd00000000000000e500000000",
            INIT_4A => X"000000b800000000000000bd00000000000000c1000000000000008c00000000",
            INIT_4B => X"000000c400000000000000c000000000000000c400000000000000ca00000000",
            INIT_4C => X"000000c600000000000000d000000000000000ca00000000000000c700000000",
            INIT_4D => X"000000c800000000000000bc00000000000000e000000000000000d700000000",
            INIT_4E => X"000000e300000000000000ed00000000000000ee00000000000000e600000000",
            INIT_4F => X"000000d300000000000000ca00000000000000ba00000000000000bc00000000",
            INIT_50 => X"000000f400000000000000f300000000000000ee00000000000000ea00000000",
            INIT_51 => X"0000009c00000000000000a900000000000000a000000000000000df00000000",
            INIT_52 => X"000000ac00000000000000b300000000000000b1000000000000008600000000",
            INIT_53 => X"000000b700000000000000b400000000000000ae00000000000000ae00000000",
            INIT_54 => X"000000be00000000000000bc00000000000000be00000000000000bb00000000",
            INIT_55 => X"000000c400000000000000d000000000000000dc00000000000000cd00000000",
            INIT_56 => X"000000f400000000000000f600000000000000e600000000000000d900000000",
            INIT_57 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_58 => X"000000f200000000000000f200000000000000e600000000000000d300000000",
            INIT_59 => X"0000009700000000000000be00000000000000b600000000000000d800000000",
            INIT_5A => X"000000a00000000000000093000000000000006e000000000000006a00000000",
            INIT_5B => X"000000aa00000000000000a6000000000000009f000000000000009e00000000",
            INIT_5C => X"000000a6000000000000009e00000000000000a300000000000000a900000000",
            INIT_5D => X"000000af00000000000000c600000000000000bd00000000000000ad00000000",
            INIT_5E => X"000000f300000000000000f800000000000000e000000000000000b700000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e100000000000000e900000000000000da00000000000000c400000000",
            INIT_61 => X"0000009f00000000000000c300000000000000b400000000000000bd00000000",
            INIT_62 => X"000000a0000000000000008d000000000000005c000000000000005d00000000",
            INIT_63 => X"0000008c000000000000008f00000000000000a800000000000000ba00000000",
            INIT_64 => X"000000a700000000000000920000000000000089000000000000008b00000000",
            INIT_65 => X"00000096000000000000008f0000000000000083000000000000009800000000",
            INIT_66 => X"000000f400000000000000f300000000000000e300000000000000bc00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c100000000000000d300000000000000c700000000000000c300000000",
            INIT_69 => X"0000008900000000000000a2000000000000009500000000000000a400000000",
            INIT_6A => X"000000a600000000000000b200000000000000aa000000000000009600000000",
            INIT_6B => X"0000009200000000000000a600000000000000cd00000000000000bd00000000",
            INIT_6C => X"000000d300000000000000c000000000000000ac000000000000009900000000",
            INIT_6D => X"0000008a0000000000000080000000000000008000000000000000af00000000",
            INIT_6E => X"000000d300000000000000bf00000000000000b100000000000000a000000000",
            INIT_6F => X"000000f300000000000000f300000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a200000000000000c800000000000000cf00000000000000c200000000",
            INIT_71 => X"00000089000000000000008e0000000000000088000000000000009c00000000",
            INIT_72 => X"0000009f00000000000000b100000000000000b200000000000000a200000000",
            INIT_73 => X"0000008b000000000000009500000000000000a3000000000000009600000000",
            INIT_74 => X"0000009300000000000000920000000000000092000000000000008d00000000",
            INIT_75 => X"00000085000000000000007f000000000000007c000000000000008600000000",
            INIT_76 => X"000000a600000000000000ad00000000000000a3000000000000009500000000",
            INIT_77 => X"000000f400000000000000f300000000000000f500000000000000cc00000000",
            INIT_78 => X"0000006e00000000000000ad00000000000000d000000000000000c300000000",
            INIT_79 => X"000000b900000000000000b4000000000000008b000000000000007100000000",
            INIT_7A => X"00000057000000000000007f000000000000009a000000000000008500000000",
            INIT_7B => X"0000005f0000000000000059000000000000004c000000000000004900000000",
            INIT_7C => X"00000058000000000000005e0000000000000060000000000000005c00000000",
            INIT_7D => X"0000006700000000000000630000000000000056000000000000005600000000",
            INIT_7E => X"0000009b000000000000008f0000000000000074000000000000006d00000000",
            INIT_7F => X"000000f500000000000000f500000000000000e800000000000000af00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "sampleifmap_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006500000000000000a100000000000000aa00000000000000b700000000",
            INIT_01 => X"000000a100000000000000b50000000000000088000000000000006000000000",
            INIT_02 => X"0000008700000000000000810000000000000084000000000000008000000000",
            INIT_03 => X"0000006a000000000000007d000000000000007d000000000000008c00000000",
            INIT_04 => X"00000027000000000000002c000000000000002b000000000000003500000000",
            INIT_05 => X"0000002800000000000000230000000000000047000000000000004d00000000",
            INIT_06 => X"0000009700000000000000910000000000000050000000000000002000000000",
            INIT_07 => X"000000f300000000000000f600000000000000db00000000000000a700000000",
            INIT_08 => X"0000007c00000000000000c200000000000000c100000000000000ca00000000",
            INIT_09 => X"0000004900000000000000990000000000000092000000000000007800000000",
            INIT_0A => X"0000009400000000000000830000000000000087000000000000006900000000",
            INIT_0B => X"0000008300000000000000a9000000000000009f00000000000000b800000000",
            INIT_0C => X"0000007a00000000000000840000000000000076000000000000006600000000",
            INIT_0D => X"00000073000000000000006f00000000000000aa00000000000000af00000000",
            INIT_0E => X"000000b500000000000000b20000000000000091000000000000006f00000000",
            INIT_0F => X"000000f400000000000000f200000000000000c500000000000000bb00000000",
            INIT_10 => X"0000007200000000000000b800000000000000c800000000000000d800000000",
            INIT_11 => X"000000240000000000000082000000000000009d000000000000007300000000",
            INIT_12 => X"0000006300000000000000810000000000000095000000000000004f00000000",
            INIT_13 => X"00000084000000000000009d0000000000000081000000000000006f00000000",
            INIT_14 => X"000000b900000000000000b700000000000000c100000000000000b100000000",
            INIT_15 => X"000000bd00000000000000ba00000000000000c100000000000000c800000000",
            INIT_16 => X"0000009700000000000000b600000000000000c700000000000000b500000000",
            INIT_17 => X"000000f600000000000000e800000000000000a2000000000000009400000000",
            INIT_18 => X"0000007100000000000000bb00000000000000cc00000000000000d900000000",
            INIT_19 => X"0000003d0000000000000071000000000000008b000000000000006000000000",
            INIT_1A => X"0000005d00000000000000730000000000000070000000000000004e00000000",
            INIT_1B => X"0000007d000000000000005e0000000000000053000000000000005500000000",
            INIT_1C => X"0000008a000000000000007f000000000000009f00000000000000bf00000000",
            INIT_1D => X"0000008f000000000000008c000000000000009500000000000000a000000000",
            INIT_1E => X"00000063000000000000009f00000000000000bd000000000000008a00000000",
            INIT_1F => X"000000f700000000000000e2000000000000009a000000000000007300000000",
            INIT_20 => X"0000007500000000000000c700000000000000d000000000000000d500000000",
            INIT_21 => X"000000540000000000000063000000000000005c000000000000004900000000",
            INIT_22 => X"0000006900000000000000610000000000000041000000000000004b00000000",
            INIT_23 => X"0000005f00000000000000670000000000000057000000000000005f00000000",
            INIT_24 => X"00000097000000000000009900000000000000a2000000000000008600000000",
            INIT_25 => X"0000008f00000000000000890000000000000090000000000000009600000000",
            INIT_26 => X"0000006f000000000000008f0000000000000099000000000000009300000000",
            INIT_27 => X"000000f700000000000000de0000000000000092000000000000007300000000",
            INIT_28 => X"0000008300000000000000cc00000000000000ce00000000000000cc00000000",
            INIT_29 => X"0000005a000000000000005c0000000000000051000000000000006500000000",
            INIT_2A => X"000000450000000000000039000000000000002d000000000000004600000000",
            INIT_2B => X"00000057000000000000007d000000000000006f000000000000006200000000",
            INIT_2C => X"0000006700000000000000700000000000000066000000000000004a00000000",
            INIT_2D => X"0000007d000000000000005e0000000000000065000000000000006200000000",
            INIT_2E => X"0000009500000000000000710000000000000052000000000000007300000000",
            INIT_2F => X"000000f800000000000000d40000000000000089000000000000009a00000000",
            INIT_30 => X"0000007500000000000000ce00000000000000d000000000000000d100000000",
            INIT_31 => X"0000005e0000000000000056000000000000007a000000000000006900000000",
            INIT_32 => X"0000002f00000000000000330000000000000036000000000000005600000000",
            INIT_33 => X"0000006300000000000000ad0000000000000083000000000000006600000000",
            INIT_34 => X"00000082000000000000009e0000000000000064000000000000002d00000000",
            INIT_35 => X"000000ab000000000000007c000000000000008a000000000000007900000000",
            INIT_36 => X"000000ab000000000000005f000000000000004b00000000000000bb00000000",
            INIT_37 => X"000000fa00000000000000cf0000000000000075000000000000009800000000",
            INIT_38 => X"0000006800000000000000cc00000000000000d600000000000000dd00000000",
            INIT_39 => X"0000008000000000000000720000000000000074000000000000003b00000000",
            INIT_3A => X"0000003000000000000000340000000000000041000000000000007c00000000",
            INIT_3B => X"0000004b000000000000006c0000000000000046000000000000003800000000",
            INIT_3C => X"0000008f00000000000000a6000000000000005f000000000000003000000000",
            INIT_3D => X"000000af000000000000008f00000000000000a7000000000000009100000000",
            INIT_3E => X"000000620000000000000048000000000000004a00000000000000af00000000",
            INIT_3F => X"000000fb00000000000000d60000000000000068000000000000005400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006300000000000000c900000000000000d400000000000000d700000000",
            INIT_41 => X"000000b000000000000000800000000000000044000000000000002f00000000",
            INIT_42 => X"0000002d00000000000000380000000000000050000000000000008700000000",
            INIT_43 => X"0000002f000000000000002b0000000000000027000000000000002800000000",
            INIT_44 => X"0000006e0000000000000050000000000000003c000000000000003700000000",
            INIT_45 => X"0000008b00000000000000900000000000000093000000000000007d00000000",
            INIT_46 => X"0000004300000000000000460000000000000043000000000000005c00000000",
            INIT_47 => X"000000fb00000000000000d9000000000000006d000000000000004500000000",
            INIT_48 => X"0000009d00000000000000cb00000000000000cf00000000000000cf00000000",
            INIT_49 => X"000000aa00000000000000850000000000000075000000000000007300000000",
            INIT_4A => X"0000003000000000000000480000000000000065000000000000007e00000000",
            INIT_4B => X"0000002d00000000000000290000000000000029000000000000002800000000",
            INIT_4C => X"000000c000000000000000530000000000000027000000000000003200000000",
            INIT_4D => X"000000c900000000000000c700000000000000dc00000000000000da00000000",
            INIT_4E => X"0000003f00000000000000380000000000000034000000000000006b00000000",
            INIT_4F => X"000000f700000000000000d2000000000000007e000000000000005a00000000",
            INIT_50 => X"000000d800000000000000ce00000000000000c000000000000000bc00000000",
            INIT_51 => X"000000a10000000000000086000000000000009a00000000000000bf00000000",
            INIT_52 => X"0000003e00000000000000680000000000000073000000000000007900000000",
            INIT_53 => X"0000002900000000000000230000000000000022000000000000002100000000",
            INIT_54 => X"000000b300000000000000550000000000000031000000000000003300000000",
            INIT_55 => X"000000bb00000000000000be00000000000000c000000000000000c700000000",
            INIT_56 => X"0000004200000000000000260000000000000027000000000000006000000000",
            INIT_57 => X"000000f500000000000000d10000000000000085000000000000006f00000000",
            INIT_58 => X"000000c600000000000000cd00000000000000c600000000000000bf00000000",
            INIT_59 => X"000000a00000000000000084000000000000009e00000000000000b500000000",
            INIT_5A => X"00000046000000000000006f0000000000000076000000000000007200000000",
            INIT_5B => X"00000031000000000000002c0000000000000026000000000000002700000000",
            INIT_5C => X"0000007e0000000000000069000000000000005d000000000000004400000000",
            INIT_5D => X"000000a600000000000000ad0000000000000096000000000000008700000000",
            INIT_5E => X"00000047000000000000002a0000000000000028000000000000004800000000",
            INIT_5F => X"000000f200000000000000cf0000000000000082000000000000007100000000",
            INIT_60 => X"000000b800000000000000c600000000000000d100000000000000ce00000000",
            INIT_61 => X"00000085000000000000008200000000000000a300000000000000ab00000000",
            INIT_62 => X"0000004d0000000000000068000000000000006f000000000000006b00000000",
            INIT_63 => X"000000390000000000000035000000000000002f000000000000003200000000",
            INIT_64 => X"0000006800000000000000570000000000000048000000000000003f00000000",
            INIT_65 => X"000000b000000000000000a80000000000000091000000000000007800000000",
            INIT_66 => X"0000004700000000000000300000000000000028000000000000004500000000",
            INIT_67 => X"000000ee00000000000000d4000000000000007e000000000000006600000000",
            INIT_68 => X"000000bd00000000000000c200000000000000c200000000000000c700000000",
            INIT_69 => X"00000065000000000000008600000000000000a600000000000000b200000000",
            INIT_6A => X"0000004f00000000000000600000000000000069000000000000006300000000",
            INIT_6B => X"0000003e000000000000003b0000000000000036000000000000003e00000000",
            INIT_6C => X"00000057000000000000004e0000000000000045000000000000004100000000",
            INIT_6D => X"0000008f00000000000000810000000000000074000000000000006400000000",
            INIT_6E => X"00000047000000000000002c0000000000000027000000000000005700000000",
            INIT_6F => X"000000e800000000000000df0000000000000085000000000000005900000000",
            INIT_70 => X"000000bc00000000000000be00000000000000bc00000000000000c100000000",
            INIT_71 => X"00000050000000000000009000000000000000bc00000000000000bd00000000",
            INIT_72 => X"0000004600000000000000580000000000000063000000000000005a00000000",
            INIT_73 => X"0000004e000000000000004a0000000000000045000000000000004900000000",
            INIT_74 => X"0000005d0000000000000056000000000000004e000000000000004e00000000",
            INIT_75 => X"00000072000000000000006d0000000000000066000000000000006100000000",
            INIT_76 => X"0000004a00000000000000300000000000000030000000000000005e00000000",
            INIT_77 => X"000000e700000000000000e800000000000000ad000000000000006400000000",
            INIT_78 => X"000000cd00000000000000d000000000000000c700000000000000c400000000",
            INIT_79 => X"0000005500000000000000a500000000000000bb00000000000000c800000000",
            INIT_7A => X"00000054000000000000004e000000000000004c000000000000004c00000000",
            INIT_7B => X"0000006300000000000000620000000000000059000000000000005400000000",
            INIT_7C => X"0000007c00000000000000720000000000000063000000000000005e00000000",
            INIT_7D => X"0000007f00000000000000800000000000000081000000000000007d00000000",
            INIT_7E => X"000000600000000000000054000000000000005b000000000000007000000000",
            INIT_7F => X"000000df00000000000000e100000000000000cc000000000000009400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "samplegold_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000009000000000000000a0000000000000010000000000000001000000000",
            INIT_01 => X"0000000d000000000000000c0000000000000008000000000000000600000000",
            INIT_02 => X"0000000f0000000000000014000000000000000b000000000000000500000000",
            INIT_03 => X"0000000000000000000000010000000000000002000000000000000700000000",
            INIT_04 => X"0000000a000000000000000b0000000000000009000000000000000300000000",
            INIT_05 => X"0000002900000000000000050000000000000003000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000001f000000000000000f0000000000000000000000000000000500000000",
            INIT_08 => X"0000004c000000000000000c000000000000000a000000000000000800000000",
            INIT_09 => X"0000000000000000000000000000000000000013000000000000002c00000000",
            INIT_0A => X"0000000000000000000000000000000000000012000000000000002100000000",
            INIT_0B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000030000000000000000000000000000000300000000",
            INIT_0D => X"0000002d00000000000000290000000000000001000000000000000800000000",
            INIT_0E => X"000000000000000000000000000000000000001c000000000000002400000000",
            INIT_0F => X"0000000e00000000000000110000000000000000000000000000002700000000",
            INIT_10 => X"000000130000000000000033000000000000000a000000000000000000000000",
            INIT_11 => X"0000000b00000000000000110000000000000000000000000000000d00000000",
            INIT_12 => X"0000006900000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000007f000000000000003a0000000000000027000000000000002b00000000",
            INIT_14 => X"0000000000000000000000140000000000000025000000000000007c00000000",
            INIT_15 => X"0000000e000000000000003c0000000000000053000000000000000000000000",
            INIT_16 => X"0000002a000000000000005e0000000000000000000000000000000300000000",
            INIT_17 => X"0000001a000000000000001e0000000000000013000000000000002e00000000",
            INIT_18 => X"000000000000000000000017000000000000002c000000000000004f00000000",
            INIT_19 => X"0000000000000000000000010000000000000013000000000000005600000000",
            INIT_1A => X"00000007000000000000003b0000000000000058000000000000000200000000",
            INIT_1B => X"00000080000000000000003b000000000000000b000000000000000000000000",
            INIT_1C => X"0000004d000000000000001e000000000000002c000000000000005000000000",
            INIT_1D => X"000000200000000000000025000000000000000f000000000000002300000000",
            INIT_1E => X"0000000e0000000000000041000000000000004f000000000000005f00000000",
            INIT_1F => X"0000000000000000000000320000000000000069000000000000001300000000",
            INIT_20 => X"0000004800000000000000350000000000000012000000000000000100000000",
            INIT_21 => X"0000007100000000000000000000000000000003000000000000001500000000",
            INIT_22 => X"0000002e000000000000000c0000000000000040000000000000005e00000000",
            INIT_23 => X"000000170000000000000000000000000000001b000000000000002400000000",
            INIT_24 => X"0000000000000000000000000000000000000035000000000000004b00000000",
            INIT_25 => X"000000540000000000000035000000000000000f000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_27 => X"00000000000000000000003c0000000000000072000000000000002200000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000004c00000000000000670000000000000056000000000000000100000000",
            INIT_2A => X"00000047000000000000008700000000000000c4000000000000002100000000",
            INIT_2B => X"0000000c00000000000000110000000000000027000000000000004800000000",
            INIT_2C => X"0000001e00000000000000170000000000000014000000000000001500000000",
            INIT_2D => X"0000006d00000000000000510000000000000044000000000000001000000000",
            INIT_2E => X"000000130000000000000016000000000000001500000000000000a300000000",
            INIT_2F => X"0000000700000000000000060000000000000007000000000000000f00000000",
            INIT_30 => X"00000023000000000000000e000000000000002a000000000000001f00000000",
            INIT_31 => X"000000390000000000000090000000000000004d000000000000000a00000000",
            INIT_32 => X"000000160000000000000010000000000000000f000000000000001500000000",
            INIT_33 => X"00000024000000000000002c000000000000001f000000000000001400000000",
            INIT_34 => X"000000180000000000000029000000000000004a000000000000000b00000000",
            INIT_35 => X"0000002600000000000000240000000000000050000000000000001c00000000",
            INIT_36 => X"0000000b000000000000000c000000000000001c000000000000003100000000",
            INIT_37 => X"0000001b0000000000000003000000000000001a000000000000001b00000000",
            INIT_38 => X"00000080000000000000007c000000000000007a000000000000001f00000000",
            INIT_39 => X"00000081000000000000007c0000000000000080000000000000008000000000",
            INIT_3A => X"0000006100000000000000710000000000000087000000000000008b00000000",
            INIT_3B => X"0000007000000000000000710000000000000069000000000000006400000000",
            INIT_3C => X"0000008200000000000000870000000000000083000000000000008100000000",
            INIT_3D => X"000000740000000000000072000000000000007b000000000000008300000000",
            INIT_3E => X"0000002d0000000000000025000000000000003c000000000000004e00000000",
            INIT_3F => X"00000060000000000000006b000000000000005d000000000000004600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008700000000000000850000000000000082000000000000006700000000",
            INIT_41 => X"000000310000000000000035000000000000003e000000000000007100000000",
            INIT_42 => X"0000001700000000000000190000000000000017000000000000002f00000000",
            INIT_43 => X"0000005c00000000000000140000000000000059000000000000003e00000000",
            INIT_44 => X"0000005900000000000000720000000000000088000000000000007200000000",
            INIT_45 => X"0000003b000000000000001b0000000000000025000000000000003500000000",
            INIT_46 => X"0000001f000000000000000e0000000000000023000000000000001400000000",
            INIT_47 => X"00000059000000000000003d0000000000000000000000000000005500000000",
            INIT_48 => X"0000001a000000000000003d0000000000000043000000000000008700000000",
            INIT_49 => X"00000024000000000000003e0000000000000016000000000000001900000000",
            INIT_4A => X"0000004200000000000000140000000000000022000000000000001800000000",
            INIT_4B => X"0000005f000000000000004d0000000000000022000000000000000400000000",
            INIT_4C => X"0000002000000000000000180000000000000028000000000000003600000000",
            INIT_4D => X"0000000c0000000000000014000000000000005c000000000000000d00000000",
            INIT_4E => X"00000009000000000000001b0000000000000016000000000000002600000000",
            INIT_4F => X"0000005500000000000000500000000000000044000000000000000300000000",
            INIT_50 => X"0000000b00000000000000170000000000000020000000000000004300000000",
            INIT_51 => X"0000001e00000000000000110000000000000001000000000000004600000000",
            INIT_52 => X"00000000000000000000000c0000000000000020000000000000001f00000000",
            INIT_53 => X"0000004500000000000000520000000000000035000000000000002c00000000",
            INIT_54 => X"0000004b0000000000000016000000000000001a000000000000000a00000000",
            INIT_55 => X"000000240000000000000024000000000000000d000000000000001100000000",
            INIT_56 => X"0000000000000000000000050000000000000001000000000000003d00000000",
            INIT_57 => X"0000001c00000000000000200000000000000031000000000000002300000000",
            INIT_58 => X"0000003100000000000000270000000000000033000000000000002000000000",
            INIT_59 => X"00000066000000000000003c0000000000000024000000000000000d00000000",
            INIT_5A => X"000000190000000000000000000000000000000d000000000000000d00000000",
            INIT_5B => X"0000000f00000000000000300000000000000033000000000000001000000000",
            INIT_5C => X"00000014000000000000000a0000000000000028000000000000002c00000000",
            INIT_5D => X"0000000f00000000000000680000000000000062000000000000003400000000",
            INIT_5E => X"0000000000000000000000470000000000000000000000000000000f00000000",
            INIT_5F => X"000000000000000000000000000000000000001f000000000000001600000000",
            INIT_60 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"000000000000000000000000000000000000003b000000000000000200000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000110000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "samplegold_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_03 => X"0000000000000000000000170000000000000016000000000000000000000000",
            INIT_04 => X"0000000f000000000000000b0000000000000025000000000000000000000000",
            INIT_05 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000021000000000000001200000000",
            INIT_08 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_0A => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_0C => X"000000000000000000000000000000000000000b000000000000002300000000",
            INIT_0D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_0E => X"0000003c00000000000000320000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000005000000000000000700000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_12 => X"00000020000000000000002f000000000000002e000000000000000000000000",
            INIT_13 => X"000000000000000000000000000000000000001c000000000000000b00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000170000000000000022000000000000002c000000000000003500000000",
            INIT_17 => X"0000003600000000000000180000000000000016000000000000002c00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_19 => X"00000041000000000000001b000000000000001b000000000000000600000000",
            INIT_1A => X"0000006200000000000000320000000000000028000000000000003600000000",
            INIT_1B => X"0000002000000000000000290000000000000025000000000000003000000000",
            INIT_1C => X"00000025000000000000001e000000000000001b000000000000001800000000",
            INIT_1D => X"0000002900000000000000260000000000000029000000000000002500000000",
            INIT_1E => X"0000001a00000000000000380000000000000057000000000000002000000000",
            INIT_1F => X"0000001600000000000000140000000000000014000000000000001900000000",
            INIT_20 => X"0000002d000000000000002a0000000000000027000000000000002000000000",
            INIT_21 => X"0000002a00000000000000230000000000000035000000000000003200000000",
            INIT_22 => X"0000001a000000000000001a000000000000001b000000000000005800000000",
            INIT_23 => X"0000002600000000000000200000000000000019000000000000001800000000",
            INIT_24 => X"000000390000000000000037000000000000002c000000000000003100000000",
            INIT_25 => X"0000003c000000000000001e000000000000002a000000000000003000000000",
            INIT_26 => X"00000017000000000000001e0000000000000019000000000000001300000000",
            INIT_27 => X"0000002000000000000000260000000000000023000000000000001a00000000",
            INIT_28 => X"00000011000000000000002e0000000000000042000000000000002d00000000",
            INIT_29 => X"0000001000000000000000150000000000000015000000000000001a00000000",
            INIT_2A => X"0000000a000000000000000a000000000000000f000000000000001900000000",
            INIT_2B => X"0000001800000000000000150000000000000011000000000000000b00000000",
            INIT_2C => X"0000000e000000000000000b0000000000000006000000000000000a00000000",
            INIT_2D => X"0000005000000000000000190000000000000013000000000000001100000000",
            INIT_2E => X"0000003800000000000000110000000000000010000000000000000e00000000",
            INIT_2F => X"0000000f0000000000000014000000000000001c000000000000003700000000",
            INIT_30 => X"0000000f00000000000000160000000000000011000000000000000b00000000",
            INIT_31 => X"000000350000000000000041000000000000000d000000000000001000000000",
            INIT_32 => X"00000070000000000000006b000000000000001c000000000000001900000000",
            INIT_33 => X"0000001d00000000000000050000000000000030000000000000006600000000",
            INIT_34 => X"00000011000000000000000c000000000000001d000000000000002b00000000",
            INIT_35 => X"0000003d000000000000004d0000000000000033000000000000001b00000000",
            INIT_36 => X"000000460000000000000079000000000000005e000000000000004100000000",
            INIT_37 => X"000000840000000000000012000000000000000f000000000000004800000000",
            INIT_38 => X"0000009e000000000000003d0000000000000022000000000000006a00000000",
            INIT_39 => X"000000380000000000000053000000000000007e000000000000007600000000",
            INIT_3A => X"0000004600000000000000460000000000000079000000000000005400000000",
            INIT_3B => X"000000b000000000000000980000000000000000000000000000002a00000000",
            INIT_3C => X"000000a100000000000000c1000000000000002c000000000000003d00000000",
            INIT_3D => X"000000780000000000000038000000000000005b00000000000000a100000000",
            INIT_3E => X"00000049000000000000004c000000000000005d000000000000009b00000000",
            INIT_3F => X"0000003600000000000000a300000000000000a3000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac00000000000000970000000000000059000000000000001c00000000",
            INIT_41 => X"00000095000000000000008f0000000000000051000000000000008700000000",
            INIT_42 => X"0000004000000000000000580000000000000047000000000000005300000000",
            INIT_43 => X"00000036000000000000004400000000000000c900000000000000b800000000",
            INIT_44 => X"0000007800000000000000af00000000000000af000000000000003b00000000",
            INIT_45 => X"000000550000000000000094000000000000007f000000000000005b00000000",
            INIT_46 => X"000000dc00000000000000430000000000000058000000000000004d00000000",
            INIT_47 => X"0000004b0000000000000080000000000000008200000000000000d700000000",
            INIT_48 => X"00000055000000000000005a0000000000000061000000000000006e00000000",
            INIT_49 => X"00000036000000000000004a000000000000004d000000000000004000000000",
            INIT_4A => X"000000d800000000000000e80000000000000021000000000000004300000000",
            INIT_4B => X"0000004e0000000000000067000000000000008f000000000000009f00000000",
            INIT_4C => X"0000005a000000000000004f0000000000000090000000000000007d00000000",
            INIT_4D => X"000000290000000000000026000000000000001a000000000000004000000000",
            INIT_4E => X"0000009f00000000000000c900000000000000d0000000000000001e00000000",
            INIT_4F => X"000000a5000000000000006e00000000000000e100000000000000d400000000",
            INIT_50 => X"000000380000000000000043000000000000007d00000000000000c800000000",
            INIT_51 => X"00000053000000000000005f000000000000005a000000000000004c00000000",
            INIT_52 => X"000000f700000000000000ba00000000000000e200000000000000a600000000",
            INIT_53 => X"00000084000000000000008500000000000000a200000000000000e500000000",
            INIT_54 => X"00000089000000000000007d0000000000000072000000000000007a00000000",
            INIT_55 => X"000000940000000000000099000000000000009a000000000000009900000000",
            INIT_56 => X"000000bb00000000000000f900000000000000d7000000000000009700000000",
            INIT_57 => X"0000007b000000000000007c000000000000007f000000000000008900000000",
            INIT_58 => X"0000009d000000000000009a0000000000000090000000000000008000000000",
            INIT_59 => X"0000008a00000000000000a800000000000000ba00000000000000a400000000",
            INIT_5A => X"0000008e000000000000009100000000000000fa00000000000000a600000000",
            INIT_5B => X"000000910000000000000085000000000000007b000000000000008800000000",
            INIT_5C => X"000000b200000000000000a200000000000000a2000000000000009b00000000",
            INIT_5D => X"00000089000000000000009f00000000000000ac00000000000000af00000000",
            INIT_5E => X"0000008d000000000000007f0000000000000073000000000000009300000000",
            INIT_5F => X"00000092000000000000009f0000000000000091000000000000008e00000000",
            INIT_60 => X"0000009600000000000000c800000000000000ba000000000000009700000000",
            INIT_61 => X"0000006f000000000000006c000000000000006d000000000000007100000000",
            INIT_62 => X"0000007c00000000000000710000000000000062000000000000007100000000",
            INIT_63 => X"000000620000000000000068000000000000006e000000000000007700000000",
            INIT_64 => X"0000006d000000000000006a0000000000000062000000000000005f00000000",
            INIT_65 => X"0000006c0000000000000073000000000000006c000000000000006800000000",
            INIT_66 => X"0000007500000000000000670000000000000061000000000000003c00000000",
            INIT_67 => X"00000046000000000000002a000000000000001d000000000000003a00000000",
            INIT_68 => X"00000076000000000000006d0000000000000062000000000000005c00000000",
            INIT_69 => X"0000008f00000000000000770000000000000076000000000000007200000000",
            INIT_6A => X"0000000d00000000000000260000000000000058000000000000007f00000000",
            INIT_6B => X"0000003a000000000000002c0000000000000028000000000000002900000000",
            INIT_6C => X"0000006800000000000000030000000000000038000000000000005100000000",
            INIT_6D => X"00000026000000000000004c0000000000000067000000000000006e00000000",
            INIT_6E => X"0000004f0000000000000022000000000000002c000000000000002800000000",
            INIT_6F => X"00000037000000000000002f0000000000000048000000000000003d00000000",
            INIT_70 => X"0000003900000000000000650000000000000000000000000000003000000000",
            INIT_71 => X"00000036000000000000003d0000000000000003000000000000000000000000",
            INIT_72 => X"0000002f0000000000000023000000000000000c000000000000003e00000000",
            INIT_73 => X"0000004300000000000000260000000000000028000000000000002400000000",
            INIT_74 => X"000000650000000000000076000000000000006a000000000000002a00000000",
            INIT_75 => X"0000002f0000000000000030000000000000003e000000000000005800000000",
            INIT_76 => X"0000002800000000000000570000000000000051000000000000000000000000",
            INIT_77 => X"0000003a00000000000000310000000000000012000000000000002b00000000",
            INIT_78 => X"000000250000000000000037000000000000007b000000000000006200000000",
            INIT_79 => X"00000000000000000000003e0000000000000040000000000000004900000000",
            INIT_7A => X"0000001b00000000000000270000000000000036000000000000005c00000000",
            INIT_7B => X"0000001c000000000000002f000000000000002b000000000000002900000000",
            INIT_7C => X"0000007800000000000000190000000000000025000000000000004900000000",
            INIT_7D => X"0000005d0000000000000024000000000000004d000000000000005c00000000",
            INIT_7E => X"0000005200000000000000380000000000000023000000000000004700000000",
            INIT_7F => X"0000002000000000000000460000000000000022000000000000003400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "samplegold_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003000000000000000510000000000000066000000000000003b00000000",
            INIT_01 => X"00000070000000000000004c0000000000000055000000000000001a00000000",
            INIT_02 => X"0000005200000000000000400000000000000035000000000000003800000000",
            INIT_03 => X"0000002d0000000000000004000000000000004c000000000000003100000000",
            INIT_04 => X"0000002400000000000000130000000000000024000000000000003300000000",
            INIT_05 => X"00000002000000000000002b0000000000000065000000000000006000000000",
            INIT_06 => X"000000300000000000000025000000000000006d000000000000003600000000",
            INIT_07 => X"0000000000000000000000030000000000000000000000000000005800000000",
            INIT_08 => X"0000002b000000000000003f000000000000004b000000000000000000000000",
            INIT_09 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"000000280000000000000037000000000000001e000000000000002800000000",
            INIT_0B => X"000000380000000000000074000000000000009d000000000000000000000000",
            INIT_0C => X"00000002000000000000000c000000000000001f000000000000003700000000",
            INIT_0D => X"0000000400000000000000000000000000000000000000000000000200000000",
            INIT_0E => X"0000004e00000000000000180000000000000016000000000000000000000000",
            INIT_0F => X"0000000700000000000000040000000000000004000000000000008800000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_11 => X"0000000400000000000000000000000000000005000000000000000000000000",
            INIT_12 => X"00000032000000000000008b0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_14 => X"0000000700000000000000090000000000000002000000000000000000000000",
            INIT_15 => X"000000000000000000000005000000000000001c000000000000000000000000",
            INIT_16 => X"0000001400000000000000230000000000000043000000000000000500000000",
            INIT_17 => X"0000000000000000000000000000000000000009000000000000001900000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000001300000000000000030000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_20 => X"000000120000000000000000000000000000000d000000000000000500000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_22 => X"00000000000000000000000a0000000000000005000000000000003e00000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000009000000000000000a00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000001c0000000000000000000000000000000d000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000016000000000000000c00000000",
            INIT_36 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000300000000000000000000000000000000000000000",
            INIT_39 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000007000000000000002600000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000f000000000000002a0000000000000031000000000000000000000000",
            INIT_3E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000007000000000000002e0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001d00000000000000480000000000000004000000000000000700000000",
            INIT_43 => X"00000031000000000000002e0000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000070000000000000019000000000000001c00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000260000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000004f00000000000000140000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_4E => X"0000000300000000000000490000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000014000000000000000c00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_52 => X"0000000200000000000000000000000000000000000000000000000600000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000030000000000000009000000000000000000000000",
            INIT_55 => X"0000000600000000000000010000000000000001000000000000000000000000",
            INIT_56 => X"00000000000000000000001d000000000000000d000000000000000000000000",
            INIT_57 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000120000000000000004000000000000000000000000",
            INIT_59 => X"0000000000000000000000030000000000000039000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000007000000000000000900000000",
            INIT_5B => X"0000000000000000000000000000000000000051000000000000000b00000000",
            INIT_5C => X"00000000000000000000001f000000000000000a000000000000000000000000",
            INIT_5D => X"00000000000000000000000c0000000000000000000000000000006500000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000006800000000",
            INIT_60 => X"0000001d00000000000000000000000000000055000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000066000000000000000000000000",
            INIT_62 => X"0000009400000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000080000000000000000000000000000001e00000000",
            INIT_65 => X"0000000000000000000000000000000000000068000000000000001e00000000",
            INIT_66 => X"0000000000000000000001010000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000056000000000000006100000000",
            INIT_6A => X"00000000000000000000000000000000000000cb000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000015000000000000000400000000",
            INIT_6C => X"0000004300000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000005f00000000",
            INIT_6E => X"0000002100000000000000000000000000000000000000000000008000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000090000000000000000000000000000002f000000000000000000000000",
            INIT_71 => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_72 => X"00000020000000000000001f0000000000000000000000000000000e00000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_74 => X"0000003900000000000000080000000000000000000000000000005500000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000002e000000000000002d000000000000000000000000",
            INIT_77 => X"000000dc00000000000000000000000000000000000000000000005e00000000",
            INIT_78 => X"00000000000000000000004b0000000000000000000000000000000000000000",
            INIT_79 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000004e0000000000000000000000000000000a000000000000000d00000000",
            INIT_7B => X"0000000000000000000000960000000000000000000000000000004100000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000500000000000000060000000000000002000000000000000000000000",
            INIT_7E => X"0000005200000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000008500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "samplegold_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000400000000000000000000000000000005000000000000000800000000",
            INIT_02 => X"000000ac00000000000000000000000000000000000000000000000e00000000",
            INIT_03 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000040000000000000006000000000000000000000000",
            INIT_05 => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_06 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000080000000000000016000000000000000000000000",
            INIT_08 => X"0000000400000000000000000000000000000000000000000000000c00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000008000000000000001c00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000001b0000000000000022000000000000000b000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000018000000000000002800000000",
            INIT_15 => X"0000000000000000000000000000000000000007000000000000001b00000000",
            INIT_16 => X"0000001500000000000000050000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000060000000000000000000000000000001700000000",
            INIT_18 => X"000000340000000000000000000000000000000d000000000000000d00000000",
            INIT_19 => X"0000002700000000000000000000000000000000000000000000002900000000",
            INIT_1A => X"0000000f00000000000000160000000000000005000000000000001500000000",
            INIT_1B => X"0000002000000000000000150000000000000017000000000000001100000000",
            INIT_1C => X"00000010000000000000001a0000000000000000000000000000002600000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000024000000000000002a0000000000000016000000000000000a00000000",
            INIT_1F => X"0000002600000000000000140000000000000007000000000000000100000000",
            INIT_20 => X"00000000000000000000000e000000000000002b000000000000002e00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000300000000000000150000000000000018000000000000000f00000000",
            INIT_23 => X"000000170000000000000021000000000000001c000000000000001c00000000",
            INIT_24 => X"0000000000000000000000170000000000000032000000000000002100000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000f00000000000000000000000000000000000000000000000100000000",
            INIT_27 => X"0000002a00000000000000000000000000000000000000000000001500000000",
            INIT_28 => X"00000000000000000000000e0000000000000022000000000000002a00000000",
            INIT_29 => X"0000001600000000000000120000000000000000000000000000000000000000",
            INIT_2A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000001900000000000000090000000000000000000000000000000000000000",
            INIT_2C => X"0000000e0000000000000010000000000000002f000000000000002800000000",
            INIT_2D => X"000000000000000000000011000000000000002e000000000000001900000000",
            INIT_2E => X"00000000000000000000001c000000000000001e000000000000000000000000",
            INIT_2F => X"0000001c0000000000000016000000000000001c000000000000000000000000",
            INIT_30 => X"0000002f00000000000000590000000000000066000000000000004e00000000",
            INIT_31 => X"000000620000000000000041000000000000002c000000000000001700000000",
            INIT_32 => X"0000003b00000000000000420000000000000068000000000000007200000000",
            INIT_33 => X"0000001f000000000000002d0000000000000027000000000000003e00000000",
            INIT_34 => X"00000041000000000000003b0000000000000020000000000000000000000000",
            INIT_35 => X"0000007c0000000000000079000000000000006c000000000000005b00000000",
            INIT_36 => X"0000009500000000000000830000000000000081000000000000008700000000",
            INIT_37 => X"000000320000000000000000000000000000002f000000000000004000000000",
            INIT_38 => X"0000007500000000000000710000000000000073000000000000007600000000",
            INIT_39 => X"000000840000000000000096000000000000008f000000000000008100000000",
            INIT_3A => X"0000008c000000000000009d00000000000000a7000000000000008500000000",
            INIT_3B => X"0000007c0000000000000058000000000000001b000000000000003900000000",
            INIT_3C => X"0000008600000000000000790000000000000076000000000000007e00000000",
            INIT_3D => X"000000a7000000000000008e0000000000000083000000000000008800000000",
            INIT_3E => X"0000006e0000000000000095000000000000009a000000000000007400000000",
            INIT_3F => X"0000006700000000000000650000000000000060000000000000004800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000085000000000000008e0000000000000082000000000000007800000000",
            INIT_41 => X"0000009700000000000000a600000000000000a2000000000000008900000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"000000000000000000000005000000000000003f000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "samplegold_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000130000000000000036000000000000001d000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000001a00000000000000220000000000000022000000000000004800000000",
            INIT_05 => X"0000004300000000000000140000000000000001000000000000000000000000",
            INIT_06 => X"0000001e00000000000000000000000000000002000000000000000100000000",
            INIT_07 => X"00000021000000000000001c0000000000000021000000000000003700000000",
            INIT_08 => X"0000000400000000000000030000000000000007000000000000000b00000000",
            INIT_09 => X"000000030000000000000068000000000000003e000000000000000800000000",
            INIT_0A => X"000000100000000000000057000000000000007d000000000000003d00000000",
            INIT_0B => X"0000003b00000000000000470000000000000000000000000000000e00000000",
            INIT_0C => X"0000000000000000000000190000000000000022000000000000001f00000000",
            INIT_0D => X"000000000000000000000000000000000000002d000000000000001c00000000",
            INIT_0E => X"00000023000000000000002e0000000000000007000000000000000000000000",
            INIT_0F => X"00000000000000000000000d000000000000007f000000000000001300000000",
            INIT_10 => X"000000330000000000000029000000000000001e000000000000001900000000",
            INIT_11 => X"0000001300000000000000000000000000000000000000000000001c00000000",
            INIT_12 => X"000000090000000000000025000000000000001b000000000000004c00000000",
            INIT_13 => X"0000002100000000000000170000000000000009000000000000006000000000",
            INIT_14 => X"00000034000000000000003d000000000000001d000000000000003800000000",
            INIT_15 => X"0000003c000000000000003e000000000000001b000000000000003000000000",
            INIT_16 => X"0000002c00000000000000010000000000000000000000000000000000000000",
            INIT_17 => X"00000009000000000000001d0000000000000003000000000000000f00000000",
            INIT_18 => X"000000120000000000000041000000000000003c000000000000000000000000",
            INIT_19 => X"0000000700000000000000000000000000000021000000000000003600000000",
            INIT_1A => X"00000000000000000000000d0000000000000032000000000000002700000000",
            INIT_1B => X"0000001d00000000000000180000000000000000000000000000000000000000",
            INIT_1C => X"0000005300000000000000140000000000000038000000000000002400000000",
            INIT_1D => X"000000560000000000000038000000000000000b000000000000001500000000",
            INIT_1E => X"0000000900000000000000000000000000000000000000000000001500000000",
            INIT_1F => X"0000004400000000000000000000000000000024000000000000003400000000",
            INIT_20 => X"00000097000000000000009b0000000000000007000000000000003900000000",
            INIT_21 => X"0000000700000000000000040000000000000051000000000000007700000000",
            INIT_22 => X"0000004800000000000000600000000000000045000000000000001d00000000",
            INIT_23 => X"00000028000000000000000e000000000000002c000000000000003000000000",
            INIT_24 => X"000000000000000000000000000000000000008e000000000000004300000000",
            INIT_25 => X"00000034000000000000001e0000000000000004000000000000000100000000",
            INIT_26 => X"00000047000000000000004a000000000000003d000000000000003c00000000",
            INIT_27 => X"0000005100000000000000180000000000000046000000000000004000000000",
            INIT_28 => X"00000035000000000000003a0000000000000000000000000000002400000000",
            INIT_29 => X"0000005100000000000000460000000000000039000000000000003400000000",
            INIT_2A => X"0000006500000000000000420000000000000041000000000000005600000000",
            INIT_2B => X"0000000000000000000000330000000000000044000000000000004100000000",
            INIT_2C => X"0000003900000000000000420000000000000040000000000000002400000000",
            INIT_2D => X"0000003700000000000000400000000000000043000000000000003b00000000",
            INIT_2E => X"0000003d000000000000001d0000000000000062000000000000004000000000",
            INIT_2F => X"0000001e0000000000000000000000000000003a000000000000004400000000",
            INIT_30 => X"0000005100000000000000370000000000000023000000000000002300000000",
            INIT_31 => X"0000007d00000000000000450000000000000041000000000000005400000000",
            INIT_32 => X"0000007b000000000000007d0000000000000037000000000000006000000000",
            INIT_33 => X"0000007900000000000000830000000000000083000000000000008000000000",
            INIT_34 => X"0000006c00000000000000850000000000000091000000000000008900000000",
            INIT_35 => X"000000710000000000000064000000000000005a000000000000005700000000",
            INIT_36 => X"0000008700000000000000880000000000000082000000000000006c00000000",
            INIT_37 => X"0000008b00000000000000750000000000000082000000000000008800000000",
            INIT_38 => X"0000001f0000000000000023000000000000004d000000000000007200000000",
            INIT_39 => X"0000006900000000000000510000000000000036000000000000002900000000",
            INIT_3A => X"0000008a00000000000000860000000000000056000000000000005600000000",
            INIT_3B => X"0000002f00000000000000490000000000000076000000000000008b00000000",
            INIT_3C => X"00000010000000000000001d0000000000000012000000000000001400000000",
            INIT_3D => X"00000030000000000000004c0000000000000029000000000000001800000000",
            INIT_3E => X"0000007700000000000000860000000000000085000000000000003300000000",
            INIT_3F => X"0000000d0000000000000019000000000000003c000000000000004a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000009000000000000001f000000000000002c000000000000001800000000",
            INIT_41 => X"0000003a000000000000001e0000000000000032000000000000000900000000",
            INIT_42 => X"0000005800000000000000570000000000000060000000000000008200000000",
            INIT_43 => X"00000008000000000000000c000000000000001c000000000000003d00000000",
            INIT_44 => X"0000000900000000000000110000000000000029000000000000003700000000",
            INIT_45 => X"0000007e00000000000000290000000000000022000000000000002100000000",
            INIT_46 => X"0000003c0000000000000038000000000000001c000000000000006300000000",
            INIT_47 => X"000000410000000000000007000000000000001a000000000000002f00000000",
            INIT_48 => X"0000000b000000000000000c0000000000000010000000000000001c00000000",
            INIT_49 => X"000000690000000000000055000000000000002c000000000000002200000000",
            INIT_4A => X"0000003000000000000000410000000000000033000000000000002f00000000",
            INIT_4B => X"0000001b00000000000000320000000000000015000000000000002000000000",
            INIT_4C => X"000000290000000000000021000000000000000c000000000000000e00000000",
            INIT_4D => X"0000003600000000000000560000000000000037000000000000002400000000",
            INIT_4E => X"0000001d00000000000000210000000000000039000000000000003300000000",
            INIT_4F => X"00000006000000000000001e0000000000000028000000000000002e00000000",
            INIT_50 => X"000000210000000000000026000000000000003b000000000000002100000000",
            INIT_51 => X"0000002600000000000000430000000000000013000000000000002000000000",
            INIT_52 => X"00000053000000000000001a0000000000000020000000000000002b00000000",
            INIT_53 => X"0000002600000000000000080000000000000011000000000000002100000000",
            INIT_54 => X"0000001e00000000000000250000000000000024000000000000006100000000",
            INIT_55 => X"0000001c000000000000001f0000000000000028000000000000000b00000000",
            INIT_56 => X"0000000a00000000000000190000000000000031000000000000002e00000000",
            INIT_57 => X"00000072000000000000005b0000000000000009000000000000000000000000",
            INIT_58 => X"0000000c0000000000000025000000000000002e000000000000000900000000",
            INIT_59 => X"0000000e000000000000000b0000000000000025000000000000003000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000038000000000000003f000000000000001f000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000044000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"00000000000000000000000b0000000000000011000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_71 => X"0000000a000000000000001b0000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000002f0000000000000014000000000000000000000000",
            INIT_73 => X"0000000200000000000000560000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_75 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000001400000000000000000000000000000035000000000000000000000000",
            INIT_79 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_7E => X"0000000d000000000000006b000000000000001a000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "samplegold_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_01 => X"0000002100000000000000060000000000000000000000000000000000000000",
            INIT_02 => X"000000030000000000000000000000000000003a000000000000000000000000",
            INIT_03 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000280000000000000012000000000000000f000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000021000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000017000000000000000800000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000003000000000000005c00000000",
            INIT_0B => X"0000002300000000000000240000000000000031000000000000001300000000",
            INIT_0C => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_0E => X"0000002100000000000000060000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000006000000000000001f00000000",
            INIT_10 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_13 => X"0000000300000000000000150000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000025000000000000008800000000",
            INIT_15 => X"00000041000000000000004d000000000000004a000000000000005800000000",
            INIT_16 => X"0000000600000000000000000000000000000001000000000000000e00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000001f000000000000001c0000000000000008000000000000006c00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000700000000000000000000000000000000000000000000000700000000",
            INIT_1C => X"000000000000000000000000000000000000002e000000000000007000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000030000000000000016000000000000000800000000",
            INIT_1F => X"0000001f00000000000000010000000000000000000000000000003f00000000",
            INIT_20 => X"0000001d0000000000000024000000000000001c000000000000005a00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000300000000000000000000000000000000000000000000000300000000",
            INIT_24 => X"0000000200000000000000050000000000000000000000000000000500000000",
            INIT_25 => X"000000000000000000000009000000000000000b000000000000000500000000",
            INIT_26 => X"00000000000000000000000b000000000000000a000000000000000000000000",
            INIT_27 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_28 => X"000000190000000000000014000000000000002e000000000000000000000000",
            INIT_29 => X"000000000000000000000015000000000000000a000000000000000000000000",
            INIT_2A => X"00000000000000000000002e0000000000000006000000000000000000000000",
            INIT_2B => X"0000000000000000000000010000000000000003000000000000000300000000",
            INIT_2C => X"0000000000000000000000000000000000000005000000000000003400000000",
            INIT_2D => X"0000000000000000000000300000000000000000000000000000001c00000000",
            INIT_2E => X"0000000b0000000000000000000000000000005c000000000000000000000000",
            INIT_2F => X"000000090000000000000000000000000000001f000000000000000000000000",
            INIT_30 => X"000000390000000000000000000000000000000e000000000000002400000000",
            INIT_31 => X"00000000000000000000002c0000000000000021000000000000001200000000",
            INIT_32 => X"0000000000000000000000410000000000000000000000000000003e00000000",
            INIT_33 => X"0000003a00000000000000380000000000000026000000000000000000000000",
            INIT_34 => X"0000004d00000000000000000000000000000000000000000000002400000000",
            INIT_35 => X"0000005b00000000000000000000000000000027000000000000000000000000",
            INIT_36 => X"0000000000000000000000500000000000000050000000000000000000000000",
            INIT_37 => X"00000046000000000000001b000000000000002a000000000000001200000000",
            INIT_38 => X"00000000000000000000004a000000000000005c000000000000000000000000",
            INIT_39 => X"0000002d000000000000004d000000000000001e000000000000001100000000",
            INIT_3A => X"0000000000000000000000000000000000000042000000000000000700000000",
            INIT_3B => X"00000000000000000000003b0000000000000030000000000000000100000000",
            INIT_3C => X"0000000000000000000000000000000000000038000000000000005100000000",
            INIT_3D => X"000000300000000000000000000000000000004d000000000000002600000000",
            INIT_3E => X"0000006700000000000000000000000000000000000000000000001100000000",
            INIT_3F => X"0000002c0000000000000000000000000000001e000000000000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000400000000000000030000000000000000000000000000003c00000000",
            INIT_41 => X"0000000000000000000000980000000000000000000000000000004100000000",
            INIT_42 => X"0000000f000000000000000b0000000000000000000000000000005100000000",
            INIT_43 => X"000000440000000000000000000000000000002b000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000003800000000000000000000000000000075000000000000000000000000",
            INIT_46 => X"0000003700000000000000030000000000000000000000000000002200000000",
            INIT_47 => X"0000000000000000000000000000000000000038000000000000001600000000",
            INIT_48 => X"0000000200000000000000000000000000000011000000000000000000000000",
            INIT_49 => X"00000033000000000000005f0000000000000000000000000000006100000000",
            INIT_4A => X"00000024000000000000004c000000000000000f000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000300000000000000000000000000000000000000000000000c00000000",
            INIT_4D => X"00000000000000000000003f00000000000000a3000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_4F => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000003000000000000000000000000000000000000000000000001f00000000",
            INIT_51 => X"0000000000000000000000050000000000000000000000000000007500000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000001f000000000000003e0000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000002000000000000000d000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000002b0000000000000028000000000000000000000000",
            INIT_58 => X"0000000000000000000000110000000000000000000000000000000c00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000001200000000000000000000000000000000000000000000000f00000000",
            INIT_5B => X"0000006f00000000000000700000000000000065000000000000003100000000",
            INIT_5C => X"00000074000000000000006b000000000000006b000000000000006f00000000",
            INIT_5D => X"000000460000000000000051000000000000006b000000000000007900000000",
            INIT_5E => X"0000005f0000000000000064000000000000005d000000000000004f00000000",
            INIT_5F => X"0000007100000000000000730000000000000077000000000000006e00000000",
            INIT_60 => X"0000005e000000000000006a000000000000007b000000000000006c00000000",
            INIT_61 => X"000000280000000000000024000000000000002a000000000000003a00000000",
            INIT_62 => X"00000044000000000000005a0000000000000047000000000000003200000000",
            INIT_63 => X"0000006e0000000000000075000000000000006f000000000000004600000000",
            INIT_64 => X"0000001e00000000000000250000000000000041000000000000005400000000",
            INIT_65 => X"0000002000000000000000250000000000000025000000000000002600000000",
            INIT_66 => X"00000038000000000000002d0000000000000050000000000000002000000000",
            INIT_67 => X"0000003e0000000000000063000000000000006e000000000000006800000000",
            INIT_68 => X"0000001900000000000000190000000000000020000000000000003e00000000",
            INIT_69 => X"00000018000000000000001c0000000000000022000000000000003800000000",
            INIT_6A => X"00000064000000000000003e0000000000000023000000000000003700000000",
            INIT_6B => X"00000041000000000000004f0000000000000066000000000000004a00000000",
            INIT_6C => X"0000003a000000000000001d000000000000001b000000000000002e00000000",
            INIT_6D => X"0000001f000000000000001f0000000000000023000000000000002e00000000",
            INIT_6E => X"00000048000000000000006a0000000000000033000000000000000f00000000",
            INIT_6F => X"0000003600000000000000530000000000000041000000000000003300000000",
            INIT_70 => X"0000002300000000000000360000000000000021000000000000002b00000000",
            INIT_71 => X"0000001c0000000000000022000000000000001c000000000000001c00000000",
            INIT_72 => X"0000003500000000000000610000000000000046000000000000003000000000",
            INIT_73 => X"0000002b00000000000000350000000000000039000000000000004000000000",
            INIT_74 => X"0000001a0000000000000024000000000000002d000000000000002000000000",
            INIT_75 => X"000000350000000000000027000000000000002b000000000000001c00000000",
            INIT_76 => X"000000310000000000000026000000000000004a000000000000002600000000",
            INIT_77 => X"00000034000000000000002c0000000000000026000000000000003100000000",
            INIT_78 => X"0000002700000000000000150000000000000024000000000000003100000000",
            INIT_79 => X"0000001c00000000000000270000000000000028000000000000004800000000",
            INIT_7A => X"000000300000000000000021000000000000002f000000000000002b00000000",
            INIT_7B => X"0000001c000000000000003a0000000000000023000000000000002900000000",
            INIT_7C => X"0000005e000000000000003e0000000000000019000000000000001c00000000",
            INIT_7D => X"0000001a00000000000000280000000000000025000000000000002a00000000",
            INIT_7E => X"0000003a000000000000002a0000000000000023000000000000002600000000",
            INIT_7F => X"000000080000000000000014000000000000001f000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "samplegold_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001500000000000000570000000000000053000000000000002200000000",
            INIT_01 => X"0000004800000000000000280000000000000026000000000000002800000000",
            INIT_02 => X"0000000f0000000000000014000000000000000f000000000000002000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_04 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000000c0000000000000037000000000000002400000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_19 => X"0000000100000000000000090000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_1C => X"0000000000000000000000030000000000000018000000000000000000000000",
            INIT_1D => X"0000002200000000000000250000000000000031000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_20 => X"00000014000000000000000a000000000000000b000000000000000600000000",
            INIT_21 => X"00000015000000000000001a0000000000000023000000000000003b00000000",
            INIT_22 => X"000000230000000000000021000000000000000c000000000000000000000000",
            INIT_23 => X"0000001800000000000000220000000000000015000000000000000000000000",
            INIT_24 => X"00000032000000000000000e000000000000000e000000000000002000000000",
            INIT_25 => X"0000000000000000000000140000000000000006000000000000002500000000",
            INIT_26 => X"00000000000000000000004b0000000000000037000000000000000000000000",
            INIT_27 => X"0000002f0000000000000044000000000000006b000000000000000500000000",
            INIT_28 => X"00000032000000000000004b0000000000000000000000000000001500000000",
            INIT_29 => X"000000000000000000000013000000000000001f000000000000001800000000",
            INIT_2A => X"00000000000000000000000e000000000000003d000000000000003800000000",
            INIT_2B => X"000000290000000000000047000000000000003f000000000000003100000000",
            INIT_2C => X"000000110000000000000031000000000000005a000000000000000e00000000",
            INIT_2D => X"00000042000000000000000b0000000000000023000000000000001900000000",
            INIT_2E => X"0000001b0000000000000000000000000000000a000000000000004d00000000",
            INIT_2F => X"0000001a0000000000000038000000000000003e000000000000005800000000",
            INIT_30 => X"0000002300000000000000140000000000000039000000000000004700000000",
            INIT_31 => X"0000006300000000000000530000000000000010000000000000002400000000",
            INIT_32 => X"0000003c000000000000000d0000000000000039000000000000001e00000000",
            INIT_33 => X"0000001000000000000000220000000000000019000000000000002100000000",
            INIT_34 => X"0000001600000000000000180000000000000015000000000000002200000000",
            INIT_35 => X"0000002d00000000000000650000000000000069000000000000000000000000",
            INIT_36 => X"000000360000000000000017000000000000001c000000000000004a00000000",
            INIT_37 => X"0000001400000000000000260000000000000013000000000000002d00000000",
            INIT_38 => X"000000000000000000000009000000000000000e000000000000000700000000",
            INIT_39 => X"0000007000000000000000330000000000000058000000000000006f00000000",
            INIT_3A => X"0000005f00000000000000510000000000000016000000000000003c00000000",
            INIT_3B => X"0000001c00000000000000100000000000000011000000000000002700000000",
            INIT_3C => X"00000074000000000000001d000000000000002b000000000000002200000000",
            INIT_3D => X"000000670000000000000082000000000000004c000000000000007a00000000",
            INIT_3E => X"0000003c000000000000004a000000000000004b000000000000005000000000",
            INIT_3F => X"00000052000000000000004a0000000000000043000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000066000000000000004d0000000000000050000000000000005300000000",
            INIT_41 => X"00000044000000000000004c0000000000000071000000000000007600000000",
            INIT_42 => X"0000004500000000000000400000000000000041000000000000004100000000",
            INIT_43 => X"0000005c00000000000000550000000000000050000000000000004e00000000",
            INIT_44 => X"00000073000000000000004b0000000000000058000000000000006000000000",
            INIT_45 => X"00000042000000000000004b0000000000000046000000000000007500000000",
            INIT_46 => X"00000055000000000000004d0000000000000047000000000000003f00000000",
            INIT_47 => X"000000650000000000000061000000000000005a000000000000005d00000000",
            INIT_48 => X"0000005a000000000000004f0000000000000056000000000000005600000000",
            INIT_49 => X"0000004b0000000000000053000000000000004d000000000000003f00000000",
            INIT_4A => X"00000054000000000000004c0000000000000050000000000000004c00000000",
            INIT_4B => X"0000003800000000000000490000000000000062000000000000006600000000",
            INIT_4C => X"000000380000000000000039000000000000003a000000000000003800000000",
            INIT_4D => X"0000003b00000000000000490000000000000042000000000000003500000000",
            INIT_4E => X"0000002b00000000000000270000000000000020000000000000002600000000",
            INIT_4F => X"00000043000000000000003a000000000000002c000000000000003100000000",
            INIT_50 => X"000000170000000000000038000000000000003c000000000000003d00000000",
            INIT_51 => X"00000000000000000000001e000000000000002d000000000000003100000000",
            INIT_52 => X"0000002100000000000000080000000000000000000000000000000000000000",
            INIT_53 => X"0000004100000000000000320000000000000011000000000000002800000000",
            INIT_54 => X"0000001000000000000000230000000000000040000000000000004200000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000003f000000000000003b0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000013000000000000002400000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_5B => X"00000000000000000000001e0000000000000027000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000026000000000000002500000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "samplegold_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000008000000000000000800000000000000080000000000000008200000000",
            INIT_05 => X"0000008100000000000000820000000000000082000000000000008100000000",
            INIT_06 => X"0000008000000000000000810000000000000080000000000000008200000000",
            INIT_07 => X"0000008500000000000000800000000000000080000000000000008000000000",
            INIT_08 => X"0000008200000000000000820000000000000082000000000000008200000000",
            INIT_09 => X"0000008000000000000000810000000000000082000000000000008200000000",
            INIT_0A => X"00000082000000000000007e000000000000008b000000000000009300000000",
            INIT_0B => X"00000087000000000000008a0000000000000081000000000000008100000000",
            INIT_0C => X"0000008300000000000000810000000000000082000000000000008300000000",
            INIT_0D => X"0000008300000000000000a1000000000000008b000000000000008600000000",
            INIT_0E => X"0000008300000000000000830000000000000088000000000000007400000000",
            INIT_0F => X"0000007f000000000000007a0000000000000073000000000000008300000000",
            INIT_10 => X"0000008100000000000000860000000000000085000000000000008300000000",
            INIT_11 => X"0000001f0000000000000038000000000000004d000000000000007c00000000",
            INIT_12 => X"00000081000000000000007f000000000000007f000000000000003f00000000",
            INIT_13 => X"0000008a000000000000008100000000000000b400000000000000b400000000",
            INIT_14 => X"00000078000000000000005f0000000000000078000000000000008700000000",
            INIT_15 => X"000000b500000000000000a10000000000000080000000000000006e00000000",
            INIT_16 => X"0000000d000000000000008100000000000000a700000000000000ba00000000",
            INIT_17 => X"00000096000000000000009c0000000000000054000000000000000b00000000",
            INIT_18 => X"000000b500000000000000cb00000000000000d400000000000000d100000000",
            INIT_19 => X"00000011000000000000001c000000000000003e000000000000007c00000000",
            INIT_1A => X"000000bb00000000000000b1000000000000007d000000000000001a00000000",
            INIT_1B => X"0000004c0000000000000052000000000000005e000000000000009800000000",
            INIT_1C => X"0000008a000000000000001b0000000000000000000000000000000f00000000",
            INIT_1D => X"000000b000000000000000b800000000000000c600000000000000b400000000",
            INIT_1E => X"0000004c0000000000000000000000000000002a00000000000000ab00000000",
            INIT_1F => X"000000000000000000000012000000000000006e000000000000006100000000",
            INIT_20 => X"00000044000000000000007c000000000000009a000000000000006000000000",
            INIT_21 => X"0000002a0000000000000009000000000000000c000000000000001800000000",
            INIT_22 => X"0000002c000000000000000f000000000000003c000000000000000000000000",
            INIT_23 => X"0000008a0000000000000098000000000000008e000000000000006900000000",
            INIT_24 => X"0000007c000000000000006e000000000000006f000000000000004e00000000",
            INIT_25 => X"0000004e0000000000000086000000000000009e000000000000009000000000",
            INIT_26 => X"000000a300000000000000ac00000000000000ab00000000000000b200000000",
            INIT_27 => X"0000005b000000000000005b0000000000000076000000000000008f00000000",
            INIT_28 => X"0000002f00000000000000500000000000000056000000000000005400000000",
            INIT_29 => X"0000003b000000000000003d000000000000003b000000000000003400000000",
            INIT_2A => X"000000930000000000000080000000000000006d000000000000005400000000",
            INIT_2B => X"0000006e000000000000007d0000000000000090000000000000009500000000",
            INIT_2C => X"000000110000000000000022000000000000003a000000000000005300000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000001b000000000000003b000000000000002d000000000000000000000000",
            INIT_31 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_32 => X"00000091000000000000002f0000000000000000000000000000000000000000",
            INIT_33 => X"0000005b000000000000007a000000000000006d000000000000006e00000000",
            INIT_34 => X"0000000000000000000000220000000000000014000000000000000e00000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"00000062000000000000003b0000000000000000000000000000000000000000",
            INIT_37 => X"0000001e00000000000000000000000000000000000000000000002300000000",
            INIT_38 => X"000000000000000000000002000000000000003e000000000000002600000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"00000028000000000000001e0000000000000021000000000000001100000000",
            INIT_3C => X"0000000e000000000000000e000000000000000d000000000000003c00000000",
            INIT_3D => X"0000000e000000000000000e000000000000000e000000000000000e00000000",
            INIT_3E => X"0000000b000000000000000e0000000000000010000000000000000e00000000",
            INIT_3F => X"0000000e000000000000000e000000000000000e000000000000000d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000d000000000000000d000000000000000d000000000000000c00000000",
            INIT_41 => X"0000000e000000000000000e000000000000000d000000000000000d00000000",
            INIT_42 => X"0000000e00000000000000050000000000000000000000000000000c00000000",
            INIT_43 => X"0000000d000000000000000d000000000000000d000000000000000d00000000",
            INIT_44 => X"0000000e000000000000000d000000000000000e000000000000000e00000000",
            INIT_45 => X"000000000000000000000001000000000000000d000000000000000d00000000",
            INIT_46 => X"0000000c000000000000000f000000000000000e000000000000000000000000",
            INIT_47 => X"000000070000000000000007000000000000000d000000000000000e00000000",
            INIT_48 => X"00000000000000000000000e000000000000000f000000000000000c00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_4A => X"0000000a0000000000000007000000000000001b000000000000000000000000",
            INIT_4B => X"0000000e00000000000000000000000000000000000000000000000c00000000",
            INIT_4C => X"000000170000000000000003000000000000000e000000000000000e00000000",
            INIT_4D => X"000000000000000000000001000000000000000c000000000000000800000000",
            INIT_4E => X"00000009000000000000000e0000000000000000000000000000000000000000",
            INIT_4F => X"0000000c000000000000000f0000000000000011000000000000000a00000000",
            INIT_50 => X"0000000300000000000000010000000000000000000000000000000c00000000",
            INIT_51 => X"0000000500000000000000000000000000000000000000000000000300000000",
            INIT_52 => X"00000000000000000000000a0000000000000021000000000000000000000000",
            INIT_53 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_54 => X"0000002100000000000000040000000000000000000000000000000000000000",
            INIT_55 => X"0000000300000000000000000000000000000001000000000000000800000000",
            INIT_56 => X"0000001300000000000000060000000000000008000000000000000000000000",
            INIT_57 => X"000000050000000000000001000000000000001b000000000000000500000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_59 => X"0000000600000000000000040000000000000000000000000000000000000000",
            INIT_5A => X"0000001300000000000000040000000000000050000000000000001200000000",
            INIT_5B => X"000000010000000000000000000000000000000c000000000000001700000000",
            INIT_5C => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000002c000000000000000c000000000000000f000000000000000000000000",
            INIT_66 => X"000000170000000000000013000000000000000f000000000000000b00000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_68 => X"00000010000000000000000f0000000000000014000000000000000100000000",
            INIT_69 => X"0000001a000000000000001f0000000000000014000000000000002000000000",
            INIT_6A => X"0000004d000000000000001a0000000000000018000000000000001400000000",
            INIT_6B => X"0000002300000000000000340000000000000036000000000000002300000000",
            INIT_6C => X"0000002300000000000000240000000000000028000000000000001c00000000",
            INIT_6D => X"0000001a0000000000000020000000000000001e000000000000000000000000",
            INIT_6E => X"0000005a0000000000000052000000000000001e000000000000001d00000000",
            INIT_6F => X"00000036000000000000003c0000000000000038000000000000005200000000",
            INIT_70 => X"00000004000000000000001d0000000000000022000000000000002200000000",
            INIT_71 => X"00000020000000000000001f0000000000000023000000000000002400000000",
            INIT_72 => X"0000003d00000000000000320000000000000036000000000000001f00000000",
            INIT_73 => X"0000002300000000000000220000000000000030000000000000004500000000",
            INIT_74 => X"000000540000000000000054000000000000001b000000000000002100000000",
            INIT_75 => X"0000005400000000000000540000000000000054000000000000005400000000",
            INIT_76 => X"0000005400000000000000520000000000000053000000000000005400000000",
            INIT_77 => X"0000005400000000000000540000000000000054000000000000005600000000",
            INIT_78 => X"0000005500000000000000550000000000000056000000000000005400000000",
            INIT_79 => X"0000005500000000000000550000000000000055000000000000005500000000",
            INIT_7A => X"0000004f00000000000000560000000000000056000000000000005400000000",
            INIT_7B => X"0000005500000000000000550000000000000055000000000000005600000000",
            INIT_7C => X"0000005500000000000000550000000000000054000000000000005300000000",
            INIT_7D => X"0000005700000000000000550000000000000057000000000000005500000000",
            INIT_7E => X"0000004b000000000000003e000000000000004d000000000000005500000000",
            INIT_7F => X"0000005b00000000000000560000000000000055000000000000005600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "samplegold_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005600000000000000550000000000000056000000000000005900000000",
            INIT_01 => X"000000430000000000000052000000000000004d000000000000005600000000",
            INIT_02 => X"0000005b000000000000004a000000000000003b000000000000004300000000",
            INIT_03 => X"0000004900000000000000460000000000000057000000000000005800000000",
            INIT_04 => X"0000005700000000000000570000000000000052000000000000005200000000",
            INIT_05 => X"0000005900000000000000510000000000000057000000000000004b00000000",
            INIT_06 => X"0000004c0000000000000049000000000000004a000000000000005400000000",
            INIT_07 => X"00000047000000000000002b000000000000002c000000000000005800000000",
            INIT_08 => X"00000047000000000000004f000000000000004d000000000000004900000000",
            INIT_09 => X"000000480000000000000058000000000000004f000000000000004a00000000",
            INIT_0A => X"0000005900000000000000360000000000000032000000000000003b00000000",
            INIT_0B => X"0000003b000000000000004e000000000000003d000000000000003800000000",
            INIT_0C => X"0000001f0000000000000012000000000000001a000000000000004c00000000",
            INIT_0D => X"0000004600000000000000500000000000000055000000000000003f00000000",
            INIT_0E => X"00000000000000000000004a000000000000003e000000000000004500000000",
            INIT_0F => X"0000004a000000000000002b000000000000000d000000000000000d00000000",
            INIT_10 => X"0000003f0000000000000039000000000000002a000000000000003400000000",
            INIT_11 => X"0000002400000000000000290000000000000033000000000000004100000000",
            INIT_12 => X"0000004600000000000000000000000000000033000000000000003100000000",
            INIT_13 => X"00000057000000000000004d0000000000000039000000000000002f00000000",
            INIT_14 => X"0000003d0000000000000035000000000000004e000000000000005b00000000",
            INIT_15 => X"000000370000000000000037000000000000003d000000000000003f00000000",
            INIT_16 => X"0000004e0000000000000047000000000000001a000000000000003900000000",
            INIT_17 => X"0000005200000000000000580000000000000054000000000000005700000000",
            INIT_18 => X"0000003300000000000000330000000000000045000000000000004400000000",
            INIT_19 => X"0000001b0000000000000018000000000000001f000000000000002900000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000002300000000000000200000000000000009000000000000000000000000",
            INIT_1C => X"0000000d0000000000000013000000000000001a000000000000001f00000000",
            INIT_1D => X"00000000000000000000000d000000000000000f000000000000000c00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000000000000000000000b000000000000000200000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002300000000000000090000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000011d0000000000000027000000000000000f000000000000000200000000",
            INIT_2D => X"0000011c000000000000011c000000000000011c000000000000011c00000000",
            INIT_2E => X"0000011b000000000000011c000000000000011d000000000000011d00000000",
            INIT_2F => X"0000011c000000000000011c000000000000011f000000000000011c00000000",
            INIT_30 => X"0000011d000000000000011e000000000000011d000000000000011c00000000",
            INIT_31 => X"0000011c000000000000011c000000000000011d000000000000011d00000000",
            INIT_32 => X"000001040000000000000117000000000000011c000000000000011d00000000",
            INIT_33 => X"0000011d000000000000011d0000000000000119000000000000010d00000000",
            INIT_34 => X"0000011f000000000000011d000000000000011d000000000000011e00000000",
            INIT_35 => X"0000011d000000000000011d000000000000011e000000000000011e00000000",
            INIT_36 => X"000000e100000000000000ef00000000000000fe000000000000010f00000000",
            INIT_37 => X"00000120000000000000011e000000000000011e000000000000011b00000000",
            INIT_38 => X"0000011f000000000000011c000000000000011b000000000000011700000000",
            INIT_39 => X"0000011300000000000001140000000000000113000000000000012000000000",
            INIT_3A => X"000000fb00000000000000e800000000000000f5000000000000010000000000",
            INIT_3B => X"000000cf0000000000000121000000000000011f000000000000011f00000000",
            INIT_3C => X"0000011e000000000000011b000000000000011d00000000000000e100000000",
            INIT_3D => X"0000011a000000000000011a0000000000000109000000000000011800000000",
            INIT_3E => X"000000e900000000000000fb000000000000010a000000000000011d00000000",
            INIT_3F => X"000000ee00000000000000e30000000000000124000000000000010b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000e1000000000000010e00000000000000f100000000000000fb00000000",
            INIT_41 => X"00000122000000000000011b000000000000010500000000000000f800000000",
            INIT_42 => X"000000e600000000000000d900000000000000ed00000000000000ff00000000",
            INIT_43 => X"000000e700000000000000ca00000000000000ba000000000000011e00000000",
            INIT_44 => X"0000007f000000000000009400000000000000f1000000000000010000000000",
            INIT_45 => X"00000108000000000000010f00000000000000da00000000000000aa00000000",
            INIT_46 => X"0000010100000000000000f100000000000000f700000000000000f900000000",
            INIT_47 => X"000000cb000000000000009a00000000000000a3000000000000006e00000000",
            INIT_48 => X"000000de00000000000000e700000000000000ea000000000000010600000000",
            INIT_49 => X"000000a400000000000000b200000000000000d200000000000000de00000000",
            INIT_4A => X"0000007f00000000000000ce00000000000000c400000000000000a900000000",
            INIT_4B => X"0000010a00000000000000e700000000000000dc00000000000000f000000000",
            INIT_4C => X"000000eb00000000000000ff0000000000000110000000000000011100000000",
            INIT_4D => X"000000d700000000000000de00000000000000f300000000000000de00000000",
            INIT_4E => X"000000dd00000000000000a600000000000000d300000000000000d600000000",
            INIT_4F => X"000000ea00000000000000ea00000000000000e700000000000000e200000000",
            INIT_50 => X"000000b400000000000000c300000000000000c700000000000000e100000000",
            INIT_51 => X"00000092000000000000009200000000000000a100000000000000ac00000000",
            INIT_52 => X"00000047000000000000004a000000000000002700000000000000a700000000",
            INIT_53 => X"00000089000000000000006f0000000000000056000000000000004d00000000",
            INIT_54 => X"000000750000000000000081000000000000008f000000000000008e00000000",
            INIT_55 => X"0000009300000000000000870000000000000089000000000000007400000000",
            INIT_56 => X"0000000200000000000000300000000000000011000000000000000000000000",
            INIT_57 => X"0000004800000000000000670000000000000000000000000000000000000000",
            INIT_58 => X"0000007500000000000000650000000000000051000000000000004a00000000",
            INIT_59 => X"0000000000000000000000950000000000000090000000000000007d00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000009300000000000000ab000000000000003b000000000000000000000000",
            INIT_5C => X"00000062000000000000006a0000000000000066000000000000007e00000000",
            INIT_5D => X"00000000000000000000000400000000000000b0000000000000008000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000001a0000000000000004000000000000000e000000000000000000000000",
            INIT_60 => X"000000920000000000000079000000000000004e000000000000002900000000",
            INIT_61 => X"000000000000000000000000000000000000001700000000000000c500000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000660000000000000037000000000000000a000000000000000000000000",
            INIT_64 => X"000000cf00000000000000a30000000000000084000000000000007500000000",
            INIT_65 => X"0000003c000000000000003c000000000000003c000000000000003d00000000",
            INIT_66 => X"0000003d000000000000003d000000000000003d000000000000003c00000000",
            INIT_67 => X"0000003d000000000000003b000000000000003e000000000000003e00000000",
            INIT_68 => X"0000003f000000000000003c000000000000003c000000000000003d00000000",
            INIT_69 => X"0000003e000000000000003e000000000000003d000000000000003d00000000",
            INIT_6A => X"00000042000000000000003f000000000000003e000000000000003e00000000",
            INIT_6B => X"0000003d0000000000000038000000000000004e000000000000005e00000000",
            INIT_6C => X"000000400000000000000043000000000000003d000000000000003d00000000",
            INIT_6D => X"0000003f000000000000003b000000000000003e000000000000003e00000000",
            INIT_6E => X"0000005500000000000000650000000000000052000000000000004000000000",
            INIT_6F => X"0000003f000000000000003f0000000000000040000000000000003600000000",
            INIT_70 => X"0000003d00000000000000390000000000000032000000000000003e00000000",
            INIT_71 => X"0000003f0000000000000053000000000000003d000000000000003f00000000",
            INIT_72 => X"00000000000000000000000c0000000000000019000000000000004800000000",
            INIT_73 => X"0000003f000000000000003f000000000000003f000000000000000300000000",
            INIT_74 => X"0000004400000000000000470000000000000075000000000000008500000000",
            INIT_75 => X"0000003a00000000000000250000000000000044000000000000004100000000",
            INIT_76 => X"00000079000000000000005a0000000000000039000000000000002900000000",
            INIT_77 => X"000000000000000000000041000000000000005a000000000000008000000000",
            INIT_78 => X"0000005c000000000000005b000000000000001d000000000000000000000000",
            INIT_79 => X"00000062000000000000007c0000000000000089000000000000008500000000",
            INIT_7A => X"0000000000000000000000000000000000000016000000000000004900000000",
            INIT_7B => X"00000077000000000000007f0000000000000039000000000000000000000000",
            INIT_7C => X"0000004b0000000000000034000000000000002a000000000000005800000000",
            INIT_7D => X"0000003f00000000000000000000000000000000000000000000001000000000",
            INIT_7E => X"000000710000000000000070000000000000007c000000000000006500000000",
            INIT_7F => X"0000003d0000000000000000000000000000000c000000000000005e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "samplegold_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000003f000000000000003200000000",
            INIT_01 => X"00000037000000000000005c000000000000006d000000000000003100000000",
            INIT_02 => X"0000000000000000000000000000000000000001000000000000001200000000",
            INIT_03 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_04 => X"0000004f0000000000000056000000000000004e000000000000001f00000000",
            INIT_05 => X"0000003d000000000000002c0000000000000028000000000000001600000000",
            INIT_06 => X"0000000e000000000000005c000000000000006a000000000000005100000000",
            INIT_07 => X"0000004d00000000000000540000000000000058000000000000006200000000",
            INIT_08 => X"0000002500000000000000260000000000000036000000000000004300000000",
            INIT_09 => X"00000011000000000000002c0000000000000027000000000000002600000000",
            INIT_0A => X"00000044000000000000004e000000000000001c000000000000001700000000",
            INIT_0B => X"0000006700000000000000650000000000000058000000000000004800000000",
            INIT_0C => X"00000042000000000000004b0000000000000051000000000000005800000000",
            INIT_0D => X"0000000000000000000000050000000000000020000000000000003300000000",
            INIT_0E => X"00000011000000000000000d0000000000000031000000000000001300000000",
            INIT_0F => X"00000000000000000000000f0000000000000015000000000000000e00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000013000000000000002e0000000000000008000000000000000000000000",
            INIT_12 => X"0000003700000000000000360000000000000021000000000000001d00000000",
            INIT_13 => X"0000002600000000000000000000000000000019000000000000002100000000",
            INIT_14 => X"0000005800000000000000560000000000000026000000000000000b00000000",
            INIT_15 => X"0000003e00000000000000170000000000000019000000000000001c00000000",
            INIT_16 => X"00000018000000000000001c0000000000000019000000000000001700000000",
            INIT_17 => X"0000004b00000000000000130000000000000000000000000000001800000000",
            INIT_18 => X"0000003100000000000000030000000000000000000000000000003700000000",
            INIT_19 => X"000000180000000000000054000000000000002a000000000000002800000000",
            INIT_1A => X"0000001000000000000000110000000000000016000000000000001600000000",
            INIT_1B => X"0000000000000000000000000000000000000019000000000000000a00000000",
            INIT_1C => X"00000028000000000000002d000000000000003d000000000000002a00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000000000000000000004000000000000000d000000000000000f00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000900000000000000460000000000000046000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000000000000000000002e0000000000000042000000000000003300000000",
            INIT_30 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000005d00000000000000710000000000000055000000000000000c00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000003200000000",
            INIT_33 => X"0000006000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000031000000000000006100000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000004d00000000000000450000000000000029000000000000000000000000",
            INIT_37 => X"00000000000000000000001d0000000000000030000000000000003f00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"00000004000000000000001e0000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000013000000000000000f0000000000000000000000000000001800000000",
            INIT_3E => X"00000025000000000000003f000000000000003c000000000000001f00000000",
            INIT_3F => X"0000004e0000000000000052000000000000005a000000000000002c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000019000000000000002c000000000000003c00000000",
            INIT_41 => X"0000001400000000000000140000000000000000000000000000000700000000",
            INIT_42 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000006800000000000000520000000000000034000000000000002800000000",
            INIT_44 => X"00000059000000000000006a0000000000000072000000000000007400000000",
            INIT_45 => X"0000000000000000000000190000000000000032000000000000004a00000000",
            INIT_46 => X"00000016000000000000000e0000000000000000000000000000000000000000",
            INIT_47 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000002e00000000000000040000000000000000000000000000000000000000",
            INIT_4B => X"0000004100000000000000010000000000000008000000000000001c00000000",
            INIT_4C => X"0000003500000000000000190000000000000011000000000000003c00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_4E => X"0000000500000000000000040000000000000000000000000000000000000000",
            INIT_4F => X"0000002d00000000000000020000000000000002000000000000000200000000",
            INIT_50 => X"000000000000000000000000000000000000000e000000000000003600000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"00000042000000000000002b0000000000000000000000000000000000000000",
            INIT_60 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_63 => X"0000000000000000000000390000000000000000000000000000000000000000",
            INIT_64 => X"0000002f00000000000000040000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000004e00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_67 => X"0000005d00000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000140000000000000000000000000000000500000000",
            INIT_69 => X"0000001e00000000000000000000000000000008000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000002f000000000000002000000000",
            INIT_6B => X"0000000800000000000000620000000000000000000000000000000000000000",
            INIT_6C => X"0000002c000000000000001a0000000000000042000000000000000600000000",
            INIT_6D => X"0000003900000000000000160000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000005800000000",
            INIT_6F => X"0000006500000000000000410000000000000000000000000000000900000000",
            INIT_70 => X"0000000000000000000000620000000000000000000000000000003c00000000",
            INIT_71 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_72 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"00000000000000000000011a0000000000000018000000000000000500000000",
            INIT_74 => X"0000000000000000000000100000000000000013000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000300000000000000080000000000000000000000000000000b00000000",
            INIT_77 => X"0000001000000000000000070000000000000068000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000009000000000000000700000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000001e000000000000000a0000000000000002000000000000000000000000",
            INIT_7B => X"0000000800000000000000000000000000000027000000000000000000000000",
            INIT_7C => X"000000140000000000000018000000000000002b000000000000001900000000",
            INIT_7D => X"0000000f00000000000000000000000000000000000000000000000500000000",
            INIT_7E => X"0000000000000000000000200000000000000003000000000000002000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000004e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "samplegold_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000007d000000000000001b00000000",
            INIT_01 => X"00000009000000000000000b0000000000000013000000000000000000000000",
            INIT_02 => X"0000001c0000000000000000000000000000002d000000000000000300000000",
            INIT_03 => X"0000000600000000000000000000000000000000000000000000001000000000",
            INIT_04 => X"000000000000000000000000000000000000000100000000000000de00000000",
            INIT_05 => X"0000002300000000000000120000000000000008000000000000000000000000",
            INIT_06 => X"0000000700000000000000000000000000000000000000000000003b00000000",
            INIT_07 => X"0000006700000000000000020000000000000000000000000000000000000000",
            INIT_08 => X"0000001c000000000000000a0000000000000000000000000000001400000000",
            INIT_09 => X"0000003500000000000000290000000000000008000000000000002600000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000001b00000000000000220000000000000001000000000000000000000000",
            INIT_0C => X"000000020000000000000009000000000000003d000000000000001700000000",
            INIT_0D => X"0000000f000000000000002f0000000000000022000000000000001800000000",
            INIT_0E => X"0000000f000000000000000f000000000000000f000000000000000f00000000",
            INIT_0F => X"0000000d000000000000000d000000000000000f000000000000000f00000000",
            INIT_10 => X"0000000f000000000000000f0000000000000014000000000000001000000000",
            INIT_11 => X"0000000f000000000000000e000000000000000f000000000000000f00000000",
            INIT_12 => X"0000000e000000000000000e000000000000000e000000000000000f00000000",
            INIT_13 => X"00000000000000000000000e000000000000000d000000000000000e00000000",
            INIT_14 => X"0000000f000000000000000f000000000000000d000000000000000200000000",
            INIT_15 => X"0000000e000000000000000a0000000000000009000000000000000f00000000",
            INIT_16 => X"0000000f000000000000000e000000000000000e000000000000000e00000000",
            INIT_17 => X"0000001100000000000000200000000000000001000000000000000700000000",
            INIT_18 => X"0000000f000000000000000d000000000000000e000000000000000b00000000",
            INIT_19 => X"0000000c0000000000000011000000000000001c000000000000001e00000000",
            INIT_1A => X"0000002000000000000000070000000000000004000000000000000d00000000",
            INIT_1B => X"00000038000000000000005c0000000000000056000000000000004100000000",
            INIT_1C => X"0000000000000000000000120000000000000015000000000000001600000000",
            INIT_1D => X"0000000b00000000000000050000000000000004000000000000000000000000",
            INIT_1E => X"00000024000000000000001a000000000000001b000000000000001b00000000",
            INIT_1F => X"0000000000000000000000000000000000000009000000000000002400000000",
            INIT_20 => X"0000006800000000000000720000000000000012000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_22 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000004000000000000000620000000000000061000000000000005000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_25 => X"000000470000000000000041000000000000002f000000000000002d00000000",
            INIT_26 => X"00000000000000000000000c0000000000000040000000000000005e00000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000001c000000000000005f000000000000003b00000000",
            INIT_29 => X"0000002000000000000000720000000000000068000000000000002300000000",
            INIT_2A => X"0000004800000000000000320000000000000011000000000000000000000000",
            INIT_2B => X"0000007a0000000000000043000000000000005c000000000000005000000000",
            INIT_2C => X"000000280000000000000046000000000000005d000000000000004b00000000",
            INIT_2D => X"0000004b00000000000000260000000000000007000000000000001000000000",
            INIT_2E => X"00000012000000000000002a000000000000003b000000000000003300000000",
            INIT_2F => X"0000000800000000000000200000000000000012000000000000000400000000",
            INIT_30 => X"0000002b000000000000001e0000000000000014000000000000001000000000",
            INIT_31 => X"00000048000000000000003d0000000000000043000000000000003b00000000",
            INIT_32 => X"0000003f000000000000004e0000000000000042000000000000003c00000000",
            INIT_33 => X"000000100000000000000017000000000000000b000000000000003600000000",
            INIT_34 => X"0000000f00000000000000000000000000000000000000000000000300000000",
            INIT_35 => X"0000003600000000000000280000000000000020000000000000001800000000",
            INIT_36 => X"0000002f000000000000004b0000000000000052000000000000004100000000",
            INIT_37 => X"0000003d000000000000003b0000000000000029000000000000002000000000",
            INIT_38 => X"0000009800000000000000810000000000000030000000000000003000000000",
            INIT_39 => X"00000066000000000000007b0000000000000082000000000000008500000000",
            INIT_3A => X"0000002e00000000000000290000000000000021000000000000002300000000",
            INIT_3B => X"00000021000000000000000d0000000000000000000000000000001200000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_3D => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000002500000000000000270000000000000027000000000000002300000000",
            INIT_3F => X"0000002600000000000000250000000000000023000000000000002100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000001a0000000000000015000000000000001f000000000000002600000000",
            INIT_42 => X"0000002d000000000000002c000000000000001e000000000000001d00000000",
            INIT_43 => X"000000180000000000000032000000000000002e000000000000002e00000000",
            INIT_44 => X"00000008000000000000001d0000000000000026000000000000000000000000",
            INIT_45 => X"0000002300000000000000200000000000000018000000000000000f00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000004900000000000000490000000000000049000000000000000000000000",
            INIT_7F => X"0000004900000000000000490000000000000049000000000000004900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "samplegold_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004900000000000000480000000000000049000000000000004800000000",
            INIT_01 => X"0000004a00000000000000490000000000000049000000000000004a00000000",
            INIT_02 => X"0000004800000000000000490000000000000049000000000000004700000000",
            INIT_03 => X"0000004900000000000000480000000000000048000000000000004800000000",
            INIT_04 => X"00000049000000000000002f000000000000001a000000000000004500000000",
            INIT_05 => X"00000041000000000000004a0000000000000049000000000000004900000000",
            INIT_06 => X"0000004b00000000000000490000000000000048000000000000004400000000",
            INIT_07 => X"00000010000000000000002e0000000000000047000000000000004500000000",
            INIT_08 => X"00000048000000000000003e000000000000002a000000000000001400000000",
            INIT_09 => X"000000510000000000000056000000000000004a000000000000004900000000",
            INIT_0A => X"0000002f00000000000000480000000000000048000000000000004c00000000",
            INIT_0B => X"00000075000000000000006c000000000000003d000000000000004500000000",
            INIT_0C => X"0000004e000000000000004d000000000000007b000000000000008600000000",
            INIT_0D => X"0000003a00000000000000000000000000000000000000000000004d00000000",
            INIT_0E => X"0000006100000000000000460000000000000045000000000000004100000000",
            INIT_0F => X"000000180000000000000045000000000000005e000000000000004f00000000",
            INIT_10 => X"0000004c000000000000001f0000000000000000000000000000000000000000",
            INIT_11 => X"00000015000000000000005500000000000000a1000000000000009400000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_13 => X"0000008d00000000000000750000000000000048000000000000001a00000000",
            INIT_14 => X"0000000000000000000000500000000000000094000000000000008000000000",
            INIT_15 => X"0000004800000000000000530000000000000002000000000000000000000000",
            INIT_16 => X"0000008c000000000000007d0000000000000049000000000000001500000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_18 => X"00000084000000000000002c000000000000000f000000000000000000000000",
            INIT_19 => X"0000009500000000000000400000000000000030000000000000001800000000",
            INIT_1A => X"0000000e0000000000000000000000000000003c00000000000000b700000000",
            INIT_1B => X"0000007d000000000000006a0000000000000055000000000000003000000000",
            INIT_1C => X"00000088000000000000005c00000000000000b3000000000000006e00000000",
            INIT_1D => X"0000001e000000000000002d0000000000000052000000000000007900000000",
            INIT_1E => X"0000002f000000000000002f000000000000004a000000000000002000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_21 => X"0000002100000000000000130000000000000004000000000000000000000000",
            INIT_22 => X"0000000c0000000000000010000000000000001c000000000000002000000000",
            INIT_23 => X"00000000000000000000002e0000000000000028000000000000002700000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002f00000000000000060000000000000000000000000000000000000000",
            INIT_27 => X"0000001200000000000000000000000000000039000000000000003f00000000",
            INIT_28 => X"0000000300000000000000010000000000000010000000000000001900000000",
            INIT_29 => X"0000006900000000000000670000000000000087000000000000008800000000",
            INIT_2A => X"0000001700000000000000280000000000000067000000000000007700000000",
            INIT_2B => X"000000000000000000000000000000000000000a000000000000004f00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000005c00000000000000470000000000000031000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_31 => X"0000004f00000000000000420000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000004f0000000000000042000000000000002f00000000",
            INIT_33 => X"0000001500000000000000140000000000000019000000000000001b00000000",
            INIT_34 => X"0000003d00000000000000000000000000000012000000000000001900000000",
            INIT_35 => X"0000003d00000000000000290000000000000030000000000000005400000000",
            INIT_36 => X"0000004300000000000000440000000000000058000000000000004b00000000",
            INIT_37 => X"0000004300000000000000430000000000000043000000000000004300000000",
            INIT_38 => X"0000004200000000000000440000000000000044000000000000004300000000",
            INIT_39 => X"0000004300000000000000430000000000000043000000000000003e00000000",
            INIT_3A => X"0000004300000000000000430000000000000044000000000000004300000000",
            INIT_3B => X"0000004300000000000000430000000000000043000000000000004300000000",
            INIT_3C => X"0000002400000000000000390000000000000043000000000000004400000000",
            INIT_3D => X"0000004300000000000000430000000000000044000000000000003900000000",
            INIT_3E => X"0000004400000000000000440000000000000042000000000000004100000000",
            INIT_3F => X"0000003f000000000000003f0000000000000043000000000000004400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000026000000000000001b0000000000000015000000000000002700000000",
            INIT_41 => X"0000003600000000000000440000000000000044000000000000004400000000",
            INIT_42 => X"0000004400000000000000450000000000000043000000000000003d00000000",
            INIT_43 => X"00000023000000000000003c0000000000000033000000000000004500000000",
            INIT_44 => X"0000003e00000000000000370000000000000024000000000000002300000000",
            INIT_45 => X"0000000900000000000000080000000000000042000000000000004000000000",
            INIT_46 => X"0000004000000000000000430000000000000043000000000000002000000000",
            INIT_47 => X"00000033000000000000003a000000000000003f000000000000004400000000",
            INIT_48 => X"0000001300000000000000170000000000000018000000000000002400000000",
            INIT_49 => X"000000440000000000000021000000000000001a000000000000003c00000000",
            INIT_4A => X"0000000b0000000000000025000000000000002d000000000000003a00000000",
            INIT_4B => X"00000026000000000000002b0000000000000019000000000000001000000000",
            INIT_4C => X"0000003b00000000000000280000000000000028000000000000002800000000",
            INIT_4D => X"00000014000000000000000a0000000000000000000000000000000000000000",
            INIT_4E => X"0000000b0000000000000000000000000000000c000000000000003100000000",
            INIT_4F => X"0000001d00000000000000290000000000000037000000000000002600000000",
            INIT_50 => X"000000000000000000000012000000000000001b000000000000001000000000",
            INIT_51 => X"00000022000000000000001f000000000000001f000000000000000600000000",
            INIT_52 => X"0000001c000000000000003a000000000000002a000000000000001f00000000",
            INIT_53 => X"00000014000000000000000c0000000000000010000000000000001300000000",
            INIT_54 => X"0000002900000000000000000000000000000021000000000000001600000000",
            INIT_55 => X"0000002f000000000000002c000000000000002f000000000000001e00000000",
            INIT_56 => X"000000030000000000000009000000000000000c000000000000002300000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000040000000000000017000000000000000d00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000003000000000000000320000000000000024000000000000000500000000",
            INIT_66 => X"0000001b00000000000000160000000000000014000000000000002300000000",
            INIT_67 => X"000000000000000000000000000000000000000a000000000000001f00000000",
            INIT_68 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000001600000000000000160000000000000041000000000000004d00000000",
            INIT_6A => X"00000021000000000000001d0000000000000020000000000000002200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_6C => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"00000020000000000000002b0000000000000025000000000000000e00000000",
            INIT_6E => X"0000000000000000000000250000000000000022000000000000001e00000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000003000000000000002c00000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"000000380000000000000017000000000000003a000000000000000b00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000009b00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000030000000000000020000000000000008b00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "samplegold_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007c00000000000000640000000000000030000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000005500000000",
            INIT_02 => X"0000007c00000000000000260000000000000036000000000000000200000000",
            INIT_03 => X"0000000000000000000000470000000000000071000000000000008a00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000005200000000000000ab00000000000000a4000000000000000400000000",
            INIT_06 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000004500000000000000150000000000000000000000000000000000000000",
            INIT_08 => X"0000005b00000000000000670000000000000054000000000000006500000000",
            INIT_09 => X"0000003d00000000000000220000000000000000000000000000002300000000",
            INIT_0A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000010000000000000034000000000000005b00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000031000000000000001b00000000",
            INIT_0F => X"0000004f00000000000000230000000000000004000000000000000e00000000",
            INIT_10 => X"0000007f00000000000000620000000000000048000000000000006e00000000",
            INIT_11 => X"00000053000000000000006e000000000000007e000000000000008600000000",
            INIT_12 => X"00000011000000000000002e0000000000000026000000000000003d00000000",
            INIT_13 => X"00000011000000000000000c0000000000000024000000000000003c00000000",
            INIT_14 => X"00000070000000000000005c0000000000000064000000000000001100000000",
            INIT_15 => X"0000009e00000000000000aa00000000000000a4000000000000008f00000000",
            INIT_16 => X"0000004b00000000000000680000000000000079000000000000009100000000",
            INIT_17 => X"000000000000000000000000000000000000000b000000000000003200000000",
            INIT_18 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_1C => X"000000000000000000000016000000000000003d000000000000001e00000000",
            INIT_1D => X"000000050000000000000022000000000000009b000000000000000000000000",
            INIT_1E => X"0000000000000000000000370000000000000054000000000000001600000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_21 => X"0000000a00000000000000380000000000000029000000000000004000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000f000000000000000f0000000000000025000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000290000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000020000000000000000000000000000001a00000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000001800000000000000260000000000000016000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_3A => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_3C => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_3E => X"0000007f00000000000000230000000000000000000000000000000000000000",
            INIT_3F => X"0000000700000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000e00000000000000000000000000000022000000000000001c00000000",
            INIT_41 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_43 => X"0000000d00000000000000010000000000000008000000000000004200000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000001c0000000000000000000000000000000f000000000000000000000000",
            INIT_47 => X"0000002200000000000000000000000000000011000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000002000000000000000a00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_4A => X"0000000000000000000000030000000000000004000000000000000000000000",
            INIT_4B => X"0000000000000000000000090000000000000002000000000000001e00000000",
            INIT_4C => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000009000000000000001900000000",
            INIT_4E => X"0000000e00000000000000060000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000001600000000000000000000000000000024000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000017000000000000002b00000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_53 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_54 => X"0000001500000000000000000000000000000004000000000000004a00000000",
            INIT_55 => X"0000001600000000000000000000000000000006000000000000000c00000000",
            INIT_56 => X"00000000000000000000002e0000000000000031000000000000001c00000000",
            INIT_57 => X"0000008000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000400000000000000070000000000000001000000000000000600000000",
            INIT_59 => X"0000003600000000000000150000000000000000000000000000000100000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000f00000000000000580000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000003000000000000000400000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000003300000000000000330000000000000033000000000000000000000000",
            INIT_60 => X"0000003300000000000000330000000000000033000000000000003300000000",
            INIT_61 => X"0000003000000000000000310000000000000035000000000000003500000000",
            INIT_62 => X"0000003300000000000000330000000000000033000000000000003300000000",
            INIT_63 => X"0000003300000000000000330000000000000033000000000000003300000000",
            INIT_64 => X"0000003400000000000000320000000000000033000000000000003300000000",
            INIT_65 => X"0000002e000000000000001b0000000000000024000000000000003000000000",
            INIT_66 => X"0000003200000000000000330000000000000033000000000000003300000000",
            INIT_67 => X"0000003400000000000000330000000000000034000000000000003300000000",
            INIT_68 => X"0000000e0000000000000028000000000000002d000000000000003400000000",
            INIT_69 => X"000000320000000000000020000000000000000b000000000000000e00000000",
            INIT_6A => X"0000002900000000000000230000000000000032000000000000003300000000",
            INIT_6B => X"0000003500000000000000360000000000000034000000000000002e00000000",
            INIT_6C => X"000000210000000000000022000000000000002f000000000000002800000000",
            INIT_6D => X"0000002a0000000000000028000000000000001f000000000000002300000000",
            INIT_6E => X"0000001d00000000000000000000000000000000000000000000002e00000000",
            INIT_6F => X"0000002f00000000000000330000000000000033000000000000003200000000",
            INIT_70 => X"0000000e0000000000000025000000000000002d000000000000003000000000",
            INIT_71 => X"0000002800000000000000040000000000000000000000000000000000000000",
            INIT_72 => X"00000021000000000000002e000000000000002f000000000000002700000000",
            INIT_73 => X"0000000200000000000000000000000000000000000000000000002200000000",
            INIT_74 => X"0000002900000000000000210000000000000020000000000000000b00000000",
            INIT_75 => X"0000000000000000000000250000000000000023000000000000003000000000",
            INIT_76 => X"00000022000000000000001e0000000000000008000000000000000000000000",
            INIT_77 => X"0000002300000000000000150000000000000000000000000000000600000000",
            INIT_78 => X"0000000d000000000000000e0000000000000016000000000000002500000000",
            INIT_79 => X"0000002100000000000000000000000000000006000000000000000d00000000",
            INIT_7A => X"000000320000000000000023000000000000001d000000000000001600000000",
            INIT_7B => X"0000000e000000000000000c0000000000000021000000000000003300000000",
            INIT_7C => X"0000001d00000000000000150000000000000013000000000000001000000000",
            INIT_7D => X"0000002a00000000000000280000000000000014000000000000001500000000",
            INIT_7E => X"0000000c00000000000000190000000000000021000000000000002d00000000",
            INIT_7F => X"000000020000000000000000000000000000000f000000000000000a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "samplegold_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000000a000000000000001a000000000000001600000000",
            INIT_09 => X"00000007000000000000000e000000000000001a000000000000001e00000000",
            INIT_0A => X"000000190000000000000013000000000000001f000000000000001a00000000",
            INIT_0B => X"00000029000000000000002b0000000000000031000000000000002700000000",
            INIT_0C => X"0000001500000000000000040000000000000016000000000000002200000000",
            INIT_0D => X"00000020000000000000000c000000000000000c000000000000001500000000",
            INIT_0E => X"0000005400000000000000800000000000000098000000000000008f00000000",
            INIT_0F => X"000000190000000000000020000000000000002f000000000000003b00000000",
            INIT_10 => X"00000010000000000000000e000000000000000d000000000000001700000000",
            INIT_11 => X"000000cf000000000000003a000000000000000d000000000000000d00000000",
            INIT_12 => X"0000002d000000000000003f000000000000005d00000000000000a300000000",
            INIT_13 => X"0000001300000000000000130000000000000016000000000000001f00000000",
            INIT_14 => X"00000011000000000000000c000000000000000e000000000000001400000000",
            INIT_15 => X"00000043000000000000004d0000000000000017000000000000000d00000000",
            INIT_16 => X"000000180000000000000018000000000000002d000000000000003a00000000",
            INIT_17 => X"0000008200000000000000810000000000000015000000000000001700000000",
            INIT_18 => X"0000008200000000000000820000000000000082000000000000008200000000",
            INIT_19 => X"0000008200000000000000820000000000000081000000000000008300000000",
            INIT_1A => X"0000008200000000000000820000000000000082000000000000008400000000",
            INIT_1B => X"0000008300000000000000830000000000000082000000000000008300000000",
            INIT_1C => X"0000008300000000000000820000000000000083000000000000008200000000",
            INIT_1D => X"0000008c0000000000000076000000000000007f000000000000008200000000",
            INIT_1E => X"0000008300000000000000820000000000000082000000000000008600000000",
            INIT_1F => X"0000008300000000000000840000000000000083000000000000008400000000",
            INIT_20 => X"0000007b00000000000000860000000000000081000000000000008300000000",
            INIT_21 => X"000000940000000000000078000000000000006f000000000000007f00000000",
            INIT_22 => X"0000008400000000000000850000000000000084000000000000008300000000",
            INIT_23 => X"0000008300000000000000830000000000000084000000000000008300000000",
            INIT_24 => X"0000007000000000000000760000000000000089000000000000007900000000",
            INIT_25 => X"00000087000000000000007a0000000000000061000000000000006600000000",
            INIT_26 => X"00000087000000000000007b0000000000000086000000000000008600000000",
            INIT_27 => X"0000007c00000000000000840000000000000084000000000000009600000000",
            INIT_28 => X"0000008100000000000000810000000000000080000000000000007b00000000",
            INIT_29 => X"0000009b00000000000000800000000000000087000000000000008500000000",
            INIT_2A => X"00000075000000000000005f0000000000000058000000000000008c00000000",
            INIT_2B => X"00000091000000000000007a0000000000000084000000000000007600000000",
            INIT_2C => X"0000006b0000000000000087000000000000009c000000000000009300000000",
            INIT_2D => X"0000008b000000000000006e000000000000004c000000000000005d00000000",
            INIT_2E => X"00000079000000000000007d0000000000000084000000000000007000000000",
            INIT_2F => X"0000004c0000000000000040000000000000002c000000000000006800000000",
            INIT_30 => X"0000008300000000000000850000000000000081000000000000006600000000",
            INIT_31 => X"0000004800000000000000920000000000000081000000000000008600000000",
            INIT_32 => X"0000007d00000000000000720000000000000048000000000000004200000000",
            INIT_33 => X"000000760000000000000064000000000000005c000000000000005500000000",
            INIT_34 => X"000000490000000000000044000000000000004d000000000000006800000000",
            INIT_35 => X"0000006c0000000000000047000000000000005d000000000000005100000000",
            INIT_36 => X"00000084000000000000007e0000000000000064000000000000005500000000",
            INIT_37 => X"0000006e00000000000000690000000000000075000000000000008a00000000",
            INIT_38 => X"0000007a0000000000000076000000000000006e000000000000007a00000000",
            INIT_39 => X"0000007f000000000000007b000000000000006a000000000000006f00000000",
            INIT_3A => X"0000006d000000000000007a000000000000007f000000000000007f00000000",
            INIT_3B => X"0000005700000000000000510000000000000063000000000000005f00000000",
            INIT_3C => X"0000005300000000000000490000000000000047000000000000004d00000000",
            INIT_3D => X"00000038000000000000002d0000000000000034000000000000001b00000000",
            INIT_3E => X"0000005c000000000000005b0000000000000053000000000000004200000000",
            INIT_3F => X"0000004000000000000000430000000000000049000000000000005600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000480000000000000039000000000000004300000000",
            INIT_41 => X"0000000000000000000000000000000000000006000000000000001100000000",
            INIT_42 => X"000000100000000000000000000000000000002d000000000000000000000000",
            INIT_43 => X"000000380000000000000021000000000000001b000000000000001400000000",
            INIT_44 => X"0000000000000000000000000000000000000046000000000000004000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000001f0000000000000021000000000000002f000000000000003d00000000",
            INIT_47 => X"0000003b00000000000000240000000000000031000000000000002900000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000005600000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000006500000000000000470000000000000034000000000000001a00000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000340000000000000027000000000000000f000000000000000000000000",
            INIT_4F => X"000000000000000000000067000000000000004e000000000000003e00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001500000000000000150000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000009000000000000000e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "samplegold_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000001f00000000000000650000000000000085000000000000003500000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000007c0000000000000066000000000000005c000000000000005d00000000",
            INIT_09 => X"0000008000000000000000830000000000000084000000000000007c00000000",
            INIT_0A => X"00000088000000000000009a0000000000000089000000000000007c00000000",
            INIT_0B => X"0000006600000000000000870000000000000080000000000000008800000000",
            INIT_0C => X"0000007d00000000000000810000000000000073000000000000006400000000",
            INIT_0D => X"0000008200000000000000850000000000000086000000000000008500000000",
            INIT_0E => X"0000009000000000000000860000000000000092000000000000009200000000",
            INIT_0F => X"0000006e000000000000006e000000000000008b000000000000008a00000000",
            INIT_10 => X"0000007d0000000000000077000000000000007c000000000000007400000000",
            INIT_11 => X"0000008d00000000000000960000000000000094000000000000007800000000",
            INIT_12 => X"0000008c000000000000009600000000000000a1000000000000006400000000",
            INIT_13 => X"00000082000000000000006c000000000000007f000000000000008b00000000",
            INIT_14 => X"0000007e0000000000000080000000000000008b000000000000009100000000",
            INIT_15 => X"0000004200000000000000780000000000000089000000000000005b00000000",
            INIT_16 => X"000000a90000000000000092000000000000009e000000000000008800000000",
            INIT_17 => X"00000079000000000000006d000000000000006b000000000000007e00000000",
            INIT_18 => X"00000079000000000000008c0000000000000091000000000000008c00000000",
            INIT_19 => X"00000008000000000000002d000000000000002c000000000000004800000000",
            INIT_1A => X"00000000000000000000005f0000000000000040000000000000002800000000",
            INIT_1B => X"00000000000000000000000e0000000000000015000000000000000900000000",
            INIT_1C => X"00000027000000000000003a0000000000000023000000000000000c00000000",
            INIT_1D => X"0000001300000000000000000000000000000001000000000000001600000000",
            INIT_1E => X"0000002600000000000000140000000000000039000000000000002e00000000",
            INIT_1F => X"0000002c00000000000000350000000000000017000000000000002c00000000",
            INIT_20 => X"000000000000000000000000000000000000000d000000000000001c00000000",
            INIT_21 => X"00000057000000000000005e0000000000000066000000000000001900000000",
            INIT_22 => X"0000000000000000000000000000000000000010000000000000006500000000",
            INIT_23 => X"000000490000000000000040000000000000002d000000000000000500000000",
            INIT_24 => X"0000006200000000000000690000000000000067000000000000005600000000",
            INIT_25 => X"0000000000000000000000290000000000000056000000000000005800000000",
            INIT_26 => X"0000005b00000000000000550000000000000066000000000000004800000000",
            INIT_27 => X"0000004e000000000000006d000000000000007a000000000000006c00000000",
            INIT_28 => X"0000003b00000000000000070000000000000026000000000000003b00000000",
            INIT_29 => X"0000002000000000000000620000000000000048000000000000004f00000000",
            INIT_2A => X"0000004e000000000000005a0000000000000032000000000000000200000000",
            INIT_2B => X"0000007200000000000000620000000000000040000000000000003400000000",
            INIT_2C => X"0000006e000000000000005c000000000000004c000000000000005000000000",
            INIT_2D => X"0000003d000000000000003f0000000000000047000000000000006500000000",
            INIT_2E => X"00000067000000000000006b000000000000005c000000000000004700000000",
            INIT_2F => X"000000570000000000000027000000000000004b000000000000005100000000",
            INIT_30 => X"0000002200000000000000390000000000000061000000000000007300000000",
            INIT_31 => X"00000042000000000000004d000000000000002b000000000000001500000000",
            INIT_32 => X"0000006600000000000000270000000000000011000000000000003000000000",
            INIT_33 => X"0000003200000000000000310000000000000028000000000000003800000000",
            INIT_34 => X"000000000000000000000006000000000000000a000000000000002500000000",
            INIT_35 => X"0000004200000000000000640000000000000061000000000000003600000000",
            INIT_36 => X"0000001600000000000000270000000000000042000000000000004600000000",
            INIT_37 => X"00000007000000000000000d0000000000000027000000000000002a00000000",
            INIT_38 => X"0000002200000000000000000000000000000000000000000000000f00000000",
            INIT_39 => X"0000000d000000000000000a0000000000000012000000000000002400000000",
            INIT_3A => X"00000000000000000000000c0000000000000014000000000000001500000000",
            INIT_3B => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000001100000000000000090000000000000001000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"000000070000000000000007000000000000000a000000000000000000000000",
            INIT_43 => X"0000000d00000000000000050000000000000007000000000000000d00000000",
            INIT_44 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_45 => X"0000000500000000000000080000000000000007000000000000000400000000",
            INIT_46 => X"0000001100000000000000160000000000000000000000000000000c00000000",
            INIT_47 => X"0000000000000000000000130000000000000009000000000000000a00000000",
            INIT_48 => X"00000012000000000000000c0000000000000011000000000000000f00000000",
            INIT_49 => X"00000017000000000000000f0000000000000005000000000000000f00000000",
            INIT_4A => X"0000000900000000000000120000000000000025000000000000000000000000",
            INIT_4B => X"0000001c00000000000000000000000000000019000000000000001100000000",
            INIT_4C => X"0000001d000000000000001a000000000000001c000000000000001900000000",
            INIT_4D => X"000000000000000000000000000000000000000b000000000000001100000000",
            INIT_4E => X"0000001600000000000000190000000000000000000000000000000000000000",
            INIT_4F => X"0000000400000000000000030000000000000000000000000000002700000000",
            INIT_50 => X"000000070000000000000011000000000000000e000000000000001100000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000001d000000000000000a0000000000000024000000000000001400000000",
            INIT_53 => X"000000070000000000000000000000000000000a000000000000000100000000",
            INIT_54 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_55 => X"0000001a00000000000000170000000000000000000000000000000000000000",
            INIT_56 => X"00000000000000000000000a000000000000001b000000000000000800000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000700000000000000170000000000000018000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000002900000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000000000000000000013000000000000001b000000000000000e00000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000001b00000000000000000000000000000002000000000000000000000000",
            INIT_61 => X"00000013000000000000000d0000000000000007000000000000001100000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000002000000000000000100000000",
            INIT_6A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000600000000000000060000000000000000000000000000000900000000",
            INIT_71 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000002000000000000000400000000",
            INIT_73 => X"0000000400000000000000020000000000000000000000000000000e00000000",
            INIT_74 => X"0000000b000000000000000a0000000000000008000000000000000400000000",
            INIT_75 => X"000000090000000000000009000000000000000a000000000000000d00000000",
            INIT_76 => X"0000001700000000000000030000000000000005000000000000000800000000",
            INIT_77 => X"0000000900000000000000060000000000000006000000000000000000000000",
            INIT_78 => X"0000003f00000000000000550000000000000002000000000000000a00000000",
            INIT_79 => X"00000058000000000000005f000000000000005e000000000000005a00000000",
            INIT_7A => X"0000005f0000000000000057000000000000005c000000000000005b00000000",
            INIT_7B => X"0000005d0000000000000059000000000000005a000000000000005600000000",
            INIT_7C => X"0000005100000000000000380000000000000050000000000000005900000000",
            INIT_7D => X"00000055000000000000004d0000000000000055000000000000005200000000",
            INIT_7E => X"0000004300000000000000590000000000000055000000000000005900000000",
            INIT_7F => X"00000052000000000000005d0000000000000057000000000000005900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "samplegold_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000450000000000000043000000000000002d000000000000004900000000",
            INIT_01 => X"00000046000000000000004c0000000000000046000000000000004a00000000",
            INIT_02 => X"0000004c00000000000000320000000000000045000000000000004800000000",
            INIT_03 => X"0000003a000000000000004e000000000000004e000000000000004d00000000",
            INIT_04 => X"0000003c00000000000000350000000000000034000000000000001a00000000",
            INIT_05 => X"0000002c00000000000000320000000000000041000000000000003700000000",
            INIT_06 => X"0000003d00000000000000200000000000000013000000000000003300000000",
            INIT_07 => X"0000000f000000000000001d000000000000002d000000000000003900000000",
            INIT_08 => X"000000260000000000000023000000000000001d000000000000001d00000000",
            INIT_09 => X"00000016000000000000001e0000000000000039000000000000002d00000000",
            INIT_0A => X"0000001600000000000000000000000000000002000000000000000c00000000",
            INIT_0B => X"0000000900000000000000040000000000000001000000000000001100000000",
            INIT_0C => X"00000026000000000000001b0000000000000018000000000000000100000000",
            INIT_0D => X"00000002000000000000000f0000000000000012000000000000002800000000",
            INIT_0E => X"0000000300000000000000230000000000000007000000000000001900000000",
            INIT_0F => X"0000000e000000000000000f0000000000000009000000000000001000000000",
            INIT_10 => X"0000002a00000000000000350000000000000031000000000000002f00000000",
            INIT_11 => X"0000002a000000000000001a0000000000000023000000000000002400000000",
            INIT_12 => X"000000200000000000000000000000000000000d000000000000003100000000",
            INIT_13 => X"0000003f000000000000002d0000000000000026000000000000001c00000000",
            INIT_14 => X"0000003d000000000000003f0000000000000049000000000000004600000000",
            INIT_15 => X"0000002600000000000000240000000000000017000000000000002c00000000",
            INIT_16 => X"0000002a00000000000000330000000000000000000000000000000900000000",
            INIT_17 => X"00000049000000000000004f000000000000004a000000000000003200000000",
            INIT_18 => X"00000025000000000000002d0000000000000036000000000000004000000000",
            INIT_19 => X"0000001d00000000000000280000000000000022000000000000001300000000",
            INIT_1A => X"00000033000000000000002b0000000000000026000000000000001b00000000",
            INIT_1B => X"000000330000000000000038000000000000003a000000000000003a00000000",
            INIT_1C => X"0000002d000000000000002f0000000000000026000000000000003000000000",
            INIT_1D => X"000000000000000000000010000000000000001d000000000000002f00000000",
            INIT_1E => X"0000003100000000000000380000000000000039000000000000002f00000000",
            INIT_1F => X"0000001600000000000000330000000000000032000000000000002c00000000",
            INIT_20 => X"0000001800000000000000210000000000000028000000000000000900000000",
            INIT_21 => X"0000002000000000000000000000000000000000000000000000000300000000",
            INIT_22 => X"000000150000000000000018000000000000002e000000000000003100000000",
            INIT_23 => X"0000000000000000000000050000000000000028000000000000002100000000",
            INIT_24 => X"0000000000000000000000000000000000000004000000000000000d00000000",
            INIT_25 => X"0000001b00000000000000110000000000000000000000000000000000000000",
            INIT_26 => X"0000000600000000000000020000000000000005000000000000001a00000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000010500000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000012d0000000000000123000000000000012100000000000000ef00000000",
            INIT_32 => X"0000012200000000000001270000000000000129000000000000012300000000",
            INIT_33 => X"00000125000000000000012c0000000000000123000000000000012e00000000",
            INIT_34 => X"000000e600000000000001000000000000000126000000000000012c00000000",
            INIT_35 => X"0000011100000000000001210000000000000115000000000000011700000000",
            INIT_36 => X"00000109000000000000011c0000000000000125000000000000011a00000000",
            INIT_37 => X"0000012a0000000000000122000000000000012600000000000000fc00000000",
            INIT_38 => X"0000010500000000000000d500000000000000f9000000000000012500000000",
            INIT_39 => X"000001010000000000000105000000000000010c000000000000010800000000",
            INIT_3A => X"000000cd00000000000000ea000000000000010600000000000000f500000000",
            INIT_3B => X"0000011900000000000001150000000000000117000000000000011600000000",
            INIT_3C => X"000000f800000000000000e500000000000000c300000000000000e400000000",
            INIT_3D => X"000000d500000000000000ef00000000000000f500000000000000f400000000",
            INIT_3E => X"0000007d000000000000007f00000000000000a000000000000000b100000000",
            INIT_3F => X"0000009400000000000000e700000000000000eb00000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a0000000000000008e000000000000008b000000000000008100000000",
            INIT_41 => X"0000009e00000000000000b700000000000000b800000000000000a700000000",
            INIT_42 => X"0000008700000000000000810000000000000083000000000000008a00000000",
            INIT_43 => X"0000006b000000000000006e000000000000007e00000000000000aa00000000",
            INIT_44 => X"00000086000000000000008d0000000000000079000000000000007e00000000",
            INIT_45 => X"0000008a000000000000008b000000000000009f00000000000000a500000000",
            INIT_46 => X"000000a7000000000000009200000000000000be000000000000009300000000",
            INIT_47 => X"0000007900000000000000790000000000000081000000000000006700000000",
            INIT_48 => X"000000be00000000000000c000000000000000b4000000000000008800000000",
            INIT_49 => X"000000b300000000000000a900000000000000a800000000000000b400000000",
            INIT_4A => X"0000006f000000000000007a00000000000000c700000000000000d200000000",
            INIT_4B => X"000000c600000000000000b000000000000000a400000000000000a000000000",
            INIT_4C => X"000000e300000000000000f100000000000000ed00000000000000e100000000",
            INIT_4D => X"000000b600000000000000a900000000000000ba00000000000000e300000000",
            INIT_4E => X"000000ae000000000000006a000000000000008800000000000000bd00000000",
            INIT_4F => X"000000ee00000000000000ee00000000000000c800000000000000b200000000",
            INIT_50 => X"000000be00000000000000d000000000000000e100000000000000eb00000000",
            INIT_51 => X"000000bb00000000000000b500000000000000a100000000000000bb00000000",
            INIT_52 => X"000000a700000000000000a500000000000000a300000000000000a800000000",
            INIT_53 => X"000000cf00000000000000da00000000000000d000000000000000c900000000",
            INIT_54 => X"000000cd00000000000000bf00000000000000c300000000000000cf00000000",
            INIT_55 => X"00000081000000000000009f00000000000000bc00000000000000c600000000",
            INIT_56 => X"000000c700000000000000ca00000000000000cd000000000000006900000000",
            INIT_57 => X"000000ba00000000000000d700000000000000b700000000000000b900000000",
            INIT_58 => X"000000a500000000000000a9000000000000007c000000000000008300000000",
            INIT_59 => X"00000038000000000000004f0000000000000064000000000000008e00000000",
            INIT_5A => X"0000008500000000000000af00000000000000c100000000000000a400000000",
            INIT_5B => X"0000008100000000000000a9000000000000009a000000000000008300000000",
            INIT_5C => X"0000005900000000000000610000000000000077000000000000007500000000",
            INIT_5D => X"00000086000000000000001f0000000000000031000000000000004000000000",
            INIT_5E => X"00000074000000000000007a0000000000000094000000000000009a00000000",
            INIT_5F => X"00000056000000000000005c0000000000000065000000000000006f00000000",
            INIT_60 => X"00000034000000000000003c0000000000000043000000000000005800000000",
            INIT_61 => X"0000003c000000000000003b000000000000001a000000000000002200000000",
            INIT_62 => X"00000040000000000000003f000000000000003b000000000000003a00000000",
            INIT_63 => X"000000390000000000000049000000000000003e000000000000004500000000",
            INIT_64 => X"0000001d00000000000000210000000000000025000000000000003200000000",
            INIT_65 => X"0000001e00000000000000160000000000000017000000000000001d00000000",
            INIT_66 => X"00000031000000000000002e000000000000002a000000000000002300000000",
            INIT_67 => X"0000001e0000000000000039000000000000003e000000000000002900000000",
            INIT_68 => X"00000005000000000000001f000000000000001a000000000000001d00000000",
            INIT_69 => X"000000230000000000000015000000000000000d000000000000001f00000000",
            INIT_6A => X"0000003d0000000000000034000000000000002e000000000000002600000000",
            INIT_6B => X"0000003d00000000000000480000000000000039000000000000003100000000",
            INIT_6C => X"0000003100000000000000330000000000000038000000000000003b00000000",
            INIT_6D => X"0000003a00000000000000370000000000000027000000000000001e00000000",
            INIT_6E => X"0000003800000000000000430000000000000042000000000000003f00000000",
            INIT_6F => X"0000004500000000000000390000000000000048000000000000006500000000",
            INIT_70 => X"0000002a000000000000003d000000000000003b000000000000004400000000",
            INIT_71 => X"0000004600000000000000440000000000000041000000000000003200000000",
            INIT_72 => X"0000007d000000000000004f0000000000000056000000000000004d00000000",
            INIT_73 => X"0000005300000000000000590000000000000051000000000000002600000000",
            INIT_74 => X"00000045000000000000002e0000000000000051000000000000004100000000",
            INIT_75 => X"00000054000000000000004b0000000000000059000000000000005300000000",
            INIT_76 => X"0000003f00000000000000710000000000000074000000000000004500000000",
            INIT_77 => X"0000006600000000000000630000000000000065000000000000007100000000",
            INIT_78 => X"000000630000000000000064000000000000005b000000000000006a00000000",
            INIT_79 => X"0000006300000000000000690000000000000073000000000000007500000000",
            INIT_7A => X"00000000000000000000001d0000000000000020000000000000003400000000",
            INIT_7B => X"0000000100000000000000590000000000000051000000000000001300000000",
            INIT_7C => X"00000000000000000000000f000000000000001c000000000000000100000000",
            INIT_7D => X"0000001d0000000000000020000000000000000a000000000000000300000000",
            INIT_7E => X"0000002700000000000000000000000000000000000000000000001a00000000",
            INIT_7F => X"0000002100000000000000060000000000000036000000000000002f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "samplegold_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000f00000000000000120000000000000006000000000000002800000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000003e000000000000004d000000000000003d000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_04 => X"0000000e00000000000000030000000000000000000000000000000000000000",
            INIT_05 => X"0000004b0000000000000050000000000000002c000000000000001d00000000",
            INIT_06 => X"00000000000000000000003a000000000000003b000000000000003e00000000",
            INIT_07 => X"00000015000000000000001d000000000000003a000000000000001300000000",
            INIT_08 => X"00000033000000000000003f0000000000000039000000000000002100000000",
            INIT_09 => X"000000230000000000000000000000000000001c000000000000001700000000",
            INIT_0A => X"00000008000000000000004e0000000000000031000000000000003300000000",
            INIT_0B => X"0000002200000000000000230000000000000000000000000000000000000000",
            INIT_0C => X"0000004700000000000000390000000000000016000000000000000b00000000",
            INIT_0D => X"00000059000000000000003c0000000000000028000000000000003100000000",
            INIT_0E => X"0000000d0000000000000012000000000000004f000000000000006500000000",
            INIT_0F => X"0000003a0000000000000038000000000000002f000000000000001700000000",
            INIT_10 => X"0000003d00000000000000190000000000000047000000000000004300000000",
            INIT_11 => X"0000003d0000000000000049000000000000005f000000000000005e00000000",
            INIT_12 => X"0000003300000000000000230000000000000009000000000000003400000000",
            INIT_13 => X"000000470000000000000005000000000000000c000000000000002700000000",
            INIT_14 => X"000000410000000000000039000000000000002c000000000000003000000000",
            INIT_15 => X"0000002b000000000000002a0000000000000029000000000000004100000000",
            INIT_16 => X"00000034000000000000004a000000000000003d000000000000001800000000",
            INIT_17 => X"0000002300000000000000300000000000000049000000000000004400000000",
            INIT_18 => X"00000022000000000000002c000000000000003f000000000000003800000000",
            INIT_19 => X"000000380000000000000018000000000000001e000000000000003200000000",
            INIT_1A => X"0000002900000000000000240000000000000031000000000000003a00000000",
            INIT_1B => X"0000000e000000000000002f0000000000000033000000000000003300000000",
            INIT_1C => X"00000020000000000000001f0000000000000027000000000000001c00000000",
            INIT_1D => X"0000001900000000000000200000000000000016000000000000001500000000",
            INIT_1E => X"0000001300000000000000150000000000000018000000000000001a00000000",
            INIT_1F => X"00000037000000000000001d000000000000002b000000000000001e00000000",
            INIT_20 => X"000000140000000000000018000000000000001b000000000000001900000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000120000000000000003000000000000000700000000",
            INIT_2C => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_2D => X"000000000000000000000003000000000000000b000000000000000700000000",
            INIT_2E => X"00000036000000000000001d0000000000000000000000000000000000000000",
            INIT_2F => X"0000002700000000000000600000000000000031000000000000000000000000",
            INIT_30 => X"0000003200000000000000260000000000000046000000000000002000000000",
            INIT_31 => X"0000003400000000000000430000000000000045000000000000003e00000000",
            INIT_32 => X"0000000000000000000000000000000000000007000000000000003400000000",
            INIT_33 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000000000000000000000000000e000000000000000600000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000900000000000000010000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_3F => X"0000000000000000000000210000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000002000000000000000c0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_46 => X"00000000000000000000001c000000000000002a000000000000002000000000",
            INIT_47 => X"00000026000000000000000f0000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000030000000000000000000000000000001600000000",
            INIT_49 => X"000000170000000000000025000000000000002a000000000000001b00000000",
            INIT_4A => X"0000000000000000000000000000000000000015000000000000001200000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000700000000000000000000000000000009000000000000002e00000000",
            INIT_4D => X"0000000600000000000000000000000000000012000000000000001400000000",
            INIT_4E => X"0000003e000000000000002b0000000000000016000000000000000900000000",
            INIT_4F => X"00000007000000000000001b000000000000001c000000000000001f00000000",
            INIT_50 => X"0000000300000000000000160000000000000017000000000000000000000000",
            INIT_51 => X"000000000000000000000002000000000000000f000000000000000300000000",
            INIT_52 => X"00000009000000000000000f000000000000001c000000000000001600000000",
            INIT_53 => X"00000005000000000000000b0000000000000014000000000000000d00000000",
            INIT_54 => X"0000000100000000000000090000000000000000000000000000000000000000",
            INIT_55 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000007000000000000000c0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000002000000000000000300000000",
            INIT_59 => X"000000220000000000000000000000000000000f000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_5B => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_5D => X"0000001f000000000000001f0000000000000000000000000000000300000000",
            INIT_5E => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_5F => X"0000003c00000000000000000000000000000006000000000000000000000000",
            INIT_60 => X"0000000d00000000000000000000000000000000000000000000001600000000",
            INIT_61 => X"0000000000000000000000240000000000000016000000000000000000000000",
            INIT_62 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000002f000000000000007f0000000000000000000000000000001f00000000",
            INIT_64 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000150000000000000012000000000000001c00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_67 => X"0000007000000000000000110000000000000012000000000000000000000000",
            INIT_68 => X"0000000f00000000000000000000000000000021000000000000000800000000",
            INIT_69 => X"0000001500000000000000090000000000000022000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_6B => X"00000000000000000000002b0000000000000010000000000000000500000000",
            INIT_6C => X"0000000000000000000000130000000000000020000000000000000f00000000",
            INIT_6D => X"0000000700000000000000000000000000000003000000000000001a00000000",
            INIT_6E => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000220000000000000000000000000000002200000000",
            INIT_70 => X"0000003d00000000000000000000000000000000000000000000000f00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_72 => X"0000000a000000000000003c0000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"000000080000000000000014000000000000000e000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000001c000000000000002b000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000019000000000000003500000000",
            INIT_79 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_7B => X"0000001000000000000000260000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_7D => X"0000000000000000000000050000000000000011000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000002d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "samplegold_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000002a000000000000000f00000000",
            INIT_01 => X"000000000000000000000000000000000000000d000000000000003d00000000",
            INIT_02 => X"0000004e00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000b00000000000000000000000000000000000000000000003500000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_0A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_0B => X"0000000400000000000000040000000000000004000000000000000d00000000",
            INIT_0C => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_0D => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_0E => X"0000000600000000000000040000000000000008000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000002000000000000000300000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000004a00000000",
            INIT_11 => X"0000005900000000000000000000000000000008000000000000000000000000",
            INIT_12 => X"00000037000000000000003d000000000000004b000000000000004f00000000",
            INIT_13 => X"0000001b000000000000001f000000000000001e000000000000002a00000000",
            INIT_14 => X"0000001800000000000000110000000000000008000000000000001600000000",
            INIT_15 => X"0000003400000000000000410000000000000015000000000000001800000000",
            INIT_16 => X"00000012000000000000001b0000000000000021000000000000002d00000000",
            INIT_17 => X"0000000000000000000000130000000000000010000000000000000c00000000",
            INIT_18 => X"0000000b000000000000000c000000000000000b000000000000000100000000",
            INIT_19 => X"00000014000000000000001f0000000000000029000000000000000c00000000",
            INIT_1A => X"0000000600000000000000080000000000000005000000000000000f00000000",
            INIT_1B => X"0000000700000000000000070000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"000000000000000000000000000000000000000f000000000000000900000000",
            INIT_1E => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000160000000000000011000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000003a000000000000000b0000000000000000000000000000000000000000",
            INIT_23 => X"0000001e0000000000000050000000000000003e000000000000004600000000",
            INIT_24 => X"0000004b00000000000000560000000000000000000000000000000400000000",
            INIT_25 => X"0000005300000000000000540000000000000049000000000000004300000000",
            INIT_26 => X"0000005000000000000000490000000000000050000000000000005300000000",
            INIT_27 => X"000000040000000000000025000000000000004d000000000000005e00000000",
            INIT_28 => X"00000041000000000000003c0000000000000050000000000000001e00000000",
            INIT_29 => X"0000006e000000000000005e000000000000004b000000000000004800000000",
            INIT_2A => X"0000003a0000000000000068000000000000007a000000000000007800000000",
            INIT_2B => X"000000050000000000000000000000000000000e000000000000000100000000",
            INIT_2C => X"0000008100000000000000800000000000000074000000000000007000000000",
            INIT_2D => X"0000004f00000000000000610000000000000065000000000000006e00000000",
            INIT_2E => X"000000000000000000000000000000000000001a000000000000003900000000",
            INIT_2F => X"0000004e000000000000005c0000000000000030000000000000000e00000000",
            INIT_30 => X"0000004c00000000000000510000000000000049000000000000003400000000",
            INIT_31 => X"0000003f00000000000000400000000000000039000000000000003d00000000",
            INIT_32 => X"0000001d00000000000000250000000000000040000000000000004c00000000",
            INIT_33 => X"0000007700000000000000750000000000000000000000000000001900000000",
            INIT_34 => X"0000005b00000000000000560000000000000048000000000000006200000000",
            INIT_35 => X"0000002c00000000000000190000000000000026000000000000004a00000000",
            INIT_36 => X"0000000000000000000000010000000000000019000000000000002900000000",
            INIT_37 => X"0000005500000000000000630000000000000062000000000000000700000000",
            INIT_38 => X"0000003000000000000000340000000000000029000000000000003e00000000",
            INIT_39 => X"0000000800000000000000140000000000000033000000000000002d00000000",
            INIT_3A => X"0000001800000000000000270000000000000019000000000000001300000000",
            INIT_3B => X"0000004a000000000000004a000000000000004d000000000000004d00000000",
            INIT_3C => X"0000003500000000000000270000000000000040000000000000005900000000",
            INIT_3D => X"0000002b0000000000000022000000000000002a000000000000002f00000000",
            INIT_3E => X"0000003c000000000000002d000000000000002b000000000000003100000000",
            INIT_3F => X"000000240000000000000030000000000000002a000000000000002900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002600000000000000380000000000000034000000000000002000000000",
            INIT_41 => X"0000002e00000000000000310000000000000033000000000000002900000000",
            INIT_42 => X"000000240000000000000021000000000000003c000000000000003800000000",
            INIT_43 => X"0000002900000000000000300000000000000035000000000000002f00000000",
            INIT_44 => X"0000003f00000000000000480000000000000031000000000000002f00000000",
            INIT_45 => X"0000003d00000000000000370000000000000031000000000000003200000000",
            INIT_46 => X"0000003a00000000000000360000000000000031000000000000003800000000",
            INIT_47 => X"0000003b00000000000000420000000000000041000000000000003b00000000",
            INIT_48 => X"0000003200000000000000350000000000000028000000000000002b00000000",
            INIT_49 => X"00000020000000000000003b000000000000003a000000000000003600000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "samplegold_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000063000000000000005c000000000000004c000000000000000000000000",
            INIT_03 => X"0000004f000000000000004d0000000000000054000000000000005500000000",
            INIT_04 => X"0000003d000000000000004b0000000000000053000000000000004800000000",
            INIT_05 => X"000000530000000000000050000000000000004e000000000000005000000000",
            INIT_06 => X"0000004600000000000000530000000000000051000000000000004000000000",
            INIT_07 => X"00000040000000000000003a000000000000003f000000000000004800000000",
            INIT_08 => X"0000004e000000000000002c0000000000000019000000000000004c00000000",
            INIT_09 => X"00000035000000000000004b0000000000000042000000000000004300000000",
            INIT_0A => X"0000004000000000000000400000000000000048000000000000004000000000",
            INIT_0B => X"000000290000000000000018000000000000002d000000000000003b00000000",
            INIT_0C => X"0000002b000000000000002b0000000000000039000000000000000000000000",
            INIT_0D => X"0000002900000000000000130000000000000042000000000000003100000000",
            INIT_0E => X"0000002b00000000000000190000000000000015000000000000001600000000",
            INIT_0F => X"000000000000000000000000000000000000002f000000000000002100000000",
            INIT_10 => X"0000000300000000000000000000000000000000000000000000000e00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002900000000000000260000000000000019000000000000000000000000",
            INIT_14 => X"00000000000000000000000a000000000000003d000000000000004500000000",
            INIT_15 => X"0000003e000000000000002c0000000000000047000000000000004300000000",
            INIT_16 => X"000000250000000000000047000000000000004f000000000000006000000000",
            INIT_17 => X"0000008b000000000000006b000000000000003c000000000000002f00000000",
            INIT_18 => X"0000003900000000000000180000000000000034000000000000004000000000",
            INIT_19 => X"0000004000000000000000460000000000000014000000000000002600000000",
            INIT_1A => X"0000007f000000000000006d0000000000000060000000000000005500000000",
            INIT_1B => X"00000019000000000000002b0000000000000069000000000000006f00000000",
            INIT_1C => X"0000006600000000000000590000000000000000000000000000000000000000",
            INIT_1D => X"00000063000000000000006d0000000000000085000000000000008300000000",
            INIT_1E => X"0000000300000000000000300000000000000042000000000000005b00000000",
            INIT_1F => X"0000003000000000000000280000000000000024000000000000000a00000000",
            INIT_20 => X"0000002d000000000000000a0000000000000027000000000000007b00000000",
            INIT_21 => X"0000002700000000000000240000000000000034000000000000004500000000",
            INIT_22 => X"000000680000000000000049000000000000004b000000000000003a00000000",
            INIT_23 => X"000000010000000000000026000000000000002d000000000000003e00000000",
            INIT_24 => X"0000002f00000000000000570000000000000072000000000000004200000000",
            INIT_25 => X"0000001a0000000000000049000000000000005a000000000000003f00000000",
            INIT_26 => X"0000001a00000000000000360000000000000033000000000000001600000000",
            INIT_27 => X"0000004100000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000900000000000000190000000000000038000000000000004800000000",
            INIT_29 => X"000000320000000000000003000000000000001b000000000000002400000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_2B => X"0000003200000000000000400000000000000000000000000000000200000000",
            INIT_2C => X"0000003e00000000000000410000000000000020000000000000002000000000",
            INIT_2D => X"00000010000000000000001f0000000000000015000000000000000000000000",
            INIT_2E => X"00000009000000000000000e0000000000000006000000000000000500000000",
            INIT_2F => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_30 => X"0000001000000000000000000000000000000000000000000000000300000000",
            INIT_31 => X"0000000f00000000000000000000000000000004000000000000001c00000000",
            INIT_32 => X"00000014000000000000000d0000000000000000000000000000001100000000",
            INIT_33 => X"0000000f00000000000000030000000000000000000000000000000000000000",
            INIT_34 => X"0000000b000000000000000a0000000000000007000000000000000c00000000",
            INIT_35 => X"0000000d0000000000000009000000000000001a000000000000003500000000",
            INIT_36 => X"0000000c00000000000000120000000000000017000000000000000d00000000",
            INIT_37 => X"00000024000000000000001f000000000000001b000000000000001700000000",
            INIT_38 => X"0000001e0000000000000002000000000000001a000000000000002600000000",
            INIT_39 => X"00000012000000000000000c000000000000000f000000000000000000000000",
            INIT_3A => X"0000000100000000000000030000000000000000000000000000001700000000",
            INIT_3B => X"0000002c0000000000000021000000000000001b000000000000000d00000000",
            INIT_3C => X"0000003c00000000000000370000000000000039000000000000003500000000",
            INIT_3D => X"0000003f00000000000000410000000000000040000000000000004000000000",
            INIT_3E => X"0000002100000000000000110000000000000015000000000000003f00000000",
            INIT_3F => X"0000003800000000000000380000000000000033000000000000002e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000025000000000000003e000000000000003c000000000000003500000000",
            INIT_41 => X"0000004200000000000000430000000000000047000000000000004100000000",
            INIT_42 => X"0000003d000000000000002e000000000000001d000000000000002200000000",
            INIT_43 => X"00000034000000000000003d000000000000003d000000000000004300000000",
            INIT_44 => X"0000002e000000000000000e000000000000002f000000000000003200000000",
            INIT_45 => X"0000002600000000000000420000000000000044000000000000004300000000",
            INIT_46 => X"0000004b00000000000000390000000000000034000000000000001f00000000",
            INIT_47 => X"0000001a000000000000002f0000000000000042000000000000004000000000",
            INIT_48 => X"0000000600000000000000100000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000041000000000000003700000000",
            INIT_4A => X"0000001a00000000000000190000000000000011000000000000000a00000000",
            INIT_4B => X"000000000000000000000000000000000000000a000000000000001100000000",
            INIT_4C => X"0000002f00000000000000210000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000001f0000000000000021000000000000003d000000000000002100000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000003700000000000000170000000000000003000000000000000000000000",
            INIT_54 => X"000000000000000000000002000000000000003c000000000000003000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000002b00000000000000260000000000000010000000000000001000000000",
            INIT_58 => X"0000000000000000000000000000000000000016000000000000001c00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"00000011000000000000000d0000000000000001000000000000000000000000",
            INIT_5B => X"0000001b000000000000001d0000000000000025000000000000001d00000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_5D => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"00000016000000000000000c0000000000000000000000000000000700000000",
            INIT_5F => X"000000000000000000000007000000000000000f000000000000001700000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000020000000000000002000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_76 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000200000000000000000000000000000000000000000000000600000000",
            INIT_78 => X"0000001f00000000000000000000000000000002000000000000000700000000",
            INIT_79 => X"0000000000000000000000000000000000000001000000000000003000000000",
            INIT_7A => X"0000000c00000000000000100000000000000000000000000000000000000000",
            INIT_7B => X"0000000400000000000000000000000000000001000000000000000000000000",
            INIT_7C => X"0000003700000000000000120000000000000025000000000000003b00000000",
            INIT_7D => X"0000000b0000000000000010000000000000000a000000000000003400000000",
            INIT_7E => X"000000210000000000000027000000000000000e000000000000001300000000",
            INIT_7F => X"000000000000000000000008000000000000000b000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "samplegold_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a30000000000000054000000000000004f000000000000005f00000000",
            INIT_01 => X"00000066000000000000004b000000000000003d000000000000007d00000000",
            INIT_02 => X"0000007000000000000000770000000000000060000000000000005600000000",
            INIT_03 => X"00000003000000000000003f0000000000000055000000000000007000000000",
            INIT_04 => X"0000000a00000000000000000000000000000011000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000000000004a000000000000000900000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_08 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000f00000000000000040000000000000007000000000000000000000000",
            INIT_0A => X"000000000000000000000000000000000000000a000000000000000a00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000900000000000000370000000000000000000000000000001900000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000001600000000000000430000000000000027000000000000001300000000",
            INIT_10 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000001400000000000000090000000000000026000000000000004200000000",
            INIT_12 => X"0000000000000000000000020000000000000028000000000000002c00000000",
            INIT_13 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000032000000000000000000000000",
            INIT_15 => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_16 => X"000000060000000000000032000000000000001f000000000000000000000000",
            INIT_17 => X"00000041000000000000003a000000000000000b000000000000000100000000",
            INIT_18 => X"0000000500000000000000000000000000000005000000000000003900000000",
            INIT_19 => X"00000015000000000000002c0000000000000048000000000000001c00000000",
            INIT_1A => X"0000004700000000000000320000000000000016000000000000002600000000",
            INIT_1B => X"0000001f00000000000000160000000000000020000000000000003a00000000",
            INIT_1C => X"00000012000000000000000e0000000000000011000000000000002400000000",
            INIT_1D => X"0000000700000000000000270000000000000018000000000000000000000000",
            INIT_1E => X"000000220000000000000020000000000000001a000000000000001700000000",
            INIT_1F => X"0000002f00000000000000070000000000000012000000000000000800000000",
            INIT_20 => X"00000040000000000000002b000000000000003e000000000000003f00000000",
            INIT_21 => X"000000280000000000000007000000000000000f000000000000004000000000",
            INIT_22 => X"0000000f00000000000000110000000000000004000000000000002700000000",
            INIT_23 => X"0000003200000000000000390000000000000000000000000000000300000000",
            INIT_24 => X"0000002000000000000000140000000000000011000000000000001c00000000",
            INIT_25 => X"0000000000000000000000000000000000000013000000000000001d00000000",
            INIT_26 => X"0000000000000000000000010000000000000008000000000000000d00000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000080000000000000000000000000000001b000000000000001100000000",
            INIT_2A => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_2C => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_2E => X"0000001600000000000000000000000000000000000000000000000500000000",
            INIT_2F => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_31 => X"0000000e00000000000000000000000000000000000000000000004500000000",
            INIT_32 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_33 => X"0000000100000000000000000000000000000005000000000000000000000000",
            INIT_34 => X"0000007300000000000000000000000000000000000000000000000f00000000",
            INIT_35 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_36 => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_37 => X"0000000200000000000000000000000000000001000000000000000000000000",
            INIT_38 => X"00000000000000000000000b0000000000000042000000000000002a00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_3A => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_3B => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000010000000000000000d00000000",
            INIT_3D => X"00000000000000000000000d0000000000000022000000000000000000000000",
            INIT_3E => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_3F => X"0000000000000000000000110000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007200000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000150000000000000000000000000000004a000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000002600000000000000120000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000006f00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000410000000000000000000000000000001900000000",
            INIT_48 => X"0000000000000000000000530000000000000003000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000001000000000000000e00000000",
            INIT_4A => X"0000000000000000000000000000000000000006000000000000000800000000",
            INIT_4B => X"000000010000000000000000000000000000000e000000000000000000000000",
            INIT_4C => X"000000040000000000000000000000000000001a000000000000000100000000",
            INIT_4D => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_4F => X"00000023000000000000001c0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000006000000000000002900000000",
            INIT_51 => X"0000000000000000000000000000000000000017000000000000000500000000",
            INIT_52 => X"000000000000000000000000000000000000001e000000000000003200000000",
            INIT_53 => X"00000009000000000000001a0000000000000016000000000000001700000000",
            INIT_54 => X"0000002800000000000000000000000000000000000000000000001c00000000",
            INIT_55 => X"0000001e00000000000000000000000000000000000000000000000300000000",
            INIT_56 => X"0000001700000000000000000000000000000000000000000000001700000000",
            INIT_57 => X"00000010000000000000000f0000000000000011000000000000000300000000",
            INIT_58 => X"0000000e000000000000000c000000000000000d000000000000000000000000",
            INIT_59 => X"0000000400000000000000000000000000000000000000000000000700000000",
            INIT_5A => X"00000000000000000000000a0000000000000000000000000000000f00000000",
            INIT_5B => X"0000000900000000000000040000000000000001000000000000001a00000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_5E => X"00000005000000000000000b0000000000000001000000000000002d00000000",
            INIT_5F => X"0000000000000000000000020000000000000007000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000003700000000000000000000000000000012000000000000000200000000",
            INIT_62 => X"0000000000000000000000000000000000000005000000000000000300000000",
            INIT_63 => X"0000000f00000000000000010000000000000009000000000000002d00000000",
            INIT_64 => X"0000002900000000000000240000000000000020000000000000001400000000",
            INIT_65 => X"0000002c000000000000002e0000000000000029000000000000002e00000000",
            INIT_66 => X"000000300000000000000031000000000000002e000000000000002f00000000",
            INIT_67 => X"00000022000000000000001a000000000000000a000000000000001200000000",
            INIT_68 => X"0000002e000000000000002e000000000000002a000000000000002a00000000",
            INIT_69 => X"0000003100000000000000170000000000000025000000000000002b00000000",
            INIT_6A => X"0000001d00000000000000330000000000000035000000000000003200000000",
            INIT_6B => X"0000003200000000000000300000000000000023000000000000001200000000",
            INIT_6C => X"0000002000000000000000220000000000000031000000000000002f00000000",
            INIT_6D => X"00000030000000000000001e0000000000000008000000000000002200000000",
            INIT_6E => X"0000002000000000000000260000000000000033000000000000003500000000",
            INIT_6F => X"000000390000000000000040000000000000003b000000000000003300000000",
            INIT_70 => X"0000000000000000000000020000000000000027000000000000003500000000",
            INIT_71 => X"0000002d00000000000000080000000000000000000000000000000000000000",
            INIT_72 => X"0000000a00000000000000010000000000000004000000000000002f00000000",
            INIT_73 => X"0000000b00000000000000100000000000000015000000000000000a00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_75 => X"000000130000000000000035000000000000001e000000000000001700000000",
            INIT_76 => X"0000000600000000000000090000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000003000000000000000f00000000",
            INIT_78 => X"00000033000000000000000b0000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000160000000000000033000000000000003a00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000700000000000000040000000000000001000000000000000100000000",
            INIT_7C => X"00000039000000000000002d000000000000001b000000000000000b00000000",
            INIT_7D => X"0000000b00000000000000000000000000000011000000000000002600000000",
            INIT_7E => X"000000030000000000000008000000000000000a000000000000000e00000000",
            INIT_7F => X"0000000e00000000000000030000000000000001000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "samplegold_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000029000000000000002a0000000000000027000000000000001200000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000003600000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000230000000000000020000000000000000d000000000000000100000000",
            INIT_04 => X"000000220000000000000021000000000000001e000000000000002300000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000200000000000000060000000000000000000000000000000000000000",
            INIT_07 => X"0000001b00000000000000180000000000000010000000000000000000000000",
            INIT_08 => X"0000000000000000000000060000000000000008000000000000000b00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_0C => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000200000000000000030000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000030000000000000001000000000000000000000000",
            INIT_1B => X"0000007900000000000000790000000000000008000000000000000000000000",
            INIT_1C => X"0000008a0000000000000090000000000000008e000000000000009100000000",
            INIT_1D => X"0000008e000000000000008b0000000000000086000000000000008c00000000",
            INIT_1E => X"0000008a0000000000000085000000000000008d000000000000008a00000000",
            INIT_1F => X"0000008c00000000000000740000000000000076000000000000008900000000",
            INIT_20 => X"00000084000000000000007f000000000000008b000000000000008300000000",
            INIT_21 => X"0000008400000000000000780000000000000087000000000000008b00000000",
            INIT_22 => X"00000089000000000000008a0000000000000083000000000000008d00000000",
            INIT_23 => X"000000780000000000000082000000000000006a000000000000007100000000",
            INIT_24 => X"0000007c00000000000000740000000000000077000000000000007f00000000",
            INIT_25 => X"000000930000000000000078000000000000005d000000000000008600000000",
            INIT_26 => X"0000006800000000000000870000000000000083000000000000008000000000",
            INIT_27 => X"000000700000000000000075000000000000006e000000000000005a00000000",
            INIT_28 => X"00000059000000000000005b000000000000006c000000000000007000000000",
            INIT_29 => X"00000082000000000000004f0000000000000047000000000000004e00000000",
            INIT_2A => X"0000004800000000000000510000000000000078000000000000007500000000",
            INIT_2B => X"0000005d00000000000000570000000000000053000000000000004b00000000",
            INIT_2C => X"0000004100000000000000470000000000000059000000000000006200000000",
            INIT_2D => X"0000004300000000000000410000000000000032000000000000004300000000",
            INIT_2E => X"0000003200000000000000310000000000000032000000000000003e00000000",
            INIT_2F => X"0000004d00000000000000370000000000000039000000000000003800000000",
            INIT_30 => X"0000004500000000000000400000000000000045000000000000004900000000",
            INIT_31 => X"0000001e00000000000000530000000000000025000000000000004f00000000",
            INIT_32 => X"0000004900000000000000360000000000000039000000000000004100000000",
            INIT_33 => X"0000004d00000000000000560000000000000057000000000000005b00000000",
            INIT_34 => X"0000006400000000000000550000000000000046000000000000004400000000",
            INIT_35 => X"0000004700000000000000220000000000000033000000000000004c00000000",
            INIT_36 => X"0000006900000000000000570000000000000048000000000000004300000000",
            INIT_37 => X"00000072000000000000006c0000000000000073000000000000007000000000",
            INIT_38 => X"000000510000000000000058000000000000005d000000000000005600000000",
            INIT_39 => X"0000006300000000000000560000000000000016000000000000002300000000",
            INIT_3A => X"0000007b0000000000000078000000000000007a000000000000006c00000000",
            INIT_3B => X"00000048000000000000005c0000000000000067000000000000007600000000",
            INIT_3C => X"000000450000000000000054000000000000004e000000000000004300000000",
            INIT_3D => X"00000065000000000000004e0000000000000047000000000000005200000000",
            INIT_3E => X"000000630000000000000064000000000000006d000000000000006900000000",
            INIT_3F => X"0000005b00000000000000640000000000000068000000000000005f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000034000000000000003d000000000000004f000000000000005400000000",
            INIT_41 => X"0000005d00000000000000630000000000000065000000000000006e00000000",
            INIT_42 => X"0000003d00000000000000560000000000000077000000000000006700000000",
            INIT_43 => X"000000460000000000000058000000000000005b000000000000004300000000",
            INIT_44 => X"0000006300000000000000190000000000000025000000000000003000000000",
            INIT_45 => X"0000004000000000000000420000000000000053000000000000006400000000",
            INIT_46 => X"0000003d000000000000003e0000000000000051000000000000005400000000",
            INIT_47 => X"0000001900000000000000300000000000000031000000000000003b00000000",
            INIT_48 => X"00000055000000000000004e0000000000000008000000000000001500000000",
            INIT_49 => X"0000004000000000000000440000000000000042000000000000005000000000",
            INIT_4A => X"0000002f000000000000002f000000000000002d000000000000003200000000",
            INIT_4B => X"0000000c0000000000000014000000000000001d000000000000001d00000000",
            INIT_4C => X"0000002000000000000000230000000000000022000000000000000700000000",
            INIT_4D => X"0000002600000000000000240000000000000022000000000000002100000000",
            INIT_4E => X"0000001600000000000000120000000000000023000000000000001e00000000",
            INIT_4F => X"000000070000000000000009000000000000000b000000000000000d00000000",
            INIT_50 => X"0000000e000000000000000c0000000000000008000000000000000600000000",
            INIT_51 => X"0000001000000000000000180000000000000013000000000000001100000000",
            INIT_52 => X"00000008000000000000000b0000000000000010000000000000002900000000",
            INIT_53 => X"000000000000000000000000000000000000000c000000000000000800000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "samplegold_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000510000000000000054000000000000005b000000000000004500000000",
            INIT_0D => X"0000005000000000000000510000000000000053000000000000005700000000",
            INIT_0E => X"0000005400000000000000510000000000000050000000000000004c00000000",
            INIT_0F => X"0000004f000000000000006a0000000000000056000000000000004f00000000",
            INIT_10 => X"0000007e00000000000000740000000000000064000000000000006900000000",
            INIT_11 => X"000000a7000000000000009e00000000000000a700000000000000a600000000",
            INIT_12 => X"00000073000000000000009f00000000000000a500000000000000a400000000",
            INIT_13 => X"0000006600000000000000510000000000000078000000000000007900000000",
            INIT_14 => X"0000003400000000000000480000000000000086000000000000007400000000",
            INIT_15 => X"0000003a000000000000003e0000000000000043000000000000004900000000",
            INIT_16 => X"0000007200000000000000830000000000000052000000000000004300000000",
            INIT_17 => X"000000570000000000000063000000000000004b000000000000007800000000",
            INIT_18 => X"0000003e0000000000000050000000000000004b000000000000004000000000",
            INIT_19 => X"0000005200000000000000590000000000000058000000000000004800000000",
            INIT_1A => X"000000790000000000000075000000000000005d000000000000004800000000",
            INIT_1B => X"0000005d00000000000000600000000000000060000000000000004d00000000",
            INIT_1C => X"0000005a000000000000005d0000000000000061000000000000005c00000000",
            INIT_1D => X"0000005800000000000000590000000000000061000000000000006800000000",
            INIT_1E => X"000000590000000000000077000000000000006d000000000000006600000000",
            INIT_1F => X"000000400000000000000060000000000000008f000000000000006d00000000",
            INIT_20 => X"0000004d000000000000004d0000000000000045000000000000004100000000",
            INIT_21 => X"00000071000000000000005c0000000000000048000000000000004800000000",
            INIT_22 => X"00000051000000000000005c000000000000006f000000000000006e00000000",
            INIT_23 => X"0000008400000000000000b5000000000000008a000000000000002b00000000",
            INIT_24 => X"0000007000000000000000720000000000000073000000000000007100000000",
            INIT_25 => X"0000007900000000000000750000000000000075000000000000007300000000",
            INIT_26 => X"0000004e000000000000006f000000000000005f000000000000007e00000000",
            INIT_27 => X"000000a400000000000000890000000000000025000000000000000000000000",
            INIT_28 => X"0000006e00000000000000770000000000000079000000000000008200000000",
            INIT_29 => X"00000070000000000000006c000000000000006c000000000000007000000000",
            INIT_2A => X"0000006d00000000000000780000000000000077000000000000006200000000",
            INIT_2B => X"000000ac00000000000000510000000000000011000000000000003c00000000",
            INIT_2C => X"0000006f000000000000008100000000000000a100000000000000c300000000",
            INIT_2D => X"0000006100000000000000760000000000000075000000000000007200000000",
            INIT_2E => X"0000007e0000000000000080000000000000007a000000000000007800000000",
            INIT_2F => X"00000020000000000000000d000000000000000f000000000000001600000000",
            INIT_30 => X"000000c000000000000000ce00000000000000a2000000000000005e00000000",
            INIT_31 => X"0000007700000000000000640000000000000079000000000000009500000000",
            INIT_32 => X"0000000000000000000000000000000000000063000000000000007a00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000ca00000000000000c400000000000000a8000000000000006500000000",
            INIT_36 => X"0000008100000000000000ba00000000000000d100000000000000cc00000000",
            INIT_37 => X"00000083000000000000008900000000000000a9000000000000008900000000",
            INIT_38 => X"000000970000000000000094000000000000007d000000000000007a00000000",
            INIT_39 => X"000000270000000000000028000000000000002f000000000000002c00000000",
            INIT_3A => X"0000004200000000000000290000000000000027000000000000002400000000",
            INIT_3B => X"0000007100000000000000690000000000000063000000000000005e00000000",
            INIT_3C => X"0000003b000000000000007f000000000000007f000000000000007c00000000",
            INIT_3D => X"0000001e00000000000000290000000000000038000000000000003c00000000",
            INIT_3E => X"0000000c00000000000000150000000000000016000000000000001900000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000010000000000000002a00000000",
            INIT_45 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_47 => X"0000000400000000000000060000000000000006000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_49 => X"0000001c0000000000000017000000000000001d000000000000002000000000",
            INIT_4A => X"0000001a0000000000000016000000000000001a000000000000001800000000",
            INIT_4B => X"0000000700000000000000000000000000000000000000000000000a00000000",
            INIT_4C => X"0000001d00000000000000080000000000000000000000000000000000000000",
            INIT_4D => X"0000002100000000000000310000000000000023000000000000002e00000000",
            INIT_4E => X"00000013000000000000001f0000000000000023000000000000001f00000000",
            INIT_4F => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_50 => X"00000018000000000000001d0000000000000017000000000000000000000000",
            INIT_51 => X"000000110000000000000018000000000000001c000000000000001900000000",
            INIT_52 => X"0000000000000000000000200000000000000013000000000000002000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"00000006000000000000000e0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_5F => X"00000019000000000000000f0000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000020000000000000011000000000000000000000000",
            INIT_63 => X"0000001d00000000000000190000000000000000000000000000000000000000",
            INIT_64 => X"000000000000000000000000000000000000000c000000000000001700000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000010000000000000004000000000000001500000000",
            INIT_67 => X"0000001d000000000000001f0000000000000018000000000000000000000000",
            INIT_68 => X"0000000c00000000000000100000000000000007000000000000001800000000",
            INIT_69 => X"0000001400000000000000000000000000000001000000000000000c00000000",
            INIT_6A => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000001200000000000000340000000000000010000000000000000000000000",
            INIT_6C => X"0000002c00000000000000110000000000000013000000000000001300000000",
            INIT_6D => X"0000000000000000000000140000000000000003000000000000000f00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000001000000000000000400000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000400000000000000020000000000000016000000000000000000000000",
            INIT_72 => X"0000000b000000000000000c000000000000000c000000000000000700000000",
            INIT_73 => X"0000000000000000000000020000000000000000000000000000000900000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000016000000000000000f000000000000000e000000000000001b00000000",
            INIT_76 => X"0000001b00000000000000180000000000000019000000000000001800000000",
            INIT_77 => X"0000001d0000000000000020000000000000001c000000000000001d00000000",
            INIT_78 => X"000000230000000000000029000000000000001e000000000000001d00000000",
            INIT_79 => X"0000001d000000000000001f000000000000001a000000000000001a00000000",
            INIT_7A => X"0000001f0000000000000023000000000000001d000000000000002000000000",
            INIT_7B => X"0000002400000000000000250000000000000021000000000000002000000000",
            INIT_7C => X"0000005600000000000000390000000000000006000000000000002800000000",
            INIT_7D => X"0000004500000000000000400000000000000035000000000000004500000000",
            INIT_7E => X"00000041000000000000003e0000000000000041000000000000004200000000",
            INIT_7F => X"0000004d00000000000000450000000000000044000000000000004400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "samplegold_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004f0000000000000053000000000000003e000000000000004e00000000",
            INIT_01 => X"00000023000000000000001f000000000000001b000000000000001b00000000",
            INIT_02 => X"0000002b00000000000000260000000000000023000000000000001f00000000",
            INIT_03 => X"000000540000000000000051000000000000004c000000000000002a00000000",
            INIT_04 => X"0000002e0000000000000048000000000000004f000000000000003a00000000",
            INIT_05 => X"000000210000000000000010000000000000001c000000000000002100000000",
            INIT_06 => X"0000002900000000000000250000000000000029000000000000002900000000",
            INIT_07 => X"0000003b00000000000000510000000000000053000000000000003f00000000",
            INIT_08 => X"00000027000000000000001c0000000000000042000000000000004e00000000",
            INIT_09 => X"0000002a000000000000001e0000000000000024000000000000002800000000",
            INIT_0A => X"0000003800000000000000290000000000000026000000000000002900000000",
            INIT_0B => X"0000004c000000000000003f0000000000000056000000000000004f00000000",
            INIT_0C => X"0000003e000000000000003d0000000000000049000000000000005200000000",
            INIT_0D => X"0000004000000000000000440000000000000040000000000000003d00000000",
            INIT_0E => X"00000052000000000000004c0000000000000047000000000000003b00000000",
            INIT_0F => X"00000045000000000000004d0000000000000045000000000000005400000000",
            INIT_10 => X"0000004700000000000000440000000000000048000000000000004a00000000",
            INIT_11 => X"0000004500000000000000460000000000000049000000000000004b00000000",
            INIT_12 => X"0000005200000000000000500000000000000052000000000000004800000000",
            INIT_13 => X"0000002800000000000000270000000000000043000000000000004700000000",
            INIT_14 => X"0000005700000000000000520000000000000047000000000000003b00000000",
            INIT_15 => X"00000051000000000000004f0000000000000050000000000000005400000000",
            INIT_16 => X"0000004a00000000000000550000000000000052000000000000005100000000",
            INIT_17 => X"0000000000000000000000190000000000000050000000000000005400000000",
            INIT_18 => X"00000053000000000000004d000000000000003f000000000000002100000000",
            INIT_19 => X"00000051000000000000004f000000000000004e000000000000005200000000",
            INIT_1A => X"0000005200000000000000480000000000000054000000000000005100000000",
            INIT_1B => X"0000000000000000000000130000000000000051000000000000005300000000",
            INIT_1C => X"0000003c00000000000000350000000000000026000000000000000000000000",
            INIT_1D => X"0000005100000000000000540000000000000054000000000000004900000000",
            INIT_1E => X"00000053000000000000004f0000000000000045000000000000005300000000",
            INIT_1F => X"0000000000000000000000000000000000000016000000000000005000000000",
            INIT_20 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000004e000000000000003d0000000000000030000000000000002d00000000",
            INIT_22 => X"0000004c00000000000000540000000000000054000000000000004500000000",
            INIT_23 => X"0000000400000000000000000000000000000000000000000000002300000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_25 => X"00000033000000000000004a000000000000002b000000000000001300000000",
            INIT_26 => X"00000038000000000000003a000000000000003b000000000000003f00000000",
            INIT_27 => X"000000470000000000000028000000000000001f000000000000003700000000",
            INIT_28 => X"0000003e0000000000000040000000000000003c000000000000004000000000",
            INIT_29 => X"0000000f0000000000000002000000000000004f000000000000004e00000000",
            INIT_2A => X"0000000000000000000000000000000000000005000000000000000c00000000",
            INIT_2B => X"0000000500000000000000090000000000000002000000000000000000000000",
            INIT_2C => X"0000000800000000000000090000000000000007000000000000000400000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000de00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000e000000000000000d300000000000000e8000000000000010000000000",
            INIT_36 => X"000000df00000000000000de00000000000000e100000000000000e700000000",
            INIT_37 => X"000000eb00000000000000e300000000000000e400000000000000e200000000",
            INIT_38 => X"0000010800000000000000e7000000000000010400000000000000fa00000000",
            INIT_39 => X"000000db00000000000000be00000000000000b7000000000000010100000000",
            INIT_3A => X"000000e000000000000000dd00000000000000db00000000000000d600000000",
            INIT_3B => X"00000108000000000000010a00000000000000e300000000000000e400000000",
            INIT_3C => X"00000100000000000000010400000000000000e3000000000000010d00000000",
            INIT_3D => X"0000009c00000000000000a100000000000000b100000000000000c300000000",
            INIT_3E => X"000000b900000000000000b300000000000000b200000000000000ab00000000",
            INIT_3F => X"00000111000000000000010a00000000000000fd00000000000000c400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009c00000000000000dd000000000000010200000000000000e200000000",
            INIT_41 => X"000000a900000000000000a600000000000000b900000000000000b000000000",
            INIT_42 => X"000000bb00000000000000b200000000000000b400000000000000ba00000000",
            INIT_43 => X"000000ef000000000000010e000000000000010900000000000000d100000000",
            INIT_44 => X"000000d400000000000000e400000000000000fe00000000000000fe00000000",
            INIT_45 => X"000000df00000000000000db00000000000000d900000000000000d200000000",
            INIT_46 => X"000000fd00000000000000eb00000000000000d300000000000000d900000000",
            INIT_47 => X"000000f700000000000000fc000000000000010e000000000000010800000000",
            INIT_48 => X"000000f100000000000000f2000000000000010b00000000000000f000000000",
            INIT_49 => X"000000f500000000000000f800000000000000fc00000000000000f700000000",
            INIT_4A => X"00000107000000000000010800000000000000fd00000000000000f300000000",
            INIT_4B => X"000000a700000000000000f60000000000000100000000000000010c00000000",
            INIT_4C => X"0000010e000000000000011200000000000000e7000000000000009000000000",
            INIT_4D => X"0000010900000000000001090000000000000110000000000000011100000000",
            INIT_4E => X"0000010e000000000000010a0000000000000109000000000000010900000000",
            INIT_4F => X"000000b400000000000001010000000000000116000000000000010600000000",
            INIT_50 => X"0000011700000000000000ff00000000000000a9000000000000005400000000",
            INIT_51 => X"0000010600000000000001030000000000000106000000000000010c00000000",
            INIT_52 => X"0000010800000000000001090000000000000106000000000000010700000000",
            INIT_53 => X"0000008100000000000001080000000000000113000000000000011600000000",
            INIT_54 => X"000000e100000000000000a30000000000000064000000000000004700000000",
            INIT_55 => X"00000109000000000000010c000000000000010d00000000000000ff00000000",
            INIT_56 => X"0000010c0000000000000104000000000000010d000000000000010700000000",
            INIT_57 => X"00000023000000000000008b0000000000000100000000000000011200000000",
            INIT_58 => X"00000058000000000000004b0000000000000048000000000000003b00000000",
            INIT_59 => X"0000010500000000000000e900000000000000b8000000000000007c00000000",
            INIT_5A => X"00000110000000000000010e0000000000000102000000000000010f00000000",
            INIT_5B => X"00000043000000000000006200000000000000b000000000000000fc00000000",
            INIT_5C => X"00000069000000000000006a0000000000000097000000000000007000000000",
            INIT_5D => X"000000f000000000000000ce000000000000008b000000000000005600000000",
            INIT_5E => X"000000d900000000000000dd00000000000000e300000000000000d400000000",
            INIT_5F => X"000000cd00000000000000b600000000000000cd00000000000000d700000000",
            INIT_60 => X"000000d800000000000000d500000000000000d300000000000000df00000000",
            INIT_61 => X"0000007d00000000000000e600000000000000e300000000000000da00000000",
            INIT_62 => X"0000007300000000000000790000000000000082000000000000008a00000000",
            INIT_63 => X"00000087000000000000007e0000000000000071000000000000007200000000",
            INIT_64 => X"0000008c00000000000000850000000000000083000000000000008200000000",
            INIT_65 => X"0000004800000000000000430000000000000082000000000000008a00000000",
            INIT_66 => X"000000310000000000000033000000000000003e000000000000004700000000",
            INIT_67 => X"00000024000000000000002e0000000000000030000000000000002f00000000",
            INIT_68 => X"0000002500000000000000240000000000000023000000000000002200000000",
            INIT_69 => X"000000270000000000000027000000000000002a000000000000004500000000",
            INIT_6A => X"00000029000000000000002d0000000000000023000000000000002300000000",
            INIT_6B => X"000000200000000000000027000000000000002c000000000000002900000000",
            INIT_6C => X"00000050000000000000004b0000000000000030000000000000001d00000000",
            INIT_6D => X"0000001a000000000000001f0000000000000011000000000000001300000000",
            INIT_6E => X"0000001d0000000000000022000000000000001e000000000000001b00000000",
            INIT_6F => X"00000020000000000000001e000000000000001e000000000000001c00000000",
            INIT_70 => X"0000001300000000000000230000000000000013000000000000001300000000",
            INIT_71 => X"0000002a0000000000000034000000000000001d000000000000001c00000000",
            INIT_72 => X"0000003e0000000000000039000000000000004c000000000000003f00000000",
            INIT_73 => X"0000002100000000000000370000000000000040000000000000004000000000",
            INIT_74 => X"0000001f00000000000000170000000000000028000000000000002a00000000",
            INIT_75 => X"00000000000000000000000c0000000000000021000000000000002300000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_77 => X"0000002900000000000000210000000000000000000000000000000000000000",
            INIT_78 => X"0000002800000000000000190000000000000010000000000000002800000000",
            INIT_79 => X"0000001a00000000000000160000000000000019000000000000001200000000",
            INIT_7A => X"00000025000000000000002c0000000000000020000000000000001100000000",
            INIT_7B => X"0000002a000000000000002d0000000000000011000000000000001d00000000",
            INIT_7C => X"00000022000000000000001a0000000000000019000000000000001500000000",
            INIT_7D => X"0000001b00000000000000240000000000000027000000000000002300000000",
            INIT_7E => X"000000120000000000000025000000000000002c000000000000002400000000",
            INIT_7F => X"0000002000000000000000240000000000000020000000000000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "samplegold_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000001a0000000000000040000000000000002400000000",
            INIT_01 => X"0000000400000000000000030000000000000000000000000000000000000000",
            INIT_02 => X"0000002500000000000000100000000000000008000000000000000700000000",
            INIT_03 => X"000000250000000000000024000000000000001f000000000000002400000000",
            INIT_04 => X"00000031000000000000005a0000000000000056000000000000002c00000000",
            INIT_05 => X"00000021000000000000001f000000000000001d000000000000001d00000000",
            INIT_06 => X"0000002a00000000000000270000000000000026000000000000002200000000",
            INIT_07 => X"0000001800000000000000220000000000000022000000000000002b00000000",
            INIT_08 => X"0000004a0000000000000047000000000000001c000000000000000100000000",
            INIT_09 => X"00000025000000000000002b0000000000000029000000000000003100000000",
            INIT_0A => X"0000002000000000000000220000000000000021000000000000002500000000",
            INIT_0B => X"0000002d000000000000002e000000000000002c000000000000002300000000",
            INIT_0C => X"00000073000000000000004c0000000000000027000000000000004900000000",
            INIT_0D => X"0000001d000000000000002a000000000000004f000000000000007000000000",
            INIT_0E => X"0000002700000000000000250000000000000028000000000000002300000000",
            INIT_0F => X"0000008700000000000000400000000000000030000000000000002f00000000",
            INIT_10 => X"0000003900000000000000240000000000000028000000000000003000000000",
            INIT_11 => X"00000071000000000000008a0000000000000075000000000000006700000000",
            INIT_12 => X"0000002900000000000000280000000000000025000000000000004400000000",
            INIT_13 => X"0000000000000000000000000000000000000039000000000000002d00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000007e00000000000000700000000000000062000000000000001d00000000",
            INIT_17 => X"00000047000000000000007a0000000000000085000000000000008200000000",
            INIT_18 => X"00000037000000000000003d0000000000000057000000000000004100000000",
            INIT_19 => X"0000003c000000000000003a000000000000002d000000000000002d00000000",
            INIT_1A => X"0000001800000000000000120000000000000015000000000000002200000000",
            INIT_1B => X"000000230000000000000019000000000000001f000000000000001d00000000",
            INIT_1C => X"0000004c00000000000000490000000000000042000000000000003f00000000",
            INIT_1D => X"00000053000000000000005c0000000000000058000000000000005300000000",
            INIT_1E => X"000000490000000000000047000000000000004d000000000000004e00000000",
            INIT_1F => X"0000003d000000000000003d000000000000003b000000000000004100000000",
            INIT_20 => X"0000002e00000000000000300000000000000034000000000000003b00000000",
            INIT_21 => X"0000002a0000000000000037000000000000000d000000000000002d00000000",
            INIT_22 => X"0000001a000000000000002d0000000000000027000000000000002600000000",
            INIT_23 => X"0000001a000000000000001f000000000000001b000000000000001900000000",
            INIT_24 => X"000000060000000000000025000000000000002e000000000000002100000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000005900000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000001d000000000000001c0000000000000023000000000000000000000000",
            INIT_2B => X"000000180000000000000023000000000000001c000000000000002000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000005d000000000000002d0000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000000000000000000002b0000000000000069000000000000006600000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000000c0000000000000015000000000000001600000000",
            INIT_49 => X"0000008600000000000000650000000000000028000000000000000000000000",
            INIT_4A => X"000000000000000000000000000000000000001f000000000000006700000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000005f000000000000005a0000000000000000000000000000000000000000",
            INIT_4F => X"0000007100000000000000740000000000000070000000000000006900000000",
            INIT_50 => X"000000300000000000000048000000000000003a000000000000004a00000000",
            INIT_51 => X"0000002d000000000000001e0000000000000027000000000000003000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_53 => X"0000000400000000000000020000000000000000000000000000000000000000",
            INIT_54 => X"00000032000000000000002d0000000000000023000000000000001200000000",
            INIT_55 => X"0000003c000000000000003e000000000000003d000000000000003700000000",
            INIT_56 => X"0000000e00000000000000180000000000000019000000000000000d00000000",
            INIT_57 => X"000000050000000000000007000000000000000c000000000000000d00000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000600000000000000350000000000000017000000000000000000000000",
            INIT_5E => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_61 => X"000000000000000000000011000000000000002f000000000000000000000000",
            INIT_62 => X"0000000000000000000000090000000000000010000000000000000000000000",
            INIT_63 => X"0000000100000000000000040000000000000000000000000000001200000000",
            INIT_64 => X"0000000000000000000000000000000000000015000000000000001d00000000",
            INIT_65 => X"000000000000000000000000000000000000000d000000000000002b00000000",
            INIT_66 => X"0000001600000000000000000000000000000001000000000000000000000000",
            INIT_67 => X"0000001900000000000000040000000000000000000000000000000000000000",
            INIT_68 => X"0000001b00000000000000000000000000000000000000000000002200000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000c00000000000000010000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"000000000000000000000000000000000000001f000000000000000100000000",
            INIT_70 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_74 => X"0000000700000000000000000000000000000000000000000000001300000000",
            INIT_75 => X"0000000000000000000000000000000000000023000000000000005500000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000090000000000000058000000000000006400000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_7C => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000001d000000000000003e0000000000000041000000000000003a00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_7F => X"0000000000000000000000000000000000000021000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "samplegold_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000490000000000000000000000000000000b000000000000000e00000000",
            INIT_02 => X"0000000900000000000000270000000000000044000000000000003a00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_04 => X"0000005000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000002e00000000000000080000000000000012000000000000005f00000000",
            INIT_07 => X"0000001000000000000000070000000000000002000000000000000400000000",
            INIT_08 => X"00000000000000000000003c0000000000000010000000000000000000000000",
            INIT_09 => X"0000000a0000000000000001000000000000000a000000000000000000000000",
            INIT_0A => X"0000000000000000000000020000000000000007000000000000000100000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000500000000000000000000000000000015000000000000000400000000",
            INIT_0D => X"00000000000000000000000c000000000000000d000000000000000200000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_11 => X"0000003500000000000000040000000000000000000000000000000000000000",
            INIT_12 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000050000000000000000000000000000000a000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"000000340000000000000000000000000000001e000000000000002000000000",
            INIT_16 => X"0000002a00000000000000260000000000000044000000000000004600000000",
            INIT_17 => X"00000030000000000000002d000000000000002b000000000000003000000000",
            INIT_18 => X"00000032000000000000002b000000000000002b000000000000002d00000000",
            INIT_19 => X"00000042000000000000003b000000000000002b000000000000002c00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000002500000000000000200000000000000000000000000000000000000000",
            INIT_1D => X"0000002f00000000000000430000000000000039000000000000002600000000",
            INIT_1E => X"000000030000000000000013000000000000000f000000000000000000000000",
            INIT_1F => X"0000001e000000000000001a000000000000001c000000000000000c00000000",
            INIT_20 => X"00000029000000000000002a0000000000000015000000000000001300000000",
            INIT_21 => X"0000000a00000000000000250000000000000046000000000000003f00000000",
            INIT_22 => X"0000000d0000000000000014000000000000001a000000000000000c00000000",
            INIT_23 => X"0000000800000000000000000000000000000000000000000000000a00000000",
            INIT_24 => X"00000043000000000000002b0000000000000028000000000000001700000000",
            INIT_25 => X"0000002d00000000000000370000000000000046000000000000004400000000",
            INIT_26 => X"00000028000000000000002e000000000000002e000000000000002600000000",
            INIT_27 => X"0000003800000000000000310000000000000028000000000000002c00000000",
            INIT_28 => X"0000003300000000000000370000000000000034000000000000003200000000",
            INIT_29 => X"0000005200000000000000550000000000000046000000000000001e00000000",
            INIT_2A => X"0000004c000000000000004e000000000000004d000000000000004f00000000",
            INIT_2B => X"000000330000000000000033000000000000003c000000000000004800000000",
            INIT_2C => X"00000033000000000000004b000000000000002e000000000000003500000000",
            INIT_2D => X"0000003600000000000000280000000000000000000000000000000000000000",
            INIT_2E => X"0000003000000000000000330000000000000036000000000000003600000000",
            INIT_2F => X"0000002b000000000000002a000000000000002f000000000000003100000000",
            INIT_30 => X"0000005f00000000000000480000000000000038000000000000002a00000000",
            INIT_31 => X"0000002500000000000000000000000000000000000000000000001a00000000",
            INIT_32 => X"00000031000000000000002e000000000000002a000000000000002a00000000",
            INIT_33 => X"0000002500000000000000380000000000000036000000000000003500000000",
            INIT_34 => X"0000002d000000000000002e0000000000000026000000000000002600000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_36 => X"0000003100000000000000340000000000000026000000000000000400000000",
            INIT_37 => X"0000001d000000000000001d0000000000000034000000000000002f00000000",
            INIT_38 => X"0000000700000000000000080000000000000012000000000000002200000000",
            INIT_39 => X"0000000000000000000000020000000000000012000000000000000e00000000",
            INIT_3A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000230000000000000025000000000000001e000000000000002e00000000",
            INIT_3C => X"00000062000000000000007e0000000000000073000000000000003000000000",
            INIT_3D => X"000000740000000000000075000000000000006e000000000000006800000000",
            INIT_3E => X"00000029000000000000003f0000000000000053000000000000006700000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000300000000000000080000000000000000000000000000000000000000",
            INIT_41 => X"00000025000000000000001c0000000000000016000000000000000300000000",
            INIT_42 => X"0000002000000000000000170000000000000019000000000000002300000000",
            INIT_43 => X"00000029000000000000002f0000000000000036000000000000003200000000",
            INIT_44 => X"000000140000000000000021000000000000002c000000000000002b00000000",
            INIT_45 => X"0000000200000000000000050000000000000009000000000000000d00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000600000000000000000000000000000001000000000000000000000000",
            INIT_48 => X"00000010000000000000000c0000000000000008000000000000000900000000",
            INIT_49 => X"0000001d00000000000000150000000000000013000000000000001200000000",
            INIT_4A => X"0000001b000000000000001a0000000000000010000000000000004f00000000",
            INIT_4B => X"0000002400000000000000270000000000000016000000000000001700000000",
            INIT_4C => X"0000001b00000000000000240000000000000022000000000000002000000000",
            INIT_4D => X"00000004000000000000004a0000000000000030000000000000001700000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "samplegold_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000004500000000000000540000000000000051000000000000000000000000",
            INIT_07 => X"0000004700000000000000490000000000000040000000000000003b00000000",
            INIT_08 => X"0000004a000000000000004a000000000000004c000000000000004900000000",
            INIT_09 => X"0000005000000000000000560000000000000053000000000000004600000000",
            INIT_0A => X"000000000000000000000044000000000000004d000000000000005000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000004b0000000000000048000000000000003f000000000000003e00000000",
            INIT_0E => X"0000001b0000000000000005000000000000002e000000000000004d00000000",
            INIT_0F => X"0000003d000000000000002e000000000000001b000000000000003400000000",
            INIT_10 => X"00000034000000000000003b000000000000003a000000000000003b00000000",
            INIT_11 => X"0000004e000000000000004f0000000000000049000000000000004600000000",
            INIT_12 => X"0000002a0000000000000025000000000000002a000000000000002200000000",
            INIT_13 => X"000000100000000000000024000000000000002a000000000000002d00000000",
            INIT_14 => X"000000410000000000000041000000000000002d000000000000001a00000000",
            INIT_15 => X"0000004a000000000000004f0000000000000050000000000000004400000000",
            INIT_16 => X"0000003500000000000000310000000000000034000000000000003400000000",
            INIT_17 => X"00000036000000000000002a000000000000002f000000000000003600000000",
            INIT_18 => X"0000004a00000000000000480000000000000051000000000000004600000000",
            INIT_19 => X"0000004b0000000000000019000000000000003b000000000000005000000000",
            INIT_1A => X"0000005f00000000000000650000000000000067000000000000006600000000",
            INIT_1B => X"00000059000000000000005e000000000000005f000000000000005f00000000",
            INIT_1C => X"000000510000000000000051000000000000004a000000000000004600000000",
            INIT_1D => X"000000000000000000000000000000000000003e000000000000005000000000",
            INIT_1E => X"0000004b000000000000004b000000000000004a000000000000003100000000",
            INIT_1F => X"0000004100000000000000420000000000000044000000000000004600000000",
            INIT_20 => X"0000005000000000000000530000000000000040000000000000003d00000000",
            INIT_21 => X"00000000000000000000001e000000000000007a000000000000005900000000",
            INIT_22 => X"0000003d000000000000003f000000000000003a000000000000000e00000000",
            INIT_23 => X"0000004800000000000000490000000000000046000000000000004500000000",
            INIT_24 => X"00000048000000000000004a0000000000000050000000000000004c00000000",
            INIT_25 => X"0000000000000000000000120000000000000009000000000000004200000000",
            INIT_26 => X"0000003600000000000000070000000000000000000000000000000000000000",
            INIT_27 => X"0000004700000000000000430000000000000045000000000000004900000000",
            INIT_28 => X"0000002000000000000000440000000000000044000000000000004d00000000",
            INIT_29 => X"0000001400000000000000060000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_2B => X"000000490000000000000041000000000000001c000000000000000000000000",
            INIT_2C => X"0000008d000000000000003d0000000000000044000000000000004400000000",
            INIT_2D => X"000000a400000000000000a0000000000000007c000000000000009600000000",
            INIT_2E => X"00000099000000000000008300000000000000a8000000000000007c00000000",
            INIT_2F => X"0000000000000000000000000000000000000047000000000000006800000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000000e000000000000000f000000000000000100000000",
            INIT_33 => X"0000002200000000000000220000000000000025000000000000000000000000",
            INIT_34 => X"000000180000000000000018000000000000001e000000000000001e00000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000c00000000000000090000000000000005000000000000000200000000",
            INIT_3A => X"00000009000000000000005f000000000000001c000000000000000c00000000",
            INIT_3B => X"0000001100000000000000130000000000000011000000000000000f00000000",
            INIT_3C => X"0000002700000000000000280000000000000025000000000000002400000000",
            INIT_3D => X"0000003c0000000000000012000000000000001d000000000000002800000000",
            INIT_3E => X"0000000c00000000000000090000000000000005000000000000005f00000000",
            INIT_3F => X"0000001e0000000000000017000000000000001c000000000000001b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002500000000000000240000000000000021000000000000002300000000",
            INIT_41 => X"0000002800000000000000220000000000000024000000000000002400000000",
            INIT_42 => X"0000001400000000000000080000000000000004000000000000002700000000",
            INIT_43 => X"000000390000000000000033000000000000003b000000000000004500000000",
            INIT_44 => X"0000002f00000000000000330000000000000036000000000000003000000000",
            INIT_45 => X"0000002700000000000000260000000000000020000000000000002900000000",
            INIT_46 => X"00000029000000000000001a0000000000000006000000000000000500000000",
            INIT_47 => X"0000002e0000000000000032000000000000002a000000000000002d00000000",
            INIT_48 => X"0000002e000000000000002c000000000000002a000000000000002800000000",
            INIT_49 => X"0000000800000000000000240000000000000025000000000000001700000000",
            INIT_4A => X"00000037000000000000004a0000000000000021000000000000000600000000",
            INIT_4B => X"0000003e000000000000003a000000000000003c000000000000003600000000",
            INIT_4C => X"000000340000000000000037000000000000003c000000000000004300000000",
            INIT_4D => X"00000008000000000000000e000000000000001f000000000000002100000000",
            INIT_4E => X"0000000e000000000000000c0000000000000017000000000000000c00000000",
            INIT_4F => X"00000014000000000000000f0000000000000013000000000000000c00000000",
            INIT_50 => X"0000001b000000000000001d0000000000000011000000000000001700000000",
            INIT_51 => X"0000000a00000000000000140000000000000016000000000000001a00000000",
            INIT_52 => X"0000001600000000000000130000000000000016000000000000000100000000",
            INIT_53 => X"0000001a00000000000000170000000000000017000000000000001800000000",
            INIT_54 => X"0000001d000000000000001f0000000000000019000000000000001b00000000",
            INIT_55 => X"0000001d0000000000000029000000000000001b000000000000001d00000000",
            INIT_56 => X"0000001d000000000000001b0000000000000008000000000000000000000000",
            INIT_57 => X"0000001b000000000000001c000000000000001f000000000000001f00000000",
            INIT_58 => X"0000001f000000000000001b000000000000001d000000000000001b00000000",
            INIT_59 => X"00000029000000000000002b0000000000000022000000000000001e00000000",
            INIT_5A => X"00000024000000000000001c0000000000000000000000000000000000000000",
            INIT_5B => X"0000001c000000000000001d0000000000000020000000000000002100000000",
            INIT_5C => X"0000002800000000000000240000000000000017000000000000001c00000000",
            INIT_5D => X"00000008000000000000002b000000000000002e000000000000002c00000000",
            INIT_5E => X"0000000a00000000000000000000000000000008000000000000001200000000",
            INIT_5F => X"0000001c000000000000001e000000000000001f000000000000001100000000",
            INIT_60 => X"0000002c000000000000002f0000000000000027000000000000001800000000",
            INIT_61 => X"000000000000000000000000000000000000001b000000000000003000000000",
            INIT_62 => X"00000000000000000000000e0000000000000013000000000000000800000000",
            INIT_63 => X"00000017000000000000000a0000000000000000000000000000000000000000",
            INIT_64 => X"0000002c000000000000002a0000000000000028000000000000002100000000",
            INIT_65 => X"000000160000000000000017000000000000002d000000000000002400000000",
            INIT_66 => X"00000029000000000000001a000000000000002c000000000000002b00000000",
            INIT_67 => X"000000090000000000000023000000000000002b000000000000001800000000",
            INIT_68 => X"0000000200000000000000040000000000000008000000000000000800000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"000000020000000000000005000000000000000d000000000000000000000000",
            INIT_70 => X"000000030000000000000005000000000000000b000000000000000400000000",
            INIT_71 => X"0000000400000000000000070000000000000007000000000000000500000000",
            INIT_72 => X"0000000100000000000000010000000000000002000000000000000300000000",
            INIT_73 => X"0000000400000000000000010000000000000003000000000000000c00000000",
            INIT_74 => X"0000000c000000000000000a0000000000000003000000000000000600000000",
            INIT_75 => X"00000009000000000000000b000000000000000d000000000000000f00000000",
            INIT_76 => X"0000000000000000000000110000000000000004000000000000000200000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000600000000000000040000000000000000000000000000000000000000",
            INIT_7B => X"0000004b000000000000002c0000000000000012000000000000000000000000",
            INIT_7C => X"0000003f0000000000000041000000000000003a000000000000004100000000",
            INIT_7D => X"000000010000000000000000000000000000002c000000000000003a00000000",
            INIT_7E => X"0000001a00000000000000010000000000000007000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "samplegold_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_02 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000040000000000000004000000000000000000000000",
            INIT_06 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000b00000000000000050000000000000006000000000000000f00000000",
            INIT_08 => X"0000000000000000000000040000000000000006000000000000000700000000",
            INIT_09 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000150000000000000071000000000000008700000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000700000000000000080000000000000001000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000005000000000000004e0000000000000083000000000000001100000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000007a00000000000000a50000000000000069000000000000001200000000",
            INIT_17 => X"0000000000000000000000000000000000000010000000000000003700000000",
            INIT_18 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_19 => X"0000002c0000000000000006000000000000000a000000000000000000000000",
            INIT_1A => X"0000007900000000000000250000000000000000000000000000001300000000",
            INIT_1B => X"0000002b000000000000007200000000000000b000000000000000bf00000000",
            INIT_1C => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000008d0000000000000086000000000000007b000000000000007500000000",
            INIT_21 => X"0000005900000000000000410000000000000061000000000000009600000000",
            INIT_22 => X"0000002400000000000000450000000000000031000000000000006800000000",
            INIT_23 => X"00000000000000000000004d0000000000000057000000000000004300000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000003000000000000000230000000000000000000000000000000000000000",
            INIT_26 => X"0000005600000000000000500000000000000046000000000000003d00000000",
            INIT_27 => X"000000410000000000000035000000000000005c000000000000005b00000000",
            INIT_28 => X"000000220000000000000024000000000000002a000000000000003700000000",
            INIT_29 => X"00000008000000000000000d000000000000001a000000000000001d00000000",
            INIT_2A => X"0000000000000000000000030000000000000003000000000000000600000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000500000000000000220000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000570000000000000000000000000000000000000000",
            INIT_34 => X"0000000e00000000000000030000000000000013000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000006000000000000000500000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000080000000000000036000000000000000900000000",
            INIT_38 => X"0000000200000000000000000000000000000000000000000000001200000000",
            INIT_39 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_3A => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000001700000000000000000000000000000000000000000000002e00000000",
            INIT_3C => X"00000000000000000000001d000000000000000a000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"000000000000000000000000000000000000000a000000000000000900000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000001000000000000005000000000",
            INIT_47 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000050000000000000005b00000000",
            INIT_4B => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000000000000000000000000000000000000d000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000b500000000000000310000000000000000000000000000000000000000",
            INIT_52 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000006b00000000000000050000000000000015000000000000000000000000",
            INIT_56 => X"0000001f00000000000000070000000000000000000000000000000000000000",
            INIT_57 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_58 => X"0000000f000000000000000f0000000000000000000000000000000000000000",
            INIT_59 => X"0000000200000000000000100000000000000008000000000000000e00000000",
            INIT_5A => X"00000000000000000000000e0000000000000002000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_5C => X"00000008000000000000000b0000000000000003000000000000000000000000",
            INIT_5D => X"0000000000000000000000060000000000000009000000000000000a00000000",
            INIT_5E => X"00000005000000000000000b0000000000000007000000000000001300000000",
            INIT_5F => X"00000014000000000000000a000000000000000f000000000000000400000000",
            INIT_60 => X"0000000800000000000000000000000000000004000000000000000300000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000010000000000000000000000000000000800000000",
            INIT_63 => X"00000005000000000000001a0000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_66 => X"0000000000000000000000000000000000000003000000000000000800000000",
            INIT_67 => X"0000002000000000000000160000000000000010000000000000002000000000",
            INIT_68 => X"0000002800000000000000250000000000000024000000000000002800000000",
            INIT_69 => X"0000002800000000000000280000000000000028000000000000002600000000",
            INIT_6A => X"00000027000000000000002c0000000000000027000000000000002600000000",
            INIT_6B => X"00000061000000000000001e000000000000000d000000000000000c00000000",
            INIT_6C => X"00000062000000000000005f0000000000000062000000000000006500000000",
            INIT_6D => X"0000004b000000000000005c000000000000005d000000000000006500000000",
            INIT_6E => X"0000000d00000000000000280000000000000028000000000000003300000000",
            INIT_6F => X"0000006700000000000000630000000000000020000000000000000900000000",
            INIT_70 => X"0000005e000000000000006c000000000000006d000000000000006300000000",
            INIT_71 => X"000000330000000000000059000000000000005e000000000000005f00000000",
            INIT_72 => X"0000000c00000000000000110000000000000026000000000000002500000000",
            INIT_73 => X"000000590000000000000058000000000000007c000000000000003100000000",
            INIT_74 => X"00000067000000000000005e0000000000000061000000000000005c00000000",
            INIT_75 => X"000000200000000000000047000000000000005a000000000000006100000000",
            INIT_76 => X"00000014000000000000000f000000000000001a000000000000001e00000000",
            INIT_77 => X"000000190000000000000019000000000000001c000000000000002400000000",
            INIT_78 => X"000000210000000000000020000000000000001e000000000000002300000000",
            INIT_79 => X"0000001c000000000000001d000000000000002a000000000000001d00000000",
            INIT_7A => X"0000001d00000000000000080000000000000014000000000000001d00000000",
            INIT_7B => X"0000002900000000000000250000000000000020000000000000002100000000",
            INIT_7C => X"0000002100000000000000230000000000000022000000000000002700000000",
            INIT_7D => X"0000001e000000000000001f0000000000000022000000000000001f00000000",
            INIT_7E => X"00000006000000000000000b0000000000000025000000000000002500000000",
            INIT_7F => X"0000002700000000000000270000000000000025000000000000001d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "samplegold_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001f00000000000000210000000000000023000000000000002600000000",
            INIT_01 => X"00000022000000000000001e000000000000001e000000000000001f00000000",
            INIT_02 => X"00000007000000000000001c0000000000000043000000000000002b00000000",
            INIT_03 => X"0000002600000000000000290000000000000028000000000000001400000000",
            INIT_04 => X"0000002000000000000000210000000000000022000000000000002500000000",
            INIT_05 => X"0000002800000000000000270000000000000024000000000000001a00000000",
            INIT_06 => X"00000010000000000000001d0000000000000033000000000000003000000000",
            INIT_07 => X"00000022000000000000001d000000000000000f000000000000000700000000",
            INIT_08 => X"0000001c000000000000001f0000000000000024000000000000002800000000",
            INIT_09 => X"0000002c0000000000000029000000000000002a000000000000002900000000",
            INIT_0A => X"00000024000000000000001a0000000000000012000000000000002700000000",
            INIT_0B => X"000000020000000000000000000000000000000a000000000000001b00000000",
            INIT_0C => X"000000220000000000000023000000000000001a000000000000000b00000000",
            INIT_0D => X"0000004700000000000000360000000000000028000000000000002b00000000",
            INIT_0E => X"000000420000000000000034000000000000002f000000000000004500000000",
            INIT_0F => X"0000002900000000000000320000000000000037000000000000003700000000",
            INIT_10 => X"0000000e00000000000000060000000000000026000000000000002e00000000",
            INIT_11 => X"0000000700000000000000030000000000000006000000000000000700000000",
            INIT_12 => X"000000080000000000000008000000000000000a000000000000000800000000",
            INIT_13 => X"00000008000000000000000b000000000000000c000000000000000a00000000",
            INIT_14 => X"0000001c000000000000001e0000000000000016000000000000000b00000000",
            INIT_15 => X"0000001600000000000000180000000000000017000000000000001900000000",
            INIT_16 => X"0000000e00000000000000100000000000000012000000000000001400000000",
            INIT_17 => X"0000000d0000000000000011000000000000000d000000000000000c00000000",
            INIT_18 => X"0000001500000000000000150000000000000016000000000000001200000000",
            INIT_19 => X"0000001500000000000000140000000000000013000000000000001500000000",
            INIT_1A => X"0000001200000000000000120000000000000013000000000000001500000000",
            INIT_1B => X"0000001a0000000000000003000000000000000d000000000000001300000000",
            INIT_1C => X"0000001600000000000000160000000000000017000000000000001600000000",
            INIT_1D => X"0000001d000000000000001d000000000000001f000000000000001c00000000",
            INIT_1E => X"0000000900000000000000150000000000000018000000000000001c00000000",
            INIT_1F => X"00000078000000000000006a0000000000000000000000000000000000000000",
            INIT_20 => X"0000006500000000000000670000000000000057000000000000006000000000",
            INIT_21 => X"00000061000000000000005e0000000000000061000000000000006100000000",
            INIT_22 => X"0000006c00000000000000650000000000000061000000000000006200000000",
            INIT_23 => X"0000007500000000000000830000000000000071000000000000007500000000",
            INIT_24 => X"00000059000000000000005e000000000000004d000000000000003f00000000",
            INIT_25 => X"0000005e0000000000000060000000000000005a000000000000005800000000",
            INIT_26 => X"0000007c000000000000007b000000000000007c000000000000006500000000",
            INIT_27 => X"000000430000000000000075000000000000007f000000000000007100000000",
            INIT_28 => X"000000320000000000000025000000000000002b000000000000003600000000",
            INIT_29 => X"0000004a000000000000003e0000000000000033000000000000003600000000",
            INIT_2A => X"0000006b000000000000007e000000000000007d000000000000007800000000",
            INIT_2B => X"000000400000000000000032000000000000005f000000000000007d00000000",
            INIT_2C => X"000000490000000000000041000000000000003b000000000000004500000000",
            INIT_2D => X"0000005b00000000000000470000000000000043000000000000004100000000",
            INIT_2E => X"0000007b000000000000006c0000000000000080000000000000007c00000000",
            INIT_2F => X"0000006100000000000000600000000000000060000000000000007500000000",
            INIT_30 => X"0000006100000000000000640000000000000061000000000000006200000000",
            INIT_31 => X"0000007a0000000000000071000000000000006d000000000000006100000000",
            INIT_32 => X"0000007900000000000000730000000000000075000000000000008000000000",
            INIT_33 => X"0000006a00000000000000670000000000000068000000000000007c00000000",
            INIT_34 => X"0000006b00000000000000690000000000000069000000000000006c00000000",
            INIT_35 => X"0000007d000000000000007a000000000000007d000000000000007300000000",
            INIT_36 => X"00000054000000000000003c0000000000000064000000000000007900000000",
            INIT_37 => X"0000007d000000000000007e0000000000000089000000000000008a00000000",
            INIT_38 => X"0000007b000000000000007b0000000000000078000000000000007c00000000",
            INIT_39 => X"0000007e0000000000000081000000000000007d000000000000007c00000000",
            INIT_3A => X"00000019000000000000002b000000000000006a000000000000007e00000000",
            INIT_3B => X"0000007a00000000000000840000000000000090000000000000006a00000000",
            INIT_3C => X"0000007a00000000000000780000000000000078000000000000007800000000",
            INIT_3D => X"00000081000000000000007e000000000000007d000000000000007900000000",
            INIT_3E => X"00000020000000000000000d0000000000000073000000000000007f00000000",
            INIT_3F => X"0000008300000000000000840000000000000069000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007b00000000000000790000000000000078000000000000008200000000",
            INIT_41 => X"0000007f000000000000007c000000000000007c000000000000007f00000000",
            INIT_42 => X"00000017000000000000000f0000000000000020000000000000006f00000000",
            INIT_43 => X"0000005b00000000000000330000000000000023000000000000001900000000",
            INIT_44 => X"0000007f00000000000000860000000000000089000000000000007900000000",
            INIT_45 => X"00000068000000000000007e000000000000007c000000000000007c00000000",
            INIT_46 => X"0000002300000000000000040000000000000000000000000000002900000000",
            INIT_47 => X"000000080000000000000011000000000000000a000000000000002300000000",
            INIT_48 => X"0000007800000000000000700000000000000058000000000000003a00000000",
            INIT_49 => X"0000007d000000000000007a000000000000007b000000000000007d00000000",
            INIT_4A => X"000000730000000000000070000000000000005f000000000000006b00000000",
            INIT_4B => X"0000006c0000000000000067000000000000006b000000000000006600000000",
            INIT_4C => X"0000003800000000000000330000000000000074000000000000007100000000",
            INIT_4D => X"0000002e000000000000002e0000000000000030000000000000003100000000",
            INIT_4E => X"000000460000000000000043000000000000003e000000000000003000000000",
            INIT_4F => X"0000004f0000000000000051000000000000004c000000000000004800000000",
            INIT_50 => X"000000230000000000000027000000000000001c000000000000004e00000000",
            INIT_51 => X"0000001600000000000000150000000000000016000000000000001f00000000",
            INIT_52 => X"0000000c000000000000000d0000000000000013000000000000001700000000",
            INIT_53 => X"0000001e000000000000000d000000000000000a000000000000000b00000000",
            INIT_54 => X"000000080000000000000009000000000000000b000000000000000400000000",
            INIT_55 => X"000000090000000000000006000000000000000a000000000000000800000000",
            INIT_56 => X"0000000700000000000000030000000000000004000000000000000700000000",
            INIT_57 => X"00000000000000000000002f000000000000001c000000000000001700000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "samplegold_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000001f00000000000000210000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_19 => X"0000000d000000000000000a0000000000000000000000000000000000000000",
            INIT_1A => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_1E => X"00000019000000000000000c0000000000000034000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000017000000000000001e000000000000001b000000000000002200000000",
            INIT_23 => X"000000000000000000000000000000000000001f000000000000000000000000",
            INIT_24 => X"000000020000000000000000000000000000001a000000000000000f00000000",
            INIT_25 => X"0000002b00000000000000000000000000000018000000000000001100000000",
            INIT_26 => X"0000000000000000000000000000000000000009000000000000002600000000",
            INIT_27 => X"0000001e0000000000000028000000000000001e000000000000002c00000000",
            INIT_28 => X"00000027000000000000002d0000000000000010000000000000000f00000000",
            INIT_29 => X"0000000b00000000000000340000000000000013000000000000001c00000000",
            INIT_2A => X"000000080000000000000000000000000000000e000000000000000f00000000",
            INIT_2B => X"0000001b00000000000000270000000000000005000000000000002400000000",
            INIT_2C => X"000000170000000000000000000000000000001c000000000000002300000000",
            INIT_2D => X"0000002e0000000000000024000000000000001c000000000000003b00000000",
            INIT_2E => X"0000002f00000000000000370000000000000000000000000000000000000000",
            INIT_2F => X"0000003600000000000000220000000000000015000000000000003d00000000",
            INIT_30 => X"00000034000000000000003e000000000000003b000000000000002200000000",
            INIT_31 => X"0000000f00000000000000000000000000000050000000000000005e00000000",
            INIT_32 => X"0000001c000000000000000b000000000000001b000000000000003c00000000",
            INIT_33 => X"0000004200000000000000230000000000000030000000000000005000000000",
            INIT_34 => X"0000002800000000000000320000000000000038000000000000003700000000",
            INIT_35 => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000004f00000000000000400000000000000045000000000000001e00000000",
            INIT_38 => X"0000000b00000000000000250000000000000034000000000000003f00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000002500000000000000060000000000000019000000000000000000000000",
            INIT_3B => X"0000001c000000000000003e0000000000000052000000000000004e00000000",
            INIT_3C => X"0000001e00000000000000220000000000000034000000000000003400000000",
            INIT_3D => X"00000000000000000000002a0000000000000077000000000000004b00000000",
            INIT_3E => X"0000006a00000000000000360000000000000015000000000000000000000000",
            INIT_3F => X"000000380000000000000041000000000000003c000000000000006b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000110000000000000032000000000000001f00000000",
            INIT_41 => X"0000000000000000000000280000000000000059000000000000003200000000",
            INIT_42 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_43 => X"000000480000000000000046000000000000003e000000000000004100000000",
            INIT_44 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000390000000000000049000000000000000000000000",
            INIT_46 => X"00000044000000000000002c0000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000040000000000000006300000000",
            INIT_48 => X"0000002c00000000000000210000000000000020000000000000000000000000",
            INIT_49 => X"00000026000000000000003e0000000000000004000000000000001d00000000",
            INIT_4A => X"00000017000000000000002e000000000000002f000000000000003100000000",
            INIT_4B => X"0000002800000000000000310000000000000006000000000000004900000000",
            INIT_4C => X"0000001a0000000000000020000000000000002c000000000000001f00000000",
            INIT_4D => X"00000039000000000000001c0000000000000031000000000000000800000000",
            INIT_4E => X"0000005000000000000000170000000000000031000000000000002300000000",
            INIT_4F => X"0000001c000000000000001d000000000000003e000000000000000700000000",
            INIT_50 => X"0000000c00000000000000170000000000000020000000000000002000000000",
            INIT_51 => X"0000002200000000000000290000000000000039000000000000003a00000000",
            INIT_52 => X"000000140000000000000052000000000000002a000000000000001200000000",
            INIT_53 => X"0000003800000000000000100000000000000025000000000000002900000000",
            INIT_54 => X"00000042000000000000002e0000000000000013000000000000002100000000",
            INIT_55 => X"0000001400000000000000420000000000000013000000000000002c00000000",
            INIT_56 => X"000000240000000000000018000000000000004e000000000000004200000000",
            INIT_57 => X"00000004000000000000003d0000000000000018000000000000000000000000",
            INIT_58 => X"0000000d00000000000000300000000000000043000000000000002600000000",
            INIT_59 => X"0000003a00000000000000460000000000000032000000000000004800000000",
            INIT_5A => X"0000000000000000000000200000000000000029000000000000004600000000",
            INIT_5B => X"0000000c000000000000001f000000000000003d000000000000001300000000",
            INIT_5C => X"0000003800000000000000380000000000000034000000000000003c00000000",
            INIT_5D => X"0000005900000000000000290000000000000030000000000000003200000000",
            INIT_5E => X"000000170000000000000000000000000000001d000000000000002700000000",
            INIT_5F => X"00000032000000000000001f000000000000002c000000000000003500000000",
            INIT_60 => X"00000035000000000000003c000000000000003c000000000000004100000000",
            INIT_61 => X"00000024000000000000003f000000000000003a000000000000003900000000",
            INIT_62 => X"0000002d00000000000000180000000000000000000000000000003100000000",
            INIT_63 => X"0000003c00000000000000210000000000000027000000000000002900000000",
            INIT_64 => X"00000041000000000000003a0000000000000045000000000000003b00000000",
            INIT_65 => X"0000002c00000000000000210000000000000038000000000000004200000000",
            INIT_66 => X"000000210000000000000030000000000000002a000000000000000000000000",
            INIT_67 => X"00000041000000000000001f000000000000003c000000000000002100000000",
            INIT_68 => X"0000003b00000000000000360000000000000039000000000000003600000000",
            INIT_69 => X"0000000b0000000000000028000000000000002e000000000000003b00000000",
            INIT_6A => X"0000002b00000000000000160000000000000019000000000000002800000000",
            INIT_6B => X"000000320000000000000032000000000000003e000000000000001a00000000",
            INIT_6C => X"000000320000000000000033000000000000002f000000000000003900000000",
            INIT_6D => X"00000006000000000000003a0000000000000022000000000000001500000000",
            INIT_6E => X"00000038000000000000002b0000000000000022000000000000003100000000",
            INIT_6F => X"00000027000000000000002f0000000000000045000000000000001c00000000",
            INIT_70 => X"0000002b00000000000000300000000000000032000000000000002c00000000",
            INIT_71 => X"0000004100000000000000330000000000000024000000000000003100000000",
            INIT_72 => X"0000003b0000000000000011000000000000003d000000000000002c00000000",
            INIT_73 => X"0000002600000000000000310000000000000034000000000000003400000000",
            INIT_74 => X"0000003b00000000000000370000000000000038000000000000003700000000",
            INIT_75 => X"0000003000000000000000410000000000000031000000000000002000000000",
            INIT_76 => X"000000330000000000000036000000000000002f000000000000003f00000000",
            INIT_77 => X"00000034000000000000002d0000000000000039000000000000002b00000000",
            INIT_78 => X"00000025000000000000003e000000000000002b000000000000002d00000000",
            INIT_79 => X"0000003b00000000000000460000000000000042000000000000001100000000",
            INIT_7A => X"00000027000000000000003d000000000000003b000000000000003c00000000",
            INIT_7B => X"0000003200000000000000320000000000000032000000000000004800000000",
            INIT_7C => X"000000180000000000000028000000000000003e000000000000001200000000",
            INIT_7D => X"0000003a00000000000000540000000000000059000000000000002400000000",
            INIT_7E => X"0000003700000000000000370000000000000039000000000000003900000000",
            INIT_7F => X"000000260000000000000025000000000000002f000000000000003800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "samplegold_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000057000000000000002c00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000300000000000000010000000000000000000000000000000000000000",
            INIT_13 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_1B => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000000000000000000000c0000000000000000000000000000000400000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_24 => X"000000000000000000000006000000000000000b000000000000000300000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000c00000000000000070000000000000000000000000000000000000000",
            INIT_28 => X"000000000000000000000000000000000000000d000000000000001100000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000f000000000000000e0000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_2D => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_2F => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000b000000000000002f000000000000001a000000000000000d00000000",
            INIT_3A => X"0000003400000000000000230000000000000023000000000000000500000000",
            INIT_3B => X"0000003d0000000000000044000000000000003c000000000000004300000000",
            INIT_3C => X"00000027000000000000004d000000000000002d000000000000001700000000",
            INIT_3D => X"000000000000000000000006000000000000003b000000000000003300000000",
            INIT_3E => X"00000033000000000000003d000000000000001f000000000000001e00000000",
            INIT_3F => X"0000002800000000000000600000000000000048000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000430000000000000043000000000000003e000000000000004600000000",
            INIT_41 => X"00000021000000000000000c0000000000000005000000000000003300000000",
            INIT_42 => X"00000041000000000000001b0000000000000048000000000000002500000000",
            INIT_43 => X"00000064000000000000005a0000000000000089000000000000005200000000",
            INIT_44 => X"0000003400000000000000360000000000000034000000000000002000000000",
            INIT_45 => X"000000170000000000000036000000000000002a000000000000000c00000000",
            INIT_46 => X"000000580000000000000038000000000000003b000000000000002600000000",
            INIT_47 => X"0000002b000000000000005e0000000000000079000000000000009a00000000",
            INIT_48 => X"0000003c0000000000000016000000000000006b000000000000006c00000000",
            INIT_49 => X"0000003f000000000000001a0000000000000033000000000000005b00000000",
            INIT_4A => X"00000087000000000000005d0000000000000057000000000000004400000000",
            INIT_4B => X"00000063000000000000002d0000000000000047000000000000008600000000",
            INIT_4C => X"0000005900000000000000380000000000000053000000000000009700000000",
            INIT_4D => X"000000620000000000000066000000000000006c000000000000005400000000",
            INIT_4E => X"00000089000000000000007f0000000000000055000000000000005d00000000",
            INIT_4F => X"0000007c000000000000004d0000000000000031000000000000003b00000000",
            INIT_50 => X"00000056000000000000005c0000000000000065000000000000008b00000000",
            INIT_51 => X"0000006b00000000000000660000000000000062000000000000005b00000000",
            INIT_52 => X"0000004f00000000000000770000000000000077000000000000007200000000",
            INIT_53 => X"0000008700000000000000700000000000000057000000000000004700000000",
            INIT_54 => X"0000006f00000000000000680000000000000033000000000000008400000000",
            INIT_55 => X"0000008a00000000000000650000000000000067000000000000007500000000",
            INIT_56 => X"000000580000000000000032000000000000007b000000000000008400000000",
            INIT_57 => X"000000770000000000000075000000000000006b000000000000006300000000",
            INIT_58 => X"0000007c00000000000000810000000000000065000000000000009600000000",
            INIT_59 => X"00000084000000000000007e000000000000007a000000000000008400000000",
            INIT_5A => X"0000006800000000000000680000000000000043000000000000006900000000",
            INIT_5B => X"000000620000000000000064000000000000005b000000000000004400000000",
            INIT_5C => X"0000009600000000000000920000000000000093000000000000009800000000",
            INIT_5D => X"000000380000000000000061000000000000007a000000000000007e00000000",
            INIT_5E => X"00000046000000000000004f0000000000000059000000000000005400000000",
            INIT_5F => X"0000008300000000000000640000000000000053000000000000005500000000",
            INIT_60 => X"00000084000000000000008700000000000000a000000000000000ac00000000",
            INIT_61 => X"0000006800000000000000600000000000000065000000000000007800000000",
            INIT_62 => X"000000520000000000000058000000000000007f000000000000007800000000",
            INIT_63 => X"000000a2000000000000008e0000000000000067000000000000006900000000",
            INIT_64 => X"00000073000000000000008a000000000000008800000000000000a300000000",
            INIT_65 => X"0000006b00000000000000760000000000000063000000000000005a00000000",
            INIT_66 => X"0000005d000000000000006e00000000000000a800000000000000a600000000",
            INIT_67 => X"00000085000000000000006a0000000000000083000000000000006d00000000",
            INIT_68 => X"0000004d000000000000007b0000000000000089000000000000009a00000000",
            INIT_69 => X"0000001a00000000000000380000000000000060000000000000004100000000",
            INIT_6A => X"00000057000000000000007a00000000000000a6000000000000008b00000000",
            INIT_6B => X"000000890000000000000048000000000000005e000000000000005700000000",
            INIT_6C => X"000000320000000000000039000000000000006e000000000000009100000000",
            INIT_6D => X"0000000f000000000000000a0000000000000033000000000000007600000000",
            INIT_6E => X"0000006a000000000000009300000000000000b4000000000000008a00000000",
            INIT_6F => X"0000006d0000000000000071000000000000004c000000000000006500000000",
            INIT_70 => X"00000056000000000000003a0000000000000037000000000000006c00000000",
            INIT_71 => X"0000003d00000000000000240000000000000030000000000000003000000000",
            INIT_72 => X"000000390000000000000040000000000000001a000000000000004e00000000",
            INIT_73 => X"0000002800000000000000630000000000000066000000000000005800000000",
            INIT_74 => X"000000360000000000000037000000000000003f000000000000007a00000000",
            INIT_75 => X"0000004f0000000000000039000000000000004b000000000000003300000000",
            INIT_76 => X"0000004e000000000000002d0000000000000050000000000000003000000000",
            INIT_77 => X"0000006b000000000000001a0000000000000064000000000000003c00000000",
            INIT_78 => X"0000006c00000000000000670000000000000044000000000000000400000000",
            INIT_79 => X"00000018000000000000004e0000000000000044000000000000004800000000",
            INIT_7A => X"0000005e0000000000000053000000000000004c000000000000002500000000",
            INIT_7B => X"000000450000000000000061000000000000001b000000000000004c00000000",
            INIT_7C => X"0000003a00000000000000120000000000000053000000000000004600000000",
            INIT_7D => X"0000007b00000000000000310000000000000029000000000000004600000000",
            INIT_7E => X"0000002000000000000000450000000000000026000000000000007d00000000",
            INIT_7F => X"0000006f00000000000000480000000000000077000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "samplegold_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003e00000000000000530000000000000026000000000000004700000000",
            INIT_01 => X"0000000d000000000000006b000000000000004c000000000000002d00000000",
            INIT_02 => X"000000750000000000000067000000000000003e000000000000004600000000",
            INIT_03 => X"0000005d000000000000007e0000000000000052000000000000006c00000000",
            INIT_04 => X"00000025000000000000003e000000000000005a000000000000003400000000",
            INIT_05 => X"0000004d00000000000000200000000000000037000000000000004600000000",
            INIT_06 => X"00000080000000000000002f0000000000000060000000000000005700000000",
            INIT_07 => X"0000002700000000000000400000000000000074000000000000005800000000",
            INIT_08 => X"0000004800000000000000500000000000000055000000000000004f00000000",
            INIT_09 => X"0000003d000000000000004b000000000000003b000000000000003900000000",
            INIT_0A => X"0000004c000000000000006a0000000000000034000000000000002e00000000",
            INIT_0B => X"00000040000000000000003d000000000000005b000000000000006a00000000",
            INIT_0C => X"0000003c000000000000003a000000000000002d000000000000005b00000000",
            INIT_0D => X"0000002f00000000000000200000000000000038000000000000003700000000",
            INIT_0E => X"00000080000000000000005b000000000000003f000000000000003400000000",
            INIT_0F => X"0000006500000000000000610000000000000035000000000000003300000000",
            INIT_10 => X"0000003a00000000000000220000000000000036000000000000004d00000000",
            INIT_11 => X"0000003f000000000000004b0000000000000049000000000000003600000000",
            INIT_12 => X"000000430000000000000060000000000000006f000000000000006400000000",
            INIT_13 => X"0000006400000000000000540000000000000069000000000000007300000000",
            INIT_14 => X"000000390000000000000026000000000000003c000000000000004700000000",
            INIT_15 => X"000000580000000000000049000000000000003f000000000000004100000000",
            INIT_16 => X"0000003e00000000000000750000000000000031000000000000003900000000",
            INIT_17 => X"0000004d000000000000003e0000000000000037000000000000005700000000",
            INIT_18 => X"0000004e000000000000003e0000000000000041000000000000002000000000",
            INIT_19 => X"0000003a000000000000004b0000000000000048000000000000004a00000000",
            INIT_1A => X"0000005c0000000000000005000000000000001c000000000000003d00000000",
            INIT_1B => X"00000039000000000000003a000000000000005f000000000000004500000000",
            INIT_1C => X"0000002c00000000000000420000000000000049000000000000004d00000000",
            INIT_1D => X"0000007300000000000000540000000000000065000000000000004300000000",
            INIT_1E => X"0000006e000000000000007d0000000000000092000000000000007a00000000",
            INIT_1F => X"0000007c00000000000000520000000000000045000000000000007200000000",
            INIT_20 => X"0000004a0000000000000038000000000000003e000000000000006100000000",
            INIT_21 => X"0000005c00000000000000770000000000000063000000000000005100000000",
            INIT_22 => X"000000730000000000000076000000000000009a000000000000007400000000",
            INIT_23 => X"0000001300000000000000560000000000000078000000000000007600000000",
            INIT_24 => X"0000008400000000000000550000000000000043000000000000004500000000",
            INIT_25 => X"00000049000000000000006a000000000000005f000000000000004100000000",
            INIT_26 => X"00000065000000000000007d0000000000000092000000000000004800000000",
            INIT_27 => X"0000005e000000000000006e0000000000000074000000000000007000000000",
            INIT_28 => X"0000002a0000000000000034000000000000006e000000000000006b00000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_2A => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_2B => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000150000000000000007000000000000000000000000",
            INIT_2F => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_30 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_32 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000005000000000000000300000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000020000000000000000000000000",
            INIT_37 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000001500000000000000000000000000000000000000000000000b00000000",
            INIT_3C => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000800000000000000000000000000000000000000000000000e00000000",
            INIT_48 => X"000000000000000000000000000000000000000e000000000000000b00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000000000000000000017000000000000001f000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_4C => X"000000000000000000000000000000000000003c000000000000000800000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"00000000000000000000004a0000000000000021000000000000000000000000",
            INIT_57 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000034000000000000002d00000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"00000000000000000000004e0000000000000030000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_5D => X"0000000900000000000000000000000000000000000000000000002100000000",
            INIT_5E => X"0000000000000000000000340000000000000017000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"00000000000000000000000d000000000000003a000000000000002100000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000005f00000000000000000000000000000009000000000000001d00000000",
            INIT_63 => X"0000001c00000000000000070000000000000026000000000000000000000000",
            INIT_64 => X"000000410000000000000000000000000000007b000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_66 => X"00000006000000000000003e0000000000000000000000000000000800000000",
            INIT_67 => X"0000000000000000000000180000000000000000000000000000003b00000000",
            INIT_68 => X"00000000000000000000003a0000000000000000000000000000009b00000000",
            INIT_69 => X"0000000000000000000000010000000000000017000000000000000000000000",
            INIT_6A => X"0000000000000000000000180000000000000046000000000000000000000000",
            INIT_6B => X"0000008800000000000000320000000000000000000000000000002d00000000",
            INIT_6C => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_6D => X"0000000200000000000000000000000000000000000000000000006300000000",
            INIT_6E => X"0000006300000000000000000000000000000000000000000000004100000000",
            INIT_6F => X"00000000000000000000005e0000000000000034000000000000000000000000",
            INIT_70 => X"0000008a00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000200000000000000640000000000000000000000000000000000000000",
            INIT_72 => X"0000002400000000000000000000000000000053000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_74 => X"00000003000000000000008d0000000000000000000000000000000000000000",
            INIT_75 => X"00000000000000000000000f000000000000002e000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_77 => X"00000000000000000000000f0000000000000000000000000000006500000000",
            INIT_78 => X"000000000000000000000039000000000000004d000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_7A => X"0000000f0000000000000008000000000000000f000000000000000000000000",
            INIT_7B => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_7C => X"0000000500000000000000000000000000000025000000000000004000000000",
            INIT_7D => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_7E => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_7F => X"00000012000000000000000c0000000000000000000000000000000800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "samplegold_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_02 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_04 => X"000000110000000000000029000000000000000b000000000000003200000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_06 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000002a00000000000000000000000000000044000000000000000000000000",
            INIT_08 => X"0000000000000000000000630000000000000000000000000000000800000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000e00000000000000120000000000000001000000000000000000000000",
            INIT_0B => X"00000000000000000000001f0000000000000000000000000000000e00000000",
            INIT_0C => X"0000000000000000000000040000000000000034000000000000002200000000",
            INIT_0D => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_0E => X"00000064000000000000001f0000000000000000000000000000002e00000000",
            INIT_0F => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000004a0000000000000000000000000000000e00000000",
            INIT_11 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000009300000000000000450000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_14 => X"0000000600000000000000120000000000000035000000000000000000000000",
            INIT_15 => X"0000002b00000000000000590000000000000000000000000000000000000000",
            INIT_16 => X"0000008b00000000000000750000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_18 => X"0000000000000000000000060000000000000018000000000000000000000000",
            INIT_19 => X"0000002400000000000000850000000000000000000000000000000000000000",
            INIT_1A => X"00000022000000000000002b000000000000002a000000000000002900000000",
            INIT_1B => X"0000000000000000000000170000000000000019000000000000002400000000",
            INIT_1C => X"000000020000000000000011000000000000000a000000000000000000000000",
            INIT_1D => X"0000002400000000000000260000000000000020000000000000000300000000",
            INIT_1E => X"0000000a00000000000000200000000000000027000000000000001d00000000",
            INIT_1F => X"000000160000000000000016000000000000001d000000000000000b00000000",
            INIT_20 => X"00000035000000000000001b0000000000000011000000000000000e00000000",
            INIT_21 => X"0000001a00000000000000000000000000000000000000000000001f00000000",
            INIT_22 => X"000000330000000000000036000000000000001b000000000000001900000000",
            INIT_23 => X"000000120000000000000000000000000000000c000000000000001100000000",
            INIT_24 => X"0000001e000000000000001c000000000000000f000000000000001200000000",
            INIT_25 => X"0000001a000000000000001d0000000000000032000000000000001a00000000",
            INIT_26 => X"0000000000000000000000000000000000000019000000000000002a00000000",
            INIT_27 => X"00000000000000000000001c0000000000000023000000000000001900000000",
            INIT_28 => X"0000002000000000000000020000000000000014000000000000000000000000",
            INIT_29 => X"0000001b00000000000000110000000000000027000000000000001b00000000",
            INIT_2A => X"0000001b00000000000000340000000000000007000000000000000a00000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_2C => X"00000008000000000000000d0000000000000010000000000000001300000000",
            INIT_2D => X"0000000000000000000000150000000000000044000000000000001d00000000",
            INIT_2E => X"0000000000000000000000030000000000000017000000000000000800000000",
            INIT_2F => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"00000004000000000000001b0000000000000025000000000000001500000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000002100000000000000110000000000000000000000000000000000000000",
            INIT_34 => X"0000000200000000000000160000000000000015000000000000001000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_36 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_37 => X"0000002500000000000000000000000000000000000000000000000300000000",
            INIT_38 => X"0000000000000000000000020000000000000001000000000000001f00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000000000014000000000000001c000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000001900000000000000060000000000000000000000000000002e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000d0000000000000021000000000000002300000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001a00000000000000220000000000000000000000000000000000000000",
            INIT_43 => X"0000001600000000000000160000000000000030000000000000003f00000000",
            INIT_44 => X"0000000000000000000000000000000000000017000000000000000800000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_47 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000160000000000000018000000000000000000000000",
            INIT_4D => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000001b0000000000000007000000000000002100000000",
            INIT_4F => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000035000000000000002e000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "samplegold_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000004800000000000000280000000000000033000000000000000000000000",
            INIT_0B => X"00000026000000000000003a0000000000000000000000000000003500000000",
            INIT_0C => X"000000120000000000000018000000000000001c000000000000002b00000000",
            INIT_0D => X"00000033000000000000001a0000000000000000000000000000004e00000000",
            INIT_0E => X"00000036000000000000002c0000000000000041000000000000003b00000000",
            INIT_0F => X"00000039000000000000000c0000000000000018000000000000000000000000",
            INIT_10 => X"0000005c0000000000000010000000000000003a000000000000003100000000",
            INIT_11 => X"00000000000000000000003a000000000000006a000000000000002300000000",
            INIT_12 => X"0000000000000000000000160000000000000029000000000000000600000000",
            INIT_13 => X"0000002400000000000000260000000000000064000000000000005000000000",
            INIT_14 => X"0000003500000000000000660000000000000029000000000000000000000000",
            INIT_15 => X"0000006d00000000000000160000000000000035000000000000004900000000",
            INIT_16 => X"000000670000000000000033000000000000001a000000000000002d00000000",
            INIT_17 => X"0000002b000000000000003f0000000000000000000000000000001a00000000",
            INIT_18 => X"0000004400000000000000260000000000000063000000000000006100000000",
            INIT_19 => X"00000041000000000000005e0000000000000022000000000000000000000000",
            INIT_1A => X"0000000700000000000000440000000000000050000000000000000c00000000",
            INIT_1B => X"0000003500000000000000600000000000000050000000000000006500000000",
            INIT_1C => X"0000000000000000000000390000000000000033000000000000002b00000000",
            INIT_1D => X"00000056000000000000003e000000000000003e000000000000000000000000",
            INIT_1E => X"0000005b00000000000000180000000000000023000000000000006800000000",
            INIT_1F => X"00000068000000000000001c000000000000002d000000000000004300000000",
            INIT_20 => X"0000003200000000000000000000000000000039000000000000002300000000",
            INIT_21 => X"0000000e0000000000000039000000000000003b000000000000004b00000000",
            INIT_22 => X"0000000a00000000000000240000000000000030000000000000001400000000",
            INIT_23 => X"000000230000000000000039000000000000002a000000000000001500000000",
            INIT_24 => X"00000044000000000000001a0000000000000005000000000000004b00000000",
            INIT_25 => X"0000000a000000000000004d0000000000000027000000000000004b00000000",
            INIT_26 => X"00000047000000000000002f000000000000001f000000000000002100000000",
            INIT_27 => X"00000030000000000000002f000000000000002e000000000000002700000000",
            INIT_28 => X"0000001a0000000000000050000000000000004c000000000000000000000000",
            INIT_29 => X"00000029000000000000003a000000000000000c000000000000001e00000000",
            INIT_2A => X"00000015000000000000001a000000000000002c000000000000002100000000",
            INIT_2B => X"0000002000000000000000000000000000000000000000000000002500000000",
            INIT_2C => X"0000002200000000000000130000000000000009000000000000003700000000",
            INIT_2D => X"0000003f00000000000000270000000000000000000000000000002600000000",
            INIT_2E => X"0000001500000000000000200000000000000021000000000000002100000000",
            INIT_2F => X"000000000000000000000047000000000000002e000000000000000c00000000",
            INIT_30 => X"0000003a00000000000000470000000000000026000000000000004200000000",
            INIT_31 => X"0000002a00000000000000270000000000000040000000000000003b00000000",
            INIT_32 => X"0000001800000000000000160000000000000011000000000000000300000000",
            INIT_33 => X"000000a0000000000000006e000000000000005e000000000000003a00000000",
            INIT_34 => X"00000030000000000000002f0000000000000055000000000000005d00000000",
            INIT_35 => X"0000001400000000000000190000000000000015000000000000003400000000",
            INIT_36 => X"0000003800000000000000000000000000000012000000000000002d00000000",
            INIT_37 => X"0000004d00000000000000030000000000000000000000000000003700000000",
            INIT_38 => X"000000150000000000000042000000000000003c000000000000005800000000",
            INIT_39 => X"0000001c00000000000000230000000000000000000000000000000000000000",
            INIT_3A => X"0000002d00000000000000190000000000000005000000000000000e00000000",
            INIT_3B => X"0000005200000000000000040000000000000000000000000000000f00000000",
            INIT_3C => X"0000004100000000000000310000000000000050000000000000005400000000",
            INIT_3D => X"0000000000000000000000230000000000000013000000000000005100000000",
            INIT_3E => X"00000001000000000000004b0000000000000034000000000000000000000000",
            INIT_3F => X"000000490000000000000018000000000000000e000000000000002700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000080000000000000048000000000000005f000000000000006c00000000",
            INIT_41 => X"0000004800000000000000020000000000000000000000000000000000000000",
            INIT_42 => X"0000000d000000000000000e0000000000000082000000000000005d00000000",
            INIT_43 => X"0000000000000000000000020000000000000002000000000000000a00000000",
            INIT_44 => X"0000001900000000000000220000000000000009000000000000000f00000000",
            INIT_45 => X"0000000700000000000000360000000000000010000000000000001900000000",
            INIT_46 => X"0000001600000000000000200000000000000019000000000000000d00000000",
            INIT_47 => X"0000000100000000000000000000000000000007000000000000000500000000",
            INIT_48 => X"0000001900000000000000190000000000000018000000000000000d00000000",
            INIT_49 => X"0000001e00000000000000160000000000000037000000000000001400000000",
            INIT_4A => X"0000000a000000000000000a0000000000000005000000000000001600000000",
            INIT_4B => X"0000001b00000000000000190000000000000002000000000000000100000000",
            INIT_4C => X"000000230000000000000006000000000000001c000000000000000300000000",
            INIT_4D => X"0000000c00000000000000220000000000000025000000000000003f00000000",
            INIT_4E => X"00000007000000000000000b0000000000000025000000000000000b00000000",
            INIT_4F => X"0000000e000000000000000f000000000000002f000000000000002500000000",
            INIT_50 => X"000000330000000000000035000000000000002c000000000000000a00000000",
            INIT_51 => X"0000000e00000000000000120000000000000026000000000000002900000000",
            INIT_52 => X"00000031000000000000000c0000000000000020000000000000002200000000",
            INIT_53 => X"0000002f000000000000002e000000000000000b000000000000002f00000000",
            INIT_54 => X"00000026000000000000003f0000000000000039000000000000003900000000",
            INIT_55 => X"0000001f000000000000000b0000000000000018000000000000001d00000000",
            INIT_56 => X"0000002b00000000000000350000000000000031000000000000002800000000",
            INIT_57 => X"0000003d000000000000003c000000000000003d000000000000002600000000",
            INIT_58 => X"00000023000000000000001b0000000000000043000000000000003000000000",
            INIT_59 => X"0000003200000000000000220000000000000017000000000000001700000000",
            INIT_5A => X"0000004a000000000000003d0000000000000045000000000000004400000000",
            INIT_5B => X"0000004a00000000000000350000000000000036000000000000003a00000000",
            INIT_5C => X"000000180000000000000022000000000000002b000000000000003b00000000",
            INIT_5D => X"00000030000000000000002a0000000000000024000000000000001400000000",
            INIT_5E => X"0000004700000000000000470000000000000038000000000000004e00000000",
            INIT_5F => X"000000490000000000000030000000000000004e000000000000005000000000",
            INIT_60 => X"0000002b000000000000001a0000000000000023000000000000002800000000",
            INIT_61 => X"00000024000000000000003c0000000000000022000000000000002400000000",
            INIT_62 => X"0000004c000000000000004f0000000000000043000000000000004600000000",
            INIT_63 => X"00000027000000000000003c0000000000000046000000000000004a00000000",
            INIT_64 => X"0000001900000000000000210000000000000024000000000000000f00000000",
            INIT_65 => X"0000003500000000000000340000000000000017000000000000001200000000",
            INIT_66 => X"000000440000000000000049000000000000004e000000000000004000000000",
            INIT_67 => X"0000001600000000000000150000000000000030000000000000004700000000",
            INIT_68 => X"0000001500000000000000230000000000000012000000000000002400000000",
            INIT_69 => X"0000004d0000000000000034000000000000001b000000000000003100000000",
            INIT_6A => X"000000440000000000000040000000000000004a000000000000004100000000",
            INIT_6B => X"000000260000000000000025000000000000001c000000000000003d00000000",
            INIT_6C => X"0000001d000000000000002f0000000000000055000000000000005100000000",
            INIT_6D => X"00000044000000000000004d000000000000003c000000000000002e00000000",
            INIT_6E => X"00000049000000000000004b0000000000000042000000000000004100000000",
            INIT_6F => X"0000002e000000000000002d0000000000000025000000000000002500000000",
            INIT_70 => X"0000001c000000000000003f000000000000005e000000000000005500000000",
            INIT_71 => X"0000003c00000000000000220000000000000045000000000000004100000000",
            INIT_72 => X"00000022000000000000003e0000000000000049000000000000004c00000000",
            INIT_73 => X"000000250000000000000022000000000000001d000000000000002700000000",
            INIT_74 => X"00000042000000000000004c0000000000000066000000000000004c00000000",
            INIT_75 => X"0000003c000000000000003f0000000000000037000000000000002800000000",
            INIT_76 => X"000000190000000000000007000000000000002a000000000000004b00000000",
            INIT_77 => X"0000003600000000000000290000000000000008000000000000002000000000",
            INIT_78 => X"0000004e000000000000005a0000000000000063000000000000004d00000000",
            INIT_79 => X"00000028000000000000002e000000000000002e000000000000004000000000",
            INIT_7A => X"0000000000000000000000460000000000000029000000000000002a00000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_7F => X"0000001b00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "samplegold_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_01 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_02 => X"0000000000000000000000130000000000000025000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_04 => X"0000000000000000000000200000000000000015000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000002100000000000000010000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_0D => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_19 => X"000000370000000000000019000000000000001e000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_1B => X"0000001f00000000000000000000000000000000000000000000000500000000",
            INIT_1C => X"0000002000000000000000000000000000000000000000000000002300000000",
            INIT_1D => X"0000005e000000000000000d0000000000000009000000000000000500000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_21 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000700000000000000020000000000000002000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_27 => X"0000005800000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000005b00000000",
            INIT_29 => X"0000004900000000000000430000000000000018000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_2B => X"0000007f00000000000000000000000000000005000000000000001a00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000006300000000",
            INIT_2D => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"00000000000000000000001f0000000000000003000000000000000000000000",
            INIT_2F => X"0000005d00000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000004d00000000",
            INIT_31 => X"0000004b00000000000000250000000000000018000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_34 => X"0000000000000000000000090000000000000000000000000000004500000000",
            INIT_35 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000007f00000000",
            INIT_37 => X"0000005100000000000000000000000000000000000000000000001700000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"000000490000000000000000000000000000001e000000000000000000000000",
            INIT_3A => X"00000000000000000000002a0000000000000013000000000000000000000000",
            INIT_3B => X"000000000000000000000044000000000000000d000000000000000000000000",
            INIT_3C => X"000000470000000000000000000000000000001e000000000000000000000000",
            INIT_3D => X"0000000000000000000000290000000000000000000000000000000000000000",
            INIT_3E => X"0000002500000000000000000000000000000016000000000000000000000000",
            INIT_3F => X"0000002500000000000000000000000000000000000000000000002100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000120000000000000000000000000000002100000000",
            INIT_41 => X"0000005800000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"00000025000000000000003b0000000000000000000000000000002d00000000",
            INIT_43 => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000004e00000000000000830000000000000000000000000000000000000000",
            INIT_46 => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_47 => X"0000000b00000000000000000000000000000010000000000000000000000000",
            INIT_48 => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000380000000000000093000000000000000000000000",
            INIT_4A => X"00000000000000000000001d0000000000000007000000000000000000000000",
            INIT_4B => X"0000000000000000000000030000000000000002000000000000000000000000",
            INIT_4C => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000022000000000000006400000000",
            INIT_4E => X"0000000000000000000000340000000000000000000000000000000000000000",
            INIT_4F => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000007800000000000000000000000000000046000000000000000000000000",
            INIT_51 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_52 => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_53 => X"0000000f00000000000000000000000000000000000000000000000b00000000",
            INIT_54 => X"000000090000000000000043000000000000000d000000000000001400000000",
            INIT_55 => X"000000000000000000000000000000000000002f000000000000000d00000000",
            INIT_56 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_57 => X"0000003300000000000000130000000000000006000000000000001400000000",
            INIT_58 => X"0000000000000000000000470000000000000000000000000000000700000000",
            INIT_59 => X"0000002000000000000000000000000000000000000000000000002800000000",
            INIT_5A => X"0000001100000000000000100000000000000005000000000000000000000000",
            INIT_5B => X"00000000000000000000001a0000000000000003000000000000000400000000",
            INIT_5C => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_5E => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_5F => X"000000000000000000000000000000000000001d000000000000001300000000",
            INIT_60 => X"0000002500000000000000000000000000000000000000000000000100000000",
            INIT_61 => X"0000003e00000000000000000000000000000000000000000000002500000000",
            INIT_62 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"00000031000000000000000b0000000000000000000000000000003500000000",
            INIT_64 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_66 => X"0000005900000000000000360000000000000000000000000000000000000000",
            INIT_67 => X"0000000f000000000000003a0000000000000000000000000000000000000000",
            INIT_68 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000230000000000000000000000000000001200000000",
            INIT_6A => X"00000000000000000000001f0000000000000000000000000000000600000000",
            INIT_6B => X"000000000000000000000007000000000000000a000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000100000000000000000000000000000017000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000003000000000000000300000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000010000000000000007000000000000002000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_75 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_77 => X"000000000000000000000004000000000000000a000000000000000500000000",
            INIT_78 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000001000000000000000c0000000000000000000000000000000e00000000",
            INIT_7A => X"0000000700000000000000000000000000000000000000000000000900000000",
            INIT_7B => X"0000000900000000000000000000000000000003000000000000000700000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_7D => X"0000000900000000000000000000000000000007000000000000000000000000",
            INIT_7E => X"0000001000000000000000000000000000000000000000000000000100000000",
            INIT_7F => X"0000001a0000000000000032000000000000001c000000000000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "samplegold_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000010000000000000016000000000000000c000000000000000f00000000",
            INIT_01 => X"0000000600000000000000140000000000000000000000000000000100000000",
            INIT_02 => X"0000002f00000000000000070000000000000000000000000000000000000000",
            INIT_03 => X"00000037000000000000003d0000000000000045000000000000004200000000",
            INIT_04 => X"0000001100000000000000370000000000000041000000000000003c00000000",
            INIT_05 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_06 => X"0000003500000000000000420000000000000002000000000000000000000000",
            INIT_07 => X"0000005400000000000000510000000000000049000000000000003f00000000",
            INIT_08 => X"0000000200000000000000460000000000000038000000000000004800000000",
            INIT_09 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_0A => X"00000043000000000000004a0000000000000019000000000000000000000000",
            INIT_0B => X"000000460000000000000048000000000000004e000000000000004900000000",
            INIT_0C => X"00000004000000000000000d000000000000003b000000000000003e00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000004a00000000000000460000000000000018000000000000000000000000",
            INIT_0F => X"000000430000000000000043000000000000004d000000000000004c00000000",
            INIT_10 => X"000000000000000000000000000000000000000a000000000000003700000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_12 => X"000000480000000000000049000000000000002f000000000000000c00000000",
            INIT_13 => X"0000003a00000000000000480000000000000048000000000000004600000000",
            INIT_14 => X"0000003200000000000000190000000000000000000000000000000d00000000",
            INIT_15 => X"0000000900000000000000000000000000000000000000000000001500000000",
            INIT_16 => X"000000450000000000000043000000000000004e000000000000003400000000",
            INIT_17 => X"00000006000000000000003a000000000000004d000000000000005100000000",
            INIT_18 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000002600000000000000000000000000000000000000000000000800000000",
            INIT_1A => X"00000049000000000000004c0000000000000025000000000000003600000000",
            INIT_1B => X"000000000000000000000000000000000000003c000000000000005000000000",
            INIT_1C => X"0000000e00000000000000000000000000000000000000000000000500000000",
            INIT_1D => X"0000001300000000000000000000000000000000000000000000000f00000000",
            INIT_1E => X"0000004600000000000000460000000000000043000000000000001c00000000",
            INIT_1F => X"0000000300000000000000000000000000000000000000000000002300000000",
            INIT_20 => X"0000000f00000000000000000000000000000000000000000000000100000000",
            INIT_21 => X"0000000d00000000000000000000000000000000000000000000000e00000000",
            INIT_22 => X"0000001c00000000000000270000000000000029000000000000002e00000000",
            INIT_23 => X"0000000000000000000000110000000000000001000000000000000900000000",
            INIT_24 => X"0000000d0000000000000000000000000000001b000000000000000f00000000",
            INIT_25 => X"0000002c00000000000000200000000000000017000000000000000d00000000",
            INIT_26 => X"0000001700000000000000030000000000000030000000000000001500000000",
            INIT_27 => X"00000019000000000000000a0000000000000021000000000000000f00000000",
            INIT_28 => X"0000001300000000000000070000000000000000000000000000001f00000000",
            INIT_29 => X"00000016000000000000001b000000000000001d000000000000001300000000",
            INIT_2A => X"0000001f00000000000000120000000000000013000000000000003500000000",
            INIT_2B => X"00000019000000000000001e0000000000000029000000000000002200000000",
            INIT_2C => X"0000001300000000000000100000000000000009000000000000000000000000",
            INIT_2D => X"0000003a00000000000000280000000000000008000000000000003000000000",
            INIT_2E => X"0000000a0000000000000029000000000000002c000000000000003100000000",
            INIT_2F => X"00000000000000000000000f000000000000000f000000000000002300000000",
            INIT_30 => X"0000001b0000000000000009000000000000001e000000000000002300000000",
            INIT_31 => X"0000004c000000000000003a0000000000000023000000000000000e00000000",
            INIT_32 => X"0000004b000000000000000b000000000000001f000000000000003900000000",
            INIT_33 => X"0000002a00000000000000240000000000000001000000000000002400000000",
            INIT_34 => X"0000002300000000000000240000000000000009000000000000000300000000",
            INIT_35 => X"0000004200000000000000420000000000000042000000000000002d00000000",
            INIT_36 => X"0000004f000000000000004b0000000000000009000000000000000a00000000",
            INIT_37 => X"0000001000000000000000260000000000000020000000000000000d00000000",
            INIT_38 => X"00000023000000000000002b0000000000000029000000000000003300000000",
            INIT_39 => X"00000000000000000000004d000000000000003b000000000000003000000000",
            INIT_3A => X"00000041000000000000004d0000000000000031000000000000000700000000",
            INIT_3B => X"0000001d0000000000000017000000000000001e000000000000002000000000",
            INIT_3C => X"0000002400000000000000230000000000000024000000000000002000000000",
            INIT_3D => X"0000001c000000000000000a0000000000000042000000000000003500000000",
            INIT_3E => X"0000002d0000000000000042000000000000003b000000000000003800000000",
            INIT_3F => X"0000002400000000000000210000000000000029000000000000000200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002000000000000000400000000000000018000000000000001800000000",
            INIT_41 => X"0000002f00000000000000290000000000000009000000000000004000000000",
            INIT_42 => X"0000002500000000000000410000000000000042000000000000003b00000000",
            INIT_43 => X"000000300000000000000028000000000000002e000000000000002500000000",
            INIT_44 => X"000000330000000000000030000000000000002f000000000000002900000000",
            INIT_45 => X"0000002300000000000000380000000000000032000000000000001200000000",
            INIT_46 => X"00000035000000000000003e0000000000000038000000000000003500000000",
            INIT_47 => X"0000002a00000000000000330000000000000035000000000000003500000000",
            INIT_48 => X"0000002b0000000000000012000000000000001a000000000000002800000000",
            INIT_49 => X"0000003400000000000000170000000000000030000000000000002300000000",
            INIT_4A => X"0000004200000000000000470000000000000028000000000000002500000000",
            INIT_4B => X"0000002800000000000000310000000000000032000000000000003a00000000",
            INIT_4C => X"0000002c000000000000003c000000000000002a000000000000001e00000000",
            INIT_4D => X"00000036000000000000002d000000000000001a000000000000002d00000000",
            INIT_4E => X"0000004100000000000000420000000000000040000000000000003400000000",
            INIT_4F => X"0000001e0000000000000024000000000000002e000000000000002900000000",
            INIT_50 => X"0000007300000000000000440000000000000046000000000000003600000000",
            INIT_51 => X"0000003f000000000000002b000000000000002c000000000000004b00000000",
            INIT_52 => X"00000038000000000000004a000000000000002a000000000000004100000000",
            INIT_53 => X"0000002c000000000000000e0000000000000022000000000000003600000000",
            INIT_54 => X"0000006c00000000000000220000000000000011000000000000003b00000000",
            INIT_55 => X"000000330000000000000031000000000000002d000000000000005300000000",
            INIT_56 => X"000000370000000000000039000000000000001f000000000000002100000000",
            INIT_57 => X"000000410000000000000021000000000000000c000000000000001e00000000",
            INIT_58 => X"0000006800000000000000210000000000000000000000000000000f00000000",
            INIT_59 => X"00000036000000000000002e0000000000000039000000000000005b00000000",
            INIT_5A => X"0000002e00000000000000370000000000000035000000000000002300000000",
            INIT_5B => X"0000000000000000000000410000000000000018000000000000000300000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "samplegold_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000001100000000000000190000000000000000000000000000001600000000",
            INIT_15 => X"0000001000000000000000180000000000000012000000000000001400000000",
            INIT_16 => X"0000000000000000000000000000000000000003000000000000001500000000",
            INIT_17 => X"00000029000000000000000f0000000000000000000000000000000000000000",
            INIT_18 => X"000000160000000000000016000000000000001d000000000000002700000000",
            INIT_19 => X"00000009000000000000000e0000000000000011000000000000000f00000000",
            INIT_1A => X"0000000a00000000000000110000000000000000000000000000000000000000",
            INIT_1B => X"00000017000000000000002d000000000000000a000000000000000c00000000",
            INIT_1C => X"00000024000000000000001f0000000000000024000000000000001900000000",
            INIT_1D => X"00000000000000000000001a0000000000000018000000000000001500000000",
            INIT_1E => X"00000019000000000000000e0000000000000000000000000000000000000000",
            INIT_1F => X"00000028000000000000001e000000000000003f000000000000000700000000",
            INIT_20 => X"0000002f0000000000000030000000000000002e000000000000002500000000",
            INIT_21 => X"0000001800000000000000270000000000000025000000000000002300000000",
            INIT_22 => X"000000100000000000000000000000000000000a000000000000000f00000000",
            INIT_23 => X"000000260000000000000022000000000000001a000000000000003b00000000",
            INIT_24 => X"00000000000000000000001c0000000000000028000000000000002500000000",
            INIT_25 => X"00000024000000000000002e0000000000000028000000000000001700000000",
            INIT_26 => X"0000001900000000000000100000000000000014000000000000000400000000",
            INIT_27 => X"000000360000000000000027000000000000000c000000000000001f00000000",
            INIT_28 => X"0000003c0000000000000052000000000000001e000000000000001600000000",
            INIT_29 => X"00000000000000000000002a0000000000000026000000000000000b00000000",
            INIT_2A => X"000000460000000000000000000000000000000a000000000000000800000000",
            INIT_2B => X"00000034000000000000001a000000000000002f000000000000003d00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000005c00000000",
            INIT_2D => X"000000000000000000000000000000000000000b000000000000002600000000",
            INIT_2E => X"000000430000000000000016000000000000000e000000000000000700000000",
            INIT_2F => X"0000002a00000000000000370000000000000025000000000000004400000000",
            INIT_30 => X"0000001900000000000000380000000000000046000000000000003b00000000",
            INIT_31 => X"0000000200000000000000000000000000000000000000000000001100000000",
            INIT_32 => X"0000004500000000000000320000000000000012000000000000001a00000000",
            INIT_33 => X"0000006c000000000000004d000000000000005b000000000000003a00000000",
            INIT_34 => X"0000000d0000000000000077000000000000007c000000000000006800000000",
            INIT_35 => X"0000002500000000000000110000000000000005000000000000000000000000",
            INIT_36 => X"00000049000000000000003c0000000000000041000000000000001f00000000",
            INIT_37 => X"0000001a0000000000000000000000000000005b000000000000004500000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_39 => X"0000003b000000000000002b000000000000000b000000000000000600000000",
            INIT_3A => X"0000004000000000000000000000000000000045000000000000005500000000",
            INIT_3B => X"0000000b000000000000005d000000000000003f000000000000003c00000000",
            INIT_3C => X"0000002c00000000000000000000000000000000000000000000000800000000",
            INIT_3D => X"0000003c000000000000001f0000000000000045000000000000003900000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000041000000000000002a0000000000000000000000000000000000000000",
            INIT_41 => X"0000004e00000000000000290000000000000034000000000000002100000000",
            INIT_42 => X"00000001000000000000000a000000000000001f000000000000001a00000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"00000027000000000000000b0000000000000000000000000000000000000000",
            INIT_45 => X"00000038000000000000002b0000000000000040000000000000003a00000000",
            INIT_46 => X"0000000400000000000000270000000000000019000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000a00000000000000220000000000000014000000000000000000000000",
            INIT_49 => X"0000001400000000000000110000000000000017000000000000002b00000000",
            INIT_4A => X"0000001e00000000000000250000000000000036000000000000002a00000000",
            INIT_4B => X"0000001000000000000000170000000000000015000000000000000e00000000",
            INIT_4C => X"0000005f0000000000000068000000000000004a000000000000000200000000",
            INIT_4D => X"0000005b00000000000000630000000000000060000000000000006100000000",
            INIT_4E => X"0000003b0000000000000041000000000000003f000000000000005a00000000",
            INIT_4F => X"000000340000000000000046000000000000003e000000000000003800000000",
            INIT_50 => X"0000006400000000000000620000000000000059000000000000005c00000000",
            INIT_51 => X"000000650000000000000069000000000000006b000000000000006600000000",
            INIT_52 => X"00000042000000000000003d0000000000000044000000000000004d00000000",
            INIT_53 => X"000000470000000000000043000000000000003f000000000000004500000000",
            INIT_54 => X"0000006a00000000000000680000000000000065000000000000005800000000",
            INIT_55 => X"0000006300000000000000760000000000000066000000000000006800000000",
            INIT_56 => X"00000049000000000000004a0000000000000055000000000000004800000000",
            INIT_57 => X"0000005900000000000000480000000000000045000000000000004700000000",
            INIT_58 => X"0000006b000000000000006a000000000000006a000000000000006000000000",
            INIT_59 => X"0000006000000000000000660000000000000068000000000000006900000000",
            INIT_5A => X"0000004b00000000000000400000000000000049000000000000006000000000",
            INIT_5B => X"0000006200000000000000590000000000000043000000000000004700000000",
            INIT_5C => X"000000530000000000000068000000000000006b000000000000006800000000",
            INIT_5D => X"0000006100000000000000630000000000000051000000000000005500000000",
            INIT_5E => X"0000004300000000000000450000000000000047000000000000003800000000",
            INIT_5F => X"000000620000000000000064000000000000004d000000000000005e00000000",
            INIT_60 => X"0000004500000000000000330000000000000064000000000000006000000000",
            INIT_61 => X"0000002b00000000000000420000000000000052000000000000003800000000",
            INIT_62 => X"0000006800000000000000460000000000000042000000000000003f00000000",
            INIT_63 => X"0000005c000000000000004b0000000000000050000000000000005900000000",
            INIT_64 => X"000000460000000000000034000000000000003d000000000000004e00000000",
            INIT_65 => X"000000380000000000000025000000000000002a000000000000004900000000",
            INIT_66 => X"0000006400000000000000420000000000000042000000000000004100000000",
            INIT_67 => X"0000004b00000000000000560000000000000051000000000000004600000000",
            INIT_68 => X"00000037000000000000003e0000000000000050000000000000005900000000",
            INIT_69 => X"00000043000000000000003b0000000000000028000000000000002700000000",
            INIT_6A => X"000000490000000000000060000000000000004c000000000000003900000000",
            INIT_6B => X"0000003f000000000000004f0000000000000040000000000000004500000000",
            INIT_6C => X"00000015000000000000003a0000000000000042000000000000004c00000000",
            INIT_6D => X"0000001b000000000000004d0000000000000048000000000000002300000000",
            INIT_6E => X"0000000d000000000000003e0000000000000063000000000000004200000000",
            INIT_6F => X"000000530000000000000030000000000000004d000000000000005000000000",
            INIT_70 => X"0000002e000000000000002d000000000000002d000000000000003c00000000",
            INIT_71 => X"000000480000000000000007000000000000005a000000000000004a00000000",
            INIT_72 => X"0000003800000000000000040000000000000039000000000000005a00000000",
            INIT_73 => X"0000002b0000000000000050000000000000002c000000000000003000000000",
            INIT_74 => X"00000049000000000000002f000000000000002d000000000000002f00000000",
            INIT_75 => X"0000004f000000000000004a000000000000000e000000000000005b00000000",
            INIT_76 => X"000000460000000000000043000000000000003e000000000000004100000000",
            INIT_77 => X"000000230000000000000024000000000000002f000000000000005100000000",
            INIT_78 => X"0000004d000000000000003d000000000000002e000000000000001f00000000",
            INIT_79 => X"0000004d000000000000004e0000000000000058000000000000003300000000",
            INIT_7A => X"0000004a00000000000000440000000000000050000000000000004f00000000",
            INIT_7B => X"00000024000000000000002c0000000000000035000000000000003d00000000",
            INIT_7C => X"000000490000000000000036000000000000003b000000000000002d00000000",
            INIT_7D => X"0000004d00000000000000430000000000000053000000000000004800000000",
            INIT_7E => X"0000003f00000000000000550000000000000049000000000000003000000000",
            INIT_7F => X"0000004b0000000000000042000000000000003e000000000000004800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "samplegold_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004a0000000000000036000000000000004f000000000000004600000000",
            INIT_01 => X"0000004d0000000000000055000000000000004a000000000000005600000000",
            INIT_02 => X"0000004c000000000000004c0000000000000057000000000000005000000000",
            INIT_03 => X"0000004f00000000000000560000000000000054000000000000004d00000000",
            INIT_04 => X"0000000000000000000000000000000000000052000000000000004700000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000002f000000000000002e000000000000002c000000000000002100000000",
            INIT_3E => X"0000002200000000000000240000000000000020000000000000002100000000",
            INIT_3F => X"0000001500000000000000130000000000000018000000000000000c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004900000000000000520000000000000023000000000000001d00000000",
            INIT_41 => X"0000002d00000000000000330000000000000037000000000000003300000000",
            INIT_42 => X"0000000000000000000000180000000000000021000000000000001f00000000",
            INIT_43 => X"00000025000000000000002c000000000000001b000000000000001300000000",
            INIT_44 => X"0000003a000000000000004c0000000000000047000000000000001e00000000",
            INIT_45 => X"0000002d0000000000000036000000000000003f000000000000003c00000000",
            INIT_46 => X"0000001d000000000000002b0000000000000032000000000000001c00000000",
            INIT_47 => X"000000250000000000000025000000000000001d000000000000001800000000",
            INIT_48 => X"0000004400000000000000430000000000000048000000000000005d00000000",
            INIT_49 => X"0000002b00000000000000380000000000000040000000000000004700000000",
            INIT_4A => X"00000017000000000000002d000000000000003f000000000000002f00000000",
            INIT_4B => X"0000004400000000000000270000000000000017000000000000001400000000",
            INIT_4C => X"000000440000000000000046000000000000004a000000000000004e00000000",
            INIT_4D => X"0000002500000000000000470000000000000043000000000000003e00000000",
            INIT_4E => X"000000190000000000000028000000000000003f000000000000003200000000",
            INIT_4F => X"0000004e00000000000000390000000000000028000000000000002000000000",
            INIT_50 => X"0000006a000000000000003e000000000000004d000000000000004d00000000",
            INIT_51 => X"00000038000000000000004d0000000000000054000000000000006900000000",
            INIT_52 => X"00000015000000000000000a000000000000001c000000000000003400000000",
            INIT_53 => X"00000073000000000000006f0000000000000014000000000000002100000000",
            INIT_54 => X"0000007900000000000000730000000000000059000000000000006500000000",
            INIT_55 => X"0000003e0000000000000059000000000000004d000000000000006300000000",
            INIT_56 => X"0000001700000000000000120000000000000006000000000000001200000000",
            INIT_57 => X"0000006400000000000000760000000000000051000000000000002c00000000",
            INIT_58 => X"0000008e00000000000000620000000000000083000000000000008300000000",
            INIT_59 => X"000000180000000000000052000000000000008d000000000000009100000000",
            INIT_5A => X"00000039000000000000000e0000000000000031000000000000001400000000",
            INIT_5B => X"00000086000000000000004e000000000000007b000000000000005f00000000",
            INIT_5C => X"0000006d00000000000000630000000000000060000000000000008000000000",
            INIT_5D => X"000000070000000000000005000000000000003a000000000000005700000000",
            INIT_5E => X"00000059000000000000003b000000000000002e000000000000005100000000",
            INIT_5F => X"0000006e00000000000000470000000000000040000000000000009500000000",
            INIT_60 => X"00000013000000000000002e000000000000005b000000000000005c00000000",
            INIT_61 => X"0000006500000000000000090000000000000000000000000000000500000000",
            INIT_62 => X"00000083000000000000005a0000000000000046000000000000005300000000",
            INIT_63 => X"0000002100000000000000120000000000000000000000000000003a00000000",
            INIT_64 => X"0000000000000000000000000000000000000022000000000000002d00000000",
            INIT_65 => X"0000007a00000000000000550000000000000007000000000000000a00000000",
            INIT_66 => X"0000004e0000000000000064000000000000004e000000000000004900000000",
            INIT_67 => X"00000011000000000000001a000000000000001e000000000000001a00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000003c0000000000000070000000000000001b000000000000000c00000000",
            INIT_6A => X"0000003a000000000000005e000000000000004b000000000000005200000000",
            INIT_6B => X"0000001100000000000000240000000000000038000000000000003200000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"00000049000000000000003c0000000000000025000000000000000b00000000",
            INIT_6E => X"00000035000000000000003f000000000000003d000000000000004e00000000",
            INIT_6F => X"00000027000000000000002e000000000000003f000000000000003e00000000",
            INIT_70 => X"00000018000000000000001e0000000000000023000000000000002200000000",
            INIT_71 => X"0000004800000000000000420000000000000046000000000000002900000000",
            INIT_72 => X"0000003800000000000000420000000000000046000000000000004300000000",
            INIT_73 => X"0000002e000000000000002d0000000000000031000000000000003900000000",
            INIT_74 => X"00000028000000000000002b0000000000000038000000000000003a00000000",
            INIT_75 => X"00000032000000000000003e000000000000000d000000000000004400000000",
            INIT_76 => X"000000330000000000000041000000000000003d000000000000004100000000",
            INIT_77 => X"000000230000000000000024000000000000002e000000000000004600000000",
            INIT_78 => X"00000047000000000000002e0000000000000015000000000000001b00000000",
            INIT_79 => X"0000003d000000000000003c0000000000000042000000000000005900000000",
            INIT_7A => X"000000450000000000000035000000000000003d000000000000003900000000",
            INIT_7B => X"0000001d00000000000000250000000000000024000000000000002e00000000",
            INIT_7C => X"0000004700000000000000560000000000000025000000000000002a00000000",
            INIT_7D => X"0000004900000000000000430000000000000047000000000000004000000000",
            INIT_7E => X"000000220000000000000040000000000000003d000000000000004400000000",
            INIT_7F => X"0000002e0000000000000023000000000000001d000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "samplegold_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004c0000000000000042000000000000005c000000000000002100000000",
            INIT_01 => X"00000049000000000000004e000000000000004b000000000000004300000000",
            INIT_02 => X"0000003b00000000000000410000000000000040000000000000004800000000",
            INIT_03 => X"00000026000000000000001c000000000000002f000000000000004100000000",
            INIT_04 => X"0000004c0000000000000045000000000000003a000000000000004e00000000",
            INIT_05 => X"00000026000000000000003d000000000000004f000000000000004900000000",
            INIT_06 => X"0000005f0000000000000041000000000000003b000000000000003b00000000",
            INIT_07 => X"00000029000000000000002b0000000000000030000000000000002a00000000",
            INIT_08 => X"0000005e00000000000000490000000000000032000000000000004100000000",
            INIT_09 => X"0000006300000000000000500000000000000035000000000000003600000000",
            INIT_0A => X"00000024000000000000005b000000000000003e000000000000002700000000",
            INIT_0B => X"0000004a00000000000000000000000000000027000000000000002f00000000",
            INIT_0C => X"000000430000000000000033000000000000004e000000000000004c00000000",
            INIT_0D => X"0000001300000000000000000000000000000025000000000000006600000000",
            INIT_0E => X"00000025000000000000001b0000000000000036000000000000004500000000",
            INIT_0F => X"0000004e0000000000000012000000000000002b000000000000002900000000",
            INIT_10 => X"0000003700000000000000400000000000000031000000000000004c00000000",
            INIT_11 => X"00000040000000000000003f0000000000000040000000000000003800000000",
            INIT_12 => X"00000029000000000000000c0000000000000020000000000000003b00000000",
            INIT_13 => X"000000540000000000000039000000000000000e000000000000002400000000",
            INIT_14 => X"0000007200000000000000560000000000000057000000000000005900000000",
            INIT_15 => X"000000460000000000000096000000000000007e000000000000006d00000000",
            INIT_16 => X"000000340000000000000049000000000000001b000000000000000b00000000",
            INIT_17 => X"000000410000000000000074000000000000003d000000000000001300000000",
            INIT_18 => X"0000003600000000000000010000000000000066000000000000004700000000",
            INIT_19 => X"0000000b000000000000000d0000000000000013000000000000004400000000",
            INIT_1A => X"00000029000000000000002f000000000000004c000000000000000e00000000",
            INIT_1B => X"0000005c00000000000000110000000000000077000000000000005800000000",
            INIT_1C => X"0000004000000000000000790000000000000047000000000000005700000000",
            INIT_1D => X"0000001c000000000000000b000000000000002a000000000000003b00000000",
            INIT_1E => X"00000043000000000000001e000000000000003c000000000000006400000000",
            INIT_1F => X"000000000000000000000000000000000000001b000000000000001b00000000",
            INIT_20 => X"0000002500000000000000270000000000000036000000000000003600000000",
            INIT_21 => X"0000005200000000000000300000000000000023000000000000002700000000",
            INIT_22 => X"0000004b0000000000000032000000000000002f000000000000002100000000",
            INIT_23 => X"0000001a00000000000000150000000000000039000000000000003900000000",
            INIT_24 => X"0000000200000000000000080000000000000008000000000000000f00000000",
            INIT_25 => X"000000300000000000000028000000000000002a000000000000000c00000000",
            INIT_26 => X"0000004d0000000000000035000000000000003f000000000000002800000000",
            INIT_27 => X"0000001700000000000000320000000000000017000000000000001a00000000",
            INIT_28 => X"000000080000000000000000000000000000000a000000000000000c00000000",
            INIT_29 => X"0000000a00000000000000250000000000000030000000000000000700000000",
            INIT_2A => X"0000001a000000000000001c0000000000000014000000000000002900000000",
            INIT_2B => X"000000280000000000000032000000000000003a000000000000003300000000",
            INIT_2C => X"0000002d00000000000000230000000000000020000000000000001d00000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000800000000000000050000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000060000000000000005000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_41 => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001300000000000000000000000000000000000000000000001b00000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_45 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000010000000000000014000000000000000000000000",
            INIT_4D => X"0000006300000000000000470000000000000035000000000000003400000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000210000000000000005000000000000007700000000",
            INIT_51 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000001f000000000000000a000000000000000000000000",
            INIT_54 => X"00000046000000000000002d000000000000003d000000000000003e00000000",
            INIT_55 => X"00000000000000000000001e000000000000001e000000000000000400000000",
            INIT_56 => X"00000000000000000000000b0000000000000007000000000000001100000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_58 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000b0000000000000013000000000000000d000000000000000c00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000050000000000000009000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_67 => X"000000020000000000000000000000000000000a000000000000000000000000",
            INIT_68 => X"0000001900000000000000010000000000000000000000000000000400000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000011000000000000000400000000",
            INIT_6D => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000010000000000000001000000000000000100000000",
            INIT_71 => X"00000000000000000000000b0000000000000000000000000000000100000000",
            INIT_72 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000d00000000000000000000000000000003000000000000001100000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"00000002000000000000001a0000000000000000000000000000000300000000",
            INIT_78 => X"00000008000000000000000000000000000000a0000000000000000600000000",
            INIT_79 => X"00000000000000000000003a0000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_7B => X"000000120000000000000004000000000000001e000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000047000000000000008100000000",
            INIT_7D => X"0000000000000000000000000000000000000009000000000000001100000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_7F => X"000000000000000000000003000000000000000c000000000000000f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "samplegold_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003300000000000000000000000000000000000000000000008600000000",
            INIT_01 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_02 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000006900000000000000000000000000000000000000000000002300000000",
            INIT_04 => X"0000002000000000000000340000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000000d0000000000000009000000000000000000000000",
            INIT_06 => X"0000005400000000000000550000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000700000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000002f0000000000000082000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_0A => X"0000000000000000000000850000000000000047000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000049000000000000000000000000",
            INIT_0C => X"0000003600000000000000060000000000000011000000000000002b00000000",
            INIT_0D => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000096000000000000002300000000",
            INIT_0F => X"0000000000000000000000000000000000000007000000000000001000000000",
            INIT_10 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_11 => X"00000044000000000000001e0000000000000000000000000000000000000000",
            INIT_12 => X"00000000000000000000000a000000000000000f000000000000003800000000",
            INIT_13 => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_15 => X"0000000a00000000000000280000000000000009000000000000000000000000",
            INIT_16 => X"0000000000000000000000320000000000000000000000000000002d00000000",
            INIT_17 => X"0000001f00000000000000070000000000000000000000000000001600000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000000000000000000000b0000000000000000000000000000000900000000",
            INIT_1A => X"0000000300000000000000000000000000000012000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000900000000000000080000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000020000000000000015000000000000000400000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"000000000000000000000000000000000000000c000000000000001200000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_49 => X"000000020000000000000013000000000000000a000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000260000000000000027000000000000002200000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000030000000000000003000000000000000100000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "samplegold_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000000000000000000003b000000000000000c000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000000000000a0000000000000007000000000000000500000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000300000000000000000000000000000006000000000000000700000000",
            INIT_17 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000000000000000000002000000000000002a000000000000002200000000",
            INIT_19 => X"0000000500000000000000000000000000000003000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00000003000000000000000d0000000000000000000000000000000000000000",
            INIT_1E => X"0000000400000000000000000000000000000000000000000000000100000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000007000000000000001b000000000000000f000000000000000f00000000",
            INIT_22 => X"0000000000000000000000210000000000000038000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_24 => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000002600000000000000080000000000000004000000000000000100000000",
            INIT_26 => X"0000005a000000000000003a0000000000000000000000000000001800000000",
            INIT_27 => X"0000000600000000000000000000000000000000000000000000003600000000",
            INIT_28 => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000001b00000000000000350000000000000000000000000000000100000000",
            INIT_2A => X"0000001e0000000000000015000000000000001e000000000000001800000000",
            INIT_2B => X"0000003000000000000000060000000000000000000000000000000600000000",
            INIT_2C => X"00000018000000000000002f0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000220000000000000015000000000000000000000000",
            INIT_30 => X"0000000000000000000000190000000000000027000000000000000000000000",
            INIT_31 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000a00000000000000090000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000003a000000000000000e00000000",
            INIT_34 => X"0000001300000000000000000000000000000000000000000000000400000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000700000000000000000000000000000000000000000000001a00000000",
            INIT_38 => X"0000002c000000000000000d000000000000002c000000000000000600000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000700000000000000000000000000000001000000000000000000000000",
            INIT_3D => X"0000001c00000000000000220000000000000018000000000000000b00000000",
            INIT_3E => X"0000000000000000000000000000000000000010000000000000002300000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000020000000000000008000000000000000000000000",
            INIT_41 => X"0000002f00000000000000190000000000000014000000000000000e00000000",
            INIT_42 => X"000000000000000000000000000000000000001c000000000000002300000000",
            INIT_43 => X"00000012000000000000000b0000000000000000000000000000001500000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_45 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_46 => X"0000005e000000000000005e0000000000000011000000000000000000000000",
            INIT_47 => X"000000650000000000000064000000000000005d000000000000006000000000",
            INIT_48 => X"00000023000000000000003c000000000000004f000000000000005800000000",
            INIT_49 => X"0000002c00000000000000270000000000000029000000000000002400000000",
            INIT_4A => X"000000650000000000000068000000000000005f000000000000002500000000",
            INIT_4B => X"0000006e000000000000006e000000000000006c000000000000006900000000",
            INIT_4C => X"0000001f000000000000002c0000000000000054000000000000006300000000",
            INIT_4D => X"0000002d0000000000000037000000000000002f000000000000002a00000000",
            INIT_4E => X"0000006f000000000000006c0000000000000059000000000000006400000000",
            INIT_4F => X"0000007000000000000000720000000000000076000000000000007100000000",
            INIT_50 => X"0000003e00000000000000410000000000000048000000000000006500000000",
            INIT_51 => X"0000005400000000000000340000000000000033000000000000003900000000",
            INIT_52 => X"00000075000000000000006d000000000000006a000000000000006300000000",
            INIT_53 => X"0000006400000000000000670000000000000074000000000000007800000000",
            INIT_54 => X"00000031000000000000004e0000000000000066000000000000006500000000",
            INIT_55 => X"0000005a00000000000000480000000000000037000000000000003400000000",
            INIT_56 => X"0000007000000000000000760000000000000072000000000000006c00000000",
            INIT_57 => X"000000570000000000000060000000000000005a000000000000005a00000000",
            INIT_58 => X"0000003200000000000000270000000000000048000000000000005900000000",
            INIT_59 => X"0000006c0000000000000069000000000000001e000000000000003300000000",
            INIT_5A => X"0000005500000000000000560000000000000075000000000000007200000000",
            INIT_5B => X"0000004b0000000000000043000000000000003a000000000000004200000000",
            INIT_5C => X"00000030000000000000002b0000000000000021000000000000002e00000000",
            INIT_5D => X"0000006000000000000000690000000000000049000000000000003400000000",
            INIT_5E => X"0000004000000000000000520000000000000068000000000000005b00000000",
            INIT_5F => X"0000001b0000000000000041000000000000004d000000000000004600000000",
            INIT_60 => X"00000042000000000000002e000000000000002a000000000000001800000000",
            INIT_61 => X"00000058000000000000005a000000000000005f000000000000004000000000",
            INIT_62 => X"0000005400000000000000560000000000000071000000000000006a00000000",
            INIT_63 => X"00000011000000000000001a0000000000000046000000000000004f00000000",
            INIT_64 => X"00000045000000000000004a000000000000003b000000000000002f00000000",
            INIT_65 => X"0000005300000000000000460000000000000058000000000000005d00000000",
            INIT_66 => X"000000420000000000000040000000000000004f000000000000006500000000",
            INIT_67 => X"0000003300000000000000100000000000000005000000000000002400000000",
            INIT_68 => X"0000004d00000000000000460000000000000051000000000000003300000000",
            INIT_69 => X"0000004e000000000000004c0000000000000019000000000000004700000000",
            INIT_6A => X"0000000f0000000000000019000000000000005e000000000000003f00000000",
            INIT_6B => X"0000003c00000000000000350000000000000016000000000000001500000000",
            INIT_6C => X"0000003600000000000000490000000000000047000000000000005400000000",
            INIT_6D => X"0000003b00000000000000180000000000000018000000000000001800000000",
            INIT_6E => X"0000000900000000000000050000000000000011000000000000002700000000",
            INIT_6F => X"0000004d000000000000003a0000000000000034000000000000002000000000",
            INIT_70 => X"0000004a000000000000004c0000000000000040000000000000004d00000000",
            INIT_71 => X"0000000800000000000000310000000000000039000000000000002b00000000",
            INIT_72 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"000000540000000000000051000000000000002a000000000000003300000000",
            INIT_74 => X"0000004000000000000000510000000000000046000000000000005200000000",
            INIT_75 => X"0000001100000000000000220000000000000040000000000000003c00000000",
            INIT_76 => X"0000001600000000000000170000000000000001000000000000000700000000",
            INIT_77 => X"000000500000000000000041000000000000004a000000000000003200000000",
            INIT_78 => X"0000004b00000000000000410000000000000039000000000000004400000000",
            INIT_79 => X"0000003100000000000000340000000000000039000000000000004c00000000",
            INIT_7A => X"0000002e00000000000000390000000000000039000000000000003600000000",
            INIT_7B => X"0000004f000000000000004e0000000000000051000000000000004700000000",
            INIT_7C => X"0000004900000000000000540000000000000058000000000000004b00000000",
            INIT_7D => X"0000004f00000000000000490000000000000043000000000000004800000000",
            INIT_7E => X"00000000000000000000003a000000000000004a000000000000004f00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "samplegold_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000006000000000000000a00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_0D => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_11 => X"00000000000000000000001f0000000000000000000000000000000600000000",
            INIT_12 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000030000000000000038000000000000000000000000",
            INIT_14 => X"0000000000000000000000110000000000000009000000000000000100000000",
            INIT_15 => X"00000000000000000000000c0000000000000016000000000000000400000000",
            INIT_16 => X"0000000400000000000000050000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000700000000000000000000000000000001000000000000000000000000",
            INIT_19 => X"0000000800000000000000000000000000000016000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_1D => X"0000002300000000000000010000000000000000000000000000000000000000",
            INIT_1E => X"0000003c000000000000004b0000000000000003000000000000001e00000000",
            INIT_1F => X"0000000a000000000000000e000000000000005a000000000000006300000000",
            INIT_20 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000001b000000000000007d0000000000000000000000000000000000000000",
            INIT_22 => X"0000001100000000000000000000000000000000000000000000000b00000000",
            INIT_23 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_24 => X"0000001e00000000000000160000000000000000000000000000000000000000",
            INIT_25 => X"0000004700000000000000760000000000000006000000000000000000000000",
            INIT_26 => X"000000290000000000000007000000000000002d000000000000005c00000000",
            INIT_27 => X"0000000000000000000000360000000000000000000000000000000900000000",
            INIT_28 => X"00000000000000000000000a0000000000000000000000000000000600000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000000290000000000000004000000000000000a000000000000000700000000",
            INIT_2B => X"00000000000000000000000c0000000000000041000000000000001800000000",
            INIT_2C => X"00000000000000000000002b0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000180000000000000000000000000000002a000000000000000200000000",
            INIT_30 => X"00000000000000000000000b0000000000000007000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000003000000000000000f0000000000000006000000000000002000000000",
            INIT_38 => X"000000020000000000000012000000000000000e000000000000000b00000000",
            INIT_39 => X"0000001200000000000000000000000000000008000000000000002f00000000",
            INIT_3A => X"0000001300000000000000220000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000000000001000000000000000c000000000000001900000000",
            INIT_3C => X"0000002c0000000000000008000000000000001e000000000000000900000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_3E => X"0000000000000000000000340000000000000000000000000000001700000000",
            INIT_3F => X"0000000e00000000000000000000000000000001000000000000000d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003200000000000000050000000000000000000000000000001a00000000",
            INIT_41 => X"0000000000000000000000080000000000000026000000000000000000000000",
            INIT_42 => X"000000070000000000000000000000000000001d000000000000000800000000",
            INIT_43 => X"000000140000000000000012000000000000000c000000000000000000000000",
            INIT_44 => X"0000001300000000000000000000000000000000000000000000001900000000",
            INIT_45 => X"0000000100000000000000000000000000000006000000000000004000000000",
            INIT_46 => X"0000000500000000000000060000000000000000000000000000000300000000",
            INIT_47 => X"0000000000000000000000090000000000000014000000000000000200000000",
            INIT_48 => X"0000005a00000000000000070000000000000000000000000000003600000000",
            INIT_49 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_4A => X"00000015000000000000000c0000000000000000000000000000001000000000",
            INIT_4B => X"00000023000000000000000f000000000000003f000000000000000000000000",
            INIT_4C => X"00000000000000000000003b0000000000000027000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_4E => X"0000000a00000000000000000000000000000015000000000000000d00000000",
            INIT_4F => X"0000000100000000000000000000000000000016000000000000001400000000",
            INIT_50 => X"0000000000000000000000000000000000000033000000000000004c00000000",
            INIT_51 => X"0000001800000000000000000000000000000025000000000000000400000000",
            INIT_52 => X"0000002500000000000000080000000000000000000000000000000000000000",
            INIT_53 => X"0000006400000000000000000000000000000001000000000000000000000000",
            INIT_54 => X"0000004200000000000000000000000000000000000000000000004100000000",
            INIT_55 => X"0000004a00000000000000060000000000000000000000000000001800000000",
            INIT_56 => X"0000000300000000000000580000000000000000000000000000000000000000",
            INIT_57 => X"0000001500000000000000480000000000000027000000000000000300000000",
            INIT_58 => X"0000002200000000000000830000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000c00000000000000000000000000000000000000000",
            INIT_5A => X"0000006400000000000000000000000000000042000000000000000000000000",
            INIT_5B => X"00000000000000000000001a0000000000000006000000000000001c00000000",
            INIT_5C => X"00000000000000000000002b000000000000008d000000000000000000000000",
            INIT_5D => X"00000000000000000000000b0000000000000072000000000000000a00000000",
            INIT_5E => X"0000002b00000000000000340000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_60 => X"000000000000000000000009000000000000000c000000000000004e00000000",
            INIT_61 => X"0000000a0000000000000000000000000000002a000000000000002700000000",
            INIT_62 => X"0000000a00000000000000030000000000000025000000000000003300000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000200000000000000000000000000000000c00000000",
            INIT_65 => X"0000002c00000000000000000000000000000026000000000000004b00000000",
            INIT_66 => X"0000000000000000000000160000000000000014000000000000002700000000",
            INIT_67 => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000001b00000000000000170000000000000027000000000000000000000000",
            INIT_69 => X"00000000000000000000002f0000000000000000000000000000000000000000",
            INIT_6A => X"0000001100000000000000000000000000000007000000000000001900000000",
            INIT_6B => X"0000000600000000000000000000000000000000000000000000000b00000000",
            INIT_6C => X"0000000800000000000000100000000000000001000000000000001100000000",
            INIT_6D => X"0000000d00000000000000150000000000000007000000000000001500000000",
            INIT_6E => X"0000001e00000000000000130000000000000000000000000000000000000000",
            INIT_6F => X"00000079000000000000006e0000000000000070000000000000000000000000",
            INIT_70 => X"0000007c00000000000000800000000000000083000000000000008100000000",
            INIT_71 => X"0000005100000000000000430000000000000059000000000000006c00000000",
            INIT_72 => X"0000005200000000000000550000000000000051000000000000005000000000",
            INIT_73 => X"0000008200000000000000790000000000000071000000000000006c00000000",
            INIT_74 => X"0000008b000000000000008d000000000000008b000000000000008600000000",
            INIT_75 => X"0000005700000000000000490000000000000042000000000000007700000000",
            INIT_76 => X"0000006100000000000000580000000000000063000000000000006400000000",
            INIT_77 => X"000000840000000000000081000000000000007b000000000000006800000000",
            INIT_78 => X"000000870000000000000086000000000000008e000000000000008800000000",
            INIT_79 => X"00000069000000000000006a000000000000006f000000000000007000000000",
            INIT_7A => X"00000068000000000000005b0000000000000061000000000000006200000000",
            INIT_7B => X"000000910000000000000083000000000000007f000000000000007700000000",
            INIT_7C => X"00000087000000000000007d0000000000000081000000000000008f00000000",
            INIT_7D => X"00000061000000000000005f0000000000000069000000000000007e00000000",
            INIT_7E => X"0000007c000000000000006c0000000000000051000000000000006200000000",
            INIT_7F => X"00000072000000000000007f0000000000000086000000000000007d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "samplegold_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000074000000000000007c0000000000000071000000000000007900000000",
            INIT_01 => X"0000005e00000000000000590000000000000050000000000000005900000000",
            INIT_02 => X"00000078000000000000007a0000000000000072000000000000004100000000",
            INIT_03 => X"0000004b0000000000000055000000000000005b000000000000007500000000",
            INIT_04 => X"0000004300000000000000630000000000000062000000000000005800000000",
            INIT_05 => X"00000049000000000000005b0000000000000051000000000000004200000000",
            INIT_06 => X"00000064000000000000006b000000000000006d000000000000005f00000000",
            INIT_07 => X"0000005e0000000000000064000000000000005f000000000000005c00000000",
            INIT_08 => X"0000003a000000000000003c0000000000000054000000000000005b00000000",
            INIT_09 => X"0000005c00000000000000680000000000000055000000000000005000000000",
            INIT_0A => X"0000006f000000000000005f000000000000005e000000000000006c00000000",
            INIT_0B => X"0000005b000000000000005a0000000000000066000000000000007b00000000",
            INIT_0C => X"0000005900000000000000340000000000000038000000000000005b00000000",
            INIT_0D => X"0000006b00000000000000680000000000000080000000000000005100000000",
            INIT_0E => X"00000072000000000000005a0000000000000052000000000000005500000000",
            INIT_0F => X"0000003700000000000000460000000000000056000000000000005d00000000",
            INIT_10 => X"0000004f00000000000000530000000000000033000000000000002d00000000",
            INIT_11 => X"00000052000000000000005a0000000000000061000000000000008300000000",
            INIT_12 => X"0000007d000000000000006b0000000000000056000000000000002b00000000",
            INIT_13 => X"00000047000000000000003d000000000000003a000000000000007400000000",
            INIT_14 => X"0000008500000000000000530000000000000053000000000000003f00000000",
            INIT_15 => X"0000003500000000000000510000000000000053000000000000006800000000",
            INIT_16 => X"0000004c00000000000000600000000000000043000000000000002200000000",
            INIT_17 => X"0000004a000000000000003c0000000000000025000000000000003100000000",
            INIT_18 => X"0000007d000000000000007e0000000000000053000000000000004800000000",
            INIT_19 => X"0000006e000000000000006a0000000000000073000000000000005500000000",
            INIT_1A => X"0000001800000000000000230000000000000059000000000000007100000000",
            INIT_1B => X"0000004600000000000000370000000000000016000000000000001600000000",
            INIT_1C => X"0000006a00000000000000840000000000000086000000000000005300000000",
            INIT_1D => X"0000007c000000000000006b0000000000000066000000000000005800000000",
            INIT_1E => X"00000030000000000000003c0000000000000053000000000000007400000000",
            INIT_1F => X"0000004a00000000000000400000000000000034000000000000002b00000000",
            INIT_20 => X"00000063000000000000007b0000000000000072000000000000007900000000",
            INIT_21 => X"00000085000000000000007c0000000000000071000000000000005a00000000",
            INIT_22 => X"0000006b00000000000000680000000000000067000000000000006c00000000",
            INIT_23 => X"0000008200000000000000590000000000000064000000000000006800000000",
            INIT_24 => X"0000007b00000000000000830000000000000087000000000000008800000000",
            INIT_25 => X"00000076000000000000007b0000000000000080000000000000008a00000000",
            INIT_26 => X"0000007d000000000000007f000000000000007e000000000000007900000000",
            INIT_27 => X"0000000000000000000000000000000000000068000000000000007500000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000005000000000000000b000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000000000000000000000000000000000000d000000000000000400000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000040000000000000003000000000000000e00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000b00000000000000120000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000003000000000000000500000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000070000000000000008000000000000001f000000000000000000000000",
            INIT_3B => X"00000011000000000000001f0000000000000003000000000000000700000000",
            INIT_3C => X"000000000000000000000006000000000000000c000000000000001a00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000013000000000000001b0000000000000029000000000000000300000000",
            INIT_3F => X"0000000700000000000000240000000000000026000000000000001000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000000000000000000000d000000000000000700000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000002d000000000000001c000000000000001c000000000000002400000000",
            INIT_43 => X"00000031000000000000002e000000000000000b000000000000002100000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_45 => X"0000002100000000000000000000000000000000000000000000000200000000",
            INIT_46 => X"0000002e00000000000000390000000000000009000000000000001e00000000",
            INIT_47 => X"00000024000000000000002a0000000000000024000000000000000900000000",
            INIT_48 => X"0000001d00000000000000000000000000000000000000000000000c00000000",
            INIT_49 => X"0000003100000000000000220000000000000000000000000000000000000000",
            INIT_4A => X"00000007000000000000002a0000000000000039000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_4C => X"00000000000000000000002d0000000000000000000000000000000000000000",
            INIT_4D => X"00000000000000000000002e000000000000001d000000000000000000000000",
            INIT_4E => X"0000000c00000000000000050000000000000009000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000100000000000000160000000000000032000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000022000000000000000500000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000080000000000000000000000000000002b000000000000000600000000",
            INIT_55 => X"0000000000000000000000000000000000000023000000000000000500000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"00000002000000000000000e0000000000000000000000000000000400000000",
            INIT_59 => X"0000000400000000000000000000000000000004000000000000000400000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"00000033000000000000002f0000000000000032000000000000001800000000",
            INIT_61 => X"0000000d00000000000000270000000000000031000000000000003700000000",
            INIT_62 => X"0000000d000000000000000d0000000000000010000000000000000f00000000",
            INIT_63 => X"00000024000000000000001b0000000000000007000000000000000f00000000",
            INIT_64 => X"0000003900000000000000350000000000000031000000000000003500000000",
            INIT_65 => X"0000000d0000000000000025000000000000003e000000000000003f00000000",
            INIT_66 => X"0000001600000000000000180000000000000015000000000000001100000000",
            INIT_67 => X"00000031000000000000001c0000000000000013000000000000001200000000",
            INIT_68 => X"0000003e000000000000003e0000000000000033000000000000003700000000",
            INIT_69 => X"0000001300000000000000120000000000000031000000000000004400000000",
            INIT_6A => X"00000018000000000000001d0000000000000020000000000000001e00000000",
            INIT_6B => X"00000031000000000000002e000000000000001c000000000000001300000000",
            INIT_6C => X"0000003b00000000000000400000000000000045000000000000003500000000",
            INIT_6D => X"0000002100000000000000310000000000000039000000000000003800000000",
            INIT_6E => X"00000018000000000000001a000000000000001d000000000000001e00000000",
            INIT_6F => X"0000003a0000000000000032000000000000002b000000000000001c00000000",
            INIT_70 => X"0000002b000000000000001c0000000000000028000000000000003200000000",
            INIT_71 => X"000000170000000000000010000000000000002b000000000000003a00000000",
            INIT_72 => X"000000220000000000000020000000000000001a000000000000001800000000",
            INIT_73 => X"0000000600000000000000310000000000000028000000000000002000000000",
            INIT_74 => X"0000001d00000000000000190000000000000001000000000000000000000000",
            INIT_75 => X"00000016000000000000000d000000000000000a000000000000001900000000",
            INIT_76 => X"00000011000000000000001e000000000000000a000000000000001a00000000",
            INIT_77 => X"0000000f00000000000000020000000000000014000000000000001500000000",
            INIT_78 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000001700000000000000110000000000000002000000000000000000000000",
            INIT_7A => X"00000011000000000000000f0000000000000014000000000000001700000000",
            INIT_7B => X"00000000000000000000001d000000000000000a000000000000000300000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"00000023000000000000000a0000000000000005000000000000000400000000",
            INIT_7E => X"00000000000000000000000e0000000000000006000000000000001300000000",
            INIT_7F => X"00000013000000000000001c0000000000000016000000000000001b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "samplegold_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000500000000000000000000000000000009000000000000001200000000",
            INIT_01 => X"00000011000000000000002a0000000000000000000000000000000600000000",
            INIT_02 => X"0000001100000000000000030000000000000000000000000000000000000000",
            INIT_03 => X"000000070000000000000017000000000000000f000000000000001c00000000",
            INIT_04 => X"00000000000000000000000c0000000000000000000000000000000100000000",
            INIT_05 => X"00000000000000000000001a0000000000000025000000000000000000000000",
            INIT_06 => X"00000022000000000000000a0000000000000001000000000000000000000000",
            INIT_07 => X"000000000000000000000007000000000000001b000000000000002d00000000",
            INIT_08 => X"000000000000000000000009000000000000000e000000000000000700000000",
            INIT_09 => X"000000050000000000000007000000000000001d000000000000003000000000",
            INIT_0A => X"0000000b0000000000000015000000000000000b000000000000001300000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000350000000000000000000000000000001a000000000000001000000000",
            INIT_0D => X"0000001600000000000000140000000000000017000000000000002700000000",
            INIT_0E => X"0000000000000000000000120000000000000026000000000000002600000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000002e00000000000000230000000000000007000000000000001400000000",
            INIT_11 => X"0000001d00000000000000120000000000000022000000000000001e00000000",
            INIT_12 => X"0000000c00000000000000140000000000000027000000000000002800000000",
            INIT_13 => X"00000011000000000000000b0000000000000009000000000000000e00000000",
            INIT_14 => X"0000002b00000000000000250000000000000027000000000000000900000000",
            INIT_15 => X"0000002f0000000000000028000000000000001f000000000000002400000000",
            INIT_16 => X"0000002b000000000000002c000000000000002b000000000000002c00000000",
            INIT_17 => X"0000001c00000000000000210000000000000026000000000000002a00000000",
            INIT_18 => X"0000002f00000000000000270000000000000024000000000000000e00000000",
            INIT_19 => X"0000002000000000000000220000000000000027000000000000002f00000000",
            INIT_1A => X"00000006000000000000001b0000000000000036000000000000002000000000",
            INIT_1B => X"0000002700000000000000000000000000000000000000000000000300000000",
            INIT_1C => X"0000002200000000000000240000000000000023000000000000001b00000000",
            INIT_1D => X"0000000b00000000000000120000000000000013000000000000001a00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_1F => X"00000036000000000000002e0000000000000000000000000000000000000000",
            INIT_20 => X"0000000900000000000000100000000000000018000000000000001e00000000",
            INIT_21 => X"0000000000000000000000010000000000000004000000000000000800000000",
            INIT_22 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_23 => X"0000000600000000000000060000000000000007000000000000000000000000",
            INIT_24 => X"0000000000000000000000060000000000000002000000000000000500000000",
            INIT_25 => X"0000002a00000000000000020000000000000000000000000000000000000000",
            INIT_26 => X"00000009000000000000000c0000000000000000000000000000000000000000",
            INIT_27 => X"0000000d000000000000000b0000000000000007000000000000000000000000",
            INIT_28 => X"0000000900000000000000070000000000000004000000000000000800000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000005000000000000000b0000000000000009000000000000000900000000",
            INIT_2C => X"00000072000000000000001b0000000000000000000000000000000000000000",
            INIT_2D => X"000000070000000000000000000000000000000000000000000000a500000000",
            INIT_2E => X"0000000d00000000000000090000000000000000000000000000000000000000",
            INIT_2F => X"0000005800000000000000000000000000000003000000000000000d00000000",
            INIT_30 => X"00000000000000000000002e0000000000000061000000000000006d00000000",
            INIT_31 => X"000000000000000000000000000000000000000e000000000000002800000000",
            INIT_32 => X"00000000000000000000000e000000000000000f000000000000000000000000",
            INIT_33 => X"000000050000000000000000000000000000000d000000000000000000000000",
            INIT_34 => X"0000006000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000000e000000000000009a00000000",
            INIT_36 => X"0000002900000000000000080000000000000004000000000000001000000000",
            INIT_37 => X"0000000000000000000000080000000000000009000000000000002200000000",
            INIT_38 => X"00000062000000000000007f0000000000000098000000000000008400000000",
            INIT_39 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000f00000000000000000000000000000012000000000000000000000000",
            INIT_3B => X"00000073000000000000005c000000000000000c000000000000000000000000",
            INIT_3C => X"00000000000000000000000c00000000000000c700000000000000b600000000",
            INIT_3D => X"000000a8000000000000001e000000000000005b000000000000003400000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000004900000000",
            INIT_3F => X"0000008d000000000000007f000000000000005b000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007400000000000000860000000000000094000000000000003c00000000",
            INIT_41 => X"0000000000000000000000100000000000000022000000000000008400000000",
            INIT_42 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000063000000000000005e00000000",
            INIT_44 => X"000000000000000000000049000000000000004d000000000000002100000000",
            INIT_45 => X"0000000000000000000000030000000000000006000000000000000a00000000",
            INIT_46 => X"0000006500000000000000030000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000004300000000",
            INIT_48 => X"0000000000000000000000000000000000000045000000000000003a00000000",
            INIT_49 => X"00000068000000000000004e000000000000003e000000000000001400000000",
            INIT_4A => X"0000009400000000000000dd00000000000000d100000000000000b900000000",
            INIT_4B => X"0000000800000000000000000000000000000025000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_50 => X"000000c800000000000000c800000000000000c9000000000000000000000000",
            INIT_51 => X"000000aa00000000000000b000000000000000bb00000000000000ca00000000",
            INIT_52 => X"0000006d000000000000007e000000000000008d000000000000009d00000000",
            INIT_53 => X"0000005300000000000000360000000000000037000000000000006300000000",
            INIT_54 => X"000000a000000000000000a300000000000000ae00000000000000bc00000000",
            INIT_55 => X"000000820000000000000088000000000000008a000000000000009400000000",
            INIT_56 => X"0000004600000000000000710000000000000073000000000000007a00000000",
            INIT_57 => X"00000086000000000000005e000000000000004a000000000000002000000000",
            INIT_58 => X"0000007a000000000000007c000000000000007e000000000000007900000000",
            INIT_59 => X"0000007700000000000000780000000000000077000000000000007600000000",
            INIT_5A => X"00000035000000000000001a000000000000005e000000000000007400000000",
            INIT_5B => X"00000072000000000000006b0000000000000061000000000000005e00000000",
            INIT_5C => X"0000007900000000000000770000000000000074000000000000007400000000",
            INIT_5D => X"0000006e0000000000000078000000000000007b000000000000007900000000",
            INIT_5E => X"000000690000000000000050000000000000002a000000000000002000000000",
            INIT_5F => X"000000750000000000000074000000000000006c000000000000006400000000",
            INIT_60 => X"00000071000000000000007a0000000000000077000000000000007400000000",
            INIT_61 => X"0000001b00000000000000430000000000000065000000000000006900000000",
            INIT_62 => X"00000065000000000000005f0000000000000051000000000000003900000000",
            INIT_63 => X"0000007200000000000000740000000000000073000000000000007400000000",
            INIT_64 => X"00000040000000000000005b0000000000000067000000000000007000000000",
            INIT_65 => X"00000000000000000000000a0000000000000006000000000000002e00000000",
            INIT_66 => X"00000076000000000000005a0000000000000039000000000000003a00000000",
            INIT_67 => X"00000063000000000000006b000000000000006e000000000000007300000000",
            INIT_68 => X"0000000700000000000000000000000000000000000000000000002600000000",
            INIT_69 => X"000000180000000000000000000000000000001a000000000000003900000000",
            INIT_6A => X"000000700000000000000073000000000000003b000000000000002300000000",
            INIT_6B => X"0000002c0000000000000024000000000000004a000000000000006e00000000",
            INIT_6C => X"0000003700000000000000380000000000000015000000000000000e00000000",
            INIT_6D => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000003800000000000000670000000000000070000000000000003100000000",
            INIT_6F => X"0000003700000000000000170000000000000000000000000000001400000000",
            INIT_70 => X"0000000000000000000000000000000000000005000000000000002c00000000",
            INIT_71 => X"000000210000000000000036000000000000002a000000000000000000000000",
            INIT_72 => X"0000000f00000000000000000000000000000066000000000000006f00000000",
            INIT_73 => X"0000000000000000000000370000000000000027000000000000000000000000",
            INIT_74 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_75 => X"0000007600000000000000000000000000000000000000000000001300000000",
            INIT_76 => X"0000000d00000000000000000000000000000000000000000000001600000000",
            INIT_77 => X"0000000000000000000000000000000000000039000000000000002000000000",
            INIT_78 => X"0000000000000000000000190000000000000010000000000000000000000000",
            INIT_79 => X"00000017000000000000004c0000000000000000000000000000000000000000",
            INIT_7A => X"0000001a000000000000001b0000000000000000000000000000000000000000",
            INIT_7B => X"0000000c00000000000000000000000000000000000000000000002500000000",
            INIT_7C => X"0000000000000000000000000000000000000034000000000000000d00000000",
            INIT_7D => X"000000000000000000000017000000000000003e000000000000001800000000",
            INIT_7E => X"000000150000000000000006000000000000001f000000000000000000000000",
            INIT_7F => X"0000000200000000000000190000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "samplegold_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002600000000000000000000000000000015000000000000001800000000",
            INIT_01 => X"0000000000000000000000060000000000000023000000000000003a00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_03 => X"0000000300000000000000000000000000000016000000000000000000000000",
            INIT_04 => X"000000360000000000000021000000000000000c000000000000001500000000",
            INIT_05 => X"0000000f0000000000000009000000000000000a000000000000001b00000000",
            INIT_06 => X"000000140000000000000010000000000000000f000000000000000e00000000",
            INIT_07 => X"0000001d00000000000000090000000000000004000000000000002a00000000",
            INIT_08 => X"0000000000000000000000000000000000000023000000000000001e00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"000000150000000000000027000000000000000f000000000000000200000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_21 => X"00000025000000000000004c0000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000000000000000000004d0000000000000053000000000000001700000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000005f00000000000000500000000000000033000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000009000000000000005200000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000004600000000000000510000000000000052000000000000004e00000000",
            INIT_2D => X"00000020000000000000002a000000000000001b000000000000002300000000",
            INIT_2E => X"0000000000000000000000150000000000000023000000000000000000000000",
            INIT_2F => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000003600000000000000000000000000000000000000000000004700000000",
            INIT_31 => X"000000000000000000000000000000000000002a000000000000004100000000",
            INIT_32 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_33 => X"00000031000000000000004b0000000000000014000000000000000000000000",
            INIT_34 => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_36 => X"0000000c00000000000000000000000000000000000000000000000b00000000",
            INIT_37 => X"000000000000000000000027000000000000004c000000000000002b00000000",
            INIT_38 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000001900000000000000100000000000000000000000000000000000000000",
            INIT_3B => X"000000000000000000000000000000000000000b000000000000001d00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000500000000000000100000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"00000021000000000000000d0000000000000001000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000025000000000000002900000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"000000b7000000000000008f000000000000006e000000000000005200000000",
            INIT_56 => X"000000010000000000000001000000000000001700000000000000d500000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000006700000000000000460000000000000012000000000000000000000000",
            INIT_59 => X"000000ec000000000000005d0000000000000027000000000000003100000000",
            INIT_5A => X"000000000000000000000003000000000000000000000000000000a400000000",
            INIT_5B => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000004c000000000000003e000000000000002a000000000000003200000000",
            INIT_5D => X"000000b3000000000000011500000000000000a8000000000000005c00000000",
            INIT_5E => X"00000000000000000000002d0000000000000000000000000000003f00000000",
            INIT_5F => X"0000002d00000000000000420000000000000008000000000000000000000000",
            INIT_60 => X"0000011300000000000000e30000000000000052000000000000001a00000000",
            INIT_61 => X"0000003600000000000000630000000000000105000000000000012d00000000",
            INIT_62 => X"0000006d00000000000000000000000000000099000000000000004e00000000",
            INIT_63 => X"000000080000000000000009000000000000002d000000000000004d00000000",
            INIT_64 => X"000000d8000000000000010a00000000000000fb000000000000007300000000",
            INIT_65 => X"000000b9000000000000009d00000000000000d5000000000000010100000000",
            INIT_66 => X"00000097000000000000008f0000000000000019000000000000009e00000000",
            INIT_67 => X"00000071000000000000001d0000000000000000000000000000001e00000000",
            INIT_68 => X"0000002f000000000000006b00000000000000cb00000000000000f500000000",
            INIT_69 => X"0000004d00000000000000ae00000000000000e300000000000000c800000000",
            INIT_6A => X"00000015000000000000007a000000000000003f000000000000000800000000",
            INIT_6B => X"000000fc00000000000000c10000000000000044000000000000000400000000",
            INIT_6C => X"00000035000000000000000e000000000000001e000000000000009300000000",
            INIT_6D => X"000000000000000000000000000000000000005600000000000000c100000000",
            INIT_6E => X"00000049000000000000002e0000000000000078000000000000003e00000000",
            INIT_6F => X"0000008400000000000000f800000000000000bd000000000000008c00000000",
            INIT_70 => X"0000007000000000000000050000000000000032000000000000003a00000000",
            INIT_71 => X"0000002f00000000000000000000000000000000000000000000002e00000000",
            INIT_72 => X"0000007e0000000000000051000000000000003f000000000000005200000000",
            INIT_73 => X"0000004300000000000000690000000000000094000000000000008e00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_75 => X"0000001800000000000000150000000000000005000000000000000000000000",
            INIT_76 => X"0000000000000000000000010000000000000000000000000000000300000000",
            INIT_77 => X"0000002600000000000000080000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000005f0000000000000054000000000000004e000000000000002e00000000",
            INIT_7A => X"00000050000000000000004e0000000000000054000000000000006000000000",
            INIT_7B => X"0000003200000000000000440000000000000053000000000000004200000000",
            INIT_7C => X"0000004f000000000000001d0000000000000026000000000000003900000000",
            INIT_7D => X"0000003b000000000000003f0000000000000044000000000000004200000000",
            INIT_7E => X"0000002c0000000000000035000000000000002f000000000000003400000000",
            INIT_7F => X"0000002c000000000000002a000000000000001b000000000000002900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "samplegold_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004900000000000000460000000000000017000000000000000000000000",
            INIT_01 => X"0000001c0000000000000025000000000000002a000000000000003300000000",
            INIT_02 => X"0000001a000000000000001e0000000000000021000000000000001b00000000",
            INIT_03 => X"00000000000000000000000e0000000000000036000000000000001b00000000",
            INIT_04 => X"000000140000000000000014000000000000001e000000000000002000000000",
            INIT_05 => X"0000001100000000000000140000000000000013000000000000001500000000",
            INIT_06 => X"00000056000000000000001f0000000000000016000000000000001300000000",
            INIT_07 => X"00000029000000000000002b0000000000000015000000000000001e00000000",
            INIT_08 => X"000000160000000000000012000000000000000f000000000000000a00000000",
            INIT_09 => X"0000001f00000000000000230000000000000015000000000000001000000000",
            INIT_0A => X"0000000000000000000000060000000000000000000000000000000100000000",
            INIT_0B => X"0000000e000000000000001f0000000000000021000000000000001c00000000",
            INIT_0C => X"0000001200000000000000190000000000000014000000000000000f00000000",
            INIT_0D => X"0000004400000000000000020000000000000000000000000000000000000000",
            INIT_0E => X"0000002900000000000000270000000000000000000000000000006d00000000",
            INIT_0F => X"000000100000000000000010000000000000001b000000000000001600000000",
            INIT_10 => X"0000004900000000000000040000000000000013000000000000001900000000",
            INIT_11 => X"00000000000000000000005b0000000000000079000000000000007300000000",
            INIT_12 => X"0000002b0000000000000006000000000000003d000000000000000000000000",
            INIT_13 => X"0000000700000000000000150000000000000011000000000000001e00000000",
            INIT_14 => X"0000002900000000000000150000000000000031000000000000000000000000",
            INIT_15 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000080000000000000035000000000000007800000000",
            INIT_17 => X"000000320000000000000024000000000000000c000000000000001100000000",
            INIT_18 => X"0000000000000000000000000000000000000034000000000000004400000000",
            INIT_19 => X"0000006b00000000000000550000000000000048000000000000003700000000",
            INIT_1A => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000003e00000000000000100000000000000032000000000000000000000000",
            INIT_1C => X"0000002f00000000000000230000000000000000000000000000001500000000",
            INIT_1D => X"000000000000000000000001000000000000006f000000000000006600000000",
            INIT_1E => X"0000006400000000000000000000000000000046000000000000001300000000",
            INIT_1F => X"0000000000000000000000310000000000000021000000000000006500000000",
            INIT_20 => X"00000097000000000000006a0000000000000025000000000000000000000000",
            INIT_21 => X"0000005c00000000000000510000000000000047000000000000004c00000000",
            INIT_22 => X"00000017000000000000001e000000000000001f000000000000009700000000",
            INIT_23 => X"0000000000000000000000000000000000000001000000000000002e00000000",
            INIT_24 => X"000000190000000000000012000000000000007f000000000000001f00000000",
            INIT_25 => X"0000002300000000000000610000000000000035000000000000000e00000000",
            INIT_26 => X"0000001a00000000000000120000000000000014000000000000001400000000",
            INIT_27 => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000001400000000000000060000000000000000000000000000006400000000",
            INIT_29 => X"0000000b000000000000001b000000000000006b000000000000003700000000",
            INIT_2A => X"0000005c00000000000000560000000000000041000000000000001800000000",
            INIT_2B => X"0000009f00000000000000b000000000000000a8000000000000009600000000",
            INIT_2C => X"0000003b000000000000002d000000000000003d000000000000001600000000",
            INIT_2D => X"0000001a000000000000000b0000000000000014000000000000003b00000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2F => X"000000160000000000000015000000000000000d000000000000000500000000",
            INIT_30 => X"000000140000000000000015000000000000003c000000000000003b00000000",
            INIT_31 => X"0000000d00000000000000000000000000000000000000000000000f00000000",
            INIT_32 => X"000000170000000000000015000000000000001b000000000000001300000000",
            INIT_33 => X"0000000e000000000000002f000000000000000d000000000000001100000000",
            INIT_34 => X"000000010000000000000024000000000000000a000000000000000300000000",
            INIT_35 => X"0000001700000000000000130000000000000002000000000000000900000000",
            INIT_36 => X"0000000c00000000000000120000000000000012000000000000001800000000",
            INIT_37 => X"0000000000000000000000000000000000000002000000000000000700000000",
            INIT_38 => X"0000002700000000000000000000000000000000000000000000000900000000",
            INIT_39 => X"0000000b00000000000000100000000000000018000000000000002b00000000",
            INIT_3A => X"0000000000000000000000000000000000000001000000000000000200000000",
            INIT_3B => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_3C => X"00000001000000000000000c0000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000400000000000000000000000000000009000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000300000000000000060000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000000000000000000007d000000000000004800000000",
            INIT_47 => X"0000000000000000000000030000000000000000000000000000003100000000",
            INIT_48 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_49 => X"00000030000000000000003f000000000000003d000000000000003100000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000010000000000000003e00000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000000000000000000003e000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_50 => X"0000000000000000000000160000000000000025000000000000002500000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000000000000000000000000000000000000b000000000000000b00000000",
            INIT_55 => X"00000000000000000000007f000000000000003d000000000000000000000000",
            INIT_56 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_57 => X"0000000500000000000000000000000000000016000000000000007f00000000",
            INIT_58 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"00000012000000000000007c0000000000000019000000000000004700000000",
            INIT_5A => X"0000000000000000000000090000000000000062000000000000002400000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_5C => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_5D => X"0000001c0000000000000012000000000000000e000000000000000000000000",
            INIT_5E => X"0000000900000000000000000000000000000006000000000000000100000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000c000000000000002b0000000000000048000000000000000000000000",
            INIT_62 => X"0000003f0000000000000040000000000000000d000000000000000000000000",
            INIT_63 => X"000000ae00000000000000a9000000000000009e000000000000006100000000",
            INIT_64 => X"00000000000000000000001b0000000000000005000000000000008b00000000",
            INIT_65 => X"0000000000000000000000010000000000000018000000000000003200000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000000000000000000000d000000000000002a000000000000001b00000000",
            INIT_69 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_6B => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_6C => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000190000000000000007000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_75 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_77 => X"0000000700000000000000280000000000000000000000000000000a00000000",
            INIT_78 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_79 => X"0000000800000000000000090000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000110000000000000008000000000000000800000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"000000210000000000000030000000000000001b000000000000000000000000",
            INIT_7E => X"000000170000000000000000000000000000001c000000000000000700000000",
            INIT_7F => X"0000000000000000000000000000000000000032000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "samplegold_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000016000000000000002c00000000",
            INIT_02 => X"00000000000000000000006200000000000000bd000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_04 => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_05 => X"0000003000000000000000190000000000000000000000000000002000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000007400000000",
            INIT_07 => X"0000002000000000000000000000000000000036000000000000001a00000000",
            INIT_08 => X"0000002600000000000000000000000000000015000000000000000000000000",
            INIT_09 => X"000000000000000000000008000000000000008c000000000000008300000000",
            INIT_0A => X"0000004000000000000000200000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000008f0000000000000026000000000000001900000000",
            INIT_0C => X"000000e600000000000000420000000000000000000000000000001f00000000",
            INIT_0D => X"0000003500000000000000000000000000000000000000000000002700000000",
            INIT_0E => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_0F => X"000000000000000000000000000000000000001c000000000000008900000000",
            INIT_10 => X"0000000b00000000000000c80000000000000059000000000000000000000000",
            INIT_11 => X"000000d100000000000000360000000000000000000000000000000000000000",
            INIT_12 => X"0000003d00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000002600000000000000000000000000000000000000000000000f00000000",
            INIT_14 => X"00000000000000000000000000000000000000bb000000000000006200000000",
            INIT_15 => X"0000002a00000000000000a20000000000000000000000000000001100000000",
            INIT_16 => X"0000001e000000000000002c0000000000000000000000000000000000000000",
            INIT_17 => X"0000001200000000000000660000000000000000000000000000001c00000000",
            INIT_18 => X"0000004200000000000000000000000000000000000000000000005f00000000",
            INIT_19 => X"00000000000000000000006c0000000000000008000000000000000000000000",
            INIT_1A => X"0000000800000000000000210000000000000016000000000000001800000000",
            INIT_1B => X"00000025000000000000002a0000000000000049000000000000000000000000",
            INIT_1C => X"0000000000000000000000630000000000000000000000000000001400000000",
            INIT_1D => X"0000000f0000000000000000000000000000001a000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000042000000000000000000000000",
            INIT_21 => X"0000000000000000000000160000000000000004000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000006000000000000000a00000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000150000000000000045000000000000001600000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000011000000000000002300000000",
            INIT_37 => X"0000000000000000000000000000000000000035000000000000006c00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000003b000000000000003b0000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000028000000000000005c00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000008300000000000000270000000000000015000000000000001800000000",
            INIT_3E => X"00000002000000000000003f000000000000007500000000000000af00000000",
            INIT_3F => X"00000000000000000000004f000000000000002a000000000000002600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001100000000000000120000000000000000000000000000000000000000",
            INIT_41 => X"000000170000000000000044000000000000003e000000000000000d00000000",
            INIT_42 => X"00000042000000000000000e000000000000000b000000000000001c00000000",
            INIT_43 => X"0000003c00000000000000000000000000000040000000000000007000000000",
            INIT_44 => X"00000021000000000000001c000000000000002e000000000000004400000000",
            INIT_45 => X"000000000000000000000033000000000000002e000000000000003400000000",
            INIT_46 => X"0000003d0000000000000065000000000000006f000000000000000000000000",
            INIT_47 => X"0000002f00000000000000000000000000000000000000000000000900000000",
            INIT_48 => X"00000058000000000000005a0000000000000023000000000000002a00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000003700000000",
            INIT_4A => X"00000000000000000000000d000000000000001d000000000000000000000000",
            INIT_4B => X"0000003400000000000000450000000000000029000000000000000000000000",
            INIT_4C => X"0000003e000000000000004c0000000000000040000000000000004400000000",
            INIT_4D => X"0000000f0000000000000034000000000000002e000000000000002600000000",
            INIT_4E => X"00000000000000000000001a0000000000000017000000000000002d00000000",
            INIT_4F => X"0000007600000000000000550000000000000040000000000000002b00000000",
            INIT_50 => X"000000390000000000000035000000000000004e000000000000008600000000",
            INIT_51 => X"0000000400000000000000220000000000000051000000000000004300000000",
            INIT_52 => X"0000000f0000000000000000000000000000000d000000000000001400000000",
            INIT_53 => X"0000000000000000000000000000000000000008000000000000000a00000000",
            INIT_54 => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"000000180000000000000006000000000000001f000000000000001c00000000",
            INIT_56 => X"0000005200000000000000240000000000000000000000000000002200000000",
            INIT_57 => X"000000460000000000000050000000000000004e000000000000005b00000000",
            INIT_58 => X"0000000c000000000000001c0000000000000033000000000000003c00000000",
            INIT_59 => X"0000002d000000000000002b000000000000002b000000000000002100000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "samplegold_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000a00000000000000000000000000000004000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000003600000000000000490000000000000034000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000320000000000000061000000000000002a000000000000000000000000",
            INIT_27 => X"00000007000000000000008d0000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000001b00000000000000300000000000000078000000000000005800000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000001a00000000000000000000000000000017000000000000000000000000",
            INIT_2E => X"000000fc00000000000000f9000000000000009c000000000000001a00000000",
            INIT_2F => X"0000002000000000000000000000000000000000000000000000005d00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000006a00000000",
            INIT_31 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000002400000000000000360000000000000042000000000000009e00000000",
            INIT_33 => X"0000005e000000000000009c0000000000000041000000000000000000000000",
            INIT_34 => X"0000001600000000000000100000000000000094000000000000000000000000",
            INIT_35 => X"0000004700000000000000680000000000000009000000000000000000000000",
            INIT_36 => X"0000007000000000000000000000000000000000000000000000004100000000",
            INIT_37 => X"0000000000000000000000000000000000000046000000000000009100000000",
            INIT_38 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_39 => X"00000000000000000000004c0000000000000096000000000000005900000000",
            INIT_3A => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000004d00000000000000320000000000000000000000000000002a00000000",
            INIT_3D => X"0000002100000000000000000000000000000053000000000000007500000000",
            INIT_3E => X"00000000000000000000001e0000000000000015000000000000000a00000000",
            INIT_3F => X"0000002f00000000000000180000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008f000000000000009e0000000000000091000000000000002700000000",
            INIT_41 => X"0000002b000000000000003e0000000000000000000000000000004800000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_43 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_46 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_47 => X"0000002f00000000000000420000000000000031000000000000001000000000",
            INIT_48 => X"0000000d00000000000000190000000000000027000000000000003200000000",
            INIT_49 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000c800000000000000c60000000000000017000000000000000c00000000",
            INIT_4B => X"000000ab00000000000000c000000000000000cc00000000000000cb00000000",
            INIT_4C => X"000000660000000000000082000000000000009600000000000000a300000000",
            INIT_4D => X"0000000a000000000000001b000000000000004b000000000000005f00000000",
            INIT_4E => X"000000a600000000000000aa00000000000000bb000000000000003e00000000",
            INIT_4F => X"0000007600000000000000780000000000000086000000000000009500000000",
            INIT_50 => X"00000053000000000000005a0000000000000064000000000000006f00000000",
            INIT_51 => X"0000004c000000000000001c0000000000000000000000000000003e00000000",
            INIT_52 => X"00000068000000000000006b000000000000006f000000000000007300000000",
            INIT_53 => X"000000620000000000000062000000000000005e000000000000006200000000",
            INIT_54 => X"00000007000000000000002a000000000000005b000000000000005f00000000",
            INIT_55 => X"00000051000000000000004c000000000000003f000000000000002400000000",
            INIT_56 => X"0000005f000000000000005b000000000000005a000000000000005700000000",
            INIT_57 => X"00000067000000000000006b0000000000000067000000000000006100000000",
            INIT_58 => X"0000003a00000000000000000000000000000015000000000000005800000000",
            INIT_59 => X"0000005a00000000000000510000000000000050000000000000005500000000",
            INIT_5A => X"0000005e000000000000005d000000000000005b000000000000005c00000000",
            INIT_5B => X"0000005c00000000000000640000000000000060000000000000005800000000",
            INIT_5C => X"0000004a00000000000000480000000000000015000000000000000d00000000",
            INIT_5D => X"0000005a000000000000005a0000000000000059000000000000004a00000000",
            INIT_5E => X"0000003400000000000000450000000000000051000000000000005a00000000",
            INIT_5F => X"000000000000000000000002000000000000001d000000000000002a00000000",
            INIT_60 => X"0000004100000000000000330000000000000000000000000000003b00000000",
            INIT_61 => X"000000490000000000000058000000000000005b000000000000005d00000000",
            INIT_62 => X"000000000000000000000004000000000000001a000000000000003600000000",
            INIT_63 => X"0000001e00000000000000210000000000000000000000000000000000000000",
            INIT_64 => X"0000005a000000000000001f0000000000000000000000000000000c00000000",
            INIT_65 => X"0000001700000000000000380000000000000041000000000000005900000000",
            INIT_66 => X"0000002700000000000000000000000000000004000000000000000700000000",
            INIT_67 => X"000000000000000000000027000000000000002a000000000000003000000000",
            INIT_68 => X"0000004300000000000000570000000000000006000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_6A => X"0000002800000000000000310000000000000018000000000000000000000000",
            INIT_6B => X"0000000d000000000000000d0000000000000027000000000000003500000000",
            INIT_6C => X"0000001f000000000000002c0000000000000045000000000000002000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000210000000000000015000000000000001900000000",
            INIT_6F => X"0000001b0000000000000017000000000000001c000000000000000e00000000",
            INIT_70 => X"0000000000000000000000000000000000000010000000000000002e00000000",
            INIT_71 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_73 => X"0000002500000000000000030000000000000009000000000000000900000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000021000000000000001c0000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000110000000000000000000000000000000d00000000",
            INIT_78 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000170000000000000017000000000000001900000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "samplegold_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000c000000000000000e0000000000000007000000000000000000000000",
            INIT_04 => X"0000000f0000000000000002000000000000000f000000000000000c00000000",
            INIT_05 => X"0000000b00000000000000000000000000000005000000000000003c00000000",
            INIT_06 => X"0000000000000000000000020000000000000000000000000000002a00000000",
            INIT_07 => X"00000008000000000000000b000000000000000d000000000000000e00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000011000000000000002a0000000000000026000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000004000000000000000700000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000002c000000000000001c0000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000005300000000000000420000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000068000000000000005d0000000000000000000000000000000000000000",
            INIT_1B => X"0000000a00000000000000000000000000000045000000000000007900000000",
            INIT_1C => X"0000000e000000000000003d0000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000002a00000000000000220000000000000004000000000000000000000000",
            INIT_22 => X"0000001600000000000000000000000000000000000000000000003200000000",
            INIT_23 => X"0000000000000000000000000000000000000011000000000000001100000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"00000013000000000000000c000000000000000f000000000000000000000000",
            INIT_26 => X"0000006e0000000000000002000000000000001d000000000000000d00000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000006700000000",
            INIT_28 => X"0000000000000000000000b00000000000000000000000000000002300000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2A => X"0000008000000000000000590000000000000040000000000000000500000000",
            INIT_2B => X"00000073000000000000003c0000000000000023000000000000009a00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2D => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_2E => X"0000006300000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000027000000000000000e00000000",
            INIT_30 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000006400000000000000090000000000000000000000000000000000000000",
            INIT_33 => X"0000000e00000000000000000000000000000015000000000000001a00000000",
            INIT_34 => X"000000dd000000000000009e0000000000000043000000000000005300000000",
            INIT_35 => X"0000001e000000000000006700000000000000eb00000000000000e900000000",
            INIT_36 => X"0000000a00000000000000590000000000000002000000000000002000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"00000023000000000000003a0000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000001d00000000000000130000000000000025000000000000001800000000",
            INIT_3C => X"0000002600000000000000120000000000000020000000000000002400000000",
            INIT_3D => X"0000000e00000000000000160000000000000000000000000000001a00000000",
            INIT_3E => X"0000000f000000000000001a0000000000000000000000000000003600000000",
            INIT_3F => X"0000001b0000000000000022000000000000002b000000000000002100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001600000000000000190000000000000013000000000000001b00000000",
            INIT_41 => X"0000001800000000000000380000000000000000000000000000001600000000",
            INIT_42 => X"00000021000000000000001c0000000000000019000000000000000000000000",
            INIT_43 => X"000000120000000000000010000000000000001a000000000000001900000000",
            INIT_44 => X"000000060000000000000010000000000000000f000000000000001200000000",
            INIT_45 => X"0000000000000000000000100000000000000019000000000000000000000000",
            INIT_46 => X"00000010000000000000000e000000000000000e000000000000002300000000",
            INIT_47 => X"00000005000000000000000f000000000000000f000000000000001400000000",
            INIT_48 => X"000000330000000000000015000000000000000c000000000000000e00000000",
            INIT_49 => X"0000001600000000000000170000000000000014000000000000000000000000",
            INIT_4A => X"0000001600000000000000130000000000000013000000000000000e00000000",
            INIT_4B => X"0000000000000000000000000000000000000007000000000000000800000000",
            INIT_4C => X"0000000c000000000000002a000000000000002e000000000000000000000000",
            INIT_4D => X"0000001000000000000000100000000000000019000000000000001a00000000",
            INIT_4E => X"0000000000000000000000150000000000000017000000000000001400000000",
            INIT_4F => X"00000013000000000000000d0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000f30000000000000000000000000000000000000000",
            INIT_51 => X"0000001700000000000000110000000000000017000000000000002a00000000",
            INIT_52 => X"0000000400000000000000000000000000000000000000000000002100000000",
            INIT_53 => X"0000000000000000000000000000000000000038000000000000001900000000",
            INIT_54 => X"00000000000000000000005400000000000000d6000000000000000000000000",
            INIT_55 => X"00000000000000000000001a0000000000000013000000000000000e00000000",
            INIT_56 => X"000000060000000000000000000000000000000f000000000000001e00000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"000000000000000000000000000000000000006400000000000000aa00000000",
            INIT_59 => X"0000000000000000000000290000000000000000000000000000001a00000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_5B => X"000000ab00000000000000500000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000004f000000000000000000000000000000b7000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000310000000000000000000000000000005800000000",
            INIT_60 => X"0000000000000000000000000000000000000049000000000000000500000000",
            INIT_61 => X"0000000000000000000000240000000000000032000000000000005800000000",
            INIT_62 => X"00000052000000000000008a0000000000000000000000000000000000000000",
            INIT_63 => X"0000004100000000000000320000000000000000000000000000000c00000000",
            INIT_64 => X"00000000000000000000000c0000000000000000000000000000006d00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000005500000000",
            INIT_66 => X"00000013000000000000000000000000000000c5000000000000000000000000",
            INIT_67 => X"0000000b00000000000000910000000000000000000000000000000000000000",
            INIT_68 => X"0000004300000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000002a0000000000000039000000000000000000000000000000cd00000000",
            INIT_6B => X"000000000000000000000000000000000000007e000000000000000000000000",
            INIT_6C => X"00000000000000000000002b0000000000000000000000000000000000000000",
            INIT_6D => X"0000003e000000000000000c0000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000400000000000000013000000000000000000000000",
            INIT_6F => X"0000000a00000000000000000000000000000000000000000000001800000000",
            INIT_70 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_71 => X"00000000000000000000000b000000000000000a000000000000000600000000",
            INIT_72 => X"000000000000000000000000000000000000002b000000000000002300000000",
            INIT_73 => X"0000011300000000000001120000000000000120000000000000000000000000",
            INIT_74 => X"000000ea00000000000000f00000000000000102000000000000010d00000000",
            INIT_75 => X"000000a200000000000000a300000000000000c700000000000000db00000000",
            INIT_76 => X"0000008b000000000000003d0000000000000041000000000000008d00000000",
            INIT_77 => X"000000ed00000000000000f200000000000000f3000000000000010300000000",
            INIT_78 => X"000000bf00000000000000cd00000000000000cf00000000000000e000000000",
            INIT_79 => X"00000068000000000000009a00000000000000ad00000000000000b500000000",
            INIT_7A => X"000000ba000000000000009f000000000000005f000000000000003100000000",
            INIT_7B => X"000000be00000000000000c700000000000000c700000000000000c000000000",
            INIT_7C => X"000000b600000000000000b800000000000000c100000000000000bd00000000",
            INIT_7D => X"00000051000000000000002c000000000000005d00000000000000ad00000000",
            INIT_7E => X"000000b800000000000000ac000000000000009b000000000000008600000000",
            INIT_7F => X"000000c400000000000000bf00000000000000bb00000000000000ba00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "samplegold_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009b00000000000000b500000000000000c100000000000000c700000000",
            INIT_01 => X"000000a000000000000000890000000000000025000000000000002d00000000",
            INIT_02 => X"000000c000000000000000c000000000000000b500000000000000a200000000",
            INIT_03 => X"0000009c00000000000000b700000000000000c100000000000000c000000000",
            INIT_04 => X"0000002d0000000000000086000000000000009f00000000000000a600000000",
            INIT_05 => X"0000009800000000000000970000000000000084000000000000003300000000",
            INIT_06 => X"000000bb00000000000000be00000000000000c200000000000000c000000000",
            INIT_07 => X"0000003f000000000000005c000000000000008c00000000000000ad00000000",
            INIT_08 => X"00000034000000000000002e0000000000000013000000000000002200000000",
            INIT_09 => X"000000c2000000000000008c0000000000000077000000000000001800000000",
            INIT_0A => X"0000007700000000000000a700000000000000bd00000000000000c200000000",
            INIT_0B => X"0000001400000000000000040000000000000012000000000000003100000000",
            INIT_0C => X"000000100000000000000045000000000000001c000000000000000600000000",
            INIT_0D => X"000000bf00000000000000c0000000000000005f000000000000001f00000000",
            INIT_0E => X"0000002b0000000000000037000000000000006e000000000000009500000000",
            INIT_0F => X"0000002b00000000000000450000000000000030000000000000002000000000",
            INIT_10 => X"0000001700000000000000300000000000000020000000000000001e00000000",
            INIT_11 => X"0000003e00000000000000a200000000000000c0000000000000004100000000",
            INIT_12 => X"000000000000000000000000000000000000000a000000000000000e00000000",
            INIT_13 => X"0000002d000000000000001f000000000000001b000000000000002400000000",
            INIT_14 => X"0000002f00000000000000390000000000000050000000000000003e00000000",
            INIT_15 => X"000000080000000000000024000000000000007500000000000000ad00000000",
            INIT_16 => X"0000001200000000000000000000000000000001000000000000000d00000000",
            INIT_17 => X"0000003f00000000000000020000000000000006000000000000001100000000",
            INIT_18 => X"00000084000000000000001d000000000000001c000000000000002a00000000",
            INIT_19 => X"0000000a000000000000000d000000000000000d000000000000000700000000",
            INIT_1A => X"00000011000000000000000f0000000000000000000000000000000900000000",
            INIT_1B => X"0000000c00000000000000000000000000000000000000000000000100000000",
            INIT_1C => X"0000000e0000000000000071000000000000000c000000000000000a00000000",
            INIT_1D => X"0000000000000000000000080000000000000011000000000000000d00000000",
            INIT_1E => X"0000000f00000000000000200000000000000013000000000000000000000000",
            INIT_1F => X"00000012000000000000000a0000000000000000000000000000001100000000",
            INIT_20 => X"0000000400000000000000110000000000000057000000000000001d00000000",
            INIT_21 => X"00000010000000000000001b0000000000000008000000000000000d00000000",
            INIT_22 => X"00000020000000000000000b0000000000000020000000000000001000000000",
            INIT_23 => X"0000001e000000000000000b0000000000000000000000000000000a00000000",
            INIT_24 => X"0000000000000000000000000000000000000020000000000000005800000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000d000000000000000e0000000000000007000000000000000000000000",
            INIT_27 => X"0000005300000000000000110000000000000006000000000000000000000000",
            INIT_28 => X"00000000000000000000000c0000000000000008000000000000002700000000",
            INIT_29 => X"0000000e000000000000000c0000000000000008000000000000000400000000",
            INIT_2A => X"0000000c000000000000000c0000000000000009000000000000000300000000",
            INIT_2B => X"000000000000000000000000000000000000000b000000000000000c00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000300000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005200000000000000620000000000000044000000000000001c00000000",
            INIT_41 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"000000190000000000000033000000000000001f000000000000000000000000",
            INIT_44 => X"0000000d000000000000007c000000000000003e000000000000001600000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000500000000000000080000000000000010000000000000000a00000000",
            INIT_48 => X"00000000000000000000003d0000000000000080000000000000004100000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"00000013000000000000000d0000000000000020000000000000000000000000",
            INIT_4B => X"0000009300000000000000880000000000000074000000000000003200000000",
            INIT_4C => X"0000000700000000000000010000000000000000000000000000007200000000",
            INIT_4D => X"0000000000000000000000140000000000000000000000000000003f00000000",
            INIT_4E => X"0000005300000000000000060000000000000000000000000000001500000000",
            INIT_4F => X"00000095000000000000006d000000000000007f000000000000008200000000",
            INIT_50 => X"0000004000000000000000510000000000000037000000000000003e00000000",
            INIT_51 => X"0000000400000000000000320000000000000060000000000000000000000000",
            INIT_52 => X"0000007a0000000000000045000000000000000a000000000000000000000000",
            INIT_53 => X"000000950000000000000027000000000000002e000000000000005700000000",
            INIT_54 => X"00000000000000000000001f000000000000004f000000000000006b00000000",
            INIT_55 => X"0000000000000000000000000000000000000038000000000000001200000000",
            INIT_56 => X"0000002200000000000000780000000000000070000000000000002900000000",
            INIT_57 => X"0000006300000000000000340000000000000000000000000000000700000000",
            INIT_58 => X"0000001a00000000000000000000000000000000000000000000001300000000",
            INIT_59 => X"00000031000000000000001f0000000000000000000000000000003f00000000",
            INIT_5A => X"0000001c00000000000000120000000000000076000000000000006200000000",
            INIT_5B => X"00000001000000000000004f0000000000000000000000000000000000000000",
            INIT_5C => X"0000003200000000000000110000000000000000000000000000000000000000",
            INIT_5D => X"0000006a00000000000000610000000000000045000000000000002400000000",
            INIT_5E => X"0000001800000000000000290000000000000034000000000000006b00000000",
            INIT_5F => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"00000000000000000000000f000000000000000c000000000000000000000000",
            INIT_63 => X"000000c400000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"000000cf00000000000000d900000000000000d600000000000000cb00000000",
            INIT_65 => X"0000009500000000000000a900000000000000b600000000000000bf00000000",
            INIT_66 => X"000000060000000000000050000000000000006b000000000000007400000000",
            INIT_67 => X"000000b800000000000000ca000000000000004b000000000000002400000000",
            INIT_68 => X"0000009800000000000000a900000000000000ba00000000000000bd00000000",
            INIT_69 => X"0000006e000000000000007d0000000000000088000000000000009400000000",
            INIT_6A => X"0000002c0000000000000000000000000000001f000000000000005c00000000",
            INIT_6B => X"000000930000000000000092000000000000008f000000000000005800000000",
            INIT_6C => X"0000007c000000000000007c0000000000000083000000000000008c00000000",
            INIT_6D => X"00000005000000000000006f000000000000006f000000000000007500000000",
            INIT_6E => X"0000005600000000000000400000000000000010000000000000000000000000",
            INIT_6F => X"0000007600000000000000780000000000000077000000000000007400000000",
            INIT_70 => X"000000700000000000000078000000000000007e000000000000007b00000000",
            INIT_71 => X"0000000300000000000000000000000000000052000000000000006800000000",
            INIT_72 => X"000000710000000000000062000000000000005e000000000000004a00000000",
            INIT_73 => X"0000007c0000000000000079000000000000007d000000000000007b00000000",
            INIT_74 => X"00000049000000000000005f0000000000000059000000000000006600000000",
            INIT_75 => X"00000047000000000000000a0000000000000000000000000000000c00000000",
            INIT_76 => X"0000007b000000000000007a000000000000005e000000000000005e00000000",
            INIT_77 => X"0000002e000000000000006d0000000000000075000000000000007a00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000003300000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000073000000000000007b000000000000007b000000000000005500000000",
            INIT_7B => X"000000000000000000000000000000000000001f000000000000006a00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000003600000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001900000000000000490000000000000078000000000000007b00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "samplegold_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000007900000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000005900000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000000000000000000006e0000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000039000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000001b000000000000000b0000000000000009000000000000000900000000",
            INIT_1D => X"0000000900000000000000070000000000000005000000000000001200000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000140000000000000004000000000000000300000000",
            INIT_21 => X"0000000000000000000000000000000000000007000000000000000a00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"00000007000000000000000a0000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000008000000000000000f00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000e00000000000000050000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000001000000000000000180000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000020000000000000009000000000000001100000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"000000000000000000000000000000000000002e000000000000003d00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000004a00000000000000490000000000000011000000000000001300000000",
            INIT_33 => X"0000001300000000000000000000000000000000000000000000003300000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_35 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000002f0000000000000026000000000000002a000000000000002300000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000000000000000000000000000000000001d000000000000002200000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000700000000000000210000000000000000000000000000000000000000",
            INIT_3E => X"00000051000000000000007d000000000000009e000000000000003c00000000",
            INIT_3F => X"0000000000000000000000070000000000000015000000000000003a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"00000097000000000000008a0000000000000000000000000000000000000000",
            INIT_42 => X"00000043000000000000003b000000000000005e00000000000000a400000000",
            INIT_43 => X"0000000000000000000000000000000000000015000000000000000e00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000005100000000000000bc00000000000000db000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"00000018000000000000002e000000000000003f000000000000004f00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000001400000000000000050000000000000000000000000000000000000000",
            INIT_4D => X"0000002600000000000000360000000000000023000000000000000d00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000023000000000000000600000000",
            INIT_50 => X"0000002c00000000000000220000000000000007000000000000000100000000",
            INIT_51 => X"0000000300000000000000000000000000000000000000000000001100000000",
            INIT_52 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_54 => X"0000001e000000000000001a000000000000001a000000000000000000000000",
            INIT_55 => X"000000280000000000000031000000000000002c000000000000001a00000000",
            INIT_56 => X"0000001c000000000000001d000000000000001b000000000000001f00000000",
            INIT_57 => X"0000001c000000000000001e000000000000001b000000000000001900000000",
            INIT_58 => X"00000028000000000000001d0000000000000018000000000000001900000000",
            INIT_59 => X"0000003c0000000000000040000000000000004b000000000000003600000000",
            INIT_5A => X"0000002900000000000000270000000000000022000000000000002a00000000",
            INIT_5B => X"0000001a0000000000000026000000000000002a000000000000002b00000000",
            INIT_5C => X"0000003f000000000000002c000000000000001c000000000000001900000000",
            INIT_5D => X"0000004e000000000000005f000000000000005a000000000000005300000000",
            INIT_5E => X"0000002c000000000000002f000000000000002e000000000000003500000000",
            INIT_5F => X"0000001e000000000000001e0000000000000022000000000000002400000000",
            INIT_60 => X"00000056000000000000004b000000000000003b000000000000001400000000",
            INIT_61 => X"0000004c00000000000000620000000000000067000000000000005f00000000",
            INIT_62 => X"0000002500000000000000290000000000000033000000000000003d00000000",
            INIT_63 => X"00000019000000000000002e000000000000002a000000000000002e00000000",
            INIT_64 => X"0000005300000000000000540000000000000051000000000000003000000000",
            INIT_65 => X"000000650000000000000067000000000000006a000000000000005a00000000",
            INIT_66 => X"0000003f0000000000000039000000000000003d000000000000004f00000000",
            INIT_67 => X"0000002c0000000000000000000000000000001f000000000000002500000000",
            INIT_68 => X"00000050000000000000004e0000000000000059000000000000003e00000000",
            INIT_69 => X"0000006000000000000000690000000000000066000000000000006000000000",
            INIT_6A => X"00000019000000000000003a0000000000000042000000000000005100000000",
            INIT_6B => X"00000041000000000000000b0000000000000016000000000000001700000000",
            INIT_6C => X"0000005a00000000000000590000000000000046000000000000004b00000000",
            INIT_6D => X"00000052000000000000006c000000000000005d000000000000005500000000",
            INIT_6E => X"00000024000000000000001f0000000000000027000000000000003d00000000",
            INIT_6F => X"0000004d00000000000000170000000000000029000000000000002300000000",
            INIT_70 => X"0000004b000000000000005b0000000000000060000000000000004800000000",
            INIT_71 => X"0000003d00000000000000510000000000000062000000000000005a00000000",
            INIT_72 => X"0000002400000000000000260000000000000027000000000000003100000000",
            INIT_73 => X"0000003e000000000000002a0000000000000029000000000000003700000000",
            INIT_74 => X"00000056000000000000004a0000000000000059000000000000005500000000",
            INIT_75 => X"000000330000000000000048000000000000005b000000000000005b00000000",
            INIT_76 => X"00000000000000000000001a0000000000000027000000000000002d00000000",
            INIT_77 => X"0000004b000000000000004d000000000000001c000000000000003700000000",
            INIT_78 => X"000000580000000000000055000000000000004f000000000000005800000000",
            INIT_79 => X"00000011000000000000003b000000000000003c000000000000005800000000",
            INIT_7A => X"0000003d00000000000000230000000000000000000000000000000800000000",
            INIT_7B => X"00000058000000000000004c0000000000000050000000000000003f00000000",
            INIT_7C => X"000000550000000000000054000000000000004f000000000000005500000000",
            INIT_7D => X"000000000000000000000000000000000000003f000000000000004300000000",
            INIT_7E => X"0000004d0000000000000030000000000000001d000000000000000c00000000",
            INIT_7F => X"0000005300000000000000490000000000000034000000000000004c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "samplegold_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000052000000000000004e000000000000004b000000000000005200000000",
            INIT_01 => X"0000001c00000000000000170000000000000015000000000000003a00000000",
            INIT_02 => X"00000049000000000000003a0000000000000028000000000000002800000000",
            INIT_03 => X"0000004500000000000000590000000000000050000000000000003d00000000",
            INIT_04 => X"000000470000000000000052000000000000004a000000000000004c00000000",
            INIT_05 => X"0000002d000000000000002f000000000000002d000000000000002400000000",
            INIT_06 => X"000000430000000000000041000000000000003c000000000000003500000000",
            INIT_07 => X"000000460000000000000041000000000000004d000000000000004d00000000",
            INIT_08 => X"0000002b0000000000000050000000000000004c000000000000004d00000000",
            INIT_09 => X"0000004b00000000000000410000000000000038000000000000002d00000000",
            INIT_0A => X"0000004a00000000000000440000000000000043000000000000004500000000",
            INIT_0B => X"000000450000000000000046000000000000004b000000000000004800000000",
            INIT_0C => X"0000000000000000000000000000000000000048000000000000004e00000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"000000140000000000000014000000000000000a000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000100000000000000012000000000000001200000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000000000000000000000000000000000000b000000000000000900000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000001400000000000000090000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000010000000000000003000000000000002300000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000004c00000000000000400000000000000032000000000000000000000000",
            INIT_2F => X"0000000000000000000000060000000000000005000000000000003300000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000050000000000000019000000000000005c000000000000005d00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000004200000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000011000000000000003200000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000004d00000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000041000000000000004d000000000000004d000000000000004600000000",
            INIT_46 => X"00000032000000000000003d0000000000000039000000000000004000000000",
            INIT_47 => X"0000000e00000000000000190000000000000024000000000000002a00000000",
            INIT_48 => X"00000044000000000000004b0000000000000006000000000000000b00000000",
            INIT_49 => X"0000002200000000000000270000000000000032000000000000004200000000",
            INIT_4A => X"0000002700000000000000260000000000000020000000000000002d00000000",
            INIT_4B => X"00000022000000000000001c000000000000001d000000000000001e00000000",
            INIT_4C => X"0000002c00000000000000420000000000000043000000000000002200000000",
            INIT_4D => X"000000000000000000000000000000000000000b000000000000002000000000",
            INIT_4E => X"0000003d00000000000000400000000000000025000000000000000300000000",
            INIT_4F => X"0000002b00000000000000370000000000000039000000000000003f00000000",
            INIT_50 => X"00000000000000000000002f000000000000003d000000000000003a00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000003900000000000000420000000000000030000000000000000700000000",
            INIT_53 => X"0000005c00000000000000220000000000000032000000000000003f00000000",
            INIT_54 => X"00000000000000000000000a0000000000000063000000000000007000000000",
            INIT_55 => X"000000000000000000000000000000000000001e000000000000001a00000000",
            INIT_56 => X"0000003a0000000000000026000000000000000f000000000000000000000000",
            INIT_57 => X"000000a5000000000000009b000000000000002c000000000000003700000000",
            INIT_58 => X"00000019000000000000000f000000000000000a000000000000008d00000000",
            INIT_59 => X"0000000000000000000000060000000000000011000000000000002400000000",
            INIT_5A => X"00000042000000000000002a000000000000000a000000000000000000000000",
            INIT_5B => X"00000098000000000000009d000000000000009d000000000000003a00000000",
            INIT_5C => X"00000026000000000000002a000000000000000c000000000000004100000000",
            INIT_5D => X"00000000000000000000000b000000000000001c000000000000001200000000",
            INIT_5E => X"000000350000000000000039000000000000001e000000000000000000000000",
            INIT_5F => X"0000007f00000000000000920000000000000097000000000000009000000000",
            INIT_60 => X"0000000f000000000000001e0000000000000014000000000000004700000000",
            INIT_61 => X"0000000000000000000000000000000000000023000000000000002c00000000",
            INIT_62 => X"0000009d000000000000002e0000000000000021000000000000001300000000",
            INIT_63 => X"0000009c000000000000008200000000000000c600000000000000b700000000",
            INIT_64 => X"0000002900000000000000170000000000000050000000000000006300000000",
            INIT_65 => X"0000000a0000000000000000000000000000000e000000000000002a00000000",
            INIT_66 => X"0000010300000000000000e4000000000000001d000000000000001800000000",
            INIT_67 => X"0000007e000000000000008d00000000000000e100000000000000fd00000000",
            INIT_68 => X"0000002c00000000000000240000000000000028000000000000004400000000",
            INIT_69 => X"0000000900000000000000020000000000000005000000000000002100000000",
            INIT_6A => X"000000a5000000000000011c000000000000012d000000000000000100000000",
            INIT_6B => X"00000020000000000000003e0000000000000044000000000000007000000000",
            INIT_6C => X"0000002000000000000000260000000000000024000000000000001d00000000",
            INIT_6D => X"0000000000000000000000190000000000000000000000000000000900000000",
            INIT_6E => X"0000005e000000000000008b00000000000000cf00000000000000f000000000",
            INIT_6F => X"0000000e00000000000000230000000000000000000000000000001c00000000",
            INIT_70 => X"0000001a00000000000000230000000000000014000000000000000800000000",
            INIT_71 => X"000000750000000000000016000000000000001b000000000000000000000000",
            INIT_72 => X"0000004700000000000000580000000000000066000000000000006c00000000",
            INIT_73 => X"00000009000000000000001f000000000000001d000000000000001f00000000",
            INIT_74 => X"0000000d00000000000000230000000000000041000000000000002400000000",
            INIT_75 => X"00000049000000000000004b0000000000000022000000000000000700000000",
            INIT_76 => X"0000002600000000000000280000000000000033000000000000004200000000",
            INIT_77 => X"00000017000000000000000b0000000000000012000000000000001200000000",
            INIT_78 => X"0000000400000000000000060000000000000022000000000000003700000000",
            INIT_79 => X"0000001600000000000000250000000000000033000000000000000d00000000",
            INIT_7A => X"0000001800000000000000220000000000000003000000000000000100000000",
            INIT_7B => X"0000000400000000000000000000000000000000000000000000000a00000000",
            INIT_7C => X"0000000000000000000000000000000000000009000000000000000f00000000",
            INIT_7D => X"0000003900000000000000300000000000000037000000000000003500000000",
            INIT_7E => X"0000003e00000000000000480000000000000057000000000000004f00000000",
            INIT_7F => X"0000003300000000000000360000000000000034000000000000003200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "samplegold_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000036000000000000001c0000000000000020000000000000002d00000000",
            INIT_01 => X"0000005800000000000000430000000000000034000000000000003600000000",
            INIT_02 => X"00000042000000000000005f0000000000000075000000000000006f00000000",
            INIT_03 => X"0000000d00000000000000170000000000000025000000000000002f00000000",
            INIT_04 => X"00000039000000000000003b0000000000000012000000000000000800000000",
            INIT_05 => X"00000074000000000000006f000000000000004e000000000000004100000000",
            INIT_06 => X"00000022000000000000004b000000000000007e000000000000008100000000",
            INIT_07 => X"00000035000000000000002f000000000000002e000000000000002a00000000",
            INIT_08 => X"00000027000000000000002f0000000000000036000000000000003b00000000",
            INIT_09 => X"00000068000000000000006c0000000000000075000000000000003500000000",
            INIT_0A => X"0000005c00000000000000720000000000000080000000000000007100000000",
            INIT_0B => X"0000002c000000000000002c0000000000000033000000000000005800000000",
            INIT_0C => X"0000005500000000000000260000000000000000000000000000000000000000",
            INIT_0D => X"00000075000000000000005b000000000000005a000000000000006300000000",
            INIT_0E => X"0000007100000000000000860000000000000087000000000000008300000000",
            INIT_0F => X"0000002700000000000000260000000000000029000000000000003700000000",
            INIT_10 => X"0000004e000000000000003e000000000000005d000000000000003c00000000",
            INIT_11 => X"000000730000000000000087000000000000007c000000000000004500000000",
            INIT_12 => X"0000004d00000000000000800000000000000087000000000000007b00000000",
            INIT_13 => X"0000004900000000000000490000000000000037000000000000003b00000000",
            INIT_14 => X"0000006e000000000000003a0000000000000036000000000000004000000000",
            INIT_15 => X"00000071000000000000006c000000000000007f000000000000008a00000000",
            INIT_16 => X"0000004c000000000000006b000000000000007b000000000000008300000000",
            INIT_17 => X"0000003c000000000000002f000000000000003b000000000000004b00000000",
            INIT_18 => X"00000051000000000000000c000000000000002d000000000000004100000000",
            INIT_19 => X"00000084000000000000007a0000000000000072000000000000006a00000000",
            INIT_1A => X"0000002e00000000000000500000000000000076000000000000008300000000",
            INIT_1B => X"000000170000000000000004000000000000001e000000000000002c00000000",
            INIT_1C => X"0000006e0000000000000046000000000000003f000000000000004300000000",
            INIT_1D => X"00000085000000000000007d0000000000000080000000000000007e00000000",
            INIT_1E => X"0000000000000000000000530000000000000054000000000000007100000000",
            INIT_1F => X"00000074000000000000008d0000000000000055000000000000000800000000",
            INIT_20 => X"0000007b0000000000000086000000000000005a000000000000007f00000000",
            INIT_21 => X"0000007a000000000000008b000000000000007a000000000000007b00000000",
            INIT_22 => X"0000005c0000000000000043000000000000002d000000000000005a00000000",
            INIT_23 => X"000000af0000000000000095000000000000009d00000000000000a900000000",
            INIT_24 => X"00000081000000000000007e000000000000007f000000000000008900000000",
            INIT_25 => X"0000003800000000000000680000000000000088000000000000008600000000",
            INIT_26 => X"0000005f00000000000000a700000000000000aa000000000000002700000000",
            INIT_27 => X"0000005200000000000000790000000000000065000000000000004d00000000",
            INIT_28 => X"0000006100000000000000750000000000000072000000000000005200000000",
            INIT_29 => X"0000003d000000000000003b000000000000005f000000000000006e00000000",
            INIT_2A => X"00000038000000000000004b0000000000000058000000000000006100000000",
            INIT_2B => X"0000006a000000000000005b0000000000000032000000000000003b00000000",
            INIT_2C => X"0000007a0000000000000062000000000000005e000000000000005e00000000",
            INIT_2D => X"0000003e000000000000003f0000000000000040000000000000006800000000",
            INIT_2E => X"0000005500000000000000640000000000000050000000000000003500000000",
            INIT_2F => X"000000620000000000000052000000000000003f000000000000003c00000000",
            INIT_30 => X"0000006f00000000000000800000000000000088000000000000006d00000000",
            INIT_31 => X"0000005a000000000000004b000000000000003e000000000000004b00000000",
            INIT_32 => X"00000038000000000000002c0000000000000039000000000000004c00000000",
            INIT_33 => X"00000042000000000000003f0000000000000049000000000000004600000000",
            INIT_34 => X"0000003a00000000000000560000000000000059000000000000004b00000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000000000000000000001000000000000000b000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000000000000000000006000000000000000c000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000006000000000000002200000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"000000000000000000000000000000000000000e000000000000000d00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000a00000000000000020000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000015000000000000001400000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000020000000000000002000000000000000000000000",
            INIT_5B => X"0000001b00000000000000300000000000000001000000000000000000000000",
            INIT_5C => X"00000000000000000000001c000000000000000a000000000000003300000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000005000000000000000580000000000000000000000000000000000000000",
            INIT_5F => X"0000000500000000000000000000000000000002000000000000000800000000",
            INIT_60 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_61 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000120000000000000018000000000000000000000000",
            INIT_63 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000023000000000000000a0000000000000000000000000000000000000000",
            INIT_67 => X"0000000500000000000000000000000000000000000000000000001600000000",
            INIT_68 => X"00000000000000000000002b0000000000000010000000000000000100000000",
            INIT_69 => X"000000140000000000000005000000000000000a000000000000000600000000",
            INIT_6A => X"0000000000000000000000000000000000000012000000000000002300000000",
            INIT_6B => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_6C => X"0000001100000000000000170000000000000003000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000005000000000000000400000000",
            INIT_6E => X"0000000200000000000000000000000000000000000000000000001200000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000f00000000000000090000000000000006000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000004000000000000001e00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000700000000000000000000000000000000000000000000000300000000",
            INIT_7A => X"00000011000000000000000d000000000000000b000000000000000900000000",
            INIT_7B => X"0000000000000000000000000000000000000008000000000000001900000000",
            INIT_7C => X"0000000e00000000000000110000000000000000000000000000000000000000",
            INIT_7D => X"00000037000000000000000b0000000000000000000000000000000000000000",
            INIT_7E => X"0000000a00000000000000030000000000000000000000000000000500000000",
            INIT_7F => X"0000000000000000000000070000000000000005000000000000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "samplegold_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_01 => X"00000000000000000000003c0000000000000001000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_03 => X"000000000000000000000000000000000000001b000000000000001e00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000400000000000000000000000000000036000000000000000800000000",
            INIT_06 => X"0000002500000000000000000000000000000000000000000000001100000000",
            INIT_07 => X"000000070000000000000000000000000000000e000000000000000800000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_09 => X"0000001900000000000000130000000000000000000000000000001900000000",
            INIT_0A => X"0000000b00000000000000070000000000000000000000000000000000000000",
            INIT_0B => X"0000001c00000000000000120000000000000000000000000000000900000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000170000000000000000000000000000000400000000",
            INIT_0E => X"00000001000000000000001a0000000000000000000000000000000000000000",
            INIT_0F => X"00000000000000000000000e0000000000000013000000000000000000000000",
            INIT_10 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000010000000000000013000000000000000000000000",
            INIT_12 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000003000000000000000d0000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000005000000000000000f00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000001b0000000000000000000000000000002b000000000000000c00000000",
            INIT_19 => X"0000000000000000000000000000000000000009000000000000001a00000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000003900000000000000100000000000000000000000000000001c00000000",
            INIT_1D => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000030000000000000000000000000000000600000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000001400000000000000240000000000000007000000000000000000000000",
            INIT_21 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000000f000000000000001a00000000",
            INIT_24 => X"0000000700000000000000120000000000000000000000000000000000000000",
            INIT_25 => X"0000001c00000000000000000000000000000003000000000000000000000000",
            INIT_26 => X"00000000000000000000000e0000000000000017000000000000001900000000",
            INIT_27 => X"0000001900000000000000120000000000000005000000000000000000000000",
            INIT_28 => X"0000001c00000000000000190000000000000016000000000000001500000000",
            INIT_29 => X"0000001b000000000000001c0000000000000028000000000000002100000000",
            INIT_2A => X"000000000000000000000000000000000000000c000000000000001100000000",
            INIT_2B => X"0000001700000000000000070000000000000000000000000000000000000000",
            INIT_2C => X"0000002a000000000000002a0000000000000026000000000000001c00000000",
            INIT_2D => X"0000000600000000000000160000000000000015000000000000002500000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000011000000000000001b0000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000050000000000000007000000000000000b00000000",
            INIT_31 => X"00000000000000000000002d000000000000001c000000000000001600000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000003f0000000000000004000000000000000a000000000000000500000000",
            INIT_35 => X"0000000000000000000000000000000000000025000000000000004300000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000a00000000000000160000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000008000000000000001100000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000001400000000000000030000000000000002000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000900000000000000050000000000000014000000000000000f00000000",
            INIT_41 => X"0000000000000000000000000000000000000017000000000000002a00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000001200000000000000020000000000000000000000000000000000000000",
            INIT_44 => X"000000070000000000000029000000000000003f000000000000001f00000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000002700000000000000430000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000800000000000000030000000000000003000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000100000000000000060000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "samplegold_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000001f000000000000001a0000000000000020000000000000000000000000",
            INIT_17 => X"00000017000000000000001f0000000000000010000000000000001200000000",
            INIT_18 => X"0000000b00000000000000120000000000000017000000000000001300000000",
            INIT_19 => X"000000180000000000000013000000000000000a000000000000000800000000",
            INIT_1A => X"0000000a000000000000001b000000000000001c000000000000001f00000000",
            INIT_1B => X"00000017000000000000000f0000000000000007000000000000001200000000",
            INIT_1C => X"000000320000000000000026000000000000001b000000000000001000000000",
            INIT_1D => X"00000017000000000000002a0000000000000037000000000000003800000000",
            INIT_1E => X"0000000700000000000000090000000000000000000000000000001700000000",
            INIT_1F => X"0000002f0000000000000012000000000000000d000000000000001400000000",
            INIT_20 => X"000000140000000000000024000000000000002f000000000000003b00000000",
            INIT_21 => X"00000026000000000000001d0000000000000000000000000000000700000000",
            INIT_22 => X"000000240000000000000016000000000000001c000000000000002700000000",
            INIT_23 => X"00000009000000000000000e000000000000001a000000000000002700000000",
            INIT_24 => X"0000001000000000000000130000000000000008000000000000001700000000",
            INIT_25 => X"0000003b00000000000000760000000000000069000000000000001000000000",
            INIT_26 => X"0000003d0000000000000030000000000000001a000000000000000b00000000",
            INIT_27 => X"0000000f00000000000000140000000000000017000000000000002000000000",
            INIT_28 => X"0000001c000000000000001b000000000000001d000000000000001600000000",
            INIT_29 => X"0000001400000000000000110000000000000033000000000000004600000000",
            INIT_2A => X"00000018000000000000001b0000000000000048000000000000003100000000",
            INIT_2B => X"0000001a0000000000000017000000000000001c000000000000002500000000",
            INIT_2C => X"0000001e0000000000000008000000000000000b000000000000001300000000",
            INIT_2D => X"0000000b000000000000002c0000000000000027000000000000001d00000000",
            INIT_2E => X"0000002f000000000000001d000000000000000e000000000000000600000000",
            INIT_2F => X"0000000b000000000000001e0000000000000016000000000000002300000000",
            INIT_30 => X"0000003f00000000000000350000000000000000000000000000000000000000",
            INIT_31 => X"0000005200000000000000480000000000000024000000000000002b00000000",
            INIT_32 => X"0000002500000000000000330000000000000026000000000000002800000000",
            INIT_33 => X"000000120000000000000015000000000000001c000000000000001a00000000",
            INIT_34 => X"0000008b0000000000000065000000000000004a000000000000001500000000",
            INIT_35 => X"0000002a0000000000000030000000000000004b000000000000006100000000",
            INIT_36 => X"0000002800000000000000240000000000000028000000000000002100000000",
            INIT_37 => X"00000000000000000000000b0000000000000024000000000000002000000000",
            INIT_38 => X"000000080000000000000020000000000000008100000000000000a000000000",
            INIT_39 => X"0000001400000000000000180000000000000003000000000000000c00000000",
            INIT_3A => X"0000001e000000000000002a000000000000002b000000000000002e00000000",
            INIT_3B => X"0000004d00000000000000000000000000000000000000000000001b00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_3D => X"0000001e00000000000000000000000000000001000000000000000000000000",
            INIT_3E => X"0000001600000000000000190000000000000011000000000000001a00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000f0000000000000008000000000000001b000000000000000500000000",
            INIT_41 => X"0000002200000000000000110000000000000014000000000000002f00000000",
            INIT_42 => X"0000000600000000000000060000000000000025000000000000003200000000",
            INIT_43 => X"0000000a00000000000000020000000000000000000000000000000000000000",
            INIT_44 => X"0000000d00000000000000220000000000000019000000000000001b00000000",
            INIT_45 => X"0000003a000000000000003e0000000000000029000000000000001100000000",
            INIT_46 => X"0000000100000000000000000000000000000011000000000000001900000000",
            INIT_47 => X"000000000000000000000000000000000000001a000000000000001400000000",
            INIT_48 => X"000000090000000000000018000000000000000a000000000000000000000000",
            INIT_49 => X"0000001200000000000000000000000000000001000000000000000700000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000c000000000000000b0000000000000000000000000000000000000000",
            INIT_4F => X"000000250000000000000020000000000000000f000000000000000b00000000",
            INIT_50 => X"000000080000000000000008000000000000000b000000000000001f00000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_52 => X"0000000c000000000000000b000000000000000a000000000000000000000000",
            INIT_53 => X"000000320000000000000035000000000000002a000000000000001500000000",
            INIT_54 => X"00000012000000000000000d0000000000000012000000000000002e00000000",
            INIT_55 => X"0000001000000000000000100000000000000010000000000000001100000000",
            INIT_56 => X"0000000c000000000000000f0000000000000008000000000000000a00000000",
            INIT_57 => X"0000004c000000000000004a000000000000003e000000000000003100000000",
            INIT_58 => X"000000230000000000000023000000000000001f000000000000002c00000000",
            INIT_59 => X"0000000b00000000000000140000000000000016000000000000001c00000000",
            INIT_5A => X"0000003400000000000000260000000000000012000000000000000d00000000",
            INIT_5B => X"000000550000000000000059000000000000004b000000000000004200000000",
            INIT_5C => X"000000180000000000000030000000000000002d000000000000003500000000",
            INIT_5D => X"00000027000000000000001e000000000000001c000000000000001800000000",
            INIT_5E => X"0000003200000000000000350000000000000029000000000000003300000000",
            INIT_5F => X"0000005a000000000000005d000000000000005b000000000000004800000000",
            INIT_60 => X"00000031000000000000002e000000000000003f000000000000005000000000",
            INIT_61 => X"0000002c0000000000000030000000000000002e000000000000003300000000",
            INIT_62 => X"0000004f0000000000000040000000000000002c000000000000002a00000000",
            INIT_63 => X"0000005e000000000000005f0000000000000051000000000000004b00000000",
            INIT_64 => X"00000034000000000000003a000000000000003f000000000000004d00000000",
            INIT_65 => X"0000002c00000000000000260000000000000027000000000000002600000000",
            INIT_66 => X"0000004e0000000000000045000000000000002e000000000000002800000000",
            INIT_67 => X"0000005100000000000000590000000000000051000000000000004a00000000",
            INIT_68 => X"000000270000000000000020000000000000002b000000000000004400000000",
            INIT_69 => X"00000039000000000000002c0000000000000036000000000000002d00000000",
            INIT_6A => X"0000004b0000000000000053000000000000004d000000000000003700000000",
            INIT_6B => X"0000003e00000000000000540000000000000057000000000000004e00000000",
            INIT_6C => X"0000003a00000000000000330000000000000021000000000000002f00000000",
            INIT_6D => X"000000460000000000000041000000000000005f000000000000004600000000",
            INIT_6E => X"0000004a000000000000004a000000000000005d000000000000003900000000",
            INIT_6F => X"0000003700000000000000440000000000000055000000000000005300000000",
            INIT_70 => X"000000510000000000000051000000000000004b000000000000002b00000000",
            INIT_71 => X"000000470000000000000044000000000000004c000000000000003e00000000",
            INIT_72 => X"00000052000000000000004a000000000000004b000000000000005600000000",
            INIT_73 => X"0000002000000000000000330000000000000047000000000000005800000000",
            INIT_74 => X"0000003b000000000000004d000000000000004e000000000000004d00000000",
            INIT_75 => X"00000040000000000000003f0000000000000042000000000000003b00000000",
            INIT_76 => X"000000520000000000000050000000000000004d000000000000004d00000000",
            INIT_77 => X"0000002f00000000000000310000000000000030000000000000004600000000",
            INIT_78 => X"0000003a00000000000000280000000000000017000000000000002300000000",
            INIT_79 => X"000000360000000000000034000000000000002f000000000000003a00000000",
            INIT_7A => X"00000048000000000000004f0000000000000043000000000000004000000000",
            INIT_7B => X"0000001600000000000000160000000000000034000000000000003600000000",
            INIT_7C => X"0000002c00000000000000220000000000000021000000000000001a00000000",
            INIT_7D => X"0000003d00000000000000380000000000000031000000000000003700000000",
            INIT_7E => X"0000003d0000000000000048000000000000004e000000000000004300000000",
            INIT_7F => X"00000029000000000000001f0000000000000019000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "samplegold_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003200000000000000280000000000000024000000000000002800000000",
            INIT_01 => X"0000003000000000000000370000000000000038000000000000003800000000",
            INIT_02 => X"0000003500000000000000390000000000000047000000000000003f00000000",
            INIT_03 => X"0000002a00000000000000250000000000000022000000000000002000000000",
            INIT_04 => X"000000370000000000000034000000000000002e000000000000002b00000000",
            INIT_05 => X"0000003600000000000000330000000000000031000000000000003500000000",
            INIT_06 => X"00000000000000000000002e0000000000000035000000000000003500000000",
            INIT_07 => X"0000000800000000000000090000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000001400000000000000000000000000000009000000000000000200000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001500000000000000000000000000000003000000000000000000000000",
            INIT_0F => X"0000000800000000000000000000000000000002000000000000000c00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_1D => X"00000000000000000000000b0000000000000011000000000000000000000000",
            INIT_1E => X"0000000000000000000000280000000000000012000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000011000000000000000d0000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000021000000000000000200000000",
            INIT_29 => X"00000000000000000000002f0000000000000000000000000000002600000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_2B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000003a000000000000000c0000000000000000000000000000000000000000",
            INIT_2D => X"0000001800000000000000370000000000000038000000000000005200000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000000000000000000000000000000000007a000000000000008600000000",
            INIT_31 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_33 => X"0000002700000000000000000000000000000004000000000000000000000000",
            INIT_34 => X"000000000000000000000000000000000000000f000000000000002700000000",
            INIT_35 => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000210000000000000033000000000000001700000000",
            INIT_39 => X"0000002800000000000000050000000000000005000000000000000000000000",
            INIT_3A => X"0000000300000000000000070000000000000000000000000000003000000000",
            INIT_3B => X"0000001500000000000000310000000000000020000000000000000e00000000",
            INIT_3C => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_3D => X"0000001300000000000000000000000000000000000000000000000100000000",
            INIT_3E => X"000000020000000000000003000000000000000b000000000000002000000000",
            INIT_3F => X"0000000300000000000000000000000000000007000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_41 => X"0000000d00000000000000080000000000000006000000000000000900000000",
            INIT_42 => X"0000000000000000000000050000000000000000000000000000000800000000",
            INIT_43 => X"0000000400000000000000000000000000000000000000000000000800000000",
            INIT_44 => X"0000000700000000000000080000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000f000000000000000a0000000000000005000000000000000200000000",
            INIT_4A => X"0000001a00000000000000000000000000000000000000000000001300000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"00000008000000000000000c0000000000000001000000000000001300000000",
            INIT_4E => X"0000003700000000000000400000000000000000000000000000000000000000",
            INIT_4F => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000070000000000000007000000000000000000000000",
            INIT_52 => X"00000000000000000000003e0000000000000031000000000000000000000000",
            INIT_53 => X"00000000000000000000000c0000000000000005000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000010000000000000000100000000",
            INIT_56 => X"000000000000000000000000000000000000007d000000000000000000000000",
            INIT_57 => X"0000000900000000000000000000000000000000000000000000000b00000000",
            INIT_58 => X"0000000000000000000000070000000000000000000000000000000300000000",
            INIT_59 => X"0000001000000000000000000000000000000000000000000000001b00000000",
            INIT_5A => X"0000000f0000000000000000000000000000004e000000000000000000000000",
            INIT_5B => X"00000008000000000000000e0000000000000000000000000000000000000000",
            INIT_5C => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000004c00000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000001a0000000000000000000000000000004f000000000000000100000000",
            INIT_5F => X"0000000600000000000000030000000000000000000000000000000000000000",
            INIT_60 => X"000000000000000000000026000000000000000d000000000000000000000000",
            INIT_61 => X"0000000000000000000000590000000000000021000000000000000000000000",
            INIT_62 => X"0000000000000000000000260000000000000000000000000000002500000000",
            INIT_63 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_64 => X"000000250000000000000000000000000000000b000000000000002600000000",
            INIT_65 => X"00000000000000000000000a0000000000000000000000000000009b00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_67 => X"0000000000000000000000030000000000000006000000000000000200000000",
            INIT_68 => X"0000002a00000000000000160000000000000035000000000000002000000000",
            INIT_69 => X"0000000000000000000000000000000000000035000000000000000e00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_6B => X"000000320000000000000000000000000000001b000000000000000800000000",
            INIT_6C => X"0000000000000000000000000000000000000004000000000000000b00000000",
            INIT_6D => X"000000090000000000000000000000000000001d000000000000000f00000000",
            INIT_6E => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000007000000000000002400000000",
            INIT_70 => X"00000000000000000000001b0000000000000012000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_72 => X"0000001100000000000000010000000000000000000000000000000000000000",
            INIT_73 => X"0000001200000000000000190000000000000000000000000000000a00000000",
            INIT_74 => X"000000000000000000000000000000000000000e000000000000000300000000",
            INIT_75 => X"00000002000000000000000a0000000000000015000000000000001400000000",
            INIT_76 => X"00000009000000000000000f0000000000000000000000000000000000000000",
            INIT_77 => X"00000010000000000000000b000000000000000b000000000000000800000000",
            INIT_78 => X"0000001400000000000000130000000000000013000000000000001300000000",
            INIT_79 => X"0000000d000000000000000e000000000000000f000000000000001100000000",
            INIT_7A => X"000000150000000000000012000000000000000d000000000000000d00000000",
            INIT_7B => X"0000000f0000000000000010000000000000000c000000000000000a00000000",
            INIT_7C => X"000000130000000000000012000000000000000b000000000000001400000000",
            INIT_7D => X"00000023000000000000001d0000000000000017000000000000001400000000",
            INIT_7E => X"0000000800000000000000280000000000000028000000000000002400000000",
            INIT_7F => X"0000000b000000000000000b0000000000000010000000000000000a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "samplegold_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001a0000000000000015000000000000000d000000000000000c00000000",
            INIT_01 => X"00000027000000000000002a0000000000000024000000000000002600000000",
            INIT_02 => X"0000000f000000000000000c0000000000000026000000000000002500000000",
            INIT_03 => X"0000000900000000000000000000000000000014000000000000002500000000",
            INIT_04 => X"00000014000000000000001e000000000000001b000000000000001100000000",
            INIT_05 => X"0000002b000000000000002b0000000000000024000000000000001c00000000",
            INIT_06 => X"00000032000000000000002a0000000000000024000000000000003200000000",
            INIT_07 => X"0000001300000000000000070000000000000000000000000000001800000000",
            INIT_08 => X"000000160000000000000018000000000000001a000000000000001800000000",
            INIT_09 => X"0000004700000000000000470000000000000035000000000000001b00000000",
            INIT_0A => X"0000001600000000000000260000000000000022000000000000002700000000",
            INIT_0B => X"000000090000000000000007000000000000000e000000000000001000000000",
            INIT_0C => X"0000000c00000000000000170000000000000019000000000000001300000000",
            INIT_0D => X"0000001a0000000000000045000000000000004c000000000000002f00000000",
            INIT_0E => X"0000001500000000000000330000000000000024000000000000001e00000000",
            INIT_0F => X"0000000f000000000000000d000000000000000a000000000000000400000000",
            INIT_10 => X"00000021000000000000000a0000000000000015000000000000001300000000",
            INIT_11 => X"00000028000000000000001e000000000000002c000000000000003100000000",
            INIT_12 => X"00000026000000000000003e000000000000002c000000000000002c00000000",
            INIT_13 => X"0000000c000000000000000a0000000000000018000000000000002600000000",
            INIT_14 => X"00000020000000000000000f000000000000000a000000000000001000000000",
            INIT_15 => X"0000004400000000000000330000000000000027000000000000003400000000",
            INIT_16 => X"00000033000000000000003e0000000000000038000000000000003a00000000",
            INIT_17 => X"0000000c00000000000000040000000000000001000000000000002100000000",
            INIT_18 => X"0000003d000000000000001d0000000000000006000000000000000800000000",
            INIT_19 => X"0000002f000000000000002b0000000000000041000000000000004200000000",
            INIT_1A => X"0000001f0000000000000024000000000000002e000000000000001a00000000",
            INIT_1B => X"00000007000000000000000c0000000000000002000000000000000100000000",
            INIT_1C => X"0000003500000000000000490000000000000028000000000000000200000000",
            INIT_1D => X"00000000000000000000000e000000000000001f000000000000003400000000",
            INIT_1E => X"0000000b000000000000000e0000000000000008000000000000000a00000000",
            INIT_1F => X"00000012000000000000000b0000000000000011000000000000000700000000",
            INIT_20 => X"00000009000000000000000a000000000000004d000000000000003e00000000",
            INIT_21 => X"0000000000000000000000130000000000000019000000000000001900000000",
            INIT_22 => X"000000010000000000000002000000000000001b000000000000000a00000000",
            INIT_23 => X"0000004100000000000000280000000000000015000000000000000f00000000",
            INIT_24 => X"0000001b000000000000000f000000000000000d000000000000005000000000",
            INIT_25 => X"0000001800000000000000230000000000000027000000000000002500000000",
            INIT_26 => X"0000000b00000000000000000000000000000007000000000000001600000000",
            INIT_27 => X"000000470000000000000045000000000000002d000000000000000c00000000",
            INIT_28 => X"0000002b00000000000000250000000000000024000000000000001c00000000",
            INIT_29 => X"00000024000000000000002a000000000000003b000000000000003500000000",
            INIT_2A => X"0000000500000000000000000000000000000007000000000000001800000000",
            INIT_2B => X"0000002600000000000000470000000000000045000000000000001b00000000",
            INIT_2C => X"000000470000000000000044000000000000003a000000000000002f00000000",
            INIT_2D => X"000000470000000000000045000000000000003a000000000000004300000000",
            INIT_2E => X"00000039000000000000002b000000000000002b000000000000003a00000000",
            INIT_2F => X"0000001c0000000000000021000000000000004f000000000000004c00000000",
            INIT_30 => X"0000001d000000000000001f0000000000000021000000000000002300000000",
            INIT_31 => X"0000000d000000000000000f0000000000000019000000000000001500000000",
            INIT_32 => X"0000000000000000000000000000000000000005000000000000000a00000000",
            INIT_33 => X"0000001d000000000000001a0000000000000020000000000000000000000000",
            INIT_34 => X"0000001600000000000000170000000000000011000000000000001400000000",
            INIT_35 => X"00000001000000000000000a000000000000000b000000000000000e00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000012000000000000000e000000000000001c000000000000001e00000000",
            INIT_38 => X"0000000200000000000000010000000000000000000000000000000700000000",
            INIT_39 => X"0000001000000000000000110000000000000011000000000000000c00000000",
            INIT_3A => X"000000180000000000000008000000000000000f000000000000000e00000000",
            INIT_3B => X"0000000100000000000000000000000000000000000000000000001800000000",
            INIT_3C => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000f0000000000000013000000000000001f000000000000001d00000000",
            INIT_3E => X"00000024000000000000001c0000000000000000000000000000000800000000",
            INIT_3F => X"0000001100000000000000000000000000000000000000000000001400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_41 => X"00000004000000000000000e0000000000000011000000000000000d00000000",
            INIT_42 => X"00000030000000000000004a0000000000000043000000000000000000000000",
            INIT_43 => X"0000001100000000000000110000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_45 => X"00000006000000000000000c000000000000000c000000000000000a00000000",
            INIT_46 => X"00000000000000000000003e0000000000000048000000000000004a00000000",
            INIT_47 => X"000000090000000000000012000000000000001f000000000000000000000000",
            INIT_48 => X"0000000200000000000000000000000000000000000000000000000c00000000",
            INIT_49 => X"00000042000000000000000b0000000000000012000000000000000800000000",
            INIT_4A => X"000000000000000000000033000000000000003b000000000000004000000000",
            INIT_4B => X"0000001700000000000000040000000000000000000000000000000000000000",
            INIT_4C => X"0000000900000000000000000000000000000000000000000000000c00000000",
            INIT_4D => X"0000004e00000000000000450000000000000003000000000000000b00000000",
            INIT_4E => X"00000010000000000000003b000000000000001b000000000000004500000000",
            INIT_4F => X"00000014000000000000001a0000000000000001000000000000001a00000000",
            INIT_50 => X"0000000200000000000000080000000000000000000000000000000200000000",
            INIT_51 => X"00000076000000000000006c0000000000000057000000000000000000000000",
            INIT_52 => X"000000220000000000000030000000000000004c000000000000005b00000000",
            INIT_53 => X"0000000d00000000000000170000000000000015000000000000000900000000",
            INIT_54 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_55 => X"0000003f0000000000000041000000000000007f000000000000008b00000000",
            INIT_56 => X"0000000f00000000000000160000000000000029000000000000002d00000000",
            INIT_57 => X"00000000000000000000000e0000000000000014000000000000001400000000",
            INIT_58 => X"0000008400000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000230000000000000036000000000000006f00000000",
            INIT_5A => X"0000000b0000000000000000000000000000000e000000000000000000000000",
            INIT_5B => X"000000000000000000000004000000000000000d000000000000000e00000000",
            INIT_5C => X"0000003600000000000000390000000000000000000000000000000100000000",
            INIT_5D => X"00000000000000000000000f0000000000000021000000000000002d00000000",
            INIT_5E => X"0000001800000000000000080000000000000007000000000000001000000000",
            INIT_5F => X"0000000000000000000000000000000000000010000000000000001a00000000",
            INIT_60 => X"0000001a0000000000000019000000000000001d000000000000000000000000",
            INIT_61 => X"0000000000000000000000030000000000000009000000000000001100000000",
            INIT_62 => X"00000026000000000000000e0000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_64 => X"0000000000000000000000000000000000000009000000000000000f00000000",
            INIT_65 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000200000000000000040000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "samplegold_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000f00000000000000050000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000000000000000000000c000000000000000c000000000000000900000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000008000000000000001400000000",
            INIT_19 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000a00000000000000000000000000000000000000000000001400000000",
            INIT_1D => X"0000000000000000000000010000000000000014000000000000001000000000",
            INIT_1E => X"0000000000000000000000060000000000000013000000000000001500000000",
            INIT_1F => X"0000001a00000000000000210000000000000011000000000000000400000000",
            INIT_20 => X"0000003700000000000000280000000000000000000000000000000000000000",
            INIT_21 => X"00000025000000000000002a000000000000002f000000000000002500000000",
            INIT_22 => X"0000001f000000000000000f0000000000000006000000000000000e00000000",
            INIT_23 => X"0000000000000000000000390000000000000036000000000000003300000000",
            INIT_24 => X"00000021000000000000004c0000000000000024000000000000000000000000",
            INIT_25 => X"0000004a000000000000003d0000000000000043000000000000002b00000000",
            INIT_26 => X"00000041000000000000003e0000000000000000000000000000003900000000",
            INIT_27 => X"0000000000000000000000000000000000000046000000000000004200000000",
            INIT_28 => X"000000460000000000000049000000000000002d000000000000000000000000",
            INIT_29 => X"00000031000000000000006b0000000000000058000000000000004500000000",
            INIT_2A => X"000000460000000000000052000000000000005b000000000000001100000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000004100000000",
            INIT_2C => X"00000008000000000000004c000000000000005d000000000000004c00000000",
            INIT_2D => X"00000056000000000000002e0000000000000015000000000000001100000000",
            INIT_2E => X"0000007200000000000000750000000000000066000000000000004d00000000",
            INIT_2F => X"00000049000000000000003c0000000000000003000000000000002100000000",
            INIT_30 => X"0000004800000000000000580000000000000065000000000000003100000000",
            INIT_31 => X"0000004e00000000000000510000000000000039000000000000002500000000",
            INIT_32 => X"000000500000000000000057000000000000006a000000000000007100000000",
            INIT_33 => X"0000003d00000000000000400000000000000058000000000000005100000000",
            INIT_34 => X"0000000a000000000000003c0000000000000062000000000000006700000000",
            INIT_35 => X"00000072000000000000005d000000000000004c000000000000002400000000",
            INIT_36 => X"000000530000000000000052000000000000003f000000000000005200000000",
            INIT_37 => X"000000470000000000000041000000000000003c000000000000006b00000000",
            INIT_38 => X"000000360000000000000033000000000000003c000000000000003f00000000",
            INIT_39 => X"0000005a00000000000000790000000000000059000000000000004600000000",
            INIT_3A => X"0000004b000000000000005a0000000000000058000000000000003c00000000",
            INIT_3B => X"0000005400000000000000530000000000000050000000000000003900000000",
            INIT_3C => X"0000005c000000000000004f0000000000000058000000000000003200000000",
            INIT_3D => X"0000006c0000000000000084000000000000009400000000000000a200000000",
            INIT_3E => X"0000004100000000000000360000000000000048000000000000004d00000000",
            INIT_3F => X"0000003b00000000000000390000000000000034000000000000005a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002300000000000000360000000000000053000000000000004000000000",
            INIT_41 => X"0000004b00000000000000720000000000000095000000000000006500000000",
            INIT_42 => X"00000066000000000000005b000000000000004c000000000000003900000000",
            INIT_43 => X"0000000d0000000000000045000000000000007b000000000000008700000000",
            INIT_44 => X"0000001d00000000000000380000000000000054000000000000002b00000000",
            INIT_45 => X"00000054000000000000005b0000000000000056000000000000003000000000",
            INIT_46 => X"0000005c00000000000000520000000000000052000000000000005300000000",
            INIT_47 => X"0000005000000000000000620000000000000074000000000000005c00000000",
            INIT_48 => X"00000049000000000000003a0000000000000024000000000000004400000000",
            INIT_49 => X"0000004b00000000000000550000000000000062000000000000003900000000",
            INIT_4A => X"0000003f0000000000000075000000000000006e000000000000006b00000000",
            INIT_4B => X"0000001c0000000000000051000000000000005a000000000000005900000000",
            INIT_4C => X"00000031000000000000003f0000000000000040000000000000004700000000",
            INIT_4D => X"0000006800000000000000540000000000000057000000000000005c00000000",
            INIT_4E => X"0000006a00000000000000570000000000000077000000000000006d00000000",
            INIT_4F => X"0000004600000000000000310000000000000048000000000000006800000000",
            INIT_50 => X"0000005e000000000000002d0000000000000050000000000000005300000000",
            INIT_51 => X"00000054000000000000005e000000000000004d000000000000004c00000000",
            INIT_52 => X"000000510000000000000058000000000000005a000000000000001e00000000",
            INIT_53 => X"0000003500000000000000340000000000000027000000000000004100000000",
            INIT_54 => X"0000003c0000000000000069000000000000002e000000000000002900000000",
            INIT_55 => X"0000005600000000000000610000000000000062000000000000004900000000",
            INIT_56 => X"00000019000000000000003b0000000000000046000000000000006300000000",
            INIT_57 => X"0000001d00000000000000240000000000000029000000000000002e00000000",
            INIT_58 => X"0000004900000000000000570000000000000019000000000000003f00000000",
            INIT_59 => X"0000004a000000000000004a000000000000003c000000000000004200000000",
            INIT_5A => X"0000004b000000000000001e000000000000002c000000000000004d00000000",
            INIT_5B => X"000000500000000000000051000000000000004e000000000000004500000000",
            INIT_5C => X"0000003f00000000000000460000000000000040000000000000001a00000000",
            INIT_5D => X"0000003c0000000000000037000000000000002e000000000000002200000000",
            INIT_5E => X"00000037000000000000005d0000000000000010000000000000003200000000",
            INIT_5F => X"0000001a00000000000000470000000000000045000000000000003f00000000",
            INIT_60 => X"0000002600000000000000420000000000000050000000000000002800000000",
            INIT_61 => X"000000220000000000000032000000000000001f000000000000000000000000",
            INIT_62 => X"0000002d000000000000002f000000000000003a000000000000002700000000",
            INIT_63 => X"0000004600000000000000200000000000000034000000000000003300000000",
            INIT_64 => X"00000009000000000000002a000000000000002b000000000000005500000000",
            INIT_65 => X"0000003e0000000000000026000000000000001a000000000000001b00000000",
            INIT_66 => X"0000001b00000000000000220000000000000037000000000000001f00000000",
            INIT_67 => X"000000320000000000000043000000000000002d000000000000002e00000000",
            INIT_68 => X"0000001200000000000000160000000000000036000000000000001900000000",
            INIT_69 => X"0000002f000000000000002f0000000000000022000000000000000b00000000",
            INIT_6A => X"0000004100000000000000230000000000000024000000000000003800000000",
            INIT_6B => X"0000002a000000000000002c0000000000000034000000000000002f00000000",
            INIT_6C => X"00000017000000000000000a0000000000000018000000000000002f00000000",
            INIT_6D => X"000000380000000000000029000000000000002a000000000000001e00000000",
            INIT_6E => X"00000035000000000000003d0000000000000022000000000000002500000000",
            INIT_6F => X"0000001b000000000000002f000000000000002a000000000000003600000000",
            INIT_70 => X"000000170000000000000023000000000000000e000000000000001d00000000",
            INIT_71 => X"0000002c0000000000000038000000000000002c000000000000001d00000000",
            INIT_72 => X"0000003600000000000000320000000000000030000000000000002500000000",
            INIT_73 => X"00000016000000000000001d0000000000000043000000000000001b00000000",
            INIT_74 => X"00000032000000000000001f000000000000001c000000000000000f00000000",
            INIT_75 => X"000000230000000000000035000000000000003f000000000000002200000000",
            INIT_76 => X"0000002500000000000000340000000000000023000000000000003100000000",
            INIT_77 => X"0000001400000000000000180000000000000018000000000000003e00000000",
            INIT_78 => X"0000002800000000000000280000000000000042000000000000000200000000",
            INIT_79 => X"0000004600000000000000270000000000000048000000000000002700000000",
            INIT_7A => X"0000001f000000000000002b0000000000000036000000000000002a00000000",
            INIT_7B => X"0000001300000000000000110000000000000019000000000000002300000000",
            INIT_7C => X"0000003500000000000000240000000000000035000000000000001e00000000",
            INIT_7D => X"0000002b000000000000003a0000000000000030000000000000003c00000000",
            INIT_7E => X"000000250000000000000026000000000000002c000000000000002200000000",
            INIT_7F => X"000000150000000000000022000000000000002a000000000000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "samplegold_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000000000380000000000000032000000000000002100000000",
            INIT_01 => X"0000001d000000000000002f0000000000000031000000000000002400000000",
            INIT_02 => X"0000001a000000000000001a000000000000001e000000000000003800000000",
            INIT_03 => X"0000001b00000000000000210000000000000027000000000000003200000000",
            INIT_04 => X"00000029000000000000002c000000000000002c000000000000004100000000",
            INIT_05 => X"0000003b000000000000002e000000000000002d000000000000002800000000",
            INIT_06 => X"00000031000000000000002e0000000000000005000000000000001c00000000",
            INIT_07 => X"0000003800000000000000250000000000000021000000000000002a00000000",
            INIT_08 => X"0000002b0000000000000029000000000000002b000000000000002b00000000",
            INIT_09 => X"0000002200000000000000420000000000000032000000000000002d00000000",
            INIT_0A => X"0000002c000000000000002c0000000000000036000000000000001600000000",
            INIT_0B => X"0000002d0000000000000034000000000000002f000000000000002a00000000",
            INIT_0C => X"0000002d00000000000000310000000000000038000000000000002700000000",
            INIT_0D => X"0000001a00000000000000230000000000000040000000000000003200000000",
            INIT_0E => X"0000002400000000000000300000000000000024000000000000002100000000",
            INIT_0F => X"0000002c00000000000000310000000000000031000000000000003b00000000",
            INIT_10 => X"000000000000000000000000000000000000002f000000000000003700000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000700000000000000070000000000000019000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000000e000000000000000400000000",
            INIT_17 => X"00000009000000000000000c0000000000000012000000000000001900000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000070000000000000000000000000000001f000000000000002b00000000",
            INIT_1A => X"0000002600000000000000120000000000000003000000000000000b00000000",
            INIT_1B => X"0000000000000000000000210000000000000029000000000000002b00000000",
            INIT_1C => X"0000002100000000000000040000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000004000000000000003100000000",
            INIT_1E => X"0000003e000000000000002a0000000000000029000000000000000100000000",
            INIT_1F => X"00000000000000000000000e0000000000000029000000000000003600000000",
            INIT_20 => X"0000003200000000000000130000000000000004000000000000001700000000",
            INIT_21 => X"000000030000000000000000000000000000000b000000000000002900000000",
            INIT_22 => X"00000023000000000000003f000000000000002b000000000000002400000000",
            INIT_23 => X"0000001c0000000000000018000000000000001c000000000000001000000000",
            INIT_24 => X"0000001f000000000000002a0000000000000019000000000000000600000000",
            INIT_25 => X"0000001c00000000000000060000000000000005000000000000000800000000",
            INIT_26 => X"0000000a00000000000000260000000000000040000000000000003600000000",
            INIT_27 => X"00000012000000000000000d0000000000000012000000000000001700000000",
            INIT_28 => X"0000000e00000000000000230000000000000022000000000000001500000000",
            INIT_29 => X"0000002e000000000000001c0000000000000012000000000000001b00000000",
            INIT_2A => X"0000001a000000000000001a000000000000003b000000000000003f00000000",
            INIT_2B => X"0000002a000000000000001e0000000000000006000000000000001000000000",
            INIT_2C => X"000000150000000000000009000000000000002b000000000000001e00000000",
            INIT_2D => X"0000002c00000000000000200000000000000013000000000000000e00000000",
            INIT_2E => X"0000000b00000000000000190000000000000028000000000000003e00000000",
            INIT_2F => X"000000300000000000000033000000000000001a000000000000001d00000000",
            INIT_30 => X"0000000100000000000000000000000000000022000000000000002800000000",
            INIT_31 => X"00000023000000000000000a0000000000000000000000000000001300000000",
            INIT_32 => X"00000022000000000000000f0000000000000023000000000000001b00000000",
            INIT_33 => X"0000003a000000000000003b000000000000002b000000000000002600000000",
            INIT_34 => X"0000000a000000000000000d0000000000000001000000000000002a00000000",
            INIT_35 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_36 => X"000000290000000000000025000000000000001c000000000000002a00000000",
            INIT_37 => X"0000002c0000000000000021000000000000001f000000000000002e00000000",
            INIT_38 => X"000000020000000000000000000000000000000d000000000000002d00000000",
            INIT_39 => X"0000002700000000000000000000000000000009000000000000000a00000000",
            INIT_3A => X"00000034000000000000003a000000000000001e000000000000001f00000000",
            INIT_3B => X"0000001f00000000000000200000000000000019000000000000002400000000",
            INIT_3C => X"0000001100000000000000070000000000000000000000000000000600000000",
            INIT_3D => X"0000001700000000000000220000000000000000000000000000000500000000",
            INIT_3E => X"00000005000000000000002c0000000000000034000000000000001300000000",
            INIT_3F => X"0000000000000000000000150000000000000018000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000100000000000000070000000000000001000000000000000000000000",
            INIT_41 => X"00000006000000000000000a000000000000001d000000000000000000000000",
            INIT_42 => X"0000000e0000000000000003000000000000002d000000000000003300000000",
            INIT_43 => X"0000000000000000000000000000000000000002000000000000000600000000",
            INIT_44 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000002d00000000000000000000000000000005000000000000001000000000",
            INIT_46 => X"000000000000000000000004000000000000001e000000000000002d00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000006f000000000000007b000000000000007f000000000000001400000000",
            INIT_4A => X"0000007e00000000000000790000000000000071000000000000006e00000000",
            INIT_4B => X"0000009000000000000000930000000000000067000000000000003600000000",
            INIT_4C => X"0000000200000000000000000000000000000089000000000000008d00000000",
            INIT_4D => X"0000007d00000000000000ad0000000000000089000000000000006c00000000",
            INIT_4E => X"0000007100000000000000a500000000000000a0000000000000009000000000",
            INIT_4F => X"000000a300000000000000ab00000000000000bb000000000000008100000000",
            INIT_50 => X"0000005000000000000000000000000000000000000000000000009e00000000",
            INIT_51 => X"0000006900000000000000a900000000000000d8000000000000007a00000000",
            INIT_52 => X"000000a7000000000000008e000000000000008b000000000000007a00000000",
            INIT_53 => X"000000c200000000000000cb00000000000000d000000000000000cd00000000",
            INIT_54 => X"00000086000000000000006c0000000000000029000000000000001d00000000",
            INIT_55 => X"00000067000000000000008e00000000000000d300000000000000d200000000",
            INIT_56 => X"000000e500000000000000d3000000000000008d000000000000006300000000",
            INIT_57 => X"000000a500000000000000e100000000000000e500000000000000fb00000000",
            INIT_58 => X"000000ac000000000000008300000000000000ba000000000000009800000000",
            INIT_59 => X"00000072000000000000008400000000000000c000000000000000d600000000",
            INIT_5A => X"000000fd00000000000000ef00000000000000c6000000000000008d00000000",
            INIT_5B => X"000000be00000000000000c200000000000000b500000000000000c700000000",
            INIT_5C => X"000000ca00000000000000b6000000000000009b00000000000000c000000000",
            INIT_5D => X"000000940000000000000085000000000000008200000000000000b600000000",
            INIT_5E => X"000000cf000000000000010300000000000000f300000000000000b700000000",
            INIT_5F => X"0000009a00000000000000b700000000000000bb000000000000009f00000000",
            INIT_60 => X"000000a500000000000000b300000000000000a900000000000000b800000000",
            INIT_61 => X"000000b700000000000000a700000000000000a9000000000000009800000000",
            INIT_62 => X"000000bc00000000000000fd000000000000010700000000000000f100000000",
            INIT_63 => X"000000ba000000000000009300000000000000b500000000000000b700000000",
            INIT_64 => X"0000009800000000000000bc00000000000000c500000000000000c600000000",
            INIT_65 => X"000000af00000000000000b8000000000000009c00000000000000b700000000",
            INIT_66 => X"000000b500000000000000e900000000000000fa000000000000010900000000",
            INIT_67 => X"000000ea00000000000000b300000000000000b0000000000000009c00000000",
            INIT_68 => X"0000007600000000000000a400000000000000c600000000000000e100000000",
            INIT_69 => X"00000082000000000000006f00000000000000a4000000000000009900000000",
            INIT_6A => X"000000ab00000000000000ca00000000000000d200000000000000c200000000",
            INIT_6B => X"000000e400000000000000d000000000000000cd00000000000000ca00000000",
            INIT_6C => X"00000098000000000000008a00000000000000d300000000000000f500000000",
            INIT_6D => X"0000008700000000000000810000000000000083000000000000008d00000000",
            INIT_6E => X"000000d500000000000000b900000000000000db000000000000008d00000000",
            INIT_6F => X"000000c000000000000000bd00000000000000da00000000000000d600000000",
            INIT_70 => X"00000084000000000000008f00000000000000cf00000000000000d600000000",
            INIT_71 => X"00000075000000000000008a000000000000009a000000000000008600000000",
            INIT_72 => X"000000ed00000000000000ca00000000000000bf00000000000000d500000000",
            INIT_73 => X"000000c800000000000000c000000000000000c000000000000000e300000000",
            INIT_74 => X"000000900000000000000078000000000000008500000000000000bd00000000",
            INIT_75 => X"000000ca0000000000000078000000000000008d00000000000000a500000000",
            INIT_76 => X"000000c400000000000000ea00000000000000c000000000000000b200000000",
            INIT_77 => X"000000a500000000000000b600000000000000be000000000000008b00000000",
            INIT_78 => X"000000850000000000000083000000000000007d000000000000007700000000",
            INIT_79 => X"0000009e00000000000000c10000000000000078000000000000008900000000",
            INIT_7A => X"0000009800000000000000c700000000000000e700000000000000a500000000",
            INIT_7B => X"00000062000000000000007c0000000000000091000000000000009e00000000",
            INIT_7C => X"0000006b00000000000000680000000000000075000000000000006e00000000",
            INIT_7D => X"00000086000000000000009800000000000000a8000000000000008400000000",
            INIT_7E => X"0000008100000000000000b100000000000000d500000000000000e600000000",
            INIT_7F => X"000000680000000000000056000000000000005d000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "samplegold_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007c0000000000000065000000000000006b000000000000007300000000",
            INIT_01 => X"0000004700000000000000400000000000000000000000000000001500000000",
            INIT_02 => X"0000003e00000000000000450000000000000046000000000000003c00000000",
            INIT_03 => X"000000270000000000000008000000000000002e000000000000002f00000000",
            INIT_04 => X"0000001500000000000000480000000000000044000000000000003c00000000",
            INIT_05 => X"00000017000000000000003f000000000000003f000000000000000900000000",
            INIT_06 => X"00000046000000000000003d0000000000000040000000000000002e00000000",
            INIT_07 => X"0000004500000000000000400000000000000000000000000000005100000000",
            INIT_08 => X"000000130000000000000015000000000000004a000000000000004700000000",
            INIT_09 => X"000000430000000000000019000000000000002e000000000000001a00000000",
            INIT_0A => X"00000031000000000000006c0000000000000055000000000000004600000000",
            INIT_0B => X"0000003d00000000000000480000000000000051000000000000001100000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_0D => X"0000000f0000000000000032000000000000002d000000000000005700000000",
            INIT_0E => X"00000046000000000000000f0000000000000020000000000000002400000000",
            INIT_0F => X"0000005d000000000000005c0000000000000035000000000000002e00000000",
            INIT_10 => X"0000006200000000000000460000000000000010000000000000003d00000000",
            INIT_11 => X"0000004c000000000000003f000000000000003a000000000000001400000000",
            INIT_12 => X"0000003d0000000000000038000000000000001f000000000000002800000000",
            INIT_13 => X"000000570000000000000064000000000000007b000000000000005600000000",
            INIT_14 => X"00000021000000000000004e0000000000000062000000000000004d00000000",
            INIT_15 => X"00000013000000000000003a0000000000000054000000000000003c00000000",
            INIT_16 => X"0000006100000000000000470000000000000034000000000000001100000000",
            INIT_17 => X"000000560000000000000065000000000000006b000000000000007500000000",
            INIT_18 => X"0000002f000000000000003f0000000000000047000000000000006d00000000",
            INIT_19 => X"00000028000000000000002b0000000000000019000000000000003800000000",
            INIT_1A => X"0000005900000000000000600000000000000040000000000000002c00000000",
            INIT_1B => X"000000530000000000000058000000000000006e000000000000005500000000",
            INIT_1C => X"00000038000000000000003c0000000000000037000000000000001a00000000",
            INIT_1D => X"0000005300000000000000350000000000000047000000000000002200000000",
            INIT_1E => X"0000006800000000000000760000000000000079000000000000007500000000",
            INIT_1F => X"0000001500000000000000280000000000000053000000000000007600000000",
            INIT_20 => X"0000003d000000000000001c0000000000000018000000000000003a00000000",
            INIT_21 => X"00000048000000000000003b0000000000000050000000000000002900000000",
            INIT_22 => X"0000006700000000000000640000000000000092000000000000005700000000",
            INIT_23 => X"0000004900000000000000420000000000000038000000000000004100000000",
            INIT_24 => X"0000001e000000000000002c000000000000004a000000000000005800000000",
            INIT_25 => X"0000002200000000000000430000000000000055000000000000002700000000",
            INIT_26 => X"0000006200000000000000630000000000000058000000000000003900000000",
            INIT_27 => X"0000005400000000000000390000000000000038000000000000003f00000000",
            INIT_28 => X"00000052000000000000004d0000000000000048000000000000004000000000",
            INIT_29 => X"0000004b00000000000000330000000000000027000000000000004c00000000",
            INIT_2A => X"0000003500000000000000720000000000000066000000000000003f00000000",
            INIT_2B => X"0000002e000000000000004d0000000000000048000000000000003f00000000",
            INIT_2C => X"00000024000000000000005e0000000000000048000000000000003b00000000",
            INIT_2D => X"0000004200000000000000410000000000000038000000000000004300000000",
            INIT_2E => X"00000047000000000000004f000000000000007a000000000000006900000000",
            INIT_2F => X"0000005500000000000000410000000000000043000000000000006100000000",
            INIT_30 => X"0000004600000000000000390000000000000053000000000000006100000000",
            INIT_31 => X"0000006f000000000000003b0000000000000051000000000000004c00000000",
            INIT_32 => X"000000490000000000000043000000000000005c000000000000007d00000000",
            INIT_33 => X"0000005a0000000000000059000000000000004e000000000000000900000000",
            INIT_34 => X"00000046000000000000003f0000000000000036000000000000004f00000000",
            INIT_35 => X"00000073000000000000007f0000000000000035000000000000003200000000",
            INIT_36 => X"0000004f000000000000004b0000000000000043000000000000005e00000000",
            INIT_37 => X"000000320000000000000055000000000000004f000000000000006400000000",
            INIT_38 => X"0000002a00000000000000380000000000000038000000000000003e00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_42 => X"0000002f00000000000000220000000000000002000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_56 => X"00000000000000000000001a000000000000004b000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000d0000000000000038000000000000001c000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_5D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_69 => X"00000000000000000000000b000000000000000e000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_6D => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"00000003000000000000000e0000000000000011000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"000000b100000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000d00000000000000000000000000000000000000000000003400000000",
            INIT_73 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000004000000000000009400000000",
            INIT_75 => X"0000006900000000000000680000000000000000000000000000000000000000",
            INIT_76 => X"0000001000000000000000000000000000000000000000000000002100000000",
            INIT_77 => X"000000b500000000000000000000000000000000000000000000001400000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000002100000000000000a30000000000000021000000000000000000000000",
            INIT_7A => X"0000001f00000000000000000000000000000000000000000000003600000000",
            INIT_7B => X"00000013000000000000003e0000000000000017000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000005d00000000000000000000000000000062000000000000004300000000",
            INIT_7E => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000490000000000000000000000000000006900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "samplegold_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000330000000000000000000000000000001b000000000000000000000000",
            INIT_01 => X"0000000000000000000000620000000000000000000000000000000000000000",
            INIT_02 => X"0000004600000000000000100000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000045000000000000002300000000",
            INIT_04 => X"0000000000000000000000040000000000000000000000000000002600000000",
            INIT_05 => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_06 => X"0000001f00000000000000360000000000000003000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000005600000000",
            INIT_08 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000230000000000000000000000000000000a000000000000000000000000",
            INIT_0A => X"00000050000000000000001b000000000000001c000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000740000000000000000000000000000000800000000",
            INIT_0D => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000004c000000000000003a0000000000000000000000000000000400000000",
            INIT_0F => X"0000000800000000000000000000000000000008000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000030000000000000000000000000",
            INIT_11 => X"00000000000000000000003b0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000560000000000000000000000000000000000000000",
            INIT_13 => X"0000000500000000000000000000000000000000000000000000005c00000000",
            INIT_14 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_15 => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_16 => X"000000260000000000000000000000000000000f000000000000000400000000",
            INIT_17 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_18 => X"00000008000000000000002c0000000000000000000000000000000000000000",
            INIT_19 => X"0000000e00000000000000040000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_1B => X"000000000000000000000000000000000000004a000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_1D => X"0000000c00000000000000000000000000000038000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000600000000000000000000000000000000000000000000003e00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_22 => X"0000004300000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000040000000000000000000000000000000f00000000",
            INIT_24 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000400000000000000280000000000000000000000000000000000000000",
            INIT_26 => X"0000003500000000000000270000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000300000000000000040000000000000027000000000000000000000000",
            INIT_29 => X"000000290000000000000006000000000000000e000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000006000000000000000a00000000",
            INIT_2D => X"0000000700000000000000280000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_2F => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_31 => X"0000000000000000000000160000000000000025000000000000000000000000",
            INIT_32 => X"0000000000000000000000120000000000000014000000000000000000000000",
            INIT_33 => X"0000000d000000000000000b0000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000021000000000000005e000000000000005b00000000",
            INIT_36 => X"0000001300000000000000310000000000000020000000000000000000000000",
            INIT_37 => X"0000000200000000000000000000000000000006000000000000000c00000000",
            INIT_38 => X"0000001100000000000000000000000000000000000000000000000900000000",
            INIT_39 => X"0000000900000000000000000000000000000000000000000000001200000000",
            INIT_3A => X"0000000900000000000000000000000000000004000000000000000500000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_3E => X"000000190000000000000023000000000000000f000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000f000000000000000f0000000000000003000000000000000000000000",
            INIT_42 => X"0000000a000000000000000f000000000000001d000000000000001100000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000f00000000000000140000000000000006000000000000000c00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000001100000000000000040000000000000007000000000000000000000000",
            INIT_49 => X"0000000000000000000000150000000000000025000000000000002700000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000180000000000000026000000000000000200000000",
            INIT_4E => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000002000000000000000400000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000001100000000000000070000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60 : if BRAM_NAME = "samplegold_layersamples_instance60" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000001a00000000000000250000000000000005000000000000000000000000",
            INIT_1B => X"0000001f000000000000001b0000000000000019000000000000001900000000",
            INIT_1C => X"000000430000000000000013000000000000003d000000000000002b00000000",
            INIT_1D => X"00000021000000000000002a000000000000002d000000000000003e00000000",
            INIT_1E => X"0000001d000000000000000a0000000000000014000000000000000700000000",
            INIT_1F => X"00000030000000000000001b0000000000000027000000000000004900000000",
            INIT_20 => X"00000041000000000000007f0000000000000003000000000000001e00000000",
            INIT_21 => X"000000070000000000000023000000000000002c000000000000003500000000",
            INIT_22 => X"000000460000000000000035000000000000002e000000000000000800000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_24 => X"0000003e00000000000000370000000000000065000000000000003400000000",
            INIT_25 => X"0000008c000000000000006d0000000000000048000000000000004800000000",
            INIT_26 => X"0000003800000000000000300000000000000010000000000000009400000000",
            INIT_27 => X"000000420000000000000026000000000000002b000000000000005000000000",
            INIT_28 => X"00000028000000000000004d000000000000005a000000000000002f00000000",
            INIT_29 => X"0000003e00000000000000780000000000000049000000000000003400000000",
            INIT_2A => X"00000021000000000000002b0000000000000046000000000000001200000000",
            INIT_2B => X"0000003900000000000000330000000000000020000000000000000700000000",
            INIT_2C => X"00000032000000000000001f0000000000000046000000000000005f00000000",
            INIT_2D => X"0000002800000000000000280000000000000039000000000000003800000000",
            INIT_2E => X"0000001800000000000000070000000000000024000000000000004400000000",
            INIT_2F => X"0000005200000000000000380000000000000046000000000000004000000000",
            INIT_30 => X"00000033000000000000003a0000000000000039000000000000004700000000",
            INIT_31 => X"0000002f00000000000000310000000000000000000000000000003300000000",
            INIT_32 => X"00000031000000000000003d000000000000001f000000000000003600000000",
            INIT_33 => X"000000460000000000000053000000000000003e000000000000004100000000",
            INIT_34 => X"0000002600000000000000270000000000000053000000000000005100000000",
            INIT_35 => X"0000003000000000000000360000000000000047000000000000000000000000",
            INIT_36 => X"0000002900000000000000210000000000000027000000000000002900000000",
            INIT_37 => X"0000002800000000000000210000000000000000000000000000001300000000",
            INIT_38 => X"00000034000000000000002a000000000000002b000000000000004500000000",
            INIT_39 => X"0000005200000000000000670000000000000045000000000000004600000000",
            INIT_3A => X"0000002700000000000000170000000000000023000000000000001d00000000",
            INIT_3B => X"0000002e00000000000000000000000000000000000000000000002300000000",
            INIT_3C => X"0000003c0000000000000039000000000000004a000000000000003d00000000",
            INIT_3D => X"00000046000000000000002a0000000000000013000000000000002e00000000",
            INIT_3E => X"000000150000000000000000000000000000003a000000000000004d00000000",
            INIT_3F => X"0000003f000000000000000c0000000000000023000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000490000000000000043000000000000003f000000000000002d00000000",
            INIT_41 => X"0000001e0000000000000024000000000000002a000000000000001c00000000",
            INIT_42 => X"0000002a0000000000000033000000000000000f000000000000000300000000",
            INIT_43 => X"0000002800000000000000380000000000000010000000000000000e00000000",
            INIT_44 => X"0000001400000000000000290000000000000039000000000000004a00000000",
            INIT_45 => X"00000000000000000000001e0000000000000033000000000000003f00000000",
            INIT_46 => X"0000001900000000000000260000000000000018000000000000003700000000",
            INIT_47 => X"0000004100000000000000200000000000000034000000000000001500000000",
            INIT_48 => X"0000002100000000000000000000000000000003000000000000003700000000",
            INIT_49 => X"0000001d00000000000000020000000000000000000000000000001200000000",
            INIT_4A => X"0000001d00000000000000050000000000000000000000000000001200000000",
            INIT_4B => X"0000003f0000000000000039000000000000001c000000000000002a00000000",
            INIT_4C => X"00000004000000000000000a0000000000000052000000000000002500000000",
            INIT_4D => X"00000016000000000000001c0000000000000000000000000000000000000000",
            INIT_4E => X"0000000e0000000000000023000000000000001d000000000000000500000000",
            INIT_4F => X"0000002f0000000000000034000000000000002a000000000000002600000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_51 => X"0000001b00000000000000190000000000000011000000000000001b00000000",
            INIT_52 => X"0000000b0000000000000000000000000000000e000000000000002300000000",
            INIT_53 => X"00000053000000000000004d000000000000004e000000000000004b00000000",
            INIT_54 => X"0000003900000000000000480000000000000056000000000000005d00000000",
            INIT_55 => X"0000006d000000000000006c0000000000000061000000000000001600000000",
            INIT_56 => X"0000003900000000000000000000000000000000000000000000006d00000000",
            INIT_57 => X"0000003d000000000000004a000000000000002f000000000000003a00000000",
            INIT_58 => X"0000002d00000000000000350000000000000051000000000000004b00000000",
            INIT_59 => X"0000006b000000000000006a0000000000000069000000000000005f00000000",
            INIT_5A => X"0000004700000000000000280000000000000000000000000000000000000000",
            INIT_5B => X"0000003100000000000000310000000000000039000000000000002500000000",
            INIT_5C => X"0000004e0000000000000046000000000000001f000000000000003000000000",
            INIT_5D => X"00000037000000000000005d0000000000000059000000000000005500000000",
            INIT_5E => X"0000001f000000000000004d0000000000000048000000000000001500000000",
            INIT_5F => X"0000002400000000000000330000000000000039000000000000003200000000",
            INIT_60 => X"000000540000000000000043000000000000003e000000000000002700000000",
            INIT_61 => X"00000049000000000000004d000000000000004b000000000000005600000000",
            INIT_62 => X"000000340000000000000029000000000000004c000000000000005400000000",
            INIT_63 => X"00000022000000000000001b000000000000002f000000000000003900000000",
            INIT_64 => X"00000067000000000000005e0000000000000054000000000000003c00000000",
            INIT_65 => X"0000005500000000000000510000000000000054000000000000005800000000",
            INIT_66 => X"0000003700000000000000350000000000000033000000000000004800000000",
            INIT_67 => X"0000003b00000000000000240000000000000022000000000000002500000000",
            INIT_68 => X"0000006300000000000000690000000000000062000000000000004e00000000",
            INIT_69 => X"0000003a000000000000005e0000000000000057000000000000006100000000",
            INIT_6A => X"0000001b0000000000000035000000000000002e000000000000004000000000",
            INIT_6B => X"0000005200000000000000380000000000000027000000000000003400000000",
            INIT_6C => X"0000006000000000000000690000000000000061000000000000006100000000",
            INIT_6D => X"000000440000000000000035000000000000004f000000000000004e00000000",
            INIT_6E => X"0000002400000000000000330000000000000027000000000000003300000000",
            INIT_6F => X"000000450000000000000048000000000000003c000000000000004000000000",
            INIT_70 => X"00000049000000000000005f0000000000000054000000000000006300000000",
            INIT_71 => X"000000400000000000000036000000000000004c000000000000004100000000",
            INIT_72 => X"0000003d000000000000003e0000000000000039000000000000003f00000000",
            INIT_73 => X"0000004500000000000000480000000000000046000000000000003d00000000",
            INIT_74 => X"000000470000000000000050000000000000005e000000000000004b00000000",
            INIT_75 => X"0000002d000000000000003d0000000000000047000000000000004200000000",
            INIT_76 => X"0000004b0000000000000038000000000000004c000000000000003a00000000",
            INIT_77 => X"0000004b000000000000004a000000000000003e000000000000003e00000000",
            INIT_78 => X"00000050000000000000003b0000000000000054000000000000005a00000000",
            INIT_79 => X"0000003c000000000000003a000000000000004c000000000000004a00000000",
            INIT_7A => X"000000400000000000000031000000000000004e000000000000003e00000000",
            INIT_7B => X"0000005b000000000000003b0000000000000041000000000000003e00000000",
            INIT_7C => X"0000004c0000000000000045000000000000003f000000000000005400000000",
            INIT_7D => X"0000004800000000000000450000000000000046000000000000004200000000",
            INIT_7E => X"00000038000000000000003e0000000000000038000000000000004400000000",
            INIT_7F => X"0000005c000000000000005c0000000000000039000000000000004100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61 : if BRAM_NAME = "samplegold_layersamples_instance61" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000039000000000000004b0000000000000043000000000000004600000000",
            INIT_01 => X"000000390000000000000046000000000000004a000000000000004100000000",
            INIT_02 => X"00000031000000000000003a0000000000000037000000000000003500000000",
            INIT_03 => X"00000047000000000000005d000000000000005b000000000000003a00000000",
            INIT_04 => X"000000500000000000000043000000000000004a000000000000003f00000000",
            INIT_05 => X"000000350000000000000032000000000000003e000000000000004300000000",
            INIT_06 => X"0000003700000000000000300000000000000033000000000000003500000000",
            INIT_07 => X"0000003200000000000000480000000000000051000000000000004f00000000",
            INIT_08 => X"000000350000000000000040000000000000004c000000000000004500000000",
            INIT_09 => X"0000003300000000000000330000000000000026000000000000003500000000",
            INIT_0A => X"0000000000000000000000350000000000000036000000000000003300000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000003b00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000026000000000000000f0000000000000000000000000000000000000000",
            INIT_13 => X"0000002c00000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"000000000000000000000000000000000000003a000000000000004700000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_18 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_19 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_1A => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_1C => X"0000000000000000000000000000000000000006000000000000000e00000000",
            INIT_1D => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_1E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_20 => X"000000000000000000000000000000000000000a000000000000000b00000000",
            INIT_21 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_25 => X"0000000300000000000000000000000000000006000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000007e000000000000000f0000000000000007000000000000000700000000",
            INIT_28 => X"000000000000000000000000000000000000000c000000000000002500000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_2A => X"0000002800000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000007100000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"000000000000000000000000000000000000002a000000000000004f00000000",
            INIT_2D => X"0000002b00000000000000130000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000003800000000",
            INIT_31 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000000f0000000000000000000000000000000f00000000",
            INIT_33 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_36 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000001300000000000000000000000000000009000000000000000000000000",
            INIT_39 => X"000000140000000000000012000000000000000c000000000000002e00000000",
            INIT_3A => X"0000002900000000000000050000000000000009000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_3D => X"0000000c00000000000000110000000000000015000000000000001400000000",
            INIT_3E => X"0000000800000000000000000000000000000000000000000000000600000000",
            INIT_3F => X"0000001600000000000000000000000000000018000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001c00000000000000000000000000000000000000000000001400000000",
            INIT_41 => X"0000000700000000000000000000000000000009000000000000001400000000",
            INIT_42 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000800000000000000000000000000000000000000000000000100000000",
            INIT_44 => X"0000000000000000000000030000000000000000000000000000000900000000",
            INIT_45 => X"0000000000000000000000000000000000000073000000000000000e00000000",
            INIT_46 => X"0000000200000000000000070000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000e00000000000000000000000000000000000000000000002300000000",
            INIT_49 => X"0000000500000000000000000000000000000000000000000000005a00000000",
            INIT_4A => X"0000000000000000000000050000000000000008000000000000000300000000",
            INIT_4B => X"0000006500000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000080000000000000000000000000000001500000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_4F => X"0000003400000000000000110000000000000000000000000000003d00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_51 => X"00000000000000000000002a0000000000000004000000000000000000000000",
            INIT_52 => X"0000005000000000000000000000000000000000000000000000000e00000000",
            INIT_53 => X"0000004a000000000000001f0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"000000010000000000000000000000000000003e000000000000000000000000",
            INIT_56 => X"00000000000000000000002d0000000000000005000000000000000000000000",
            INIT_57 => X"0000000000000000000000140000000000000030000000000000000600000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000070000000000000003000000000000003900000000",
            INIT_5A => X"00000000000000000000000d0000000000000000000000000000003900000000",
            INIT_5B => X"00000000000000000000000c0000000000000000000000000000002d00000000",
            INIT_5C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000620000000000000000000000000000001b000000000000001d00000000",
            INIT_5E => X"00000000000000000000000d000000000000001b000000000000000000000000",
            INIT_5F => X"0000001400000000000000000000000000000000000000000000003f00000000",
            INIT_60 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_62 => X"0000003600000000000000220000000000000000000000000000000000000000",
            INIT_63 => X"0000004300000000000000000000000000000020000000000000000000000000",
            INIT_64 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_66 => X"0000005300000000000000070000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000020000000000000000000000000",
            INIT_68 => X"0000003500000000000000000000000000000000000000000000000c00000000",
            INIT_69 => X"0000003c00000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000003d000000000000000d0000000000000000000000000000000000000000",
            INIT_6B => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"00000000000000000000002c0000000000000000000000000000000c00000000",
            INIT_6D => X"0000000000000000000000170000000000000015000000000000000000000000",
            INIT_6E => X"00000000000000000000003d000000000000001a000000000000000000000000",
            INIT_6F => X"0000001400000000000000210000000000000000000000000000000500000000",
            INIT_70 => X"0000000000000000000000000000000000000014000000000000000800000000",
            INIT_71 => X"0000000a00000000000000000000000000000007000000000000004800000000",
            INIT_72 => X"0000000700000000000000000000000000000029000000000000001f00000000",
            INIT_73 => X"00000012000000000000000b0000000000000000000000000000000500000000",
            INIT_74 => X"0000002000000000000000000000000000000000000000000000001e00000000",
            INIT_75 => X"0000001f000000000000000e0000000000000013000000000000001b00000000",
            INIT_76 => X"0000001b00000000000000060000000000000000000000000000000800000000",
            INIT_77 => X"00000001000000000000000f0000000000000000000000000000000000000000",
            INIT_78 => X"0000002800000000000000110000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000002c0000000000000000000000000000003100000000",
            INIT_7A => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_7B => X"0000005d000000000000001c0000000000000011000000000000000000000000",
            INIT_7C => X"000000590000000000000050000000000000004a000000000000004f00000000",
            INIT_7D => X"0000002f000000000000003a0000000000000052000000000000005000000000",
            INIT_7E => X"0000006a0000000000000066000000000000006b000000000000005f00000000",
            INIT_7F => X"00000041000000000000004b0000000000000013000000000000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62 : if BRAM_NAME = "samplegold_layersamples_instance62" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000048000000000000003e000000000000003b000000000000003f00000000",
            INIT_01 => X"0000004f00000000000000390000000000000049000000000000004d00000000",
            INIT_02 => X"000000160000000000000062000000000000005d000000000000005900000000",
            INIT_03 => X"000000390000000000000044000000000000003b000000000000001300000000",
            INIT_04 => X"000000330000000000000030000000000000002f000000000000003d00000000",
            INIT_05 => X"0000003e00000000000000320000000000000034000000000000003300000000",
            INIT_06 => X"0000003400000000000000470000000000000049000000000000004400000000",
            INIT_07 => X"00000041000000000000002f0000000000000038000000000000004000000000",
            INIT_08 => X"0000002d0000000000000034000000000000003e000000000000004800000000",
            INIT_09 => X"0000003a00000000000000450000000000000034000000000000003700000000",
            INIT_0A => X"0000003900000000000000380000000000000040000000000000002f00000000",
            INIT_0B => X"0000003f00000000000000360000000000000030000000000000003900000000",
            INIT_0C => X"000000340000000000000029000000000000002d000000000000003700000000",
            INIT_0D => X"000000270000000000000038000000000000003f000000000000003500000000",
            INIT_0E => X"0000003d00000000000000350000000000000033000000000000003700000000",
            INIT_0F => X"00000032000000000000003b0000000000000033000000000000003400000000",
            INIT_10 => X"0000002c0000000000000030000000000000002d000000000000003600000000",
            INIT_11 => X"0000003400000000000000250000000000000035000000000000003400000000",
            INIT_12 => X"000000350000000000000045000000000000003e000000000000003700000000",
            INIT_13 => X"00000038000000000000002d0000000000000039000000000000002f00000000",
            INIT_14 => X"0000003300000000000000350000000000000030000000000000002a00000000",
            INIT_15 => X"00000034000000000000002e000000000000002e000000000000003a00000000",
            INIT_16 => X"0000003100000000000000390000000000000046000000000000005c00000000",
            INIT_17 => X"0000002f0000000000000034000000000000003c000000000000003100000000",
            INIT_18 => X"00000034000000000000002d000000000000001f000000000000003500000000",
            INIT_19 => X"0000005a000000000000002b000000000000002f000000000000002900000000",
            INIT_1A => X"0000003b00000000000000410000000000000038000000000000004800000000",
            INIT_1B => X"00000045000000000000003c0000000000000032000000000000004300000000",
            INIT_1C => X"0000002400000000000000280000000000000025000000000000004500000000",
            INIT_1D => X"0000003e000000000000003f000000000000002d000000000000002f00000000",
            INIT_1E => X"000000410000000000000033000000000000002d000000000000002f00000000",
            INIT_1F => X"0000004a00000000000000440000000000000041000000000000004900000000",
            INIT_20 => X"0000002c00000000000000330000000000000046000000000000004800000000",
            INIT_21 => X"0000003e00000000000000400000000000000031000000000000002b00000000",
            INIT_22 => X"0000004100000000000000360000000000000032000000000000003d00000000",
            INIT_23 => X"000000440000000000000044000000000000003c000000000000004500000000",
            INIT_24 => X"0000002e000000000000002a000000000000003d000000000000004300000000",
            INIT_25 => X"000000440000000000000041000000000000003b000000000000002a00000000",
            INIT_26 => X"0000004500000000000000430000000000000042000000000000004400000000",
            INIT_27 => X"000000440000000000000043000000000000003d000000000000003d00000000",
            INIT_28 => X"000000230000000000000029000000000000002a000000000000004200000000",
            INIT_29 => X"0000004700000000000000480000000000000043000000000000003700000000",
            INIT_2A => X"0000003a000000000000003e0000000000000042000000000000004100000000",
            INIT_2B => X"00000041000000000000003b0000000000000039000000000000003900000000",
            INIT_2C => X"0000003000000000000000170000000000000029000000000000002c00000000",
            INIT_2D => X"000000420000000000000049000000000000005c000000000000004500000000",
            INIT_2E => X"0000003b000000000000003a0000000000000036000000000000004000000000",
            INIT_2F => X"0000002300000000000000410000000000000039000000000000003c00000000",
            INIT_30 => X"00000038000000000000002b0000000000000012000000000000002a00000000",
            INIT_31 => X"0000003d000000000000003f000000000000003c000000000000004100000000",
            INIT_32 => X"0000003f000000000000003d0000000000000038000000000000003400000000",
            INIT_33 => X"000000190000000000000000000000000000003a000000000000003c00000000",
            INIT_34 => X"0000002500000000000000210000000000000024000000000000003100000000",
            INIT_35 => X"00000000000000000000001c0000000000000025000000000000001f00000000",
            INIT_36 => X"0000002c000000000000002b0000000000000033000000000000003600000000",
            INIT_37 => X"0000003a00000000000000040000000000000000000000000000002800000000",
            INIT_38 => X"0000003a0000000000000027000000000000003e000000000000003500000000",
            INIT_39 => X"000000420000000000000011000000000000003e000000000000004000000000",
            INIT_3A => X"000000340000000000000038000000000000003d000000000000004900000000",
            INIT_3B => X"0000002b00000000000000380000000000000000000000000000000000000000",
            INIT_3C => X"0000003a000000000000002a0000000000000031000000000000006100000000",
            INIT_3D => X"00000060000000000000004c0000000000000039000000000000003c00000000",
            INIT_3E => X"00000000000000000000004a0000000000000052000000000000005500000000",
            INIT_3F => X"0000006c000000000000002f000000000000002d000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002300000000000000190000000000000021000000000000004e00000000",
            INIT_41 => X"00000069000000000000006d000000000000005f000000000000004600000000",
            INIT_42 => X"0000003e0000000000000035000000000000006e000000000000006200000000",
            INIT_43 => X"0000006000000000000000550000000000000027000000000000004d00000000",
            INIT_44 => X"00000044000000000000002e0000000000000029000000000000004900000000",
            INIT_45 => X"0000004f00000000000000710000000000000076000000000000005f00000000",
            INIT_46 => X"0000005500000000000000540000000000000052000000000000005c00000000",
            INIT_47 => X"0000004500000000000000590000000000000053000000000000003200000000",
            INIT_48 => X"0000005600000000000000400000000000000030000000000000002c00000000",
            INIT_49 => X"00000049000000000000004f0000000000000077000000000000007e00000000",
            INIT_4A => X"0000004d0000000000000039000000000000004f000000000000005100000000",
            INIT_4B => X"000000420000000000000039000000000000004d000000000000004400000000",
            INIT_4C => X"0000007b0000000000000053000000000000004e000000000000004100000000",
            INIT_4D => X"0000004e00000000000000490000000000000069000000000000007b00000000",
            INIT_4E => X"0000004c000000000000005d000000000000001f000000000000005000000000",
            INIT_4F => X"000000580000000000000032000000000000004d000000000000005500000000",
            INIT_50 => X"0000008b0000000000000068000000000000004f000000000000004400000000",
            INIT_51 => X"000000460000000000000048000000000000006e000000000000007300000000",
            INIT_52 => X"0000005b0000000000000064000000000000004d000000000000003a00000000",
            INIT_53 => X"00000039000000000000003a0000000000000034000000000000004800000000",
            INIT_54 => X"00000062000000000000004d000000000000001b000000000000004000000000",
            INIT_55 => X"0000005600000000000000460000000000000054000000000000007300000000",
            INIT_56 => X"00000070000000000000006c0000000000000061000000000000005800000000",
            INIT_57 => X"00000034000000000000003b000000000000001f000000000000004f00000000",
            INIT_58 => X"00000043000000000000002e0000000000000029000000000000003100000000",
            INIT_59 => X"000000580000000000000065000000000000004b000000000000006200000000",
            INIT_5A => X"0000006100000000000000600000000000000047000000000000005b00000000",
            INIT_5B => X"0000003100000000000000340000000000000032000000000000005300000000",
            INIT_5C => X"00000063000000000000002a0000000000000030000000000000003b00000000",
            INIT_5D => X"0000005f00000000000000670000000000000065000000000000004f00000000",
            INIT_5E => X"0000004b00000000000000520000000000000050000000000000004b00000000",
            INIT_5F => X"0000004400000000000000390000000000000031000000000000002600000000",
            INIT_60 => X"0000004e000000000000005c0000000000000025000000000000002e00000000",
            INIT_61 => X"00000034000000000000004b0000000000000068000000000000006300000000",
            INIT_62 => X"000000260000000000000040000000000000004e000000000000005500000000",
            INIT_63 => X"0000003900000000000000370000000000000032000000000000003500000000",
            INIT_64 => X"0000005900000000000000420000000000000055000000000000002900000000",
            INIT_65 => X"0000003d000000000000002c0000000000000049000000000000006b00000000",
            INIT_66 => X"0000002c0000000000000023000000000000002b000000000000003a00000000",
            INIT_67 => X"00000031000000000000002d0000000000000020000000000000002a00000000",
            INIT_68 => X"0000007100000000000000460000000000000042000000000000004e00000000",
            INIT_69 => X"0000002f000000000000002f0000000000000043000000000000005800000000",
            INIT_6A => X"000000290000000000000027000000000000001e000000000000001900000000",
            INIT_6B => X"0000000000000000000000330000000000000024000000000000002000000000",
            INIT_6C => X"0000000000000000000000000000000000000001000000000000000200000000",
            INIT_6D => X"0000000000000000000000000000000000000003000000000000000400000000",
            INIT_6E => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000007000000000000000200000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63 : if BRAM_NAME = "samplegold_layersamples_instance63" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000006d000000000000005c0000000000000050000000000000005a00000000",
            INIT_25 => X"0000001d00000000000000320000000000000041000000000000004e00000000",
            INIT_26 => X"0000007500000000000000710000000000000072000000000000004700000000",
            INIT_27 => X"0000007a00000000000000470000000000000040000000000000004f00000000",
            INIT_28 => X"000000710000000000000091000000000000007c000000000000007700000000",
            INIT_29 => X"000000b000000000000000b40000000000000093000000000000007800000000",
            INIT_2A => X"00000080000000000000006a000000000000008200000000000000a100000000",
            INIT_2B => X"0000008b000000000000008b000000000000005c000000000000007800000000",
            INIT_2C => X"000000150000000000000020000000000000005d000000000000008e00000000",
            INIT_2D => X"0000003900000000000000220000000000000012000000000000001a00000000",
            INIT_2E => X"0000007300000000000000760000000000000061000000000000005700000000",
            INIT_2F => X"0000008d0000000000000089000000000000008a000000000000006700000000",
            INIT_30 => X"0000007100000000000000700000000000000032000000000000007a00000000",
            INIT_31 => X"0000004300000000000000480000000000000058000000000000007000000000",
            INIT_32 => X"0000005400000000000000410000000000000074000000000000008000000000",
            INIT_33 => X"0000008800000000000000aa0000000000000087000000000000008e00000000",
            INIT_34 => X"00000064000000000000008a000000000000006f000000000000003c00000000",
            INIT_35 => X"0000004c000000000000005a0000000000000074000000000000006800000000",
            INIT_36 => X"0000009400000000000000100000000000000055000000000000006c00000000",
            INIT_37 => X"0000005700000000000000500000000000000070000000000000009700000000",
            INIT_38 => X"0000006e00000000000000680000000000000050000000000000004f00000000",
            INIT_39 => X"0000006f00000000000000780000000000000087000000000000006200000000",
            INIT_3A => X"000000a0000000000000007b000000000000008a000000000000008c00000000",
            INIT_3B => X"0000004b00000000000000030000000000000053000000000000008100000000",
            INIT_3C => X"00000052000000000000003a000000000000003d000000000000005500000000",
            INIT_3D => X"000000bf00000000000000950000000000000056000000000000005200000000",
            INIT_3E => X"000000450000000000000093000000000000007f000000000000009000000000",
            INIT_3F => X"0000003300000000000000420000000000000062000000000000004500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000044000000000000005e0000000000000062000000000000003e00000000",
            INIT_41 => X"000000750000000000000063000000000000006a000000000000006100000000",
            INIT_42 => X"0000009e0000000000000025000000000000004f000000000000005300000000",
            INIT_43 => X"00000004000000000000003f0000000000000045000000000000002200000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"00000070000000000000007a000000000000003b000000000000000000000000",
            INIT_46 => X"0000003300000000000000270000000000000048000000000000005f00000000",
            INIT_47 => X"00000077000000000000005d000000000000003c000000000000003100000000",
            INIT_48 => X"0000006e00000000000000730000000000000081000000000000006e00000000",
            INIT_49 => X"0000005d0000000000000075000000000000004f000000000000006f00000000",
            INIT_4A => X"00000024000000000000000f0000000000000013000000000000000000000000",
            INIT_4B => X"000000300000000000000040000000000000001c000000000000000000000000",
            INIT_4C => X"00000011000000000000004b0000000000000009000000000000002800000000",
            INIT_4D => X"000000280000000000000077000000000000007b000000000000004700000000",
            INIT_4E => X"0000005600000000000000030000000000000000000000000000000000000000",
            INIT_4F => X"000000270000000000000061000000000000001e000000000000005400000000",
            INIT_50 => X"0000004d000000000000004a0000000000000070000000000000005100000000",
            INIT_51 => X"000000310000000000000000000000000000000c000000000000007800000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_53 => X"0000002000000000000000220000000000000000000000000000000000000000",
            INIT_54 => X"0000005b00000000000000150000000000000000000000000000002100000000",
            INIT_55 => X"00000027000000000000003a000000000000004f000000000000007b00000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_57 => X"0000000c00000000000000560000000000000080000000000000004f00000000",
            INIT_58 => X"0000005c00000000000000750000000000000036000000000000000000000000",
            INIT_59 => X"0000000f00000000000000210000000000000044000000000000003d00000000",
            INIT_5A => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000049000000000000004400000000",
            INIT_5C => X"00000011000000000000001a0000000000000019000000000000001400000000",
            INIT_5D => X"0000001f00000000000000190000000000000018000000000000001200000000",
            INIT_5E => X"0000001d000000000000001a0000000000000023000000000000002900000000",
            INIT_5F => X"0000001f000000000000002c0000000000000016000000000000001e00000000",
            INIT_60 => X"00000000000000000000000a0000000000000011000000000000001000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"00000021000000000000001e000000000000000f000000000000000000000000",
            INIT_63 => X"0000000c0000000000000032000000000000001b000000000000001b00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000017000000000000001f0000000000000019000000000000000000000000",
            INIT_67 => X"00000005000000000000000c000000000000003c000000000000001900000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000001e0000000000000014000000000000001b000000000000000000000000",
            INIT_6B => X"000000000000000000000006000000000000000f000000000000002b00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000002200000000000000040000000000000016000000000000001000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000016000000000000000d000000000000000d000000000000001700000000",
            INIT_73 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000a00000000000000060000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000000d000000000000000c000000000000000d00000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"000000220000000000000000000000000000000f000000000000001200000000",
            INIT_7B => X"0000000000000000000000080000000000000002000000000000000000000000",
            INIT_7C => X"00000000000000000000001d0000000000000011000000000000000000000000",
            INIT_7D => X"0000002200000000000000000000000000000015000000000000001000000000",
            INIT_7E => X"0000000000000000000000070000000000000000000000000000000100000000",
            INIT_7F => X"0000000900000000000000000000000000000000000000000000000200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64 : if BRAM_NAME = "samplegold_layersamples_instance64" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000600000000000000270000000000000000000000000000000000000000",
            INIT_02 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_06 => X"0000000a00000000000000000000000000000002000000000000000a00000000",
            INIT_07 => X"0000000000000000000000310000000000000000000000000000000f00000000",
            INIT_08 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_09 => X"0000000a00000000000000000000000000000000000000000000002a00000000",
            INIT_0A => X"0000000f00000000000000010000000000000000000000000000000000000000",
            INIT_0B => X"0000000700000000000000310000000000000016000000000000000e00000000",
            INIT_0C => X"00000025000000000000000f0000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001600000000000000130000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000009000000000000001400000000",
            INIT_10 => X"0000000000000000000000140000000000000018000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000080000000000000009000000000000000b000000000000000000000000",
            INIT_13 => X"0000000200000000000000000000000000000000000000000000000300000000",
            INIT_14 => X"0000003b0000000000000040000000000000001e000000000000001100000000",
            INIT_15 => X"000000270000000000000027000000000000002d000000000000004500000000",
            INIT_16 => X"0000004400000000000000350000000000000027000000000000002700000000",
            INIT_17 => X"0000002a00000000000000390000000000000040000000000000003b00000000",
            INIT_18 => X"0000005600000000000000550000000000000057000000000000001f00000000",
            INIT_19 => X"0000003d00000000000000400000000000000038000000000000003400000000",
            INIT_1A => X"00000030000000000000003f000000000000004f000000000000004800000000",
            INIT_1B => X"0000002a00000000000000320000000000000044000000000000003e00000000",
            INIT_1C => X"0000002a0000000000000059000000000000005c000000000000005c00000000",
            INIT_1D => X"0000003f0000000000000042000000000000003f000000000000003100000000",
            INIT_1E => X"00000041000000000000003c0000000000000037000000000000004100000000",
            INIT_1F => X"0000005b00000000000000200000000000000025000000000000003f00000000",
            INIT_20 => X"00000036000000000000004a000000000000004e000000000000005b00000000",
            INIT_21 => X"00000056000000000000005c0000000000000048000000000000004900000000",
            INIT_22 => X"0000004000000000000000450000000000000030000000000000004f00000000",
            INIT_23 => X"0000005b000000000000005a0000000000000009000000000000002c00000000",
            INIT_24 => X"00000044000000000000003e0000000000000042000000000000004b00000000",
            INIT_25 => X"0000004d00000000000000510000000000000050000000000000005900000000",
            INIT_26 => X"0000004c00000000000000490000000000000047000000000000005600000000",
            INIT_27 => X"0000003500000000000000590000000000000053000000000000003300000000",
            INIT_28 => X"000000410000000000000038000000000000001b000000000000002600000000",
            INIT_29 => X"0000004b000000000000003e000000000000003b000000000000003a00000000",
            INIT_2A => X"0000005b000000000000005b0000000000000056000000000000003900000000",
            INIT_2B => X"00000022000000000000002a0000000000000045000000000000004000000000",
            INIT_2C => X"0000002c0000000000000041000000000000003c000000000000002300000000",
            INIT_2D => X"0000001b00000000000000160000000000000037000000000000003100000000",
            INIT_2E => X"0000003400000000000000560000000000000052000000000000003b00000000",
            INIT_2F => X"0000002400000000000000270000000000000017000000000000001c00000000",
            INIT_30 => X"00000000000000000000000f0000000000000016000000000000001600000000",
            INIT_31 => X"0000000f00000000000000000000000000000004000000000000000000000000",
            INIT_32 => X"0000000e0000000000000039000000000000005d000000000000003700000000",
            INIT_33 => X"00000015000000000000000b000000000000001a000000000000000800000000",
            INIT_34 => X"000000000000000000000000000000000000000b000000000000001200000000",
            INIT_35 => X"0000002a000000000000000a0000000000000000000000000000000900000000",
            INIT_36 => X"0000001000000000000000150000000000000044000000000000003500000000",
            INIT_37 => X"0000000700000000000000090000000000000000000000000000000000000000",
            INIT_38 => X"0000003e000000000000003d000000000000002f000000000000001f00000000",
            INIT_39 => X"0000002200000000000000200000000000000047000000000000003700000000",
            INIT_3A => X"000000000000000000000000000000000000001f000000000000004600000000",
            INIT_3B => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_3C => X"000000170000000000000014000000000000001a000000000000000700000000",
            INIT_3D => X"0000005200000000000000150000000000000015000000000000001b00000000",
            INIT_3E => X"0000000000000000000000060000000000000002000000000000001a00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000250000000000000018000000000000001100000000",
            INIT_41 => X"0000002c000000000000004f000000000000000b000000000000000500000000",
            INIT_42 => X"0000000000000000000000030000000000000025000000000000000500000000",
            INIT_43 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000025000000000000002400000000",
            INIT_45 => X"0000002c0000000000000049000000000000004a000000000000000900000000",
            INIT_46 => X"0000000000000000000000000000000000000009000000000000002400000000",
            INIT_47 => X"0000003c000000000000000e0000000000000000000000000000000000000000",
            INIT_48 => X"0000001400000000000000000000000000000000000000000000003600000000",
            INIT_49 => X"0000001100000000000000360000000000000045000000000000004c00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_4B => X"0000001f000000000000000e0000000000000000000000000000000000000000",
            INIT_4C => X"000000fc00000000000000160000000000000000000000000000000000000000",
            INIT_4D => X"000000c800000000000000c400000000000000fb00000000000000f500000000",
            INIT_4E => X"000000ff00000000000000e500000000000000d700000000000000cd00000000",
            INIT_4F => X"000000f6000000000000010600000000000000fa000000000000010700000000",
            INIT_50 => X"00000121000000000000012300000000000000d400000000000000d500000000",
            INIT_51 => X"000000c500000000000000ba00000000000000bc000000000000011500000000",
            INIT_52 => X"000000ef00000000000000eb00000000000000d300000000000000c000000000",
            INIT_53 => X"000000dc000000000000010500000000000000ff00000000000000e700000000",
            INIT_54 => X"00000115000000000000012a000000000000012a00000000000000e600000000",
            INIT_55 => X"000000c500000000000000c500000000000000b400000000000000af00000000",
            INIT_56 => X"000000d200000000000000ab00000000000000b300000000000000bd00000000",
            INIT_57 => X"000000c400000000000000c900000000000000f0000000000000010300000000",
            INIT_58 => X"000000c6000000000000010a0000000000000124000000000000012900000000",
            INIT_59 => X"000000fa00000000000000f6000000000000010200000000000000cf00000000",
            INIT_5A => X"000000f400000000000000ca00000000000000eb00000000000000f400000000",
            INIT_5B => X"0000012900000000000000a700000000000000ca000000000000010000000000",
            INIT_5C => X"000000c900000000000000c400000000000000e0000000000000012200000000",
            INIT_5D => X"000000ec00000000000000e500000000000000ed00000000000000d800000000",
            INIT_5E => X"0000011400000000000000e200000000000000f700000000000000f400000000",
            INIT_5F => X"00000114000000000000011c00000000000000dc000000000000010600000000",
            INIT_60 => X"000000c10000000000000092000000000000009c00000000000000ea00000000",
            INIT_61 => X"000000ce00000000000000c200000000000000c000000000000000b900000000",
            INIT_62 => X"0000012c000000000000011400000000000000e100000000000000d600000000",
            INIT_63 => X"000000bb00000000000000e100000000000000f5000000000000012a00000000",
            INIT_64 => X"000000c900000000000000ba000000000000009b00000000000000b700000000",
            INIT_65 => X"0000009700000000000000bb00000000000000ac00000000000000a200000000",
            INIT_66 => X"00000134000000000000010400000000000000d8000000000000009d00000000",
            INIT_67 => X"000000a300000000000000ad000000000000009200000000000000d900000000",
            INIT_68 => X"0000006a0000000000000074000000000000009100000000000000a900000000",
            INIT_69 => X"00000063000000000000005c0000000000000069000000000000006300000000",
            INIT_6A => X"000000d4000000000000011600000000000000b9000000000000009800000000",
            INIT_6B => X"0000009200000000000000740000000000000096000000000000008400000000",
            INIT_6C => X"0000006e000000000000008800000000000000b2000000000000008c00000000",
            INIT_6D => X"0000008c0000000000000062000000000000008a000000000000007f00000000",
            INIT_6E => X"0000007b00000000000000f200000000000000f200000000000000af00000000",
            INIT_6F => X"0000006a0000000000000060000000000000004b000000000000007900000000",
            INIT_70 => X"000000b000000000000000c7000000000000008f000000000000006300000000",
            INIT_71 => X"0000009600000000000000ba00000000000000b100000000000000b900000000",
            INIT_72 => X"00000059000000000000008d00000000000000f400000000000000c500000000",
            INIT_73 => X"0000007d000000000000004c000000000000002b000000000000005200000000",
            INIT_74 => X"0000008500000000000000820000000000000091000000000000004900000000",
            INIT_75 => X"000000ad00000000000000a3000000000000006300000000000000a100000000",
            INIT_76 => X"000000810000000000000063000000000000007500000000000000f800000000",
            INIT_77 => X"00000057000000000000004d000000000000001d000000000000003500000000",
            INIT_78 => X"0000009b000000000000009e00000000000000a5000000000000004a00000000",
            INIT_79 => X"000000f700000000000000a6000000000000005e000000000000007200000000",
            INIT_7A => X"0000006400000000000000a1000000000000006100000000000000b900000000",
            INIT_7B => X"0000002e0000000000000018000000000000000d000000000000001600000000",
            INIT_7C => X"0000002d00000000000000a400000000000000d000000000000000ab00000000",
            INIT_7D => X"000000e600000000000000e50000000000000095000000000000004200000000",
            INIT_7E => X"000000390000000000000074000000000000008e00000000000000b200000000",
            INIT_7F => X"00000087000000000000003c000000000000001c000000000000000e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65 : if BRAM_NAME = "samplegold_layersamples_instance65" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003e000000000000002000000000000000a300000000000000c500000000",
            INIT_01 => X"000000b400000000000000d900000000000000e900000000000000ab00000000",
            INIT_02 => X"0000002600000000000000420000000000000065000000000000006a00000000",
            INIT_03 => X"0000007f0000000000000059000000000000003c000000000000002f00000000",
            INIT_04 => X"000000b6000000000000003e000000000000001c000000000000008a00000000",
            INIT_05 => X"0000004f00000000000000350000000000000032000000000000003500000000",
            INIT_06 => X"00000000000000000000000e0000000000000016000000000000003500000000",
            INIT_07 => X"0000004b00000000000000510000000000000049000000000000002200000000",
            INIT_08 => X"00000036000000000000004a0000000000000036000000000000003800000000",
            INIT_09 => X"0000003d000000000000005c0000000000000044000000000000003600000000",
            INIT_0A => X"0000006400000000000000600000000000000041000000000000003200000000",
            INIT_0B => X"000000530000000000000042000000000000006e000000000000007000000000",
            INIT_0C => X"0000004000000000000000410000000000000053000000000000007200000000",
            INIT_0D => X"000000000000000000000000000000000000004a000000000000004b00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000007800000000000000500000000000000034000000000000002a00000000",
            INIT_10 => X"0000004300000000000000470000000000000041000000000000006200000000",
            INIT_11 => X"0000000600000000000000000000000000000000000000000000004800000000",
            INIT_12 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000053000000000000003c000000000000004a000000000000004900000000",
            INIT_14 => X"00000040000000000000005a0000000000000047000000000000004200000000",
            INIT_15 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000004000000000000000000000000000000035000000000000002b00000000",
            INIT_18 => X"000000070000000000000018000000000000002e000000000000005500000000",
            INIT_19 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000001d00000000000000210000000000000017000000000000000000000000",
            INIT_1B => X"00000061000000000000002f000000000000003f000000000000004200000000",
            INIT_1C => X"000000000000000000000000000000000000001c000000000000004300000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000005d000000000000004a0000000000000019000000000000001900000000",
            INIT_1F => X"00000010000000000000006b000000000000003e000000000000004800000000",
            INIT_20 => X"00000000000000000000000f000000000000000d000000000000002500000000",
            INIT_21 => X"0000002200000000000000310000000000000032000000000000001600000000",
            INIT_22 => X"0000001600000000000000060000000000000025000000000000003600000000",
            INIT_23 => X"000000740000000000000008000000000000002b000000000000001c00000000",
            INIT_24 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000003400000000000000060000000000000000000000000000000000000000",
            INIT_27 => X"0000000800000000000000280000000000000031000000000000004a00000000",
            INIT_28 => X"0000003a00000000000000080000000000000018000000000000001b00000000",
            INIT_29 => X"00000025000000000000002f0000000000000038000000000000002000000000",
            INIT_2A => X"00000043000000000000002d0000000000000000000000000000003700000000",
            INIT_2B => X"0000000e00000000000000120000000000000014000000000000000000000000",
            INIT_2C => X"0000000a00000000000000120000000000000008000000000000000000000000",
            INIT_2D => X"0000000000000000000000130000000000000000000000000000000700000000",
            INIT_2E => X"0000001200000000000000640000000000000022000000000000000000000000",
            INIT_2F => X"000000360000000000000013000000000000000b000000000000000000000000",
            INIT_30 => X"0000000000000000000000380000000000000000000000000000005800000000",
            INIT_31 => X"0000000000000000000000310000000000000061000000000000001700000000",
            INIT_32 => X"0000000f00000000000000000000000000000000000000000000001100000000",
            INIT_33 => X"0000000a00000000000000110000000000000009000000000000000d00000000",
            INIT_34 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_36 => X"00000009000000000000001c0000000000000019000000000000002300000000",
            INIT_37 => X"0000000000000000000000000000000000000002000000000000001b00000000",
            INIT_38 => X"00000024000000000000004a0000000000000034000000000000002000000000",
            INIT_39 => X"0000000500000000000000130000000000000000000000000000000000000000",
            INIT_3A => X"0000001500000000000000100000000000000022000000000000000a00000000",
            INIT_3B => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"000000000000000000000011000000000000002e000000000000001000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000005d000000000000003c0000000000000037000000000000003200000000",
            INIT_43 => X"0000000000000000000000060000000000000034000000000000005d00000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_4C => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000001c00000000000000000000000000000003000000000000001d00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000001000000000000000000000000000000000000000000000001d00000000",
            INIT_52 => X"0000000000000000000000210000000000000000000000000000001600000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000009000000000000001600000000",
            INIT_55 => X"000000010000000000000000000000000000000b000000000000000000000000",
            INIT_56 => X"0000003f0000000000000018000000000000000a000000000000001e00000000",
            INIT_57 => X"0000001200000000000000040000000000000000000000000000004400000000",
            INIT_58 => X"00000000000000000000000d0000000000000000000000000000000200000000",
            INIT_59 => X"0000003500000000000000380000000000000001000000000000000000000000",
            INIT_5A => X"00000009000000000000003c0000000000000041000000000000001b00000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_5C => X"0000000000000000000000070000000000000000000000000000003c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000400000000000000000000000000000000000000000",
            INIT_60 => X"0000001e00000000000000100000000000000003000000000000002400000000",
            INIT_61 => X"0000002200000000000000280000000000000015000000000000001d00000000",
            INIT_62 => X"000000000000000000000000000000000000000e000000000000003200000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000001300000000000000000000000000000000000000000000001400000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_68 => X"00000027000000000000001b000000000000003a000000000000003900000000",
            INIT_69 => X"0000003b00000000000000150000000000000017000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000300000000000000000000000000000000000000000000000600000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000001500000000000000000000000000000003000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001c000000000000002f000000000000002b000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000002000000000000000b0000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000000000000000000002a000000000000000d000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"00000000000000000000001a0000000000000019000000000000000300000000",
            INIT_78 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000015000000000000001b0000000000000000000000000000000000000000",
            INIT_7B => X"0000000200000000000000240000000000000023000000000000000800000000",
            INIT_7C => X"0000002800000000000000000000000000000000000000000000001c00000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_7F => X"0000000c000000000000006d000000000000000c000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66 : if BRAM_NAME = "samplegold_layersamples_instance66" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000440000000000000000000000000000000000000000",
            INIT_01 => X"0000007a00000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_03 => X"0000000000000000000000550000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000018000000000000004a0000000000000000000000000000000000000000",
            INIT_06 => X"0000000f00000000000000070000000000000004000000000000000000000000",
            INIT_07 => X"00000000000000000000001f0000000000000055000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000027000000000000000000000000",
            INIT_09 => X"000000000000000000000010000000000000003d000000000000000000000000",
            INIT_0A => X"0000000900000000000000150000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000068000000000000003800000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_0E => X"0000004500000000000000000000000000000000000000000000001800000000",
            INIT_0F => X"0000000000000000000000210000000000000037000000000000004f00000000",
            INIT_10 => X"000000000000000000000000000000000000005e000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000005f000000000000001b0000000000000000000000000000000a00000000",
            INIT_13 => X"0000000000000000000000000000000000000094000000000000003f00000000",
            INIT_14 => X"0000000e00000000000000360000000000000000000000000000005300000000",
            INIT_15 => X"0000001a00000000000000000000000000000000000000000000000700000000",
            INIT_16 => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_17 => X"0000002b00000000000000000000000000000000000000000000009e00000000",
            INIT_18 => X"0000001f0000000000000000000000000000002b000000000000000000000000",
            INIT_19 => X"0000000000000000000000100000000000000000000000000000006100000000",
            INIT_1A => X"000000d000000000000000000000000000000008000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000330000000000000028000000000000000000000000",
            INIT_1D => X"0000003300000000000000000000000000000000000000000000006200000000",
            INIT_1E => X"000000000000000000000091000000000000002b000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000042000000000000000000000000",
            INIT_20 => X"0000009300000000000000000000000000000049000000000000001100000000",
            INIT_21 => X"0000000000000000000000160000000000000002000000000000000100000000",
            INIT_22 => X"00000000000000000000000000000000000000d8000000000000001700000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"000000b9000000000000002e0000000000000012000000000000000100000000",
            INIT_25 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000000400000000000000ca00000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002b00000000000000560000000000000035000000000000001500000000",
            INIT_29 => X"000000aa000000000000005c0000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000002c000000000000001a000000000000001000000000",
            INIT_2D => X"0000001700000000000000cc0000000000000046000000000000000000000000",
            INIT_2E => X"0000000f00000000000000000000000000000013000000000000001300000000",
            INIT_2F => X"0000001c00000000000000390000000000000030000000000000002a00000000",
            INIT_30 => X"0000001e00000000000000000000000000000000000000000000000600000000",
            INIT_31 => X"0000001400000000000000150000000000000012000000000000000d00000000",
            INIT_32 => X"00000011000000000000000f0000000000000005000000000000001000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000d000000000000000c000000000000000c000000000000000000000000",
            INIT_36 => X"0000008d000000000000008d0000000000000074000000000000003900000000",
            INIT_37 => X"0000000400000000000000450000000000000079000000000000009000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_39 => X"0000003600000000000000110000000000000008000000000000000c00000000",
            INIT_3A => X"0000006f00000000000000610000000000000058000000000000006600000000",
            INIT_3B => X"00000000000000000000003c0000000000000087000000000000007b00000000",
            INIT_3C => X"000000090000000000000000000000000000000e000000000000000c00000000",
            INIT_3D => X"00000061000000000000003f0000000000000000000000000000000e00000000",
            INIT_3E => X"00000067000000000000006f0000000000000054000000000000004f00000000",
            INIT_3F => X"00000014000000000000002e0000000000000066000000000000006400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000000000000000000003f000000000000002400000000",
            INIT_41 => X"0000006100000000000000420000000000000055000000000000003200000000",
            INIT_42 => X"0000005600000000000000510000000000000058000000000000006700000000",
            INIT_43 => X"0000000d00000000000000120000000000000028000000000000003d00000000",
            INIT_44 => X"0000000000000000000000000000000000000002000000000000000d00000000",
            INIT_45 => X"0000006d00000000000000700000000000000080000000000000005300000000",
            INIT_46 => X"0000003f0000000000000057000000000000006d000000000000007000000000",
            INIT_47 => X"0000000900000000000000000000000000000000000000000000001c00000000",
            INIT_48 => X"0000001d00000000000000180000000000000000000000000000000000000000",
            INIT_49 => X"0000003b000000000000004f0000000000000052000000000000004700000000",
            INIT_4A => X"00000013000000000000002d0000000000000024000000000000001d00000000",
            INIT_4B => X"000000200000000000000011000000000000002d000000000000002300000000",
            INIT_4C => X"0000005100000000000000000000000000000013000000000000002a00000000",
            INIT_4D => X"0000009a0000000000000076000000000000005d000000000000003900000000",
            INIT_4E => X"00000089000000000000009a0000000000000093000000000000009c00000000",
            INIT_4F => X"0000001a00000000000000180000000000000019000000000000005300000000",
            INIT_50 => X"00000038000000000000002e000000000000002e000000000000000100000000",
            INIT_51 => X"0000002500000000000000290000000000000020000000000000002500000000",
            INIT_52 => X"00000030000000000000001a0000000000000022000000000000001f00000000",
            INIT_53 => X"0000004000000000000000310000000000000016000000000000002700000000",
            INIT_54 => X"0000006a0000000000000034000000000000002f000000000000003900000000",
            INIT_55 => X"0000004800000000000000440000000000000033000000000000003900000000",
            INIT_56 => X"00000037000000000000005e0000000000000033000000000000005a00000000",
            INIT_57 => X"0000006a00000000000000220000000000000014000000000000002700000000",
            INIT_58 => X"0000001a00000000000000000000000000000021000000000000004900000000",
            INIT_59 => X"0000001500000000000000440000000000000025000000000000001800000000",
            INIT_5A => X"0000003c0000000000000028000000000000000f000000000000001900000000",
            INIT_5B => X"0000004c000000000000003c0000000000000060000000000000008000000000",
            INIT_5C => X"0000003c0000000000000032000000000000002e000000000000003f00000000",
            INIT_5D => X"0000002d00000000000000490000000000000058000000000000005900000000",
            INIT_5E => X"0000003700000000000000420000000000000049000000000000004100000000",
            INIT_5F => X"0000004000000000000000420000000000000030000000000000004500000000",
            INIT_60 => X"0000000f0000000000000037000000000000003f000000000000003b00000000",
            INIT_61 => X"0000003c000000000000002c000000000000002b000000000000001400000000",
            INIT_62 => X"00000052000000000000004f0000000000000045000000000000004a00000000",
            INIT_63 => X"00000040000000000000003b000000000000003a000000000000003400000000",
            INIT_64 => X"000000270000000000000038000000000000003c000000000000004100000000",
            INIT_65 => X"0000005c0000000000000039000000000000003a000000000000003600000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67 : if BRAM_NAME = "samplegold_layersamples_instance67" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000004e0000000000000062000000000000005a000000000000000000000000",
            INIT_1F => X"0000006500000000000000490000000000000034000000000000001e00000000",
            INIT_20 => X"00000043000000000000004b000000000000006d000000000000008500000000",
            INIT_21 => X"0000004d000000000000005b000000000000005b000000000000004500000000",
            INIT_22 => X"0000000000000000000000390000000000000057000000000000005600000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000004400000000000000230000000000000005000000000000000000000000",
            INIT_25 => X"0000004a000000000000004e0000000000000026000000000000003b00000000",
            INIT_26 => X"0000004700000000000000080000000000000031000000000000004800000000",
            INIT_27 => X"0000004600000000000000640000000000000069000000000000006100000000",
            INIT_28 => X"0000002e0000000000000052000000000000004a000000000000002800000000",
            INIT_29 => X"00000040000000000000004a0000000000000031000000000000000e00000000",
            INIT_2A => X"0000004600000000000000510000000000000000000000000000003200000000",
            INIT_2B => X"000000560000000000000046000000000000002d000000000000003200000000",
            INIT_2C => X"00000041000000000000003b0000000000000029000000000000003a00000000",
            INIT_2D => X"00000000000000000000003b0000000000000046000000000000002600000000",
            INIT_2E => X"0000000a000000000000001f000000000000003d000000000000000000000000",
            INIT_2F => X"000000390000000000000032000000000000002b000000000000002d00000000",
            INIT_30 => X"0000008c000000000000005c000000000000005b000000000000005700000000",
            INIT_31 => X"000000010000000000000032000000000000001c000000000000003500000000",
            INIT_32 => X"0000000d000000000000001e0000000000000029000000000000000700000000",
            INIT_33 => X"000000220000000000000008000000000000001c000000000000000700000000",
            INIT_34 => X"0000002a000000000000004b0000000000000049000000000000005700000000",
            INIT_35 => X"0000006400000000000000190000000000000000000000000000000000000000",
            INIT_36 => X"0000002c0000000000000020000000000000001a000000000000002900000000",
            INIT_37 => X"0000000000000000000000120000000000000006000000000000001900000000",
            INIT_38 => X"000000000000000000000010000000000000003e000000000000000000000000",
            INIT_39 => X"0000000f00000000000000070000000000000020000000000000003100000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_3B => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000002e000000000000000d0000000000000038000000000000004c00000000",
            INIT_3D => X"0000003000000000000000190000000000000029000000000000000000000000",
            INIT_3E => X"0000009800000000000000ae00000000000000a7000000000000005400000000",
            INIT_3F => X"00000041000000000000003d00000000000000a200000000000000ac00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000200000000000000000000000000000000000000000000003000000000",
            INIT_41 => X"0000000e00000000000000000000000000000000000000000000000400000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000003000000000000000550000000000000000000000000000000200000000",
            INIT_44 => X"00000003000000000000000e000000000000001c000000000000000000000000",
            INIT_45 => X"00000019000000000000000b000000000000005c000000000000000a00000000",
            INIT_46 => X"00000005000000000000005c000000000000001d000000000000001f00000000",
            INIT_47 => X"0000000000000000000000250000000000000059000000000000004100000000",
            INIT_48 => X"000000060000000000000012000000000000004d000000000000001600000000",
            INIT_49 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000006000000000000003300000000",
            INIT_4B => X"000000690000000000000057000000000000002b000000000000004700000000",
            INIT_4C => X"00000005000000000000000e000000000000001a000000000000001700000000",
            INIT_4D => X"0000006a000000000000008e000000000000001b000000000000000c00000000",
            INIT_4E => X"0000006f00000000000000200000000000000000000000000000002600000000",
            INIT_4F => X"0000000b00000000000000120000000000000013000000000000003d00000000",
            INIT_50 => X"00000020000000000000001b0000000000000001000000000000001300000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_52 => X"0000001f0000000000000056000000000000002d000000000000000000000000",
            INIT_53 => X"0000000c00000000000000000000000000000021000000000000002d00000000",
            INIT_54 => X"0000001e0000000000000021000000000000001f000000000000000900000000",
            INIT_55 => X"0000000900000000000000000000000000000009000000000000001600000000",
            INIT_56 => X"0000004c000000000000004a0000000000000075000000000000002900000000",
            INIT_57 => X"0000002c00000000000000270000000000000045000000000000004600000000",
            INIT_58 => X"0000004d0000000000000049000000000000003b000000000000003200000000",
            INIT_59 => X"00000058000000000000004a0000000000000047000000000000005100000000",
            INIT_5A => X"0000004a00000000000000490000000000000048000000000000004800000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_5C => X"0000004300000000000000280000000000000009000000000000000300000000",
            INIT_5D => X"00000048000000000000005c000000000000004c000000000000004600000000",
            INIT_5E => X"0000001c00000000000000420000000000000047000000000000004700000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"00000048000000000000001b0000000000000000000000000000000000000000",
            INIT_61 => X"00000047000000000000004c000000000000004e000000000000005500000000",
            INIT_62 => X"00000000000000000000000c000000000000003b000000000000004600000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"00000044000000000000002a0000000000000018000000000000000000000000",
            INIT_65 => X"000000460000000000000045000000000000004b000000000000005300000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000004a000000000000003c000000000000001c000000000000000000000000",
            INIT_69 => X"0000001300000000000000420000000000000038000000000000004a00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000004700000000000000470000000000000025000000000000000000000000",
            INIT_6D => X"0000000000000000000000210000000000000036000000000000003700000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000370000000000000036000000000000001e000000000000001300000000",
            INIT_71 => X"0000000000000000000000190000000000000004000000000000002b00000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000001a00000000000000380000000000000014000000000000000000000000",
            INIT_75 => X"000000000000000000000000000000000000000b000000000000001700000000",
            INIT_76 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"000000000000000000000002000000000000000b000000000000000800000000",
            INIT_78 => X"00000000000000000000001e0000000000000033000000000000001200000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000010000000000000016000000000000002e00000000",
            INIT_7D => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000001700000000000000020000000000000000000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68 : if BRAM_NAME = "samplegold_layersamples_instance68" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000000000000000000000000000000000000e000000000000001800000000",
            INIT_07 => X"0000000000000000000000040000000000000004000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000056000000000000004b0000000000000018000000000000000000000000",
            INIT_14 => X"00000055000000000000007f000000000000008f000000000000007000000000",
            INIT_15 => X"0000000000000000000000020000000000000000000000000000001d00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000020000000000000002c0000000000000000000000000000000000000000",
            INIT_19 => X"0000002b000000000000000b0000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000001300000000000000000000000000000000000000000000000500000000",
            INIT_1C => X"00000039000000000000001e0000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_1E => X"0000001c000000000000000b000000000000003f000000000000000000000000",
            INIT_1F => X"0000001b00000000000000180000000000000022000000000000003700000000",
            INIT_20 => X"0000000000000000000000130000000000000000000000000000001700000000",
            INIT_21 => X"0000001000000000000000190000000000000000000000000000000000000000",
            INIT_22 => X"0000001200000000000000500000000000000000000000000000000000000000",
            INIT_23 => X"00000029000000000000003b000000000000002f000000000000001400000000",
            INIT_24 => X"000000000000000000000012000000000000003f000000000000004700000000",
            INIT_25 => X"0000002f0000000000000030000000000000001c000000000000000000000000",
            INIT_26 => X"00000005000000000000000d0000000000000000000000000000000000000000",
            INIT_27 => X"0000001e000000000000001d0000000000000001000000000000000300000000",
            INIT_28 => X"00000008000000000000006b0000000000000085000000000000004a00000000",
            INIT_29 => X"000000000000000000000000000000000000003d000000000000001e00000000",
            INIT_2A => X"00000027000000000000001e0000000000000013000000000000002b00000000",
            INIT_2B => X"0000006200000000000000370000000000000053000000000000005a00000000",
            INIT_2C => X"0000000000000000000000370000000000000048000000000000006500000000",
            INIT_2D => X"0000000000000000000000530000000000000011000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000052000000000000000000000000",
            INIT_31 => X"0000001300000000000000440000000000000000000000000000004d00000000",
            INIT_32 => X"000000510000000000000045000000000000003f000000000000004d00000000",
            INIT_33 => X"00000031000000000000004c0000000000000052000000000000005800000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000003900000000",
            INIT_35 => X"000000000000000000000020000000000000000e000000000000000000000000",
            INIT_36 => X"0000000300000000000000000000000000000032000000000000000400000000",
            INIT_37 => X"0000002900000000000000000000000000000020000000000000000000000000",
            INIT_38 => X"00000000000000000000001e000000000000000b000000000000000e00000000",
            INIT_39 => X"00000020000000000000007d000000000000001a000000000000000000000000",
            INIT_3A => X"0000003f00000000000000000000000000000014000000000000004b00000000",
            INIT_3B => X"0000000d000000000000002f0000000000000070000000000000001000000000",
            INIT_3C => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_3D => X"0000000300000000000000050000000000000002000000000000000000000000",
            INIT_3E => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000001800000000000000000000000000000011000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_41 => X"0000007900000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000600000000000000000000000000000011000000000000005300000000",
            INIT_43 => X"0000000000000000000000000000000000000018000000000000001c00000000",
            INIT_44 => X"000000000000000000000000000000000000000c000000000000001d00000000",
            INIT_45 => X"0000003900000000000000130000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000060000000000000000000000000000001300000000",
            INIT_47 => X"0000003900000000000000080000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_4A => X"00000000000000000000000f0000000000000001000000000000000d00000000",
            INIT_4B => X"0000000a000000000000007d000000000000001a000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_4F => X"00000000000000000000000000000000000000c3000000000000001800000000",
            INIT_50 => X"0000000000000000000000010000000000000016000000000000000000000000",
            INIT_51 => X"0000002e00000000000000230000000000000000000000000000000000000000",
            INIT_52 => X"00000010000000000000000d0000000000000000000000000000000000000000",
            INIT_53 => X"0000004900000000000000000000000000000000000000000000009e00000000",
            INIT_54 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000001500000000000000280000000000000000000000000000000000000000",
            INIT_56 => X"00000061000000000000005c0000000000000010000000000000000000000000",
            INIT_57 => X"0000000000000000000000140000000000000002000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_5A => X"00000000000000000000008d000000000000003a000000000000002900000000",
            INIT_5B => X"0000000200000000000000070000000000000018000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000d00000000000000010000000000000023000000000000001b00000000",
            INIT_5F => X"0000000000000000000000000000000000000010000000000000001300000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_61 => X"00000000000000000000006d0000000000000016000000000000000000000000",
            INIT_62 => X"000000010000000000000014000000000000000b000000000000006500000000",
            INIT_63 => X"0000001d0000000000000000000000000000000c000000000000002d00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_65 => X"0000005f00000000000000000000000000000074000000000000002200000000",
            INIT_66 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_68 => X"0000001d00000000000000000000000000000013000000000000000000000000",
            INIT_69 => X"00000000000000000000005b000000000000000000000000000000b800000000",
            INIT_6A => X"0000001900000000000000000000000000000000000000000000002000000000",
            INIT_6B => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_6C => X"000000a400000000000000040000000000000000000000000000003b00000000",
            INIT_6D => X"000000000000000000000026000000000000001b000000000000000f00000000",
            INIT_6E => X"0000002900000000000000000000000000000078000000000000000000000000",
            INIT_6F => X"0000000000000000000000460000000000000000000000000000000100000000",
            INIT_70 => X"0000000000000000000000d60000000000000012000000000000000000000000",
            INIT_71 => X"0000000000000000000000170000000000000060000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_73 => X"000000000000000000000000000000000000007e000000000000000600000000",
            INIT_74 => X"0000000000000000000000180000000000000052000000000000000000000000",
            INIT_75 => X"0000000000000000000000040000000000000040000000000000003200000000",
            INIT_76 => X"00000070000000000000000e0000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000004f00000000",
            INIT_78 => X"00000008000000000000000b0000000000000042000000000000001900000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000004a00000000",
            INIT_7A => X"0000003400000000000000640000000000000000000000000000000000000000",
            INIT_7B => X"0000000900000000000000080000000000000000000000000000000000000000",
            INIT_7C => X"0000001c00000000000000030000000000000031000000000000003000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_7E => X"000000000000000000000041000000000000000a000000000000000000000000",
            INIT_7F => X"0000003c00000000000000330000000000000035000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69 : if BRAM_NAME = "samplegold_layersamples_instance69" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000330000000000000037000000000000002c000000000000003200000000",
            INIT_01 => X"0000002f000000000000002e0000000000000030000000000000003500000000",
            INIT_02 => X"0000002c000000000000002f0000000000000039000000000000003000000000",
            INIT_03 => X"0000001c00000000000000380000000000000035000000000000003500000000",
            INIT_04 => X"000000030000000000000003000000000000000b000000000000000e00000000",
            INIT_05 => X"00000033000000000000001c0000000000000017000000000000000a00000000",
            INIT_06 => X"000000340000000000000026000000000000002e000000000000003300000000",
            INIT_07 => X"00000010000000000000002c0000000000000036000000000000003400000000",
            INIT_08 => X"000000110000000000000018000000000000001a000000000000001c00000000",
            INIT_09 => X"0000003c00000000000000390000000000000012000000000000000d00000000",
            INIT_0A => X"0000003400000000000000340000000000000019000000000000002e00000000",
            INIT_0B => X"0000002300000000000000160000000000000027000000000000003100000000",
            INIT_0C => X"0000001500000000000000120000000000000007000000000000001900000000",
            INIT_0D => X"00000040000000000000003b000000000000001d000000000000002000000000",
            INIT_0E => X"0000001a00000000000000370000000000000035000000000000002800000000",
            INIT_0F => X"000000060000000000000006000000000000000d000000000000001200000000",
            INIT_10 => X"000000150000000000000008000000000000000d000000000000000a00000000",
            INIT_11 => X"0000004700000000000000410000000000000032000000000000002300000000",
            INIT_12 => X"0000002800000000000000320000000000000037000000000000003500000000",
            INIT_13 => X"00000006000000000000000e000000000000000d000000000000000300000000",
            INIT_14 => X"000000120000000000000005000000000000000b000000000000000600000000",
            INIT_15 => X"0000003d00000000000000350000000000000035000000000000002900000000",
            INIT_16 => X"0000001a00000000000000280000000000000032000000000000003800000000",
            INIT_17 => X"0000000c000000000000000f0000000000000011000000000000001000000000",
            INIT_18 => X"0000000e00000000000000090000000000000011000000000000000f00000000",
            INIT_19 => X"000000300000000000000049000000000000002f000000000000001300000000",
            INIT_1A => X"00000020000000000000000d0000000000000037000000000000003400000000",
            INIT_1B => X"00000007000000000000000a0000000000000016000000000000001900000000",
            INIT_1C => X"0000000c00000000000000020000000000000005000000000000000e00000000",
            INIT_1D => X"0000003600000000000000340000000000000049000000000000002500000000",
            INIT_1E => X"0000001f00000000000000190000000000000021000000000000001400000000",
            INIT_1F => X"000000420000000000000039000000000000003e000000000000003100000000",
            INIT_20 => X"0000002000000000000000280000000000000032000000000000003e00000000",
            INIT_21 => X"0000001b000000000000001e000000000000002b000000000000004200000000",
            INIT_22 => X"0000000400000000000000080000000000000013000000000000000800000000",
            INIT_23 => X"0000000c000000000000000c000000000000000a000000000000001a00000000",
            INIT_24 => X"0000003b00000000000000130000000000000011000000000000001000000000",
            INIT_25 => X"00000015000000000000001c000000000000002b000000000000002f00000000",
            INIT_26 => X"0000001400000000000000210000000000000020000000000000000c00000000",
            INIT_27 => X"0000001e000000000000002a0000000000000021000000000000002500000000",
            INIT_28 => X"00000023000000000000002e0000000000000018000000000000002400000000",
            INIT_29 => X"0000000e00000000000000220000000000000030000000000000001500000000",
            INIT_2A => X"0000001900000000000000080000000000000011000000000000000100000000",
            INIT_2B => X"0000000c0000000000000012000000000000001c000000000000002400000000",
            INIT_2C => X"00000029000000000000003f0000000000000028000000000000000800000000",
            INIT_2D => X"00000011000000000000001b0000000000000022000000000000002600000000",
            INIT_2E => X"0000003500000000000000280000000000000011000000000000001000000000",
            INIT_2F => X"0000000c00000000000000120000000000000018000000000000003900000000",
            INIT_30 => X"0000002200000000000000290000000000000027000000000000002900000000",
            INIT_31 => X"0000001500000000000000160000000000000021000000000000001900000000",
            INIT_32 => X"0000002d000000000000000f000000000000000a000000000000001300000000",
            INIT_33 => X"0000001d000000000000000b000000000000000d000000000000001400000000",
            INIT_34 => X"0000001700000000000000170000000000000029000000000000001f00000000",
            INIT_35 => X"0000001600000000000000180000000000000018000000000000001b00000000",
            INIT_36 => X"0000001a00000000000000250000000000000015000000000000001700000000",
            INIT_37 => X"0000006b000000000000006d0000000000000011000000000000001100000000",
            INIT_38 => X"000000550000000000000056000000000000004d000000000000006900000000",
            INIT_39 => X"0000007a0000000000000073000000000000005d000000000000005900000000",
            INIT_3A => X"0000005b0000000000000061000000000000007a000000000000007200000000",
            INIT_3B => X"0000007500000000000000810000000000000082000000000000005500000000",
            INIT_3C => X"0000006300000000000000640000000000000059000000000000004400000000",
            INIT_3D => X"0000007400000000000000840000000000000081000000000000007200000000",
            INIT_3E => X"000000700000000000000063000000000000007a000000000000007700000000",
            INIT_3F => X"0000002800000000000000780000000000000089000000000000008900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000043000000000000004e000000000000004d000000000000005000000000",
            INIT_41 => X"000000780000000000000076000000000000004a000000000000004400000000",
            INIT_42 => X"00000088000000000000006c0000000000000055000000000000006600000000",
            INIT_43 => X"0000006e00000000000000380000000000000075000000000000008400000000",
            INIT_44 => X"0000006f00000000000000760000000000000067000000000000008200000000",
            INIT_45 => X"0000006f0000000000000083000000000000005b000000000000006800000000",
            INIT_46 => X"00000080000000000000008a000000000000004c000000000000004900000000",
            INIT_47 => X"0000006800000000000000690000000000000043000000000000006200000000",
            INIT_48 => X"000000750000000000000072000000000000006e000000000000006c00000000",
            INIT_49 => X"0000006700000000000000810000000000000075000000000000006a00000000",
            INIT_4A => X"000000570000000000000079000000000000008a000000000000004b00000000",
            INIT_4B => X"00000050000000000000005c0000000000000055000000000000002600000000",
            INIT_4C => X"0000007000000000000000640000000000000060000000000000005c00000000",
            INIT_4D => X"0000008900000000000000890000000000000090000000000000007800000000",
            INIT_4E => X"000000380000000000000052000000000000005e000000000000007000000000",
            INIT_4F => X"0000004300000000000000550000000000000052000000000000003700000000",
            INIT_50 => X"0000005700000000000000450000000000000057000000000000004c00000000",
            INIT_51 => X"0000005e0000000000000095000000000000008f000000000000007f00000000",
            INIT_52 => X"0000004800000000000000380000000000000052000000000000003200000000",
            INIT_53 => X"0000003b000000000000002d0000000000000033000000000000003f00000000",
            INIT_54 => X"0000005c000000000000003b000000000000002a000000000000003d00000000",
            INIT_55 => X"0000001b000000000000004b000000000000009c000000000000005d00000000",
            INIT_56 => X"0000003f0000000000000041000000000000002f000000000000004500000000",
            INIT_57 => X"0000001a000000000000000c0000000000000027000000000000004b00000000",
            INIT_58 => X"0000004900000000000000290000000000000005000000000000001700000000",
            INIT_59 => X"0000004400000000000000120000000000000060000000000000009000000000",
            INIT_5A => X"0000003400000000000000280000000000000031000000000000000900000000",
            INIT_5B => X"000000580000000000000057000000000000005b000000000000004f00000000",
            INIT_5C => X"00000076000000000000003b000000000000005e000000000000005600000000",
            INIT_5D => X"0000001400000000000000180000000000000017000000000000006800000000",
            INIT_5E => X"0000000d0000000000000032000000000000002a000000000000000c00000000",
            INIT_5F => X"0000004800000000000000360000000000000030000000000000005400000000",
            INIT_60 => X"0000006a00000000000000600000000000000042000000000000002200000000",
            INIT_61 => X"0000000000000000000000220000000000000039000000000000001200000000",
            INIT_62 => X"00000034000000000000001f0000000000000037000000000000000a00000000",
            INIT_63 => X"00000021000000000000004b0000000000000041000000000000004c00000000",
            INIT_64 => X"00000026000000000000006f0000000000000067000000000000003900000000",
            INIT_65 => X"0000000000000000000000170000000000000042000000000000001600000000",
            INIT_66 => X"0000005900000000000000120000000000000005000000000000000000000000",
            INIT_67 => X"0000001d0000000000000005000000000000002b000000000000005000000000",
            INIT_68 => X"0000003e00000000000000640000000000000065000000000000005700000000",
            INIT_69 => X"000000000000000000000002000000000000002c000000000000003e00000000",
            INIT_6A => X"0000006500000000000000510000000000000018000000000000000200000000",
            INIT_6B => X"0000006200000000000000200000000000000000000000000000003100000000",
            INIT_6C => X"00000027000000000000003f000000000000005d000000000000006900000000",
            INIT_6D => X"0000000900000000000000030000000000000010000000000000002900000000",
            INIT_6E => X"0000003400000000000000410000000000000027000000000000001400000000",
            INIT_6F => X"000000000000000000000065000000000000001e000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70 : if BRAM_NAME = "samplegold_layersamples_instance70" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70;

MEM_EMPTY_36Kb : if BRAM_NAME(1 to 7) = "default" generate
    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
        BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
        DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
        DO_REG => 0,                     -- Optional output register (0 or 1)
        INIT => X"000000000000000000",   -- Initial values on output port
        INIT_FILE => "NONE",
        WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        SRVAL => X"000000000000000000",  -- Set/Reset value for port output
        WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
    )
    port map (
        DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
        ADDR => bram_addr,  -- Input address, width defined by read/write port depth
        CLK => CLK,    -- 1-bit input clock
        DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
        EN => EN,      -- 1-bit input RAM enable
        REGCE => '1', -- 1-bit input output register enable
        RST => RST,    -- 1-bit input reset
        WE => bram_wr_en       -- Input write enable, width defined by write port depth
    );
-- End of BRAM_SINGLE_MACRO_inst instantiation
end generate;


end a1;