library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (

    -- ifmap
    -- channel=0
    0, 29, 34, 34, 33, 25, 23, 34, 34, 26, 28, 29, 30, 28, 27, 6, 
    0, 6, 17, 13, 24, 0, 7, 18, 21, 0, 0, 1, 17, 14, 11, 0, 
    0, 4, 17, 19, 32, 10, 0, 6, 27, 0, 0, 0, 0, 22, 3, 0, 
    0, 0, 6, 4, 0, 0, 0, 0, 27, 0, 0, 0, 0, 10, 19, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 28, 0, 
    0, 0, 0, 52, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 17, 21, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 
    0, 17, 1, 1, 0, 3, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    
    -- channel=2
    0, 89, 98, 104, 138, 182, 172, 114, 57, 63, 70, 49, 23, 6, 0, 0, 
    0, 86, 98, 110, 172, 240, 245, 115, 52, 154, 270, 249, 122, 10, 0, 0, 
    0, 91, 95, 126, 177, 261, 279, 170, 153, 314, 510, 461, 248, 60, 0, 0, 
    187, 384, 302, 307, 391, 519, 472, 338, 276, 421, 615, 563, 314, 86, 0, 0, 
    464, 790, 625, 535, 650, 886, 809, 594, 422, 532, 700, 631, 370, 136, 0, 0, 
    671, 1060, 795, 573, 719, 1031, 1021, 819, 623, 676, 852, 719, 410, 248, 63, 0, 
    749, 1171, 821, 490, 644, 1009, 1146, 953, 743, 794, 957, 745, 453, 366, 206, 36, 
    845, 1322, 978, 566, 630, 884, 1060, 877, 660, 698, 782, 583, 391, 331, 243, 73, 
    959, 1509, 1198, 824, 703, 765, 845, 783, 624, 572, 517, 345, 244, 276, 200, 46, 
    998, 1575, 1390, 1193, 1052, 985, 915, 926, 808, 523, 312, 271, 305, 383, 305, 127, 
    954, 1548, 1549, 1542, 1538, 1312, 1114, 1103, 909, 618, 456, 495, 622, 711, 614, 365, 
    849, 1471, 1628, 1771, 1794, 1416, 1090, 1019, 884, 730, 722, 847, 971, 1041, 971, 670, 
    749, 1368, 1576, 1752, 1682, 1259, 953, 909, 864, 868, 959, 1074, 1154, 1219, 1186, 875, 
    688, 1269, 1371, 1498, 1355, 1036, 903, 906, 925, 993, 1071, 1140, 1239, 1332, 1260, 874, 
    654, 1141, 1133, 1140, 970, 823, 823, 857, 927, 1029, 1073, 1126, 1246, 1356, 1220, 763, 
    388, 622, 583, 539, 440, 397, 424, 458, 515, 586, 603, 626, 718, 809, 676, 378, 
    
    -- channel=3
    79, 52, 54, 54, 59, 67, 60, 47, 53, 56, 57, 49, 48, 45, 59, 24, 
    70, 32, 37, 35, 54, 58, 23, 5, 43, 61, 52, 28, 21, 33, 52, 15, 
    74, 36, 38, 37, 54, 64, 20, 22, 45, 72, 32, 0, 0, 14, 53, 10, 
    89, 34, 42, 45, 92, 75, 18, 4, 36, 99, 44, 13, 3, 5, 54, 11, 
    117, 15, 0, 59, 82, 32, 23, 14, 47, 105, 64, 0, 11, 27, 51, 15, 
    150, 31, 0, 52, 86, 61, 48, 1, 34, 111, 48, 0, 21, 26, 35, 8, 
    170, 38, 0, 49, 103, 76, 54, 0, 27, 109, 19, 0, 26, 35, 31, 0, 
    178, 49, 0, 16, 101, 67, 5, 0, 25, 85, 2, 0, 28, 39, 31, 0, 
    180, 42, 0, 25, 46, 56, 2, 25, 35, 47, 1, 2, 30, 49, 36, 0, 
    186, 44, 0, 59, 55, 53, 43, 51, 0, 0, 5, 21, 71, 58, 55, 0, 
    179, 44, 29, 98, 20, 0, 37, 35, 0, 2, 28, 38, 50, 18, 14, 0, 
    165, 15, 48, 136, 5, 0, 32, 18, 0, 26, 40, 62, 52, 25, 41, 0, 
    163, 49, 68, 111, 0, 0, 44, 25, 37, 67, 84, 77, 70, 72, 100, 0, 
    159, 68, 95, 47, 0, 30, 69, 59, 69, 77, 74, 74, 79, 98, 94, 0, 
    161, 66, 83, 28, 0, 72, 57, 56, 74, 72, 58, 75, 91, 74, 54, 0, 
    115, 43, 46, 23, 15, 53, 39, 46, 57, 42, 32, 61, 75, 31, 15, 0, 
    
    -- channel=4
    242, 252, 273, 277, 291, 285, 269, 285, 268, 248, 226, 223, 236, 241, 248, 97, 
    451, 561, 572, 575, 606, 594, 559, 545, 528, 463, 399, 396, 432, 473, 484, 211, 
    423, 539, 569, 584, 630, 643, 573, 483, 457, 416, 365, 339, 361, 410, 483, 216, 
    346, 455, 569, 612, 622, 582, 498, 377, 378, 441, 415, 359, 337, 359, 445, 217, 
    267, 399, 523, 610, 544, 469, 433, 346, 394, 462, 418, 380, 319, 304, 360, 193, 
    328, 483, 556, 676, 682, 640, 515, 403, 387, 426, 422, 378, 328, 286, 310, 133, 
    381, 501, 553, 660, 696, 713, 575, 486, 425, 487, 483, 394, 357, 304, 320, 127, 
    376, 443, 485, 517, 592, 665, 631, 546, 501, 565, 541, 411, 371, 380, 419, 187, 
    398, 429, 428, 425, 529, 660, 662, 539, 507, 580, 537, 438, 405, 444, 504, 241, 
    448, 487, 462, 433, 464, 510, 517, 433, 405, 449, 433, 327, 324, 394, 487, 220, 
    457, 531, 501, 490, 406, 341, 402, 396, 345, 278, 208, 113, 151, 227, 302, 96, 
    381, 483, 548, 598, 487, 397, 355, 339, 251, 106, 21, 0, 33, 74, 108, 0, 
    255, 369, 562, 644, 501, 328, 202, 151, 90, 17, 0, 0, 0, 0, 9, 0, 
    86, 192, 468, 536, 330, 149, 20, 0, 0, 0, 0, 0, 0, 0, 31, 0, 
    13, 44, 297, 345, 238, 102, 30, 23, 22, 14, 13, 44, 42, 24, 43, 0, 
    44, 59, 152, 182, 161, 103, 86, 87, 94, 93, 73, 90, 125, 123, 82, 0, 
    
    -- channel=5
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    66, 16, 0, 0, 0, 17, 0, 0, 0, 37, 21, 0, 0, 0, 0, 0, 
    67, 22, 11, 0, 30, 31, 0, 0, 11, 79, 30, 0, 0, 0, 0, 0, 
    108, 15, 0, 0, 48, 32, 0, 0, 8, 102, 59, 0, 0, 0, 0, 0, 
    152, 4, 0, 0, 74, 0, 0, 0, 0, 102, 81, 0, 0, 0, 0, 0, 
    241, 25, 0, 0, 127, 44, 0, 0, 0, 104, 74, 0, 0, 0, 0, 0, 
    276, 35, 0, 0, 130, 130, 26, 0, 0, 112, 44, 0, 0, 7, 0, 0, 
    303, 29, 0, 0, 99, 129, 29, 0, 8, 85, 10, 0, 0, 35, 0, 0, 
    328, 39, 0, 0, 82, 69, 15, 0, 4, 38, 6, 0, 0, 45, 0, 0, 
    337, 84, 0, 0, 48, 12, 24, 21, 0, 0, 0, 0, 36, 52, 0, 0, 
    326, 116, 18, 79, 12, 0, 37, 46, 0, 0, 10, 51, 79, 73, 17, 0, 
    305, 151, 113, 191, 28, 0, 72, 87, 14, 25, 74, 115, 119, 95, 70, 0, 
    289, 182, 221, 215, 0, 0, 77, 96, 84, 107, 135, 137, 131, 133, 116, 0, 
    244, 211, 253, 150, 0, 0, 94, 90, 107, 130, 135, 132, 153, 164, 128, 0, 
    204, 171, 206, 118, 25, 61, 100, 93, 116, 119, 106, 117, 170, 145, 67, 0, 
    166, 120, 126, 106, 85, 103, 110, 122, 140, 125, 103, 150, 192, 127, 52, 0, 
    
    -- channel=6
    0, 31, 23, 27, 6, 7, 66, 51, 29, 19, 25, 29, 19, 17, 14, 113, 
    0, 4, 6, 11, 0, 0, 97, 68, 0, 0, 41, 74, 60, 15, 0, 154, 
    0, 13, 0, 10, 1, 0, 68, 99, 11, 0, 82, 121, 103, 43, 0, 152, 
    0, 63, 55, 0, 5, 71, 115, 160, 74, 0, 85, 177, 125, 81, 0, 127, 
    0, 111, 163, 2, 0, 175, 178, 212, 123, 0, 93, 212, 130, 92, 33, 119, 
    0, 157, 253, 86, 0, 138, 175, 248, 178, 0, 124, 249, 124, 66, 78, 157, 
    0, 192, 278, 156, 0, 35, 187, 263, 201, 0, 132, 260, 119, 57, 96, 203, 
    0, 217, 290, 191, 12, 0, 181, 227, 176, 24, 105, 219, 107, 37, 67, 207, 
    0, 245, 319, 202, 115, 51, 104, 156, 167, 79, 97, 166, 58, 3, 26, 204, 
    0, 236, 309, 164, 192, 191, 89, 130, 218, 137, 65, 79, 25, 2, 20, 227, 
    0, 199, 270, 132, 253, 349, 138, 135, 228, 162, 80, 73, 42, 39, 45, 287, 
    0, 130, 192, 133, 348, 414, 193, 148, 195, 162, 119, 118, 120, 122, 113, 380, 
    0, 115, 91, 168, 418, 370, 212, 170, 174, 175, 163, 178, 196, 187, 177, 449, 
    0, 155, 73, 184, 402, 302, 200, 190, 168, 176, 198, 184, 183, 217, 249, 453, 
    0, 207, 121, 186, 295, 206, 159, 158, 132, 162, 209, 169, 147, 230, 298, 429, 
    55, 184, 145, 150, 177, 144, 128, 135, 125, 149, 182, 164, 144, 202, 249, 264, 
    
    -- channel=7
    44, 43, 52, 54, 54, 95, 101, 64, 40, 41, 51, 47, 34, 28, 21, 17, 
    51, 54, 46, 47, 53, 123, 139, 67, 23, 90, 157, 154, 93, 29, 0, 6, 
    72, 70, 53, 50, 80, 120, 165, 104, 80, 189, 300, 261, 164, 51, 6, 19, 
    187, 210, 145, 118, 195, 250, 244, 208, 166, 256, 404, 346, 221, 96, 8, 15, 
    347, 437, 314, 194, 330, 447, 425, 350, 251, 312, 432, 386, 239, 144, 45, 4, 
    501, 639, 445, 279, 369, 553, 545, 461, 330, 382, 515, 428, 256, 187, 116, 46, 
    567, 728, 478, 300, 303, 542, 625, 534, 395, 456, 570, 449, 279, 237, 182, 98, 
    608, 821, 573, 340, 310, 493, 598, 494, 387, 400, 472, 366, 260, 227, 182, 112, 
    654, 917, 715, 480, 424, 436, 490, 458, 397, 353, 331, 263, 180, 175, 142, 89, 
    663, 958, 809, 683, 651, 537, 503, 566, 489, 351, 250, 227, 239, 262, 233, 161, 
    654, 985, 869, 865, 900, 773, 664, 715, 641, 465, 383, 413, 473, 503, 469, 343, 
    636, 954, 934, 1034, 1122, 947, 778, 750, 682, 600, 599, 693, 762, 783, 782, 582, 
    676, 957, 1005, 1140, 1106, 898, 771, 741, 721, 753, 817, 895, 943, 981, 1009, 755, 
    690, 986, 985, 1065, 966, 826, 778, 766, 779, 838, 899, 936, 999, 1078, 1089, 754, 
    696, 989, 936, 911, 818, 746, 749, 755, 797, 873, 917, 930, 1016, 1121, 1078, 690, 
    448, 637, 571, 521, 463, 444, 457, 477, 513, 560, 575, 599, 664, 724, 649, 377, 
    
    -- channel=8
    186, 202, 233, 236, 244, 255, 258, 254, 232, 217, 205, 198, 196, 196, 201, 134, 
    299, 352, 393, 397, 418, 427, 427, 393, 356, 319, 317, 319, 314, 324, 312, 183, 
    284, 332, 379, 406, 427, 434, 423, 360, 325, 309, 306, 309, 294, 289, 300, 176, 
    269, 335, 419, 452, 474, 458, 402, 344, 306, 302, 307, 312, 288, 271, 289, 151, 
    274, 345, 432, 448, 452, 451, 389, 339, 343, 325, 340, 349, 278, 256, 255, 133, 
    272, 385, 485, 487, 458, 495, 456, 401, 388, 356, 343, 359, 284, 246, 254, 130, 
    304, 397, 498, 486, 446, 502, 513, 454, 428, 377, 372, 371, 304, 243, 281, 149, 
    302, 394, 468, 455, 444, 460, 475, 444, 434, 404, 374, 356, 302, 260, 310, 196, 
    311, 380, 461, 417, 438, 448, 456, 434, 437, 405, 362, 329, 277, 298, 363, 226, 
    317, 384, 471, 438, 449, 464, 440, 407, 410, 394, 301, 259, 270, 306, 365, 212, 
    311, 407, 491, 468, 461, 462, 397, 351, 358, 284, 210, 168, 196, 237, 279, 152, 
    240, 366, 520, 535, 474, 423, 302, 240, 234, 171, 106, 79, 118, 145, 170, 96, 
    154, 260, 477, 521, 432, 329, 204, 143, 110, 70, 50, 53, 67, 75, 88, 61, 
    65, 172, 365, 391, 310, 186, 82, 57, 49, 44, 46, 56, 68, 82, 86, 65, 
    19, 93, 230, 239, 213, 120, 64, 72, 74, 77, 81, 94, 108, 108, 109, 56, 
    0, 0, 59, 60, 66, 34, 7, 19, 16, 8, 10, 22, 15, 14, 9, 22, 
    
    -- channel=9
    0, 0, 0, 0, 0, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 0, 2, 16, 73, 61, 0, 0, 46, 90, 69, 7, 0, 0, 0, 
    0, 9, 0, 7, 38, 88, 118, 51, 25, 121, 210, 167, 71, 0, 0, 0, 
    76, 101, 72, 67, 150, 199, 173, 113, 75, 177, 311, 238, 122, 11, 0, 0, 
    190, 287, 188, 141, 267, 329, 282, 219, 140, 243, 346, 266, 137, 45, 0, 0, 
    310, 451, 299, 211, 322, 463, 424, 324, 213, 295, 399, 292, 152, 105, 0, 0, 
    352, 528, 335, 186, 288, 504, 510, 386, 281, 352, 465, 320, 182, 149, 64, 25, 
    403, 588, 392, 196, 236, 416, 489, 367, 286, 311, 400, 265, 150, 147, 84, 60, 
    472, 681, 500, 310, 291, 340, 424, 367, 283, 241, 257, 177, 102, 121, 77, 46, 
    495, 762, 596, 494, 457, 385, 387, 411, 320, 201, 144, 121, 126, 155, 101, 65, 
    482, 773, 649, 647, 670, 521, 436, 488, 399, 261, 197, 220, 265, 302, 248, 155, 
    444, 727, 732, 782, 825, 625, 516, 519, 434, 342, 331, 393, 457, 490, 447, 323, 
    427, 692, 751, 840, 815, 589, 493, 473, 446, 444, 480, 540, 571, 607, 582, 450, 
    398, 658, 684, 755, 672, 501, 462, 455, 464, 501, 540, 571, 623, 668, 631, 462, 
    381, 621, 614, 608, 519, 435, 444, 450, 479, 531, 553, 571, 639, 699, 622, 425, 
    242, 431, 396, 366, 309, 287, 304, 318, 343, 379, 384, 399, 451, 498, 431, 278, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 24, 0, 0, 34, 65, 36, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 79, 145, 83, 33, 0, 0, 
    0, 101, 32, 0, 0, 44, 64, 92, 40, 0, 78, 149, 88, 34, 5, 0, 
    0, 213, 167, 30, 0, 172, 174, 167, 67, 8, 111, 169, 101, 31, 33, 0, 
    0, 255, 205, 47, 18, 107, 170, 209, 96, 59, 161, 207, 103, 40, 59, 26, 
    0, 288, 228, 57, 0, 28, 181, 238, 119, 98, 153, 187, 93, 46, 66, 32, 
    0, 346, 257, 150, 56, 70, 156, 181, 89, 81, 110, 133, 78, 26, 43, 4, 
    0, 379, 258, 203, 116, 130, 88, 101, 128, 94, 82, 71, 44, 14, 37, 16, 
    0, 355, 253, 223, 213, 237, 159, 203, 266, 190, 102, 81, 71, 90, 114, 86, 
    0, 316, 254, 254, 361, 418, 315, 295, 303, 240, 158, 163, 205, 222, 230, 222, 
    34, 334, 242, 317, 472, 450, 325, 279, 270, 248, 251, 287, 310, 324, 350, 341, 
    46, 357, 272, 344, 486, 393, 285, 273, 255, 262, 292, 308, 319, 341, 395, 390, 
    49, 370, 318, 346, 411, 331, 280, 277, 257, 275, 310, 313, 299, 362, 429, 395, 
    53, 332, 301, 290, 270, 236, 222, 230, 237, 272, 303, 295, 292, 373, 422, 328, 
    
    -- channel=11
    57, 66, 67, 67, 68, 52, 57, 53, 65, 51, 46, 46, 51, 56, 41, 25, 
    3, 4, 6, 7, 17, 0, 0, 0, 13, 0, 0, 0, 0, 3, 0, 0, 
    12, 3, 13, 8, 18, 4, 2, 7, 3, 3, 0, 0, 0, 6, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    22, 0, 0, 29, 11, 6, 0, 0, 13, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 14, 0, 16, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 3, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 2, 0, 0, 
    0, 0, 10, 2, 0, 0, 0, 0, 0, 0, 0, 7, 25, 6, 3, 0, 
    0, 0, 15, 18, 0, 1, 0, 0, 23, 21, 20, 32, 36, 32, 23, 0, 
    46, 17, 19, 0, 0, 21, 23, 17, 30, 42, 25, 16, 22, 25, 5, 0, 
    23, 43, 6, 0, 0, 0, 0, 0, 0, 2, 12, 11, 17, 17, 5, 8, 
    20, 13, 14, 0, 0, 6, 0, 8, 7, 8, 10, 15, 18, 6, 0, 4, 
    13, 0, 0, 0, 4, 17, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 20, 8, 0, 0, 8, 10, 18, 24, 32, 34, 40, 33, 37, 44, 29, 
    
    -- channel=12
    173, 273, 278, 277, 282, 301, 303, 288, 264, 248, 231, 221, 222, 228, 224, 191, 
    246, 373, 390, 395, 405, 428, 436, 385, 337, 325, 316, 306, 292, 297, 317, 251, 
    223, 356, 393, 400, 404, 434, 429, 349, 299, 297, 338, 312, 280, 270, 288, 252, 
    226, 364, 408, 446, 454, 467, 416, 326, 256, 284, 344, 317, 272, 229, 242, 235, 
    227, 386, 448, 479, 484, 500, 455, 354, 277, 306, 351, 345, 272, 212, 217, 190, 
    219, 414, 478, 463, 457, 516, 495, 406, 338, 313, 387, 369, 270, 232, 219, 174, 
    239, 428, 467, 425, 408, 491, 516, 456, 354, 320, 409, 359, 266, 252, 262, 215, 
    254, 441, 453, 383, 382, 439, 501, 437, 350, 334, 411, 337, 268, 265, 309, 257, 
    273, 473, 443, 386, 361, 407, 456, 407, 343, 351, 360, 297, 230, 280, 342, 284, 
    285, 475, 454, 420, 436, 444, 398, 385, 381, 343, 301, 220, 188, 259, 322, 275, 
    261, 451, 473, 444, 517, 453, 353, 349, 318, 245, 184, 117, 132, 209, 249, 215, 
    185, 375, 459, 478, 550, 406, 255, 235, 204, 150, 83, 72, 91, 133, 155, 160, 
    86, 231, 366, 493, 490, 265, 136, 102, 79, 47, 39, 43, 57, 72, 75, 138, 
    5, 126, 235, 393, 338, 136, 68, 56, 48, 41, 39, 45, 67, 68, 85, 146, 
    0, 45, 137, 224, 155, 71, 49, 50, 55, 64, 65, 69, 82, 101, 112, 127, 
    0, 19, 54, 88, 46, 21, 20, 25, 34, 47, 46, 37, 47, 74, 72, 60, 
    
    -- channel=13
    68, 52, 50, 54, 66, 91, 82, 64, 31, 29, 40, 41, 34, 26, 25, 0, 
    0, 14, 12, 15, 38, 71, 46, 7, 0, 41, 106, 96, 43, 11, 0, 0, 
    0, 12, 11, 16, 20, 42, 72, 42, 40, 112, 180, 155, 87, 22, 0, 0, 
    75, 144, 104, 93, 115, 140, 156, 118, 89, 144, 222, 211, 127, 39, 2, 0, 
    166, 282, 197, 142, 181, 259, 265, 222, 141, 171, 249, 226, 143, 82, 19, 0, 
    219, 378, 254, 130, 166, 323, 350, 297, 190, 215, 290, 255, 163, 123, 80, 22, 
    235, 411, 287, 128, 130, 314, 367, 325, 227, 242, 325, 265, 169, 158, 136, 59, 
    274, 486, 360, 197, 157, 238, 306, 284, 208, 202, 253, 212, 138, 128, 135, 69, 
    303, 560, 438, 294, 223, 198, 251, 289, 207, 157, 152, 124, 101, 98, 104, 47, 
    296, 563, 495, 437, 403, 314, 320, 358, 275, 162, 117, 127, 140, 158, 140, 81, 
    286, 543, 531, 548, 568, 470, 364, 389, 355, 275, 233, 270, 279, 294, 291, 213, 
    277, 534, 555, 607, 622, 514, 412, 418, 410, 374, 371, 418, 443, 463, 491, 370, 
    268, 542, 566, 602, 575, 503, 420, 407, 419, 446, 473, 512, 532, 560, 596, 443, 
    287, 519, 524, 538, 516, 484, 448, 443, 449, 479, 506, 534, 575, 625, 620, 442, 
    307, 516, 458, 468, 462, 410, 409, 418, 446, 487, 501, 519, 572, 619, 590, 398, 
    137, 307, 257, 244, 239, 215, 223, 235, 248, 267, 276, 281, 303, 340, 327, 238, 
    
    -- channel=14
    294, 415, 413, 412, 427, 452, 437, 422, 396, 376, 350, 333, 337, 343, 359, 227, 
    395, 590, 603, 603, 644, 688, 630, 563, 518, 508, 488, 449, 440, 470, 514, 306, 
    349, 562, 597, 616, 665, 679, 597, 485, 473, 525, 490, 422, 383, 403, 494, 304, 
    319, 553, 610, 675, 717, 692, 602, 467, 440, 502, 502, 414, 352, 349, 441, 284, 
    369, 550, 599, 725, 776, 722, 590, 460, 407, 514, 538, 438, 354, 330, 363, 238, 
    383, 566, 595, 725, 765, 714, 627, 504, 459, 579, 559, 425, 363, 338, 353, 198, 
    426, 576, 546, 656, 691, 760, 705, 557, 501, 583, 545, 404, 371, 379, 400, 208, 
    447, 554, 493, 582, 674, 768, 674, 539, 524, 585, 560, 410, 390, 407, 454, 260, 
    483, 564, 472, 503, 623, 636, 597, 539, 530, 549, 520, 386, 362, 447, 528, 314, 
    493, 593, 484, 540, 587, 570, 586, 571, 496, 468, 400, 305, 340, 411, 515, 284, 
    459, 587, 538, 650, 652, 536, 533, 475, 351, 257, 240, 200, 222, 278, 357, 166, 
    357, 505, 627, 750, 615, 381, 312, 260, 184, 136, 120, 93, 107, 134, 198, 18, 
    210, 332, 600, 715, 471, 229, 144, 111, 66, 38, 28, 28, 22, 33, 103, 0, 
    68, 180, 451, 511, 284, 109, 38, 15, 22, 23, 12, 11, 20, 52, 94, 0, 
    21, 54, 239, 253, 122, 58, 35, 35, 56, 56, 31, 46, 99, 94, 69, 0, 
    13, 0, 54, 48, 29, 15, 7, 19, 37, 27, 0, 33, 65, 32, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 18, 33, 26, 0, 11, 9, 10, 12, 10, 11, 26, 22, 19, 16, 4, 
    
    -- channel=16
    127, 71, 77, 77, 92, 124, 97, 69, 61, 62, 71, 63, 60, 57, 44, 0, 
    223, 132, 134, 132, 162, 195, 151, 83, 111, 165, 166, 134, 109, 96, 101, 0, 
    241, 150, 153, 140, 169, 194, 142, 84, 137, 215, 200, 134, 105, 94, 109, 0, 
    322, 213, 179, 210, 291, 265, 167, 102, 154, 265, 224, 121, 75, 83, 112, 0, 
    394, 269, 215, 239, 336, 283, 232, 141, 159, 300, 251, 117, 74, 82, 97, 0, 
    452, 279, 180, 224, 337, 282, 258, 163, 179, 333, 285, 111, 91, 104, 106, 4, 
    495, 291, 171, 187, 346, 343, 265, 160, 186, 342, 268, 96, 106, 133, 98, 0, 
    528, 296, 179, 163, 306, 367, 260, 143, 168, 285, 212, 75, 100, 155, 116, 0, 
    569, 305, 215, 185, 274, 304, 235, 188, 182, 228, 148, 51, 93, 156, 120, 0, 
    571, 319, 254, 308, 323, 291, 280, 255, 200, 135, 120, 103, 154, 204, 171, 8, 
    558, 345, 318, 420, 365, 239, 295, 271, 170, 127, 129, 148, 216, 238, 211, 14, 
    512, 341, 380, 525, 352, 166, 206, 204, 115, 109, 171, 215, 242, 243, 248, 28, 
    454, 328, 418, 510, 280, 86, 154, 177, 152, 165, 206, 221, 229, 249, 263, 20, 
    383, 299, 402, 363, 163, 81, 159, 167, 184, 208, 214, 224, 261, 276, 256, 0, 
    355, 242, 330, 237, 78, 107, 156, 162, 207, 227, 213, 239, 294, 288, 214, 0, 
    150, 43, 84, 54, 0, 16, 37, 37, 59, 53, 34, 62, 108, 68, 0, 0, 
    
    -- channel=17
    47, 232, 194, 197, 191, 224, 277, 240, 199, 184, 193, 187, 163, 160, 169, 220, 
    0, 236, 200, 206, 181, 228, 359, 276, 178, 186, 282, 291, 236, 184, 177, 304, 
    12, 249, 197, 208, 160, 190, 362, 329, 166, 162, 331, 368, 299, 194, 149, 312, 
    79, 383, 321, 265, 277, 387, 443, 418, 180, 121, 357, 454, 353, 230, 144, 284, 
    108, 527, 484, 294, 361, 563, 520, 506, 279, 147, 423, 523, 359, 269, 190, 259, 
    88, 631, 608, 261, 233, 512, 581, 632, 411, 192, 482, 571, 338, 278, 266, 292, 
    75, 693, 699, 299, 157, 388, 617, 667, 419, 216, 512, 581, 329, 263, 325, 348, 
    96, 771, 756, 446, 222, 264, 541, 564, 350, 214, 428, 508, 277, 208, 300, 392, 
    88, 827, 769, 550, 314, 282, 431, 512, 420, 282, 348, 394, 198, 172, 269, 397, 
    58, 805, 754, 600, 569, 535, 454, 539, 567, 378, 277, 290, 226, 243, 314, 464, 
    19, 745, 722, 622, 848, 787, 466, 515, 617, 487, 361, 340, 305, 349, 412, 572, 
    0, 621, 595, 626, 963, 866, 489, 473, 557, 480, 399, 393, 416, 460, 505, 726, 
    12, 538, 464, 649, 1011, 807, 514, 457, 480, 459, 452, 487, 521, 542, 587, 865, 
    92, 491, 376, 645, 922, 688, 506, 479, 450, 462, 494, 504, 536, 590, 651, 880, 
    167, 534, 365, 569, 701, 495, 432, 436, 421, 477, 528, 493, 513, 641, 710, 821, 
    65, 306, 208, 265, 300, 220, 206, 207, 195, 244, 289, 221, 220, 349, 431, 479, 
    
    -- channel=18
    105, 107, 97, 96, 91, 95, 109, 91, 86, 71, 69, 76, 82, 88, 88, 50, 
    107, 100, 91, 90, 81, 101, 115, 79, 43, 36, 49, 52, 63, 69, 88, 52, 
    91, 88, 92, 89, 84, 72, 68, 30, 12, 33, 55, 66, 65, 67, 80, 52, 
    59, 81, 85, 64, 54, 52, 43, 47, 36, 50, 74, 63, 38, 69, 82, 46, 
    67, 107, 120, 61, 84, 78, 45, 76, 29, 25, 68, 65, 31, 59, 85, 32, 
    84, 89, 124, 33, 66, 42, 54, 79, 27, 28, 90, 66, 26, 43, 85, 51, 
    80, 81, 106, 6, 53, 30, 56, 76, 27, 37, 89, 49, 23, 59, 97, 65, 
    74, 54, 87, 21, 59, 63, 84, 60, 40, 60, 78, 56, 38, 77, 106, 55, 
    84, 50, 63, 27, 78, 57, 24, 25, 44, 58, 65, 36, 31, 75, 104, 54, 
    100, 39, 36, 4, 43, 50, 0, 31, 84, 31, 24, 13, 20, 57, 63, 44, 
    86, 28, 17, 12, 94, 73, 22, 44, 59, 0, 0, 0, 6, 15, 8, 42, 
    58, 21, 16, 55, 91, 19, 0, 0, 0, 0, 0, 1, 7, 0, 0, 69, 
    53, 9, 0, 45, 61, 0, 0, 0, 0, 0, 6, 11, 5, 0, 22, 95, 
    41, 8, 0, 36, 51, 0, 10, 9, 1, 5, 11, 0, 0, 1, 40, 84, 
    64, 11, 8, 23, 17, 0, 21, 16, 12, 25, 25, 6, 15, 36, 55, 64, 
    83, 26, 25, 19, 24, 13, 27, 27, 27, 36, 37, 35, 41, 48, 45, 27, 
    
    -- channel=19
    308, 188, 161, 157, 205, 201, 113, 112, 145, 145, 124, 113, 133, 146, 149, 0, 
    407, 279, 229, 221, 318, 277, 79, 89, 238, 268, 143, 71, 102, 189, 229, 0, 
    388, 296, 249, 225, 277, 275, 112, 59, 245, 319, 100, 15, 13, 144, 264, 0, 
    421, 258, 200, 344, 316, 213, 85, 0, 180, 356, 149, 0, 0, 104, 267, 42, 
    503, 191, 61, 377, 334, 54, 0, 0, 154, 407, 176, 0, 7, 68, 172, 61, 
    545, 150, 0, 261, 404, 200, 69, 0, 111, 386, 115, 0, 34, 101, 104, 0, 
    582, 107, 0, 169, 495, 365, 68, 0, 69, 342, 79, 0, 58, 138, 72, 0, 
    593, 61, 0, 82, 378, 336, 8, 0, 88, 286, 114, 0, 80, 177, 140, 0, 
    619, 56, 0, 37, 146, 215, 191, 92, 75, 159, 98, 0, 172, 257, 198, 0, 
    651, 75, 0, 161, 64, 89, 241, 81, 0, 0, 82, 126, 230, 214, 162, 0, 
    665, 99, 70, 277, 0, 0, 54, 29, 0, 0, 85, 123, 126, 95, 70, 0, 
    574, 197, 216, 245, 0, 0, 0, 12, 0, 0, 58, 62, 37, 34, 59, 0, 
    446, 236, 350, 143, 0, 0, 0, 12, 20, 38, 48, 21, 0, 28, 48, 0, 
    353, 155, 292, 84, 0, 0, 0, 0, 31, 27, 0, 24, 58, 15, 0, 0, 
    329, 36, 104, 54, 0, 0, 21, 32, 68, 22, 0, 58, 122, 0, 0, 0, 
    180, 6, 21, 33, 10, 31, 37, 37, 51, 18, 0, 30, 64, 0, 0, 0, 
    
    -- channel=20
    38, 36, 16, 15, 17, 32, 43, 0, 7, 13, 30, 26, 16, 10, 0, 0, 
    42, 45, 10, 8, 24, 60, 56, 0, 0, 48, 99, 70, 47, 13, 0, 0, 
    59, 56, 23, 7, 23, 47, 56, 30, 46, 119, 168, 123, 67, 28, 10, 12, 
    134, 138, 79, 13, 90, 92, 91, 78, 75, 120, 212, 146, 79, 60, 8, 22, 
    246, 247, 153, 89, 214, 218, 142, 137, 80, 147, 256, 145, 78, 73, 30, 24, 
    279, 315, 200, 87, 195, 256, 225, 187, 123, 203, 275, 162, 87, 107, 69, 28, 
    293, 327, 204, 91, 103, 259, 289, 201, 164, 206, 284, 163, 100, 136, 92, 29, 
    331, 372, 233, 143, 148, 233, 263, 165, 175, 176, 214, 153, 91, 115, 82, 34, 
    351, 432, 302, 196, 217, 158, 194, 186, 164, 123, 135, 95, 77, 99, 62, 26, 
    333, 455, 332, 276, 303, 198, 214, 272, 224, 126, 89, 110, 134, 143, 115, 79, 
    325, 469, 374, 402, 461, 332, 285, 340, 274, 199, 215, 244, 263, 278, 249, 187, 
    326, 486, 443, 482, 499, 358, 321, 350, 327, 307, 327, 372, 391, 388, 392, 285, 
    336, 479, 500, 522, 482, 326, 329, 336, 339, 373, 407, 440, 449, 472, 497, 364, 
    341, 490, 489, 508, 431, 334, 373, 367, 379, 410, 431, 441, 483, 528, 509, 355, 
    356, 495, 440, 443, 374, 339, 379, 381, 402, 434, 436, 439, 519, 546, 486, 311, 
    214, 298, 264, 235, 210, 199, 218, 228, 251, 272, 270, 284, 321, 346, 301, 175, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 101, 82, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 18, 11, 0, 58, 160, 126, 53, 0, 0, 0, 
    179, 173, 34, 0, 96, 163, 164, 132, 29, 84, 179, 139, 73, 0, 0, 0, 
    268, 280, 127, 0, 77, 218, 238, 206, 94, 134, 231, 162, 79, 56, 0, 0, 
    293, 313, 157, 0, 0, 205, 274, 239, 140, 181, 258, 168, 83, 87, 50, 0, 
    347, 411, 229, 36, 1, 170, 241, 175, 110, 105, 183, 111, 59, 57, 24, 0, 
    378, 506, 344, 191, 97, 97, 160, 151, 109, 52, 57, 42, 5, 0, 0, 0, 
    362, 531, 426, 342, 283, 164, 194, 267, 195, 65, 9, 24, 40, 43, 11, 0, 
    341, 532, 475, 481, 509, 375, 313, 367, 301, 189, 151, 209, 238, 234, 210, 118, 
    339, 509, 503, 564, 609, 479, 383, 385, 362, 339, 367, 437, 468, 475, 487, 318, 
    373, 510, 518, 577, 575, 471, 411, 417, 433, 477, 523, 574, 600, 632, 675, 459, 
    439, 541, 509, 540, 510, 486, 489, 493, 506, 544, 576, 604, 644, 686, 702, 456, 
    474, 599, 510, 468, 434, 437, 467, 477, 517, 569, 583, 595, 662, 727, 680, 409, 
    307, 402, 331, 283, 256, 260, 283, 297, 326, 363, 374, 380, 430, 470, 433, 243, 
    
    -- channel=22
    37, 77, 76, 76, 65, 66, 87, 96, 87, 90, 79, 81, 79, 72, 82, 87, 
    56, 107, 115, 115, 94, 130, 151, 148, 116, 85, 98, 109, 109, 116, 100, 126, 
    57, 116, 116, 119, 119, 153, 170, 139, 98, 91, 101, 110, 99, 90, 102, 127, 
    8, 102, 123, 114, 90, 136, 177, 135, 68, 74, 107, 133, 126, 79, 96, 122, 
    7, 89, 111, 109, 123, 120, 128, 125, 75, 63, 137, 149, 112, 86, 73, 131, 
    20, 122, 184, 130, 165, 156, 135, 151, 75, 65, 127, 145, 104, 79, 69, 98, 
    11, 141, 201, 127, 116, 127, 184, 186, 100, 88, 136, 154, 102, 80, 87, 97, 
    4, 127, 160, 151, 97, 169, 192, 186, 128, 116, 166, 153, 106, 84, 95, 126, 
    13, 117, 133, 133, 112, 161, 173, 143, 168, 139, 182, 169, 85, 80, 115, 146, 
    30, 114, 129, 79, 106, 109, 118, 133, 143, 154, 122, 81, 50, 72, 103, 153, 
    18, 116, 103, 67, 127, 125, 104, 113, 126, 85, 58, 48, 21, 53, 81, 138, 
    6, 95, 98, 110, 205, 194, 109, 115, 107, 51, 4, 0, 0, 4, 5, 98, 
    0, 55, 82, 158, 220, 150, 43, 30, 20, 0, 0, 0, 0, 0, 0, 87, 
    0, 0, 88, 150, 167, 66, 0, 0, 0, 0, 0, 0, 0, 0, 4, 121, 
    0, 0, 14, 121, 115, 25, 9, 0, 0, 0, 0, 0, 0, 0, 6, 105, 
    50, 19, 31, 71, 70, 44, 46, 49, 53, 64, 56, 38, 61, 74, 58, 73, 
    
    -- channel=23
    236, 300, 329, 328, 346, 334, 310, 317, 309, 287, 259, 253, 270, 271, 251, 99, 
    442, 621, 678, 677, 734, 736, 677, 645, 619, 561, 493, 451, 462, 512, 508, 236, 
    393, 601, 691, 698, 764, 789, 693, 578, 541, 557, 507, 462, 410, 447, 486, 242, 
    307, 492, 632, 716, 721, 687, 617, 477, 467, 555, 552, 496, 399, 370, 412, 224, 
    333, 484, 635, 800, 777, 705, 593, 459, 473, 567, 568, 497, 394, 310, 294, 152, 
    422, 634, 759, 898, 946, 945, 784, 567, 517, 584, 568, 517, 439, 328, 263, 79, 
    466, 647, 726, 830, 906, 987, 879, 697, 648, 689, 638, 568, 478, 399, 350, 119, 
    484, 598, 625, 650, 781, 939, 924, 808, 756, 787, 730, 597, 509, 489, 483, 219, 
    557, 655, 620, 582, 699, 845, 882, 745, 674, 709, 704, 558, 499, 526, 569, 283, 
    622, 756, 727, 655, 610, 636, 683, 588, 533, 544, 502, 385, 376, 438, 522, 250, 
    610, 786, 840, 797, 632, 593, 630, 609, 495, 360, 233, 144, 189, 288, 339, 104, 
    494, 719, 952, 968, 779, 657, 563, 491, 376, 195, 60, 12, 67, 141, 131, 0, 
    255, 526, 926, 985, 770, 498, 308, 194, 119, 37, 0, 0, 34, 47, 29, 0, 
    32, 257, 690, 767, 548, 271, 59, 7, 0, 0, 0, 29, 44, 38, 30, 0, 
    0, 70, 376, 443, 337, 188, 75, 75, 80, 69, 56, 107, 133, 100, 46, 0, 
    15, 85, 221, 236, 200, 148, 112, 141, 176, 184, 163, 201, 252, 244, 147, 13, 
    
    -- channel=24
    51, 94, 79, 81, 98, 133, 131, 82, 52, 57, 68, 56, 44, 35, 6, 0, 
    0, 17, 4, 3, 26, 85, 93, 0, 0, 56, 132, 117, 40, 0, 0, 0, 
    0, 34, 11, 6, 18, 89, 128, 52, 39, 165, 275, 234, 109, 0, 0, 0, 
    122, 213, 148, 115, 163, 227, 244, 176, 109, 228, 368, 332, 169, 17, 0, 0, 
    310, 457, 331, 213, 367, 502, 445, 346, 218, 262, 433, 367, 214, 70, 0, 0, 
    448, 632, 445, 224, 374, 611, 583, 487, 317, 346, 510, 409, 242, 154, 30, 5, 
    485, 696, 482, 205, 277, 569, 659, 559, 392, 423, 549, 429, 245, 227, 144, 47, 
    551, 809, 577, 304, 267, 452, 586, 489, 346, 345, 428, 331, 208, 189, 156, 67, 
    604, 945, 701, 484, 355, 370, 484, 439, 337, 264, 260, 207, 129, 148, 100, 41, 
    602, 992, 830, 719, 610, 512, 515, 551, 454, 275, 157, 165, 191, 222, 166, 107, 
    566, 980, 900, 912, 924, 767, 615, 658, 558, 384, 296, 342, 398, 427, 378, 282, 
    500, 941, 949, 1024, 1083, 853, 649, 636, 587, 505, 508, 587, 632, 666, 648, 496, 
    457, 870, 947, 1027, 1001, 796, 625, 587, 593, 626, 685, 751, 800, 836, 845, 660, 
    473, 805, 818, 914, 889, 720, 650, 645, 657, 702, 747, 798, 859, 919, 890, 665, 
    488, 787, 673, 740, 693, 605, 595, 612, 655, 715, 745, 770, 861, 931, 855, 600, 
    292, 502, 396, 383, 348, 326, 340, 364, 397, 451, 468, 467, 528, 596, 538, 389, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 24, 12, 13, 3, 26, 52, 44, 13, 22, 31, 33, 21, 10, 10, 67, 
    0, 0, 0, 0, 0, 10, 89, 55, 0, 0, 66, 97, 64, 0, 0, 29, 
    0, 11, 0, 0, 0, 24, 93, 87, 3, 32, 151, 192, 146, 50, 0, 35, 
    47, 149, 52, 12, 60, 142, 154, 157, 106, 119, 240, 286, 193, 105, 25, 30, 
    86, 327, 204, 77, 122, 300, 320, 275, 191, 174, 249, 325, 206, 123, 100, 40, 
    189, 478, 357, 204, 179, 340, 406, 375, 255, 217, 323, 358, 224, 115, 137, 82, 
    232, 563, 425, 243, 162, 284, 417, 440, 303, 274, 366, 378, 231, 143, 136, 142, 
    268, 611, 480, 301, 145, 250, 410, 408, 278, 257, 297, 311, 209, 143, 141, 136, 
    289, 646, 549, 401, 275, 302, 320, 343, 280, 270, 221, 215, 160, 97, 96, 109, 
    293, 668, 569, 479, 417, 407, 305, 351, 391, 291, 195, 162, 151, 146, 146, 162, 
    278, 652, 564, 537, 594, 587, 479, 447, 498, 397, 236, 238, 262, 283, 282, 306, 
    260, 617, 561, 666, 749, 766, 585, 512, 466, 410, 370, 409, 466, 486, 494, 515, 
    303, 627, 568, 723, 850, 732, 557, 508, 482, 484, 508, 573, 604, 626, 665, 679, 
    325, 660, 608, 726, 766, 641, 530, 521, 507, 532, 582, 603, 625, 689, 766, 705, 
    332, 709, 668, 649, 607, 543, 499, 507, 512, 565, 619, 609, 623, 743, 821, 673, 
    261, 472, 433, 394, 340, 329, 323, 326, 338, 375, 408, 405, 437, 507, 539, 391, 
    
    -- channel=27
    17, 28, 23, 21, 27, 5, 11, 13, 23, 14, 6, 11, 23, 24, 30, 0, 
    37, 48, 47, 46, 54, 24, 21, 40, 48, 19, 0, 0, 6, 35, 37, 0, 
    33, 60, 51, 49, 50, 47, 19, 12, 11, 0, 0, 0, 0, 31, 40, 0, 
    0, 0, 13, 44, 5, 0, 0, 0, 5, 19, 0, 0, 0, 3, 43, 6, 
    0, 0, 0, 47, 0, 0, 0, 0, 17, 6, 0, 0, 0, 0, 16, 2, 
    0, 0, 0, 58, 51, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 66, 9, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 17, 1, 2, 8, 7, 0, 0, 9, 12, 8, 0, 
    0, 0, 0, 0, 0, 26, 33, 0, 0, 0, 11, 9, 32, 22, 35, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 4, 0, 0, 4, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 22, 11, 12, 0, 14, 38, 37, 17, 17, 21, 21, 16, 18, 29, 67, 
    0, 7, 8, 8, 0, 4, 61, 58, 0, 2, 38, 55, 43, 17, 28, 81, 
    0, 14, 12, 11, 0, 0, 64, 51, 0, 0, 34, 71, 77, 26, 12, 86, 
    0, 54, 18, 0, 5, 7, 62, 63, 0, 0, 23, 69, 75, 46, 6, 76, 
    0, 73, 72, 0, 0, 41, 72, 95, 0, 0, 20, 85, 62, 66, 24, 52, 
    0, 45, 115, 0, 0, 0, 51, 111, 4, 0, 36, 99, 38, 50, 64, 74, 
    0, 53, 126, 3, 0, 0, 12, 100, 5, 0, 35, 105, 18, 22, 66, 95, 
    0, 57, 126, 59, 0, 0, 33, 73, 15, 0, 31, 81, 22, 0, 41, 108, 
    0, 47, 99, 61, 0, 0, 8, 63, 46, 0, 38, 45, 0, 0, 29, 102, 
    0, 13, 49, 20, 75, 25, 0, 35, 98, 61, 45, 43, 0, 14, 49, 131, 
    0, 2, 0, 0, 92, 113, 8, 29, 120, 85, 42, 25, 0, 32, 73, 168, 
    0, 0, 0, 0, 121, 125, 6, 7, 56, 39, 15, 0, 0, 0, 29, 181, 
    0, 0, 0, 0, 133, 105, 4, 7, 10, 0, 0, 0, 0, 0, 3, 177, 
    0, 0, 0, 0, 126, 47, 3, 5, 0, 0, 0, 0, 0, 0, 16, 167, 
    0, 0, 0, 0, 54, 0, 0, 0, 0, 0, 6, 0, 0, 10, 61, 158, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    0, 0, 2, 0, 1, 0, 0, 15, 8, 13, 11, 13, 16, 7, 11, 42, 
    0, 20, 26, 23, 28, 0, 10, 48, 50, 44, 43, 52, 52, 45, 47, 49, 
    0, 32, 24, 27, 25, 0, 38, 75, 83, 34, 18, 38, 49, 51, 46, 44, 
    0, 65, 20, 56, 35, 34, 60, 80, 71, 0, 3, 48, 66, 71, 53, 46, 
    0, 24, 0, 59, 0, 22, 40, 60, 91, 41, 0, 66, 78, 68, 66, 56, 
    0, 18, 8, 83, 0, 22, 38, 53, 118, 30, 0, 67, 80, 56, 84, 56, 
    0, 20, 44, 99, 0, 9, 1, 56, 105, 9, 0, 84, 89, 33, 54, 49, 
    0, 23, 86, 100, 38, 0, 0, 59, 77, 0, 0, 64, 81, 5, 36, 57, 
    0, 22, 99, 84, 35, 0, 25, 81, 59, 34, 12, 69, 78, 12, 30, 50, 
    0, 8, 87, 96, 36, 88, 72, 30, 54, 52, 55, 98, 84, 11, 36, 52, 
    0, 9, 88, 58, 0, 95, 54, 5, 83, 122, 126, 123, 81, 47, 87, 85, 
    0, 13, 76, 0, 0, 135, 97, 58, 116, 143, 126, 95, 87, 87, 118, 94, 
    0, 47, 34, 0, 47, 200, 133, 99, 116, 118, 98, 93, 94, 104, 112, 75, 
    34, 93, 23, 0, 131, 180, 103, 102, 103, 96, 95, 96, 109, 106, 110, 85, 
    37, 102, 66, 51, 154, 135, 83, 95, 86, 79, 93, 114, 87, 79, 127, 108, 
    0, 61, 58, 43, 88, 76, 49, 53, 39, 31, 53, 61, 11, 30, 94, 77, 
    
    -- channel=31
    0, 4, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 1, 6, 1, 0, 0, 0, 0, 
    0, 18, 25, 11, 0, 1, 12, 9, 9, 4, 0, 0, 0, 0, 0, 0, 
    0, 40, 26, 8, 16, 33, 0, 9, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 7, 0, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 10, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 4, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 50, 7, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end inmem_package;
