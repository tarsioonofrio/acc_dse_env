library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- ifmap
    588, 450, 35, 0, 0, 0, 0, 0, 147, 83, 222, 308, 230, 136, 14, 24, 53, 230, 0, 202, 234, 0, 0, 0, 156, 189, 471, 52, 272, 253, 210, 203, 360, 76, 192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 0, 0, 0, 297, 231, 0, 0, 0, 0, 20, 110, 0, 0, 152, 14, 259, 182, 28, 18, 47, 0, 215, 239, 332, 374, 0, 0, 0, 0, 528, 429, 287, 339, 0, 0, 0, 0, 198, 21, 191, 119, 142, 297, 0, 0, 0, 0, 0, 0, 416, 358, 19, 0, 110, 99, 0, 0, 310, 158, 41, 132, 91, 0, 811, 1065, 476, 214, 0, 0, 274, 173, 167, 174, 0, 0, 0, 0, 0, 100, 0, 0, 360, 444, 0, 194, 0, 0, 0, 0, 299, 156, 0, 0, 168, 49, 103, 0, 0, 0, 0, 0, 287, 310, 701, 156, 0, 0, 0, 0, 140, 224, 235, 328, 577, 463, 0, 0, 199, 0, 0, 0, 214, 85, 69, 0, 562, 86, 428, 192, 0, 0, 0, 0, 0, 0, 27, 0, 47, 58, 0, 0, 399, 49, 0, 0, 632, 592, 144, 141, 175, 58, 53, 0, 192, 40, 236, 0, 0, 0, 166, 0, 585, 455, 0, 0, 24, 0, 295, 80, 0, 0, 0, 0, 40, 113, 0, 0, 525, 140, 171, 182, 0, 0, 0, 0, 0, 193, 0, 0, 454, 487, 195, 0, 474, 225, 173, 166, 0, 0, 0, 0, 0, 0, 0, 0
    others => 0);
end gold_package;
