library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    64, 70, 71, 69, 68, 67, 72, 76, 68, 51, 44, 53, 59, 58, 56, 
    71, 74, 74, 69, 74, 85, 54, 55, 35, 40, 18, 15, 29, 52, 55, 
    28, 64, 72, 73, 72, 59, 34, 18, 21, 47, 14, 21, 2, 20, 58, 
    0, 56, 63, 76, 55, 58, 34, 12, 13, 46, 21, 17, 9, 0, 54, 
    6, 45, 47, 88, 68, 43, 22, 11, 3, 61, 34, 6, 21, 3, 17, 
    0, 41, 49, 45, 66, 48, 38, 22, 0, 86, 14, 4, 23, 12, 7, 
    13, 12, 43, 44, 58, 69, 36, 28, 1, 73, 11, 7, 19, 28, 12, 
    22, 29, 13, 38, 50, 59, 8, 23, 17, 62, 26, 4, 24, 23, 43, 
    20, 35, 0, 46, 23, 32, 27, 22, 38, 26, 24, 0, 19, 46, 56, 
    41, 36, 0, 46, 4, 22, 54, 31, 8, 20, 0, 5, 30, 62, 53, 
    53, 36, 0, 92, 25, 6, 30, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 27, 82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 60, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=1
    24, 23, 24, 27, 25, 24, 25, 24, 25, 26, 19, 17, 18, 20, 19, 
    24, 25, 26, 27, 27, 36, 32, 24, 10, 13, 21, 16, 11, 16, 23, 
    23, 15, 23, 25, 24, 34, 7, 10, 9, 23, 33, 26, 19, 13, 17, 
    35, 19, 29, 26, 25, 20, 37, 20, 15, 26, 23, 16, 8, 6, 13, 
    40, 53, 32, 36, 73, 41, 34, 16, 11, 1, 40, 25, 20, 17, 3, 
    26, 45, 30, 0, 21, 15, 35, 32, 23, 23, 38, 15, 23, 21, 11, 
    25, 40, 21, 22, 24, 22, 57, 27, 34, 31, 32, 19, 12, 21, 25, 
    25, 49, 30, 37, 27, 62, 34, 17, 21, 28, 21, 19, 17, 22, 16, 
    38, 46, 18, 27, 18, 8, 18, 23, 30, 16, 24, 5, 1, 16, 26, 
    37, 42, 35, 22, 45, 8, 18, 50, 25, 21, 9, 4, 22, 28, 27, 
    38, 39, 34, 45, 59, 59, 42, 43, 31, 12, 18, 20, 22, 29, 23, 
    38, 28, 48, 63, 43, 0, 5, 5, 12, 18, 20, 19, 21, 24, 23, 
    26, 23, 21, 61, 20, 18, 19, 16, 18, 20, 24, 29, 29, 24, 33, 
    27, 19, 24, 47, 19, 22, 20, 19, 17, 22, 21, 24, 18, 30, 26, 
    26, 19, 7, 33, 15, 14, 20, 20, 23, 25, 25, 20, 32, 44, 26, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 11, 0, 0, 0, 29, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 0, 0, 
    53, 0, 0, 0, 1, 0, 20, 10, 2, 0, 18, 0, 5, 8, 0, 
    65, 10, 17, 0, 58, 29, 13, 18, 0, 0, 19, 32, 4, 31, 0, 
    9, 0, 25, 0, 0, 0, 34, 23, 40, 0, 8, 15, 0, 17, 35, 
    33, 0, 0, 8, 0, 0, 0, 24, 26, 0, 21, 23, 0, 1, 17, 
    24, 21, 31, 28, 0, 0, 0, 0, 7, 0, 4, 13, 0, 0, 1, 
    21, 0, 42, 0, 8, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 50, 0, 9, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 31, 0, 127, 55, 0, 0, 23, 28, 24, 27, 5, 0, 3, 
    0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 9, 2, 0, 0, 0, 2, 5, 5, 0, 0, 12, 
    12, 2, 0, 0, 4, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 3, 12, 3, 0, 6, 16, 30, 
    
    -- channel=3
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 1, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 7, 5, 0, 0, 8, 9, 0, 
    0, 30, 0, 0, 0, 41, 0, 0, 0, 35, 5, 4, 0, 8, 18, 
    0, 20, 0, 0, 0, 2, 0, 0, 4, 50, 1, 12, 0, 0, 38, 
    0, 29, 0, 9, 3, 0, 2, 0, 4, 36, 6, 0, 5, 0, 5, 
    0, 44, 0, 0, 93, 22, 8, 0, 0, 62, 0, 0, 17, 0, 0, 
    0, 38, 12, 0, 61, 26, 36, 0, 0, 83, 0, 0, 8, 11, 0, 
    0, 28, 0, 0, 20, 61, 6, 28, 0, 61, 11, 0, 19, 22, 3, 
    4, 43, 0, 40, 0, 45, 9, 3, 17, 15, 24, 0, 21, 22, 2, 
    36, 39, 0, 54, 0, 0, 22, 13, 0, 15, 5, 3, 22, 18, 0, 
    76, 31, 0, 61, 0, 0, 42, 43, 0, 0, 0, 0, 11, 24, 5, 
    82, 66, 12, 83, 30, 16, 38, 34, 14, 15, 19, 24, 23, 23, 15, 
    12, 66, 53, 56, 0, 17, 18, 18, 15, 14, 19, 17, 25, 27, 22, 
    13, 23, 73, 53, 3, 21, 11, 15, 21, 20, 24, 30, 23, 22, 39, 
    11, 26, 32, 51, 14, 28, 29, 19, 20, 18, 14, 22, 29, 18, 5, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 7, 0, 9, 6, 8, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 5, 6, 0, 4, 6, 14, 9, 0, 
    20, 0, 0, 0, 0, 0, 7, 11, 12, 0, 5, 10, 6, 9, 0, 
    30, 0, 0, 0, 0, 0, 0, 7, 13, 0, 8, 18, 6, 9, 9, 
    27, 10, 0, 0, 0, 0, 0, 2, 15, 0, 18, 18, 11, 8, 2, 
    23, 18, 10, 0, 0, 0, 6, 7, 5, 0, 6, 20, 9, 0, 0, 
    22, 20, 29, 0, 2, 9, 11, 8, 0, 0, 9, 15, 7, 0, 0, 
    10, 13, 28, 12, 22, 1, 1, 6, 10, 1, 13, 20, 0, 0, 0, 
    14, 15, 30, 0, 6, 18, 3, 21, 25, 30, 38, 33, 34, 39, 44, 
    50, 23, 14, 0, 47, 67, 60, 62, 57, 53, 54, 56, 59, 58, 62, 
    66, 46, 16, 15, 67, 52, 52, 52, 54, 55, 58, 59, 57, 61, 62, 
    73, 62, 36, 40, 50, 52, 54, 54, 53, 57, 62, 65, 67, 68, 67, 
    70, 65, 59, 64, 56, 55, 52, 49, 48, 55, 61, 60, 53, 65, 71, 
    
    -- channel=5
    2, 1, 2, 3, 6, 2, 3, 10, 13, 14, 11, 6, 1, 0, 1, 
    6, 3, 3, 5, 3, 0, 3, 16, 13, 0, 0, 0, 0, 3, 3, 
    15, 15, 8, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 43, 1, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 5, 8, 2, 0, 0, 
    19, 29, 0, 0, 0, 0, 27, 9, 0, 0, 0, 0, 0, 0, 0, 
    30, 66, 0, 11, 97, 55, 0, 0, 0, 0, 22, 15, 8, 14, 0, 
    0, 0, 0, 0, 0, 0, 15, 16, 16, 40, 0, 0, 0, 7, 27, 
    6, 0, 0, 0, 0, 7, 0, 2, 1, 5, 0, 0, 0, 11, 17, 
    4, 6, 16, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 1, 43, 0, 0, 0, 0, 25, 16, 0, 
    0, 0, 0, 62, 104, 89, 14, 0, 0, 0, 28, 46, 16, 0, 0, 
    0, 0, 16, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 19, 0, 0, 25, 
    0, 0, 0, 0, 0, 2, 7, 0, 0, 2, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 17, 2, 0, 38, 26, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 7, 0, 0, 0, 15, 0, 0, 0, 7, 0, 
    0, 27, 0, 0, 0, 10, 0, 0, 1, 31, 0, 0, 0, 0, 13, 
    0, 26, 0, 0, 0, 22, 0, 0, 0, 34, 0, 0, 0, 0, 37, 
    0, 14, 0, 47, 12, 0, 0, 0, 0, 48, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 47, 0, 0, 0, 0, 71, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 43, 10, 0, 0, 0, 59, 0, 0, 0, 10, 0, 
    0, 2, 0, 0, 24, 24, 0, 0, 0, 26, 0, 0, 11, 0, 0, 
    0, 0, 0, 25, 0, 9, 0, 0, 26, 0, 1, 0, 7, 19, 0, 
    0, 0, 0, 37, 0, 0, 29, 0, 0, 0, 0, 9, 28, 7, 0, 
    43, 0, 0, 77, 0, 0, 0, 0, 0, 0, 8, 2, 0, 1, 0, 
    23, 20, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 8, 39, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 1, 11, 
    0, 0, 21, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 20, 0, 0, 0, 0, 2, 0, 0, 4, 25, 0, 0, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    24, 27, 27, 26, 29, 27, 29, 35, 34, 27, 22, 22, 20, 23, 24, 
    29, 31, 30, 28, 24, 10, 26, 36, 24, 0, 0, 3, 18, 14, 19, 
    35, 14, 30, 31, 33, 30, 14, 11, 0, 0, 0, 0, 0, 6, 8, 
    0, 5, 21, 32, 36, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 19, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 38, 0, 0, 0, 17, 10, 0, 
    28, 37, 0, 0, 0, 47, 14, 16, 0, 0, 0, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 11, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 19, 70, 16, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 20, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 16, 28, 0, 4, 0, 0, 4, 6, 0, 
    0, 0, 0, 0, 0, 50, 0, 0, 0, 0, 37, 31, 13, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 42, 30, 9, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 34, 6, 0, 0, 0, 0, 20, 19, 
    78, 27, 0, 0, 63, 60, 42, 39, 16, 5, 0, 0, 0, 0, 0, 
    0, 57, 4, 14, 39, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 
    0, 0, 62, 46, 4, 0, 0, 0, 0, 0, 1, 11, 0, 0, 33, 
    0, 0, 11, 50, 15, 23, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    35, 39, 36, 38, 36, 36, 37, 42, 38, 31, 23, 23, 26, 32, 34, 
    36, 41, 39, 39, 36, 40, 25, 31, 19, 4, 1, 4, 11, 22, 32, 
    29, 24, 38, 40, 42, 47, 7, 3, 0, 8, 0, 0, 5, 8, 26, 
    11, 16, 35, 37, 32, 9, 15, 0, 1, 7, 0, 4, 0, 3, 22, 
    0, 20, 17, 8, 15, 0, 0, 0, 5, 0, 0, 0, 5, 3, 6, 
    0, 2, 7, 22, 16, 0, 4, 0, 10, 8, 0, 0, 4, 0, 0, 
    0, 13, 1, 31, 33, 0, 10, 0, 4, 17, 0, 0, 0, 0, 3, 
    0, 0, 0, 15, 13, 20, 0, 0, 0, 24, 0, 0, 0, 7, 7, 
    0, 0, 0, 2, 0, 0, 0, 10, 0, 14, 16, 0, 3, 14, 32, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 2, 0, 0, 12, 29, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    64, 67, 67, 71, 69, 67, 67, 69, 69, 62, 55, 52, 59, 59, 56, 
    64, 66, 67, 72, 70, 98, 88, 66, 52, 56, 69, 54, 40, 44, 58, 
    58, 37, 68, 70, 67, 79, 75, 50, 39, 66, 99, 82, 65, 26, 44, 
    95, 31, 71, 69, 80, 70, 93, 71, 58, 52, 111, 64, 63, 30, 15, 
    140, 96, 97, 74, 157, 135, 125, 83, 52, 36, 116, 93, 61, 54, 14, 
    144, 123, 112, 67, 84, 122, 141, 100, 76, 38, 150, 95, 58, 69, 47, 
    150, 133, 73, 79, 50, 105, 145, 125, 94, 61, 142, 88, 59, 67, 73, 
    158, 156, 99, 93, 61, 111, 154, 89, 82, 69, 119, 89, 51, 70, 69, 
    176, 152, 136, 81, 96, 76, 89, 82, 67, 92, 59, 68, 30, 47, 60, 
    159, 153, 149, 83, 110, 72, 88, 132, 89, 68, 62, 23, 29, 61, 79, 
    116, 154, 148, 105, 213, 130, 107, 139, 112, 71, 48, 53, 62, 70, 75, 
    74, 125, 151, 158, 200, 103, 71, 70, 68, 64, 68, 73, 81, 87, 89, 
    91, 67, 116, 191, 149, 76, 73, 69, 70, 71, 78, 87, 89, 88, 103, 
    97, 72, 66, 171, 94, 80, 84, 70, 69, 77, 83, 82, 85, 89, 97, 
    105, 77, 69, 82, 68, 57, 68, 76, 80, 92, 88, 79, 96, 129, 96, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 17, 11, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 7, 11, 0, 2, 2, 0, 0, 
    19, 11, 0, 0, 0, 0, 0, 0, 6, 5, 5, 1, 5, 2, 0, 
    36, 20, 0, 0, 7, 0, 0, 0, 3, 15, 11, 4, 10, 9, 3, 
    31, 26, 0, 0, 0, 0, 8, 1, 5, 25, 12, 8, 11, 11, 1, 
    29, 27, 10, 0, 0, 15, 14, 7, 0, 5, 4, 8, 13, 4, 0, 
    40, 42, 24, 6, 0, 6, 0, 3, 6, 0, 0, 0, 5, 0, 0, 
    28, 38, 23, 35, 15, 3, 5, 12, 15, 0, 4, 9, 2, 0, 0, 
    38, 31, 25, 38, 26, 35, 43, 38, 28, 23, 40, 49, 61, 55, 50, 
    94, 53, 31, 40, 51, 59, 68, 68, 70, 74, 81, 86, 89, 90, 88, 
    104, 84, 45, 44, 58, 76, 77, 73, 76, 81, 91, 95, 94, 97, 103, 
    109, 96, 85, 53, 65, 81, 78, 77, 79, 87, 97, 101, 100, 111, 109, 
    104, 102, 90, 77, 76, 81, 81, 78, 81, 88, 91, 92, 98, 111, 100, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 19, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 10, 3, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 2, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 2, 6, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 8, 17, 0, 15, 8, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 18, 0, 0, 0, 2, 1, 8, 
    27, 15, 0, 0, 31, 0, 0, 0, 3, 0, 12, 8, 10, 2, 0, 
    11, 30, 0, 0, 4, 0, 10, 0, 6, 13, 10, 8, 9, 4, 4, 
    15, 5, 1, 0, 0, 18, 16, 20, 3, 13, 9, 14, 15, 15, 0, 
    20, 22, 24, 1, 0, 18, 3, 6, 0, 0, 28, 16, 16, 0, 0, 
    20, 27, 17, 12, 19, 3, 0, 0, 23, 17, 12, 9, 0, 0, 0, 
    22, 18, 19, 0, 0, 6, 28, 32, 19, 4, 17, 19, 35, 29, 26, 
    86, 33, 5, 15, 69, 63, 63, 61, 56, 52, 57, 60, 60, 65, 64, 
    76, 79, 17, 48, 50, 52, 56, 54, 54, 57, 59, 62, 68, 66, 58, 
    78, 68, 77, 52, 48, 54, 52, 58, 57, 61, 71, 78, 70, 75, 97, 
    75, 74, 73, 69, 63, 70, 67, 53, 51, 55, 68, 63, 53, 73, 71, 
    
    -- channel=16
    58, 59, 59, 58, 55, 56, 59, 55, 51, 51, 49, 48, 47, 45, 38, 
    51, 50, 59, 59, 60, 76, 60, 54, 47, 43, 43, 35, 37, 41, 41, 
    54, 51, 56, 56, 59, 89, 64, 30, 28, 74, 90, 70, 44, 31, 43, 
    31, 37, 54, 56, 55, 50, 65, 55, 52, 89, 91, 68, 48, 22, 36, 
    88, 90, 71, 78, 113, 113, 102, 64, 45, 65, 92, 62, 48, 26, 24, 
    133, 137, 86, 89, 153, 144, 117, 70, 34, 95, 136, 74, 59, 50, 24, 
    132, 130, 76, 44, 82, 124, 144, 104, 58, 115, 118, 64, 53, 61, 56, 
    153, 130, 82, 49, 70, 155, 147, 105, 66, 113, 117, 66, 60, 78, 61, 
    170, 161, 111, 93, 87, 99, 77, 68, 67, 68, 77, 58, 43, 57, 63, 
    171, 168, 113, 100, 94, 78, 89, 95, 87, 87, 51, 13, 31, 60, 60, 
    144, 158, 114, 145, 148, 94, 142, 154, 94, 37, 22, 39, 61, 73, 64, 
    132, 161, 135, 201, 200, 109, 86, 84, 72, 65, 71, 77, 83, 90, 86, 
    88, 119, 158, 209, 122, 76, 73, 69, 65, 67, 75, 85, 95, 95, 99, 
    91, 79, 147, 167, 87, 81, 74, 69, 73, 80, 89, 94, 87, 99, 117, 
    97, 84, 90, 85, 68, 76, 85, 79, 81, 87, 84, 81, 100, 117, 78, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 17, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 2, 0, 11, 11, 0, 0, 0, 0, 
    35, 31, 0, 11, 55, 37, 17, 3, 0, 21, 30, 8, 4, 0, 0, 
    28, 30, 0, 0, 21, 28, 37, 14, 0, 44, 21, 0, 2, 5, 0, 
    39, 30, 0, 0, 4, 41, 32, 24, 3, 41, 22, 7, 5, 18, 0, 
    49, 48, 8, 0, 14, 39, 6, 4, 0, 20, 22, 2, 6, 0, 0, 
    58, 55, 19, 25, 8, 1, 7, 14, 10, 0, 0, 0, 0, 0, 0, 
    49, 52, 29, 43, 14, 0, 26, 46, 1, 0, 0, 0, 0, 0, 0, 
    53, 51, 24, 77, 88, 47, 45, 31, 11, 5, 15, 29, 22, 13, 11, 
    21, 48, 48, 84, 33, 11, 17, 18, 20, 23, 28, 32, 39, 39, 37, 
    35, 22, 55, 56, 11, 32, 29, 26, 27, 32, 40, 43, 38, 42, 55, 
    40, 36, 33, 27, 26, 34, 34, 29, 31, 36, 37, 36, 40, 52, 30, 
    40, 41, 33, 11, 16, 20, 23, 31, 41, 45, 36, 37, 64, 59, 35, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 1, 0, 0, 
    0, 11, 0, 0, 0, 0, 24, 35, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 18, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 9, 0, 2, 8, 0, 0, 10, 
    0, 0, 0, 0, 0, 29, 18, 0, 0, 0, 0, 41, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 34, 21, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 4, 14, 
    0, 0, 0, 0, 0, 83, 38, 38, 25, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 86, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 26, 19, 0, 0, 0, 0, 0, 0, 1, 15, 0, 0, 
    1, 0, 0, 48, 16, 4, 4, 2, 0, 0, 0, 7, 0, 0, 19, 
    
    -- channel=19
    42, 40, 44, 43, 45, 39, 42, 46, 45, 33, 28, 30, 35, 37, 38, 
    46, 39, 43, 43, 46, 47, 39, 33, 27, 33, 25, 19, 22, 32, 36, 
    20, 38, 43, 46, 45, 19, 38, 26, 20, 17, 7, 20, 15, 19, 33, 
    12, 36, 40, 44, 39, 42, 19, 16, 17, 9, 20, 9, 17, 15, 25, 
    23, 15, 40, 50, 26, 25, 14, 16, 8, 33, 18, 15, 15, 14, 16, 
    18, 16, 40, 30, 9, 25, 21, 16, 10, 22, 14, 18, 11, 16, 19, 
    28, 2, 32, 27, 10, 32, 4, 25, 7, 12, 18, 16, 18, 17, 14, 
    24, 12, 29, 28, 22, 0, 15, 13, 16, 13, 25, 13, 12, 8, 32, 
    19, 9, 17, 21, 23, 17, 22, 16, 24, 25, 1, 12, 14, 31, 36, 
    18, 13, 13, 19, 2, 20, 32, 10, 10, 8, 12, 10, 12, 23, 31, 
    7, 13, 11, 23, 34, 6, 0, 0, 7, 15, 8, 7, 6, 17, 20, 
    0, 10, 18, 11, 0, 9, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 10, 5, 0, 15, 18, 11, 0, 0, 
    21, 0, 0, 0, 0, 0, 16, 4, 6, 2, 38, 24, 20, 11, 0, 
    22, 0, 0, 0, 9, 0, 15, 27, 15, 14, 36, 24, 12, 12, 0, 
    47, 25, 30, 1, 36, 64, 50, 32, 15, 0, 32, 38, 9, 8, 15, 
    89, 47, 42, 22, 16, 62, 39, 28, 15, 0, 76, 42, 13, 16, 14, 
    89, 51, 34, 0, 0, 32, 53, 46, 26, 5, 61, 33, 14, 10, 25, 
    95, 46, 65, 12, 0, 44, 79, 37, 20, 7, 41, 31, 13, 26, 8, 
    90, 68, 83, 18, 52, 26, 22, 16, 16, 19, 16, 28, 2, 0, 3, 
    59, 67, 64, 17, 61, 48, 22, 25, 59, 34, 22, 0, 0, 1, 10, 
    28, 70, 60, 23, 74, 70, 65, 74, 65, 23, 12, 21, 38, 40, 41, 
    57, 59, 62, 53, 113, 62, 38, 40, 38, 33, 36, 37, 39, 44, 47, 
    58, 55, 58, 90, 81, 38, 39, 35, 31, 33, 35, 45, 51, 48, 48, 
    55, 47, 72, 67, 43, 39, 40, 38, 36, 41, 45, 46, 43, 51, 68, 
    61, 43, 50, 29, 35, 34, 39, 38, 36, 41, 46, 38, 37, 64, 53, 
    
    -- channel=21
    16, 16, 13, 13, 11, 12, 17, 18, 10, 9, 12, 15, 12, 11, 10, 
    10, 16, 14, 13, 12, 0, 2, 10, 15, 0, 0, 0, 10, 15, 10, 
    9, 27, 17, 15, 16, 32, 11, 9, 0, 0, 0, 0, 0, 6, 13, 
    0, 0, 13, 12, 4, 3, 0, 0, 0, 8, 0, 0, 0, 0, 13, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 16, 43, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 7, 4, 6, 0, 0, 0, 3, 6, 
    0, 0, 0, 0, 0, 22, 7, 0, 0, 0, 23, 9, 9, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 6, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 0, 0, 3, 13, 4, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    31, 37, 32, 30, 28, 34, 32, 32, 27, 27, 31, 33, 33, 24, 21, 
    25, 33, 32, 32, 34, 39, 22, 31, 41, 35, 17, 10, 20, 31, 21, 
    21, 49, 32, 33, 30, 51, 48, 25, 16, 37, 31, 29, 7, 9, 33, 
    3, 2, 27, 33, 26, 39, 25, 14, 16, 42, 44, 29, 28, 0, 26, 
    44, 18, 27, 49, 52, 33, 47, 24, 14, 42, 41, 18, 17, 4, 0, 
    54, 63, 40, 41, 114, 94, 64, 28, 1, 42, 55, 39, 24, 18, 1, 
    59, 51, 50, 32, 47, 69, 72, 51, 22, 50, 61, 24, 19, 28, 12, 
    69, 70, 16, 30, 31, 70, 66, 56, 40, 44, 65, 27, 27, 31, 31, 
    80, 79, 39, 57, 25, 66, 48, 26, 32, 26, 43, 34, 23, 33, 21, 
    95, 79, 51, 52, 36, 26, 54, 41, 11, 48, 30, 12, 9, 21, 30, 
    88, 77, 55, 68, 60, 10, 52, 82, 45, 14, 0, 3, 9, 30, 30, 
    51, 98, 71, 78, 95, 74, 47, 47, 34, 21, 18, 22, 25, 20, 23, 
    10, 43, 93, 86, 72, 25, 20, 19, 15, 13, 16, 16, 23, 33, 28, 
    20, 18, 53, 96, 39, 22, 19, 16, 22, 20, 21, 28, 27, 22, 30, 
    20, 22, 26, 42, 16, 23, 30, 26, 22, 22, 16, 21, 28, 20, 16, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 7, 12, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 10, 0, 29, 11, 11, 15, 9, 2, 6, 19, 18, 6, 0, 
    40, 20, 21, 14, 18, 9, 20, 19, 24, 32, 41, 45, 50, 51, 48, 
    62, 32, 6, 7, 13, 39, 43, 39, 40, 44, 52, 52, 55, 56, 60, 
    66, 55, 18, 27, 26, 44, 44, 41, 44, 48, 54, 56, 59, 55, 67, 
    66, 61, 46, 41, 35, 36, 42, 44, 47, 51, 53, 54, 60, 71, 70, 
    
    -- channel=24
    72, 76, 76, 77, 75, 76, 75, 76, 74, 63, 54, 57, 63, 63, 61, 
    75, 74, 76, 77, 79, 123, 72, 66, 40, 66, 68, 51, 47, 57, 64, 
    53, 56, 77, 77, 78, 74, 61, 37, 47, 88, 79, 68, 51, 38, 65, 
    51, 83, 75, 80, 77, 73, 86, 57, 57, 74, 78, 57, 48, 35, 52, 
    82, 117, 73, 89, 142, 99, 82, 61, 43, 78, 96, 61, 61, 43, 31, 
    81, 124, 80, 71, 115, 92, 114, 71, 52, 121, 94, 53, 60, 54, 44, 
    90, 110, 68, 57, 82, 126, 114, 90, 56, 119, 85, 64, 61, 75, 61, 
    111, 112, 72, 71, 77, 127, 77, 71, 62, 104, 93, 60, 61, 66, 64, 
    124, 125, 78, 100, 78, 60, 74, 81, 78, 66, 72, 29, 43, 73, 81, 
    130, 127, 88, 101, 74, 54, 88, 110, 69, 54, 27, 23, 59, 79, 67, 
    133, 122, 83, 160, 154, 99, 108, 92, 60, 39, 50, 60, 61, 66, 60, 
    76, 113, 106, 183, 101, 56, 56, 53, 56, 53, 60, 62, 72, 74, 68, 
    68, 74, 125, 150, 51, 63, 57, 57, 58, 62, 69, 76, 70, 68, 90, 
    67, 63, 92, 102, 64, 66, 65, 58, 59, 65, 67, 67, 66, 87, 65, 
    67, 66, 66, 53, 49, 55, 57, 61, 71, 78, 66, 66, 98, 95, 56, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    57, 58, 60, 60, 61, 53, 63, 64, 61, 49, 38, 41, 47, 55, 56, 
    60, 61, 63, 62, 59, 60, 60, 53, 35, 23, 23, 25, 26, 39, 53, 
    42, 34, 61, 63, 63, 31, 36, 19, 21, 11, 13, 12, 23, 21, 41, 
    29, 33, 59, 59, 59, 29, 33, 20, 15, 2, 19, 15, 14, 22, 25, 
    8, 25, 57, 33, 37, 31, 20, 22, 15, 5, 18, 25, 17, 21, 23, 
    0, 5, 52, 47, 0, 8, 27, 21, 26, 9, 14, 11, 10, 14, 23, 
    0, 12, 28, 55, 12, 20, 11, 17, 18, 2, 9, 16, 12, 12, 23, 
    1, 3, 18, 37, 20, 9, 6, 7, 15, 16, 13, 14, 7, 13, 29, 
    0, 0, 11, 11, 29, 0, 15, 23, 10, 28, 11, 7, 10, 30, 56, 
    0, 0, 10, 0, 12, 13, 5, 21, 16, 13, 7, 6, 14, 42, 46, 
    0, 0, 4, 0, 26, 19, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 
    0, 0, 0, 0, 0, 0, 20, 0, 14, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 36, 8, 0, 0, 13, 12, 34, 0, 0, 
    78, 0, 0, 0, 3, 0, 3, 16, 3, 0, 42, 0, 30, 21, 0, 
    89, 0, 35, 0, 0, 0, 35, 29, 12, 0, 9, 49, 0, 38, 0, 
    49, 0, 50, 0, 0, 16, 39, 33, 48, 0, 44, 58, 0, 20, 21, 
    52, 17, 10, 42, 0, 0, 8, 31, 61, 0, 69, 35, 0, 0, 21, 
    34, 27, 27, 22, 0, 0, 55, 4, 35, 0, 42, 41, 0, 0, 17, 
    36, 0, 79, 0, 0, 0, 24, 0, 0, 10, 0, 47, 0, 0, 0, 
    0, 0, 94, 0, 42, 0, 0, 17, 0, 4, 45, 5, 0, 0, 7, 
    0, 0, 81, 0, 101, 22, 0, 8, 64, 26, 0, 0, 0, 0, 0, 
    0, 0, 36, 0, 89, 51, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 56, 28, 0, 9, 0, 0, 0, 0, 0, 2, 0, 2, 
    24, 0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 0, 4, 52, 
    
    -- channel=29
    55, 58, 57, 57, 57, 53, 59, 64, 57, 46, 42, 47, 49, 48, 49, 
    56, 58, 60, 58, 59, 51, 44, 47, 42, 33, 11, 14, 31, 45, 48, 
    36, 61, 60, 61, 60, 68, 41, 30, 14, 23, 9, 13, 2, 21, 47, 
    5, 29, 52, 59, 48, 45, 21, 7, 8, 27, 20, 15, 15, 1, 40, 
    4, 14, 40, 51, 27, 11, 21, 11, 10, 26, 20, 3, 14, 2, 12, 
    2, 28, 40, 35, 62, 34, 26, 16, 3, 26, 15, 14, 17, 7, 0, 
    2, 14, 41, 44, 44, 33, 31, 20, 9, 31, 18, 8, 13, 13, 7, 
    2, 24, 1, 35, 27, 32, 25, 26, 23, 37, 24, 12, 15, 20, 36, 
    7, 20, 0, 27, 11, 39, 30, 15, 22, 29, 29, 20, 21, 33, 35, 
    32, 22, 3, 21, 5, 11, 30, 15, 3, 24, 15, 7, 13, 36, 46, 
    35, 21, 13, 29, 0, 0, 0, 17, 0, 1, 0, 0, 0, 3, 0, 
    5, 24, 15, 29, 13, 9, 4, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 26, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    30, 34, 28, 33, 28, 29, 29, 32, 29, 25, 23, 22, 24, 25, 27, 
    24, 29, 27, 32, 29, 35, 25, 25, 20, 17, 11, 8, 11, 18, 25, 
    30, 21, 31, 33, 28, 42, 46, 23, 10, 9, 38, 32, 13, 0, 20, 
    39, 0, 26, 27, 30, 21, 28, 20, 16, 3, 54, 22, 35, 9, 0, 
    55, 1, 35, 4, 42, 12, 52, 38, 25, 0, 37, 31, 20, 20, 0, 
    54, 48, 51, 24, 64, 59, 68, 38, 32, 0, 64, 53, 18, 24, 6, 
    56, 49, 35, 52, 7, 32, 61, 51, 46, 0, 69, 38, 14, 18, 27, 
    55, 67, 8, 34, 0, 34, 85, 45, 54, 12, 62, 45, 13, 28, 38, 
    71, 54, 60, 25, 27, 34, 46, 31, 14, 18, 38, 51, 15, 26, 18, 
    80, 57, 78, 3, 48, 18, 21, 42, 19, 46, 38, 5, 0, 3, 27, 
    41, 54, 76, 10, 69, 17, 12, 64, 52, 15, 1, 0, 0, 6, 14, 
    15, 54, 59, 17, 101, 74, 31, 34, 32, 17, 15, 16, 22, 17, 25, 
    18, 10, 32, 75, 107, 22, 18, 17, 16, 13, 13, 17, 20, 23, 25, 
    32, 10, 0, 115, 47, 18, 22, 16, 15, 17, 19, 26, 25, 19, 33, 
    35, 19, 8, 46, 24, 19, 26, 25, 15, 22, 23, 19, 13, 34, 33, 
    
    -- channel=31
    55, 53, 55, 53, 54, 51, 57, 59, 53, 46, 43, 48, 47, 47, 47, 
    55, 55, 57, 53, 56, 49, 38, 47, 35, 30, 11, 21, 39, 49, 48, 
    38, 64, 59, 55, 60, 57, 22, 22, 25, 35, 2, 5, 1, 38, 50, 
    0, 61, 50, 58, 42, 41, 16, 8, 13, 45, 0, 17, 4, 11, 59, 
    0, 29, 30, 58, 10, 12, 0, 1, 11, 50, 5, 0, 16, 0, 41, 
    0, 16, 22, 50, 45, 10, 0, 0, 0, 76, 0, 0, 21, 4, 6, 
    0, 0, 32, 27, 56, 36, 4, 0, 0, 67, 0, 0, 17, 16, 7, 
    0, 0, 1, 19, 42, 40, 0, 14, 5, 58, 0, 0, 22, 24, 25, 
    0, 0, 0, 21, 20, 24, 7, 12, 24, 22, 28, 1, 32, 34, 45, 
    1, 2, 0, 27, 0, 23, 27, 0, 13, 18, 1, 12, 31, 52, 41, 
    29, 3, 0, 53, 0, 0, 22, 0, 0, 0, 1, 0, 0, 10, 0, 
    22, 12, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    49, 50, 50, 50, 50, 50, 50, 50, 52, 48, 49, 50, 50, 50, 51, 
    49, 50, 50, 50, 50, 50, 50, 50, 46, 21, 49, 55, 50, 50, 50, 
    50, 51, 51, 50, 52, 48, 49, 31, 21, 15, 31, 59, 49, 51, 51, 
    46, 44, 49, 52, 51, 35, 57, 36, 39, 30, 35, 50, 45, 47, 49, 
    7, 26, 61, 52, 50, 44, 53, 47, 48, 33, 15, 13, 14, 54, 50, 
    35, 46, 39, 33, 41, 4, 21, 29, 45, 36, 35, 37, 24, 56, 48, 
    0, 21, 30, 51, 19, 0, 14, 42, 55, 35, 23, 18, 28, 20, 41, 
    31, 33, 17, 53, 47, 39, 49, 12, 20, 20, 14, 22, 29, 35, 28, 
    82, 35, 40, 45, 40, 29, 28, 16, 23, 8, 18, 1, 6, 7, 14, 
    16, 1, 1, 0, 4, 6, 1, 2, 4, 0, 0, 0, 0, 5, 20, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 16, 27, 
    0, 15, 6, 0, 0, 0, 50, 0, 3, 11, 27, 25, 21, 30, 41, 
    0, 0, 7, 0, 0, 0, 70, 76, 73, 51, 32, 39, 36, 36, 43, 
    0, 0, 0, 0, 0, 0, 47, 91, 55, 49, 44, 36, 29, 35, 41, 
    0, 0, 0, 0, 0, 0, 7, 40, 42, 48, 32, 25, 32, 36, 42, 
    
    -- channel=33
    59, 59, 59, 59, 59, 59, 59, 59, 58, 60, 59, 60, 60, 59, 60, 
    59, 59, 59, 59, 58, 59, 58, 58, 58, 49, 42, 54, 59, 59, 59, 
    57, 57, 59, 59, 59, 60, 58, 55, 46, 47, 47, 48, 59, 59, 60, 
    59, 60, 61, 60, 58, 55, 51, 59, 55, 58, 52, 62, 62, 62, 61, 
    12, 22, 48, 56, 58, 65, 61, 64, 61, 62, 54, 37, 28, 38, 61, 
    70, 64, 66, 46, 47, 48, 37, 41, 45, 56, 63, 66, 55, 52, 63, 
    1, 1, 33, 45, 63, 14, 8, 21, 51, 63, 52, 38, 42, 36, 35, 
    1, 35, 24, 25, 49, 63, 72, 56, 24, 18, 20, 27, 34, 47, 52, 
    15, 78, 64, 66, 61, 55, 57, 58, 57, 56, 51, 48, 33, 24, 21, 
    28, 12, 14, 13, 12, 20, 22, 19, 23, 15, 18, 14, 20, 22, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 22, 26, 
    0, 9, 9, 2, 0, 0, 0, 17, 8, 7, 13, 32, 21, 15, 30, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 31, 43, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 27, 30, 35, 47, 
    18, 2, 0, 0, 0, 0, 0, 0, 3, 24, 30, 32, 37, 42, 50, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 15, 33, 38, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 39, 0, 0, 0, 0, 0, 0, 0, 0, 34, 47, 63, 0, 0, 
    0, 0, 0, 0, 5, 49, 2, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 71, 46, 0, 0, 0, 8, 21, 19, 30, 0, 
    0, 0, 43, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    4, 0, 23, 29, 8, 0, 37, 95, 58, 54, 51, 28, 0, 0, 0, 
    33, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 4, 0, 1, 3, 2, 0, 0, 0, 0, 21, 0, 0, 0, 0, 
    44, 26, 17, 16, 16, 16, 2, 0, 28, 2, 0, 0, 0, 0, 0, 
    
    -- channel=35
    45, 47, 47, 47, 47, 47, 47, 47, 46, 45, 48, 47, 47, 47, 47, 
    46, 47, 47, 47, 47, 47, 48, 47, 44, 44, 70, 56, 46, 47, 48, 
    49, 49, 48, 47, 48, 45, 49, 42, 49, 36, 60, 75, 47, 48, 48, 
    48, 45, 49, 48, 49, 43, 58, 30, 26, 18, 19, 47, 47, 46, 48, 
    67, 72, 78, 51, 48, 40, 48, 41, 42, 35, 49, 61, 62, 80, 54, 
    7, 19, 56, 48, 57, 51, 78, 76, 77, 46, 15, 10, 3, 45, 55, 
    68, 87, 63, 41, 36, 0, 28, 28, 37, 50, 55, 59, 64, 68, 75, 
    49, 19, 25, 72, 46, 0, 10, 33, 59, 43, 19, 15, 18, 16, 25, 
    39, 47, 9, 35, 53, 52, 57, 27, 28, 37, 46, 42, 57, 63, 51, 
    88, 69, 74, 72, 69, 61, 52, 40, 47, 23, 43, 30, 27, 31, 41, 
    20, 42, 34, 47, 56, 64, 65, 63, 55, 46, 38, 36, 35, 19, 34, 
    0, 18, 0, 0, 0, 0, 33, 0, 0, 0, 4, 2, 32, 30, 28, 
    0, 2, 19, 0, 0, 0, 95, 53, 39, 33, 45, 39, 8, 25, 34, 
    0, 0, 0, 0, 0, 0, 34, 57, 32, 24, 0, 12, 19, 26, 42, 
    0, 0, 0, 0, 0, 0, 0, 28, 0, 13, 14, 14, 20, 25, 38, 
    
    -- channel=36
    12, 11, 11, 11, 11, 11, 11, 10, 10, 12, 13, 11, 11, 11, 11, 
    12, 12, 12, 12, 12, 12, 12, 11, 15, 25, 18, 14, 12, 12, 12, 
    11, 11, 11, 12, 12, 13, 13, 20, 31, 34, 17, 8, 12, 11, 12, 
    19, 17, 12, 10, 11, 17, 10, 20, 19, 24, 24, 17, 16, 14, 12, 
    49, 39, 11, 10, 13, 15, 8, 14, 12, 19, 23, 28, 35, 20, 12, 
    5, 1, 8, 17, 15, 25, 18, 15, 13, 22, 24, 15, 19, 8, 14, 
    49, 42, 32, 11, 20, 53, 43, 38, 20, 14, 17, 20, 16, 18, 22, 
    23, 11, 23, 14, 23, 13, 0, 14, 33, 46, 48, 40, 32, 27, 20, 
    4, 12, 6, 4, 12, 22, 24, 24, 15, 19, 19, 24, 25, 33, 39, 
    10, 46, 52, 56, 55, 57, 59, 57, 52, 53, 50, 50, 42, 32, 25, 
    46, 43, 52, 50, 45, 47, 55, 56, 54, 55, 53, 46, 39, 29, 15, 
    17, 8, 7, 14, 17, 18, 12, 42, 44, 40, 27, 15, 4, 14, 8, 
    16, 13, 16, 20, 16, 14, 0, 0, 0, 0, 0, 15, 11, 4, 6, 
    18, 12, 12, 16, 13, 13, 0, 0, 0, 10, 5, 0, 5, 7, 7, 
    18, 4, 8, 9, 10, 11, 1, 6, 6, 0, 0, 5, 4, 4, 7, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 40, 51, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 5, 0, 0, 0, 0, 0, 0, 
    94, 91, 5, 0, 0, 0, 0, 0, 0, 0, 37, 72, 67, 44, 0, 
    0, 0, 0, 0, 0, 0, 0, 27, 40, 0, 0, 0, 0, 0, 0, 
    0, 66, 0, 0, 0, 92, 120, 0, 0, 0, 0, 9, 26, 50, 30, 
    93, 34, 78, 53, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 22, 23, 2, 0, 72, 103, 62, 64, 77, 77, 6, 0, 14, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 14, 13, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 38, 0, 0, 0, 
    0, 26, 20, 16, 16, 18, 9, 0, 45, 53, 6, 0, 2, 6, 2, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 9, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 5, 0, 
    0, 17, 7, 12, 0, 0, 16, 31, 11, 0, 0, 0, 0, 0, 13, 
    61, 0, 0, 21, 17, 0, 0, 0, 0, 0, 0, 3, 6, 9, 0, 
    79, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 19, 0, 4, 
    0, 31, 0, 0, 0, 6, 74, 0, 4, 9, 17, 0, 0, 2, 16, 
    0, 0, 7, 0, 0, 0, 68, 0, 0, 0, 0, 16, 9, 9, 12, 
    0, 0, 2, 1, 2, 3, 19, 0, 0, 27, 24, 2, 0, 6, 12, 
    0, 0, 1, 2, 4, 5, 0, 28, 25, 14, 0, 0, 5, 4, 7, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 3, 16, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 12, 0, 6, 18, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 22, 18, 19, 22, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 16, 17, 17, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 6, 0, 0, 0, 8, 0, 0, 2, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 29, 91, 93, 39, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 27, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 38, 19, 31, 16, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    91, 86, 18, 0, 0, 0, 0, 0, 0, 0, 35, 65, 80, 54, 0, 
    0, 0, 0, 32, 30, 94, 108, 90, 51, 0, 0, 0, 0, 0, 0, 
    108, 107, 57, 0, 0, 0, 0, 0, 0, 10, 52, 75, 69, 67, 61, 
    16, 0, 0, 23, 0, 0, 0, 0, 50, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 38, 15, 0, 19, 17, 34, 61, 71, 43, 
    54, 91, 88, 85, 72, 54, 33, 16, 23, 10, 31, 21, 7, 9, 5, 
    52, 50, 62, 88, 104, 112, 109, 102, 83, 71, 52, 29, 0, 0, 0, 
    7, 14, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 36, 21, 2, 0, 57, 17, 0, 19, 58, 35, 0, 0, 0, 
    0, 0, 2, 1, 0, 0, 13, 30, 64, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 7, 6, 1, 4, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 9, 8, 6, 7, 9, 0, 12, 0, 0, 1, 9, 0, 0, 0, 
    0, 12, 12, 10, 9, 8, 3, 8, 2, 14, 8, 0, 0, 0, 0, 
    
    -- channel=44
    212, 210, 210, 210, 210, 210, 210, 210, 209, 210, 209, 210, 210, 210, 210, 
    212, 210, 210, 210, 210, 210, 210, 211, 209, 198, 170, 196, 211, 210, 211, 
    209, 208, 211, 211, 210, 212, 207, 207, 181, 170, 145, 177, 212, 211, 212, 
    203, 211, 211, 212, 212, 211, 185, 213, 189, 192, 181, 181, 213, 213, 214, 
    121, 125, 170, 206, 210, 215, 198, 212, 208, 210, 188, 165, 148, 151, 209, 
    179, 180, 191, 177, 181, 161, 141, 153, 174, 210, 199, 191, 184, 157, 206, 
    93, 93, 134, 167, 193, 143, 81, 114, 150, 196, 181, 162, 149, 154, 148, 
    30, 108, 119, 116, 177, 189, 181, 183, 147, 143, 136, 125, 130, 149, 156, 
    35, 183, 172, 177, 190, 198, 185, 182, 163, 152, 151, 147, 126, 127, 129, 
    75, 111, 114, 117, 123, 130, 137, 123, 116, 114, 99, 94, 84, 87, 98, 
    14, 10, 19, 8, 8, 16, 32, 40, 51, 48, 44, 48, 66, 87, 94, 
    1, 0, 34, 15, 0, 0, 24, 79, 54, 53, 64, 80, 80, 92, 103, 
    15, 0, 0, 0, 0, 0, 0, 83, 79, 72, 53, 56, 72, 96, 124, 
    52, 0, 0, 0, 0, 0, 0, 0, 0, 8, 42, 71, 97, 107, 137, 
    60, 0, 0, 0, 0, 0, 0, 0, 23, 54, 89, 96, 103, 123, 147, 
    
    -- channel=45
    42, 42, 42, 42, 42, 42, 42, 41, 40, 43, 45, 42, 42, 42, 42, 
    43, 43, 43, 43, 43, 43, 43, 42, 43, 46, 47, 43, 42, 43, 43, 
    42, 41, 42, 42, 42, 42, 45, 46, 54, 53, 54, 48, 43, 43, 43, 
    53, 51, 46, 42, 42, 39, 42, 43, 51, 57, 56, 60, 50, 49, 46, 
    60, 56, 46, 40, 43, 42, 45, 43, 49, 54, 60, 58, 53, 53, 49, 
    51, 49, 51, 40, 41, 49, 50, 50, 53, 54, 54, 51, 47, 52, 52, 
    57, 57, 50, 43, 52, 47, 53, 52, 52, 48, 48, 46, 43, 49, 53, 
    41, 41, 38, 37, 44, 40, 49, 54, 50, 48, 48, 46, 48, 49, 56, 
    39, 52, 42, 45, 54, 53, 57, 50, 57, 63, 63, 63, 60, 61, 54, 
    65, 66, 74, 76, 76, 74, 75, 69, 69, 62, 68, 59, 58, 52, 48, 
    31, 36, 41, 41, 41, 48, 63, 62, 59, 57, 55, 53, 52, 41, 35, 
    2, 17, 7, 5, 4, 9, 30, 46, 49, 44, 35, 31, 24, 21, 26, 
    0, 2, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 5, 22, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 27, 41, 
    1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 4, 17, 21, 30, 42, 
    
    -- channel=46
    20, 21, 21, 21, 21, 21, 21, 20, 21, 21, 21, 21, 21, 21, 21, 
    20, 21, 21, 20, 21, 20, 21, 20, 19, 1, 18, 23, 20, 21, 21, 
    20, 21, 21, 21, 21, 20, 22, 10, 8, 3, 11, 26, 21, 21, 22, 
    22, 20, 22, 22, 21, 7, 25, 12, 9, 2, 1, 22, 22, 22, 23, 
    0, 11, 30, 21, 21, 19, 21, 20, 19, 15, 3, 0, 1, 29, 24, 
    5, 7, 9, 10, 18, 2, 12, 16, 22, 13, 11, 7, 0, 15, 23, 
    0, 0, 11, 20, 0, 0, 0, 0, 18, 15, 9, 3, 11, 0, 18, 
    0, 0, 0, 9, 17, 5, 10, 0, 0, 0, 0, 0, 0, 2, 3, 
    22, 12, 8, 13, 16, 11, 18, 8, 6, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 
    
    -- channel=47
    22, 22, 22, 22, 23, 23, 23, 22, 21, 25, 24, 22, 22, 22, 23, 
    23, 23, 23, 23, 23, 23, 23, 22, 26, 43, 35, 26, 23, 23, 23, 
    24, 24, 22, 23, 22, 25, 24, 37, 48, 41, 47, 28, 23, 23, 23, 
    27, 25, 25, 23, 23, 30, 27, 22, 18, 18, 13, 30, 27, 26, 25, 
    78, 68, 35, 23, 24, 16, 20, 19, 24, 36, 57, 64, 68, 43, 28, 
    2, 2, 29, 40, 39, 71, 67, 59, 41, 26, 15, 7, 4, 23, 30, 
    82, 70, 55, 14, 29, 30, 30, 14, 28, 42, 54, 60, 52, 57, 50, 
    23, 18, 31, 37, 23, 0, 0, 42, 51, 39, 30, 20, 16, 11, 32, 
    0, 17, 0, 8, 29, 40, 53, 36, 29, 49, 45, 56, 62, 64, 53, 
    64, 75, 81, 80, 75, 67, 60, 55, 58, 50, 62, 52, 46, 43, 35, 
    56, 52, 68, 74, 79, 83, 89, 82, 76, 69, 60, 49, 36, 29, 25, 
    15, 20, 4, 7, 12, 17, 0, 6, 16, 13, 5, 14, 25, 14, 9, 
    6, 20, 19, 12, 9, 10, 34, 0, 0, 0, 16, 5, 0, 7, 15, 
    5, 7, 7, 6, 6, 6, 0, 0, 0, 0, 0, 0, 8, 16, 23, 
    4, 0, 1, 3, 0, 1, 2, 0, 0, 0, 3, 10, 11, 14, 22, 
    
    -- channel=48
    225, 224, 224, 224, 225, 226, 226, 225, 224, 225, 225, 224, 224, 224, 225, 
    227, 226, 226, 225, 225, 225, 225, 224, 223, 211, 207, 219, 225, 225, 226, 
    227, 226, 226, 226, 226, 226, 225, 221, 204, 176, 186, 218, 226, 227, 228, 
    218, 222, 225, 228, 228, 218, 216, 206, 184, 172, 163, 200, 227, 226, 228, 
    170, 182, 215, 226, 227, 210, 212, 217, 220, 223, 220, 207, 194, 207, 229, 
    159, 172, 204, 207, 215, 211, 213, 218, 224, 210, 178, 167, 148, 182, 226, 
    151, 163, 181, 185, 183, 102, 77, 101, 169, 221, 223, 211, 200, 200, 206, 
    60, 111, 122, 161, 182, 155, 169, 192, 178, 151, 121, 106, 115, 130, 165, 
    77, 171, 160, 180, 211, 217, 219, 191, 174, 179, 182, 178, 174, 171, 154, 
    146, 170, 173, 174, 173, 168, 152, 135, 137, 121, 120, 103, 96, 104, 117, 
    30, 42, 49, 56, 68, 85, 99, 101, 98, 85, 73, 70, 77, 89, 109, 
    0, 10, 19, 0, 0, 0, 16, 22, 21, 26, 42, 74, 104, 102, 110, 
    0, 0, 0, 0, 0, 0, 67, 124, 117, 110, 99, 75, 72, 99, 137, 
    0, 0, 0, 0, 0, 0, 4, 34, 31, 15, 25, 69, 96, 116, 154, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 51, 88, 95, 105, 128, 161, 
    
    -- channel=49
    76, 76, 76, 76, 76, 76, 76, 75, 75, 75, 76, 75, 76, 76, 76, 
    76, 76, 76, 76, 76, 76, 76, 76, 73, 56, 63, 76, 76, 76, 76, 
    73, 74, 76, 76, 77, 75, 75, 65, 50, 45, 47, 70, 76, 76, 77, 
    79, 78, 76, 77, 77, 66, 71, 69, 78, 79, 82, 81, 77, 77, 77, 
    21, 29, 68, 73, 75, 73, 78, 77, 81, 74, 52, 36, 27, 54, 77, 
    79, 87, 69, 50, 53, 23, 23, 33, 57, 75, 79, 83, 76, 83, 76, 
    8, 23, 38, 69, 64, 25, 37, 64, 80, 63, 45, 31, 34, 32, 48, 
    22, 59, 24, 48, 66, 86, 93, 55, 37, 43, 46, 52, 58, 70, 64, 
    64, 67, 77, 75, 72, 62, 56, 51, 56, 47, 51, 38, 30, 25, 33, 
    32, 25, 30, 34, 39, 44, 46, 46, 44, 38, 31, 27, 29, 29, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 6, 15, 32, 35, 35, 
    0, 0, 0, 0, 0, 0, 51, 48, 38, 40, 47, 44, 28, 24, 41, 
    0, 0, 0, 0, 0, 0, 0, 17, 17, 7, 0, 3, 23, 33, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 23, 21, 33, 49, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 17, 16, 27, 38, 54, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 48, 0, 0, 0, 40, 26, 1, 0, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 0, 0, 0, 13, 38, 26, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 25, 
    0, 20, 17, 22, 22, 21, 21, 14, 0, 8, 1, 22, 0, 0, 0, 
    49, 56, 44, 54, 51, 51, 45, 41, 38, 41, 33, 22, 12, 0, 0, 
    23, 0, 0, 0, 10, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 31, 36, 24, 13, 0, 0, 0, 0, 0, 46, 0, 0, 0, 
    12, 13, 13, 20, 16, 15, 0, 0, 0, 37, 0, 0, 0, 0, 0, 
    39, 3, 5, 10, 10, 9, 0, 22, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    17, 17, 17, 17, 17, 17, 17, 16, 17, 16, 16, 17, 17, 17, 17, 
    17, 17, 17, 17, 17, 17, 17, 18, 15, 5, 15, 16, 17, 17, 17, 
    16, 16, 18, 18, 17, 15, 17, 10, 7, 6, 1, 16, 16, 17, 17, 
    15, 16, 16, 17, 17, 11, 19, 17, 22, 19, 24, 14, 17, 17, 17, 
    4, 8, 17, 17, 17, 18, 16, 16, 15, 7, 0, 4, 2, 18, 18, 
    15, 18, 6, 7, 8, 0, 0, 0, 12, 19, 24, 21, 20, 16, 16, 
    0, 3, 2, 26, 6, 22, 22, 31, 13, 2, 0, 0, 0, 0, 11, 
    15, 12, 13, 10, 21, 26, 16, 0, 7, 15, 18, 19, 20, 19, 8, 
    22, 0, 18, 5, 4, 6, 1, 6, 6, 0, 0, 0, 0, 1, 8, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 1, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 9, 
    8, 2, 7, 6, 3, 0, 25, 15, 12, 13, 16, 4, 0, 12, 18, 
    6, 7, 1, 5, 8, 7, 0, 0, 2, 0, 0, 12, 15, 16, 19, 
    11, 8, 6, 6, 8, 8, 4, 0, 0, 12, 19, 12, 18, 19, 17, 
    17, 15, 14, 12, 13, 13, 16, 12, 22, 17, 16, 21, 19, 20, 19, 
    
    -- channel=52
    98, 96, 96, 96, 96, 96, 96, 96, 95, 97, 97, 96, 95, 96, 95, 
    98, 96, 96, 96, 95, 96, 96, 95, 97, 99, 72, 87, 96, 95, 96, 
    97, 96, 95, 96, 96, 98, 95, 102, 92, 81, 79, 77, 96, 96, 96, 
    93, 98, 95, 96, 98, 96, 80, 91, 76, 76, 71, 83, 98, 96, 96, 
    67, 68, 67, 94, 97, 87, 87, 91, 94, 105, 105, 91, 86, 67, 92, 
    78, 79, 88, 95, 88, 110, 91, 91, 84, 83, 77, 75, 71, 69, 93, 
    66, 54, 71, 70, 81, 74, 20, 24, 67, 101, 105, 99, 83, 86, 76, 
    0, 36, 55, 43, 60, 67, 73, 98, 73, 60, 53, 43, 45, 51, 79, 
    7, 71, 78, 86, 97, 100, 98, 95, 86, 93, 84, 92, 80, 72, 61, 
    54, 79, 78, 82, 80, 77, 73, 66, 63, 66, 57, 50, 47, 47, 44, 
    11, 0, 19, 19, 20, 27, 42, 49, 46, 43, 35, 30, 24, 39, 40, 
    0, 0, 4, 0, 0, 0, 0, 21, 8, 10, 11, 36, 47, 35, 33, 
    0, 0, 0, 0, 0, 0, 0, 49, 53, 52, 42, 14, 22, 29, 44, 
    13, 0, 0, 0, 0, 0, 0, 18, 23, 0, 0, 19, 29, 36, 48, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 3, 26, 28, 31, 42, 54, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 36, 8, 0, 0, 0, 0, 0, 0, 0, 0, 12, 25, 20, 0, 
    0, 0, 0, 8, 9, 20, 29, 22, 9, 0, 0, 0, 0, 0, 0, 
    36, 40, 25, 0, 0, 0, 0, 0, 0, 0, 8, 18, 19, 13, 18, 
    0, 0, 0, 13, 0, 0, 0, 0, 14, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 12, 12, 
    0, 23, 22, 22, 18, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 21, 26, 36, 41, 42, 33, 31, 22, 16, 10, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 8, 0, 0, 45, 46, 26, 22, 27, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 62, 58, 33, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=54
    110, 109, 109, 109, 109, 110, 110, 110, 110, 108, 111, 109, 109, 109, 110, 
    111, 110, 110, 110, 110, 110, 110, 110, 107, 103, 116, 113, 110, 110, 110, 
    113, 112, 111, 110, 111, 109, 112, 103, 105, 92, 84, 119, 111, 111, 111, 
    106, 107, 109, 112, 113, 106, 112, 99, 82, 68, 62, 76, 108, 109, 110, 
    99, 107, 121, 114, 112, 105, 94, 106, 100, 99, 99, 104, 104, 122, 111, 
    50, 58, 77, 104, 111, 102, 120, 122, 126, 107, 75, 59, 52, 65, 106, 
    94, 112, 106, 99, 75, 42, 36, 45, 63, 97, 107, 110, 112, 103, 117, 
    48, 26, 49, 84, 99, 61, 46, 63, 99, 94, 66, 51, 46, 52, 53, 
    25, 68, 61, 71, 94, 104, 104, 97, 69, 71, 83, 75, 85, 89, 88, 
    55, 104, 101, 105, 104, 98, 87, 71, 71, 63, 57, 56, 42, 44, 57, 
    18, 37, 35, 45, 52, 65, 72, 73, 66, 59, 49, 44, 44, 33, 46, 
    0, 0, 6, 0, 0, 0, 25, 0, 0, 2, 8, 11, 39, 55, 51, 
    0, 0, 9, 0, 0, 0, 42, 109, 83, 71, 73, 73, 42, 41, 55, 
    0, 0, 0, 0, 0, 0, 14, 104, 99, 73, 27, 21, 39, 47, 65, 
    0, 0, 0, 0, 0, 0, 0, 44, 18, 11, 30, 38, 41, 49, 65, 
    
    -- channel=55
    12, 12, 12, 12, 12, 12, 12, 12, 10, 11, 13, 12, 12, 12, 12, 
    12, 12, 12, 12, 12, 11, 11, 12, 9, 11, 12, 10, 12, 12, 12, 
    11, 12, 11, 12, 12, 10, 13, 9, 13, 17, 16, 17, 12, 11, 12, 
    16, 16, 14, 11, 11, 10, 7, 15, 25, 33, 29, 17, 16, 14, 14, 
    3, 1, 7, 11, 10, 18, 13, 16, 18, 16, 22, 16, 5, 10, 15, 
    37, 34, 28, 4, 0, 7, 7, 10, 21, 27, 25, 30, 32, 13, 20, 
    4, 8, 3, 10, 30, 9, 20, 12, 5, 17, 14, 9, 10, 16, 10, 
    24, 6, 11, 0, 15, 23, 30, 29, 10, 7, 8, 10, 15, 18, 15, 
    0, 43, 23, 24, 25, 21, 13, 22, 27, 34, 32, 31, 26, 21, 14, 
    37, 20, 23, 24, 25, 26, 34, 27, 28, 22, 29, 25, 23, 22, 19, 
    0, 0, 1, 0, 0, 4, 15, 19, 21, 20, 19, 22, 24, 14, 12, 
    0, 0, 4, 0, 0, 0, 25, 29, 27, 24, 22, 13, 16, 2, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 
    
    -- channel=56
    167, 167, 167, 167, 167, 167, 167, 167, 167, 166, 166, 167, 167, 167, 168, 
    167, 167, 167, 167, 167, 167, 167, 167, 165, 141, 150, 167, 167, 167, 168, 
    164, 165, 168, 168, 169, 167, 165, 154, 129, 119, 125, 156, 167, 168, 169, 
    167, 167, 169, 169, 168, 158, 163, 154, 155, 150, 153, 170, 169, 170, 171, 
    94, 108, 167, 164, 167, 162, 168, 165, 168, 160, 135, 118, 108, 139, 172, 
    145, 158, 154, 132, 146, 99, 103, 115, 138, 160, 161, 156, 141, 168, 169, 
    68, 79, 118, 147, 142, 71, 84, 128, 165, 151, 128, 109, 112, 108, 127, 
    49, 133, 88, 125, 148, 158, 168, 130, 108, 107, 105, 111, 119, 136, 140, 
    122, 137, 146, 147, 150, 147, 145, 125, 125, 110, 117, 101, 92, 91, 99, 
    81, 77, 84, 85, 91, 97, 97, 93, 93, 80, 74, 67, 71, 74, 88, 
    8, 26, 14, 8, 10, 15, 23, 24, 33, 27, 32, 42, 68, 85, 91, 
    3, 21, 32, 12, 0, 0, 76, 72, 62, 66, 81, 90, 70, 75, 106, 
    5, 1, 0, 0, 0, 0, 45, 63, 59, 45, 28, 44, 78, 96, 128, 
    19, 0, 0, 0, 0, 0, 10, 0, 0, 11, 62, 84, 88, 106, 131, 
    22, 13, 10, 7, 6, 7, 11, 12, 51, 80, 84, 87, 100, 116, 139, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 8, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 2, 15, 21, 17, 10, 2, 17, 6, 6, 10, 16, 7, 1, 5, 
    28, 15, 8, 15, 18, 18, 0, 18, 30, 28, 13, 2, 15, 8, 2, 
    28, 20, 19, 19, 20, 20, 12, 46, 43, 24, 29, 23, 10, 3, 0, 
    19, 27, 25, 22, 23, 23, 20, 25, 35, 30, 21, 8, 7, 3, 0, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 21, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 9, 9, 1, 30, 0, 0, 
    0, 0, 0, 0, 17, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 25, 0, 6, 0, 6, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 13, 0, 11, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 25, 29, 13, 0, 0, 24, 2, 0, 0, 0, 0, 0, 0, 
    41, 0, 0, 18, 11, 0, 0, 17, 9, 11, 6, 0, 0, 0, 0, 
    93, 3, 0, 6, 2, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 
    85, 13, 3, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=61
    30, 30, 30, 30, 30, 31, 31, 31, 32, 29, 30, 31, 31, 30, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 29, 24, 38, 34, 31, 31, 31, 
    32, 32, 32, 31, 31, 30, 31, 25, 28, 22, 21, 37, 31, 31, 31, 
    26, 27, 31, 32, 31, 29, 36, 27, 15, 7, 6, 17, 28, 29, 31, 
    34, 41, 42, 33, 32, 32, 26, 29, 23, 18, 18, 28, 32, 46, 31, 
    0, 0, 19, 29, 36, 23, 36, 36, 38, 29, 14, 3, 0, 11, 29, 
    27, 37, 34, 26, 13, 0, 8, 15, 13, 23, 25, 28, 32, 29, 38, 
    15, 0, 15, 36, 35, 1, 0, 3, 30, 29, 16, 10, 8, 7, 3, 
    6, 15, 0, 7, 17, 24, 26, 15, 4, 0, 6, 2, 12, 23, 25, 
    3, 19, 19, 17, 18, 17, 12, 6, 6, 0, 3, 3, 0, 0, 10, 
    6, 13, 5, 11, 15, 16, 8, 8, 6, 2, 1, 0, 5, 0, 10, 
    0, 6, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 19, 18, 
    0, 0, 13, 9, 0, 0, 35, 44, 33, 27, 28, 39, 18, 16, 19, 
    0, 0, 0, 0, 0, 0, 5, 41, 43, 41, 18, 10, 20, 19, 24, 
    2, 0, 0, 0, 0, 0, 0, 20, 18, 12, 19, 20, 19, 19, 22, 
    
    -- channel=62
    82, 80, 80, 80, 80, 81, 81, 82, 81, 81, 81, 80, 81, 80, 80, 
    82, 81, 81, 81, 81, 81, 81, 81, 81, 88, 73, 76, 81, 81, 81, 
    83, 81, 82, 82, 80, 83, 80, 86, 83, 86, 50, 68, 83, 82, 82, 
    74, 79, 81, 82, 81, 91, 74, 93, 64, 59, 45, 41, 82, 82, 82, 
    72, 71, 77, 81, 82, 90, 61, 83, 72, 86, 83, 83, 82, 68, 82, 
    41, 32, 48, 75, 87, 84, 85, 85, 78, 90, 72, 52, 50, 21, 74, 
    65, 55, 75, 66, 70, 66, 12, 17, 27, 76, 85, 87, 86, 75, 68, 
    0, 17, 41, 35, 80, 64, 31, 54, 70, 70, 54, 38, 27, 38, 34, 
    0, 52, 41, 37, 55, 78, 82, 93, 56, 54, 63, 63, 59, 63, 68, 
    0, 67, 61, 64, 63, 62, 58, 47, 45, 49, 37, 45, 26, 26, 31, 
    19, 18, 26, 29, 33, 36, 42, 39, 40, 35, 29, 21, 19, 24, 24, 
    6, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 35, 24, 
    0, 0, 0, 4, 0, 0, 0, 59, 34, 31, 29, 37, 27, 20, 30, 
    31, 0, 0, 0, 0, 0, 0, 7, 13, 17, 6, 3, 29, 30, 40, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 34, 32, 35, 43, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 14, 0, 0, 0, 
    8, 17, 18, 0, 0, 0, 6, 0, 0, 0, 0, 0, 3, 22, 0, 
    0, 0, 4, 2, 7, 0, 13, 11, 9, 0, 0, 0, 0, 21, 0, 
    7, 20, 10, 2, 0, 0, 4, 12, 19, 0, 0, 0, 4, 5, 16, 
    19, 14, 4, 32, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 5, 
    65, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    10, 19, 6, 12, 18, 17, 3, 3, 0, 0, 0, 1, 4, 0, 11, 
    6, 37, 1, 2, 12, 23, 21, 0, 0, 0, 0, 0, 5, 9, 17, 
    4, 30, 28, 14, 17, 21, 93, 10, 9, 8, 16, 21, 17, 20, 21, 
    0, 20, 24, 20, 21, 21, 63, 45, 33, 36, 28, 29, 17, 20, 18, 
    0, 18, 20, 20, 20, 20, 34, 37, 30, 36, 20, 16, 18, 17, 16, 
    
    -- channel=64
    9, 25, 35, 31, 39, 40, 46, 42, 50, 48, 46, 54, 45, 49, 53, 
    15, 31, 44, 36, 47, 42, 45, 50, 49, 17, 54, 59, 46, 50, 56, 
    22, 32, 50, 44, 50, 45, 37, 40, 48, 0, 49, 52, 43, 53, 57, 
    26, 37, 45, 57, 52, 53, 41, 26, 0, 0, 5, 4, 52, 44, 55, 
    11, 10, 13, 22, 25, 26, 24, 4, 1, 0, 3, 24, 32, 26, 20, 
    12, 10, 0, 19, 18, 8, 5, 0, 3, 7, 35, 50, 10, 55, 0, 
    3, 0, 0, 16, 17, 10, 9, 9, 11, 13, 38, 42, 31, 14, 0, 
    5, 13, 20, 18, 18, 15, 12, 5, 15, 0, 33, 44, 34, 7, 35, 
    0, 0, 18, 17, 3, 2, 6, 14, 22, 19, 36, 29, 27, 21, 28, 
    0, 13, 9, 3, 14, 14, 13, 3, 16, 26, 26, 14, 6, 0, 8, 
    11, 2, 1, 0, 1, 19, 0, 0, 17, 12, 3, 0, 0, 0, 0, 
    15, 4, 0, 0, 4, 14, 0, 0, 5, 1, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    53, 40, 55, 57, 57, 55, 60, 62, 59, 62, 58, 61, 61, 63, 59, 
    53, 38, 54, 54, 58, 52, 54, 58, 58, 51, 36, 58, 58, 62, 54, 
    53, 37, 51, 54, 60, 52, 55, 46, 49, 44, 33, 50, 53, 56, 54, 
    43, 26, 39, 37, 49, 46, 56, 45, 15, 12, 0, 0, 24, 45, 37, 
    7, 0, 10, 10, 12, 14, 17, 33, 24, 26, 18, 30, 31, 25, 8, 
    19, 29, 29, 18, 32, 35, 32, 31, 26, 30, 34, 53, 35, 46, 30, 
    24, 13, 18, 12, 29, 30, 37, 35, 41, 45, 39, 40, 48, 39, 0, 
    34, 35, 44, 47, 48, 49, 52, 44, 41, 32, 17, 30, 36, 18, 29, 
    28, 17, 20, 36, 41, 35, 33, 37, 43, 47, 43, 39, 34, 34, 39, 
    22, 38, 40, 31, 32, 46, 48, 41, 28, 39, 37, 37, 25, 14, 5, 
    26, 36, 35, 31, 26, 27, 31, 11, 14, 34, 22, 18, 15, 14, 8, 
    25, 28, 25, 12, 19, 33, 34, 19, 13, 20, 20, 10, 11, 4, 2, 
    22, 21, 22, 12, 6, 7, 12, 19, 13, 7, 12, 10, 5, 2, 3, 
    0, 0, 3, 8, 11, 8, 5, 8, 15, 18, 4, 2, 2, 4, 5, 
    1, 1, 5, 6, 11, 13, 12, 7, 4, 9, 1, 0, 3, 4, 0, 
    
    -- channel=66
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 7, 1, 20, 9, 0, 0, 0, 7, 9, 27, 47, 0, 13, 
    0, 0, 0, 0, 0, 16, 16, 39, 44, 28, 0, 0, 11, 0, 3, 
    16, 33, 34, 20, 6, 0, 0, 0, 0, 0, 0, 0, 0, 65, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 6, 0, 0, 0, 0, 
    24, 6, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 1, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    
    -- channel=67
    35, 37, 57, 49, 53, 47, 52, 47, 55, 53, 50, 52, 41, 52, 48, 
    34, 36, 59, 42, 56, 44, 53, 59, 52, 43, 56, 59, 41, 55, 50, 
    34, 31, 56, 38, 52, 40, 47, 60, 54, 22, 64, 71, 44, 57, 55, 
    39, 26, 55, 56, 51, 46, 41, 27, 40, 32, 43, 49, 88, 63, 61, 
    49, 40, 47, 60, 57, 58, 49, 40, 17, 20, 28, 3, 34, 33, 31, 
    21, 8, 13, 19, 19, 8, 27, 19, 21, 14, 16, 26, 0, 61, 0, 
    31, 14, 16, 36, 38, 20, 22, 10, 6, 13, 33, 47, 21, 20, 0, 
    17, 11, 14, 24, 34, 33, 32, 30, 44, 30, 54, 43, 28, 0, 0, 
    30, 50, 48, 50, 43, 48, 45, 32, 27, 10, 24, 27, 31, 15, 45, 
    11, 22, 41, 42, 34, 26, 29, 33, 43, 40, 35, 29, 35, 25, 25, 
    47, 33, 32, 33, 51, 55, 29, 15, 23, 46, 41, 27, 14, 9, 15, 
    56, 35, 27, 18, 18, 42, 29, 18, 25, 21, 13, 19, 3, 7, 0, 
    42, 38, 34, 28, 34, 31, 15, 13, 19, 21, 2, 10, 4, 2, 0, 
    20, 17, 12, 12, 13, 16, 15, 9, 6, 0, 8, 4, 0, 1, 0, 
    1, 1, 1, 1, 0, 0, 4, 6, 24, 0, 7, 1, 1, 4, 0, 
    
    -- channel=68
    39, 33, 29, 29, 24, 21, 16, 17, 14, 14, 13, 10, 16, 13, 13, 
    33, 25, 19, 21, 14, 15, 14, 13, 13, 26, 20, 11, 14, 11, 11, 
    24, 20, 10, 11, 5, 11, 12, 14, 13, 32, 14, 7, 11, 5, 6, 
    17, 12, 3, 0, 1, 2, 8, 11, 37, 57, 45, 49, 16, 2, 0, 
    33, 29, 34, 25, 25, 22, 30, 37, 35, 32, 29, 18, 0, 12, 24, 
    30, 25, 23, 27, 27, 34, 34, 42, 32, 30, 14, 0, 10, 0, 23, 
    32, 35, 40, 34, 41, 42, 44, 42, 36, 29, 9, 7, 13, 11, 26, 
    37, 31, 27, 28, 33, 35, 35, 34, 30, 30, 17, 11, 14, 27, 15, 
    44, 42, 45, 41, 44, 43, 42, 37, 27, 21, 7, 15, 20, 16, 10, 
    54, 37, 32, 43, 45, 35, 26, 25, 23, 22, 21, 23, 22, 28, 26, 
    39, 45, 42, 38, 35, 33, 40, 47, 32, 23, 28, 35, 29, 26, 21, 
    34, 42, 48, 49, 42, 30, 31, 25, 27, 32, 30, 29, 31, 26, 26, 
    30, 33, 35, 30, 34, 37, 35, 27, 26, 31, 30, 22, 28, 26, 24, 
    33, 34, 31, 26, 23, 24, 30, 30, 22, 26, 26, 26, 26, 23, 21, 
    21, 21, 23, 24, 25, 22, 24, 22, 18, 32, 23, 26, 24, 22, 22, 
    
    -- channel=69
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=70
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 5, 0, 0, 
    10, 20, 3, 3, 30, 20, 2, 0, 0, 8, 49, 74, 27, 0, 0, 
    0, 0, 0, 0, 0, 7, 23, 40, 57, 47, 29, 0, 0, 0, 0, 
    31, 47, 72, 64, 32, 19, 14, 0, 0, 0, 0, 0, 0, 6, 80, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 27, 42, 0, 0, 0, 0, 
    8, 46, 11, 0, 0, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 22, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    17, 1, 0, 14, 6, 0, 0, 0, 0, 0, 25, 10, 0, 44, 0, 
    0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 8, 4, 0, 0, 7, 
    0, 0, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 12, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 20, 0, 0, 0, 0, 1, 0, 
    0, 3, 2, 2, 4, 0, 0, 0, 18, 0, 0, 0, 0, 5, 0, 
    
    -- channel=72
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=74
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 26, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 31, 23, 10, 33, 32, 3, 3, 0, 
    13, 7, 24, 22, 13, 4, 2, 0, 57, 50, 35, 88, 88, 41, 45, 
    71, 59, 60, 75, 76, 78, 63, 46, 8, 0, 5, 0, 0, 0, 49, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 29, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 22, 35, 11, 0, 0, 0, 
    14, 39, 17, 2, 11, 26, 18, 0, 0, 0, 0, 0, 0, 0, 28, 
    0, 0, 0, 8, 0, 0, 0, 22, 35, 0, 0, 10, 40, 46, 38, 
    2, 0, 0, 21, 46, 28, 6, 16, 6, 33, 48, 40, 27, 16, 20, 
    10, 5, 1, 2, 0, 6, 33, 12, 10, 15, 26, 17, 4, 10, 5, 
    28, 45, 48, 33, 37, 34, 10, 6, 26, 24, 4, 9, 11, 2, 0, 
    30, 31, 17, 11, 15, 22, 16, 8, 0, 0, 7, 5, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 17, 1, 2, 1, 0, 0, 10, 
    
    -- channel=75
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=76
    182, 155, 186, 199, 204, 204, 209, 216, 204, 215, 213, 215, 219, 218, 212, 
    185, 155, 185, 200, 201, 199, 199, 203, 204, 205, 161, 207, 219, 215, 210, 
    184, 150, 177, 197, 195, 193, 191, 169, 178, 196, 110, 180, 208, 198, 197, 
    165, 134, 155, 166, 180, 176, 183, 164, 131, 107, 79, 76, 94, 159, 158, 
    81, 74, 85, 80, 98, 102, 116, 127, 103, 91, 78, 88, 99, 129, 87, 
    64, 77, 95, 79, 102, 105, 108, 109, 93, 97, 97, 141, 150, 106, 112, 
    79, 81, 81, 74, 111, 131, 131, 131, 130, 128, 122, 151, 159, 111, 94, 
    108, 115, 118, 135, 150, 160, 164, 156, 143, 136, 99, 123, 142, 133, 98, 
    104, 100, 108, 139, 151, 145, 144, 142, 135, 147, 121, 138, 137, 129, 118, 
    112, 100, 126, 133, 136, 142, 144, 134, 118, 137, 139, 136, 111, 90, 65, 
    107, 128, 126, 116, 102, 118, 134, 94, 73, 105, 106, 95, 70, 55, 39, 
    79, 117, 119, 85, 82, 89, 110, 83, 74, 80, 68, 58, 47, 32, 23, 
    65, 85, 82, 64, 63, 62, 61, 59, 53, 52, 47, 36, 37, 20, 17, 
    25, 24, 28, 29, 35, 37, 39, 41, 40, 55, 29, 23, 20, 17, 18, 
    14, 14, 21, 24, 30, 33, 34, 29, 22, 52, 16, 16, 15, 16, 13, 
    
    -- channel=77
    76, 74, 76, 73, 66, 59, 54, 50, 53, 51, 47, 46, 49, 49, 48, 
    65, 61, 62, 55, 51, 46, 45, 45, 48, 48, 44, 44, 44, 44, 44, 
    52, 50, 47, 39, 37, 38, 37, 41, 43, 39, 47, 46, 38, 34, 40, 
    35, 32, 25, 18, 17, 23, 26, 31, 45, 44, 50, 42, 32, 24, 20, 
    33, 32, 33, 30, 22, 25, 33, 44, 48, 52, 51, 32, 30, 16, 21, 
    46, 42, 41, 41, 45, 51, 62, 61, 52, 47, 45, 32, 17, 11, 26, 
    57, 45, 46, 55, 62, 63, 70, 65, 62, 58, 44, 30, 16, 21, 11, 
    64, 55, 59, 71, 73, 76, 77, 72, 64, 47, 32, 22, 25, 19, 12, 
    71, 65, 70, 77, 80, 78, 73, 61, 54, 39, 36, 35, 36, 28, 24, 
    68, 68, 75, 74, 71, 68, 61, 55, 51, 48, 44, 38, 36, 29, 26, 
    76, 79, 73, 65, 64, 64, 58, 47, 46, 48, 45, 39, 33, 29, 23, 
    70, 70, 66, 58, 57, 60, 49, 41, 42, 40, 39, 37, 29, 26, 18, 
    59, 58, 53, 49, 47, 44, 38, 40, 40, 36, 29, 31, 25, 24, 22, 
    33, 32, 33, 34, 32, 33, 36, 31, 33, 33, 26, 23, 23, 23, 20, 
    17, 19, 24, 25, 28, 30, 32, 23, 29, 28, 22, 20, 23, 23, 12, 
    
    -- channel=78
    0, 1, 12, 11, 14, 15, 19, 16, 21, 23, 18, 25, 20, 21, 23, 
    0, 3, 17, 11, 18, 13, 17, 21, 21, 0, 25, 27, 19, 22, 24, 
    0, 3, 17, 13, 18, 14, 9, 13, 23, 0, 18, 24, 15, 21, 24, 
    0, 2, 8, 16, 13, 15, 11, 0, 0, 0, 0, 0, 21, 12, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    48, 44, 45, 45, 40, 36, 32, 28, 30, 32, 30, 25, 26, 27, 24, 
    44, 39, 38, 36, 32, 31, 33, 28, 28, 46, 32, 23, 26, 28, 24, 
    37, 33, 30, 24, 26, 23, 29, 38, 34, 40, 44, 35, 28, 25, 25, 
    32, 27, 31, 19, 18, 18, 19, 28, 55, 47, 51, 72, 50, 32, 26, 
    49, 44, 45, 48, 42, 43, 41, 46, 37, 40, 39, 12, 17, 20, 39, 
    24, 25, 29, 16, 16, 26, 39, 44, 36, 28, 11, 0, 10, 5, 21, 
    41, 37, 37, 36, 42, 33, 37, 26, 23, 26, 24, 25, 7, 32, 21, 
    33, 20, 16, 27, 36, 40, 45, 51, 50, 51, 35, 20, 16, 0, 0, 
    63, 57, 53, 53, 62, 63, 58, 41, 34, 13, 10, 19, 24, 25, 26, 
    37, 37, 45, 56, 46, 41, 42, 53, 43, 33, 30, 36, 44, 42, 34, 
    49, 52, 56, 57, 65, 49, 51, 43, 40, 51, 50, 44, 39, 30, 34, 
    55, 54, 55, 45, 36, 52, 51, 35, 37, 40, 44, 35, 33, 31, 23, 
    55, 62, 58, 51, 52, 49, 37, 37, 44, 38, 32, 33, 29, 25, 20, 
    46, 43, 38, 36, 36, 36, 36, 35, 20, 32, 27, 27, 24, 22, 23, 
    20, 19, 22, 23, 23, 25, 30, 30, 29, 29, 25, 22, 24, 21, 25, 
    
    -- channel=80
    182, 177, 209, 219, 225, 225, 230, 225, 226, 237, 233, 235, 231, 233, 232, 
    185, 178, 210, 216, 222, 217, 222, 223, 225, 216, 201, 231, 233, 233, 234, 
    186, 174, 205, 209, 214, 207, 203, 201, 214, 176, 173, 227, 225, 220, 228, 
    178, 164, 194, 201, 201, 198, 189, 173, 153, 104, 98, 120, 168, 197, 201, 
    116, 112, 113, 128, 139, 147, 149, 136, 106, 96, 91, 85, 119, 130, 121, 
    62, 78, 87, 77, 89, 95, 114, 108, 95, 87, 97, 135, 121, 116, 88, 
    86, 87, 76, 92, 120, 123, 119, 108, 104, 110, 142, 174, 144, 127, 83, 
    101, 101, 107, 134, 155, 165, 169, 168, 166, 146, 134, 146, 148, 90, 52, 
    126, 127, 136, 164, 174, 171, 161, 142, 140, 124, 123, 142, 144, 134, 135, 
    94, 107, 141, 149, 142, 144, 152, 155, 148, 150, 151, 147, 133, 104, 83, 
    130, 136, 140, 135, 140, 149, 135, 88, 93, 135, 133, 104, 76, 54, 44, 
    111, 132, 116, 82, 78, 116, 123, 92, 86, 84, 75, 58, 39, 31, 13, 
    99, 117, 103, 88, 84, 76, 64, 64, 66, 57, 40, 42, 30, 14, 8, 
    38, 36, 33, 36, 44, 44, 43, 37, 38, 41, 26, 20, 13, 10, 12, 
    7, 6, 11, 15, 19, 25, 30, 25, 43, 32, 14, 10, 9, 12, 1, 
    
    -- channel=81
    70, 70, 84, 82, 84, 78, 80, 78, 80, 81, 73, 82, 79, 82, 82, 
    65, 63, 76, 73, 75, 70, 70, 74, 77, 57, 57, 80, 76, 77, 79, 
    59, 53, 67, 66, 67, 65, 59, 50, 58, 37, 49, 62, 63, 65, 73, 
    44, 41, 45, 49, 50, 55, 51, 48, 21, 11, 18, 0, 28, 38, 39, 
    5, 10, 7, 8, 8, 13, 21, 22, 27, 25, 25, 30, 30, 25, 10, 
    26, 27, 23, 28, 48, 39, 44, 30, 27, 30, 46, 70, 37, 40, 15, 
    29, 22, 16, 38, 47, 57, 60, 61, 62, 56, 56, 46, 40, 7, 0, 
    48, 53, 68, 73, 71, 71, 68, 57, 50, 26, 25, 39, 42, 33, 46, 
    38, 29, 46, 65, 58, 49, 47, 49, 51, 49, 52, 46, 42, 34, 19, 
    45, 60, 58, 48, 54, 59, 52, 34, 32, 46, 47, 36, 17, 1, 0, 
    50, 54, 48, 35, 27, 42, 36, 15, 24, 28, 17, 6, 2, 0, 0, 
    40, 44, 35, 25, 35, 36, 18, 16, 16, 12, 2, 0, 0, 0, 0, 
    20, 15, 7, 9, 5, 5, 10, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 79, 25, 38, 6, 0, 0, 
    31, 18, 28, 7, 19, 7, 16, 13, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 25, 0, 
    0, 8, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 21, 23, 
    0, 0, 0, 0, 0, 4, 0, 42, 0, 0, 3, 29, 12, 20, 0, 
    0, 0, 4, 26, 2, 0, 0, 0, 0, 7, 0, 31, 9, 12, 25, 
    0, 0, 12, 0, 17, 34, 16, 0, 0, 27, 12, 0, 20, 13, 11, 
    25, 34, 22, 4, 0, 10, 20, 18, 2, 0, 18, 7, 16, 6, 0, 
    12, 8, 9, 8, 3, 0, 0, 8, 0, 27, 5, 12, 6, 7, 12, 
    
    -- channel=83
    2, 10, 7, 7, 8, 13, 13, 13, 14, 12, 15, 18, 18, 15, 18, 
    5, 14, 10, 12, 12, 14, 11, 14, 16, 5, 21, 17, 17, 13, 20, 
    9, 17, 15, 19, 14, 19, 9, 8, 14, 6, 9, 12, 17, 15, 19, 
    7, 16, 5, 15, 13, 17, 13, 10, 7, 8, 10, 3, 6, 8, 13, 
    0, 8, 3, 1, 4, 3, 8, 0, 6, 0, 5, 15, 11, 13, 13, 
    10, 9, 4, 17, 13, 8, 3, 0, 3, 6, 18, 18, 17, 11, 9, 
    0, 7, 3, 9, 5, 12, 5, 13, 15, 11, 13, 13, 15, 0, 18, 
    4, 9, 6, 2, 2, 4, 2, 0, 1, 0, 13, 15, 14, 30, 25, 
    0, 0, 2, 0, 0, 0, 7, 12, 8, 14, 14, 13, 13, 9, 2, 
    7, 0, 0, 0, 9, 5, 1, 0, 10, 10, 9, 1, 1, 4, 11, 
    4, 0, 0, 0, 0, 9, 3, 9, 12, 0, 1, 4, 5, 8, 0, 
    0, 2, 0, 7, 8, 0, 0, 5, 8, 5, 2, 10, 4, 6, 7, 
    0, 0, 0, 0, 1, 4, 4, 2, 1, 7, 6, 5, 4, 5, 7, 
    0, 3, 4, 2, 2, 5, 7, 6, 13, 0, 6, 4, 6, 6, 4, 
    6, 8, 8, 9, 8, 7, 4, 3, 9, 6, 3, 5, 5, 6, 0, 
    
    -- channel=84
    86, 82, 85, 98, 97, 102, 98, 95, 92, 101, 103, 95, 104, 97, 100, 
    85, 81, 82, 98, 87, 96, 92, 86, 94, 101, 80, 93, 106, 95, 101, 
    83, 83, 79, 89, 81, 87, 82, 80, 88, 86, 61, 88, 99, 83, 91, 
    79, 81, 82, 79, 78, 77, 76, 77, 74, 43, 37, 55, 41, 76, 78, 
    45, 46, 44, 48, 55, 56, 63, 59, 49, 44, 36, 40, 49, 46, 55, 
    17, 38, 40, 27, 31, 49, 53, 57, 43, 36, 36, 47, 70, 10, 55, 
    35, 44, 36, 32, 47, 54, 53, 52, 48, 46, 57, 70, 58, 75, 51, 
    51, 48, 48, 66, 75, 78, 79, 84, 73, 73, 43, 52, 63, 50, 8, 
    68, 57, 55, 69, 87, 79, 68, 56, 60, 55, 51, 64, 62, 65, 53, 
    49, 49, 64, 71, 59, 64, 71, 76, 61, 57, 66, 69, 60, 48, 33, 
    48, 64, 69, 67, 62, 52, 62, 42, 37, 52, 57, 45, 33, 21, 16, 
    31, 57, 54, 37, 29, 47, 60, 44, 33, 32, 33, 16, 15, 9, 3, 
    38, 54, 45, 39, 29, 23, 23, 27, 27, 17, 14, 13, 11, 1, 0, 
    9, 6, 5, 8, 14, 12, 9, 10, 3, 24, 5, 6, 1, 0, 0, 
    0, 0, 0, 0, 0, 5, 8, 8, 1, 21, 0, 0, 0, 0, 0, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 7, 0, 9, 6, 0, 3, 0, 
    0, 0, 8, 12, 8, 3, 0, 0, 6, 23, 5, 40, 43, 14, 21, 
    26, 15, 24, 29, 32, 30, 21, 10, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    77, 74, 93, 98, 105, 105, 109, 108, 107, 113, 114, 115, 110, 112, 114, 
    80, 78, 98, 99, 106, 104, 109, 114, 108, 101, 113, 117, 112, 115, 116, 
    83, 78, 97, 99, 100, 102, 98, 102, 108, 87, 86, 120, 112, 113, 115, 
    90, 78, 97, 113, 105, 103, 94, 78, 77, 74, 49, 65, 116, 106, 110, 
    78, 69, 72, 80, 91, 93, 93, 77, 54, 35, 40, 32, 40, 64, 65, 
    24, 22, 28, 33, 36, 30, 46, 43, 35, 31, 33, 50, 33, 74, 27, 
    28, 34, 34, 41, 55, 55, 45, 39, 27, 31, 49, 82, 82, 41, 52, 
    34, 34, 39, 41, 60, 65, 67, 64, 76, 61, 75, 81, 77, 50, 15, 
    50, 64, 68, 80, 75, 79, 73, 65, 56, 53, 42, 61, 70, 61, 65, 
    39, 36, 53, 63, 67, 53, 55, 60, 75, 71, 69, 68, 65, 57, 48, 
    62, 53, 55, 59, 62, 78, 57, 44, 36, 61, 67, 56, 35, 23, 16, 
    44, 57, 48, 37, 32, 39, 57, 40, 33, 35, 26, 25, 10, 7, 3, 
    36, 51, 50, 37, 36, 38, 32, 18, 22, 25, 11, 6, 10, 0, 0, 
    15, 18, 11, 8, 9, 13, 15, 9, 10, 0, 8, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 14, 7, 0, 0, 0, 0, 0, 
    
    -- channel=87
    46, 35, 41, 38, 32, 25, 22, 21, 20, 18, 19, 15, 16, 19, 16, 
    35, 23, 28, 22, 21, 14, 11, 17, 16, 14, 0, 12, 11, 14, 9, 
    25, 14, 16, 11, 10, 7, 8, 8, 3, 17, 0, 14, 6, 7, 6, 
    12, 0, 0, 0, 0, 0, 6, 1, 6, 1, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 15, 24, 25, 2, 9, 0, 0, 
    15, 13, 19, 13, 19, 15, 26, 29, 24, 21, 19, 23, 0, 6, 4, 
    28, 12, 14, 20, 23, 31, 38, 39, 34, 31, 14, 3, 4, 0, 0, 
    37, 31, 38, 45, 44, 43, 42, 35, 32, 19, 1, 0, 0, 6, 0, 
    30, 35, 22, 37, 39, 39, 34, 28, 20, 22, 13, 6, 7, 0, 4, 
    33, 33, 47, 37, 32, 34, 30, 21, 20, 18, 13, 7, 7, 0, 0, 
    39, 42, 34, 32, 26, 27, 27, 12, 0, 13, 11, 3, 1, 2, 1, 
    33, 33, 34, 22, 23, 19, 23, 18, 12, 6, 7, 12, 1, 2, 0, 
    22, 23, 23, 19, 16, 8, 6, 10, 10, 7, 1, 4, 4, 0, 1, 
    2, 0, 4, 5, 5, 6, 5, 4, 5, 12, 3, 0, 0, 1, 0, 
    0, 0, 0, 1, 3, 6, 6, 2, 0, 6, 2, 0, 0, 2, 0, 
    
    -- channel=88
    135, 129, 159, 157, 165, 161, 169, 167, 169, 173, 161, 175, 169, 175, 170, 
    137, 130, 158, 155, 166, 156, 161, 166, 165, 146, 140, 172, 166, 172, 170, 
    136, 121, 154, 155, 163, 153, 151, 133, 146, 114, 128, 150, 157, 161, 165, 
    118, 111, 128, 134, 138, 144, 135, 131, 85, 66, 74, 65, 111, 129, 125, 
    62, 62, 69, 74, 78, 81, 88, 84, 75, 71, 68, 84, 89, 106, 79, 
    72, 73, 73, 73, 99, 89, 94, 77, 75, 81, 101, 139, 111, 114, 61, 
    73, 68, 59, 82, 101, 106, 109, 107, 115, 114, 128, 126, 111, 72, 40, 
    90, 98, 109, 118, 124, 129, 129, 119, 113, 92, 93, 113, 112, 83, 106, 
    84, 71, 98, 119, 114, 108, 112, 115, 116, 111, 117, 113, 110, 102, 86, 
    83, 103, 105, 101, 112, 121, 117, 98, 91, 115, 114, 102, 78, 59, 54, 
    98, 103, 101, 84, 81, 103, 98, 61, 81, 93, 76, 64, 54, 43, 36, 
    90, 95, 86, 66, 77, 95, 70, 61, 66, 67, 53, 47, 42, 32, 21, 
    66, 63, 52, 50, 51, 53, 55, 55, 45, 44, 43, 38, 26, 24, 23, 
    27, 27, 32, 36, 37, 36, 39, 40, 52, 40, 30, 26, 23, 26, 26, 
    21, 24, 30, 33, 37, 38, 36, 28, 43, 29, 24, 21, 22, 26, 8, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 10, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 11, 25, 5, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 5, 4, 6, 8, 
    7, 8, 5, 5, 4, 4, 2, 3, 0, 1, 5, 6, 5, 4, 12, 
    
    -- channel=91
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=92
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 83, 0, 0, 1, 0, 0, 
    17, 0, 0, 0, 0, 0, 7, 8, 18, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 13, 5, 0, 0, 0, 1, 0, 
    0, 0, 12, 0, 0, 0, 0, 12, 0, 0, 0, 0, 46, 0, 48, 
    0, 0, 4, 0, 0, 3, 0, 7, 0, 0, 0, 0, 45, 0, 71, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 82, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 29, 0, 0, 0, 7, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 20, 0, 
    0, 0, 0, 7, 0, 0, 26, 26, 0, 0, 3, 15, 15, 10, 8, 
    0, 0, 25, 6, 0, 0, 24, 13, 0, 0, 9, 8, 9, 5, 16, 
    0, 0, 11, 0, 0, 0, 2, 0, 0, 0, 9, 0, 21, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 18, 2, 3, 5, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 8, 0, 46, 0, 3, 0, 0, 28, 
    
    -- channel=93
    1, 3, 13, 13, 18, 21, 26, 27, 28, 28, 31, 32, 27, 30, 29, 
    10, 10, 23, 20, 28, 25, 30, 34, 29, 23, 38, 35, 29, 33, 32, 
    16, 15, 29, 27, 33, 29, 30, 35, 35, 21, 25, 37, 33, 39, 35, 
    23, 18, 31, 41, 42, 37, 35, 17, 19, 28, 16, 29, 50, 40, 45, 
    27, 18, 28, 31, 38, 37, 33, 23, 5, 0, 0, 2, 10, 28, 24, 
    1, 0, 0, 6, 0, 0, 0, 0, 0, 0, 2, 6, 0, 38, 1, 
    0, 0, 3, 1, 8, 0, 0, 0, 0, 0, 5, 28, 28, 15, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 29, 30, 24, 7, 5, 
    0, 5, 10, 5, 0, 6, 11, 11, 7, 6, 4, 14, 18, 12, 27, 
    0, 0, 0, 1, 8, 0, 1, 5, 16, 17, 13, 13, 15, 18, 18, 
    1, 0, 0, 0, 7, 17, 4, 9, 8, 12, 15, 18, 7, 6, 0, 
    3, 1, 0, 0, 0, 1, 6, 0, 4, 9, 2, 7, 0, 0, 0, 
    0, 2, 6, 0, 6, 11, 4, 0, 0, 8, 1, 0, 0, 0, 0, 
    3, 5, 1, 0, 0, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    72, 44, 64, 72, 78, 76, 79, 88, 74, 85, 84, 83, 84, 84, 78, 
    76, 47, 65, 78, 80, 78, 82, 85, 75, 91, 67, 77, 87, 88, 79, 
    78, 46, 63, 79, 78, 78, 85, 71, 75, 106, 34, 74, 92, 87, 77, 
    76, 47, 63, 73, 78, 73, 80, 68, 57, 74, 20, 41, 61, 77, 69, 
    56, 37, 52, 44, 60, 57, 60, 70, 52, 33, 23, 29, 10, 62, 38, 
    11, 11, 30, 14, 19, 22, 29, 43, 28, 32, 13, 25, 47, 45, 37, 
    13, 24, 32, 6, 33, 41, 35, 31, 23, 29, 20, 54, 80, 35, 65, 
    22, 25, 19, 16, 35, 46, 55, 57, 58, 64, 42, 49, 57, 54, 20, 
    39, 39, 40, 51, 58, 61, 61, 59, 44, 57, 18, 41, 52, 54, 50, 
    37, 16, 27, 46, 54, 45, 47, 53, 48, 54, 49, 60, 54, 56, 36, 
    38, 40, 46, 51, 42, 50, 60, 46, 17, 44, 55, 58, 39, 29, 16, 
    15, 44, 51, 33, 22, 19, 60, 34, 21, 36, 33, 26, 20, 9, 12, 
    18, 41, 51, 29, 28, 35, 32, 21, 22, 25, 22, 7, 19, 4, 0, 
    14, 19, 16, 11, 12, 13, 15, 18, 7, 11, 11, 4, 5, 0, 2, 
    2, 0, 0, 0, 3, 2, 5, 12, 0, 29, 0, 2, 0, 0, 5, 
    
    -- channel=95
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 16, 5, 0, 0, 2, 
    0, 3, 9, 0, 4, 0, 0, 8, 11, 0, 34, 14, 0, 4, 7, 
    0, 10, 13, 13, 7, 8, 0, 0, 0, 0, 14, 23, 35, 14, 22, 
    11, 13, 14, 26, 20, 21, 11, 0, 0, 0, 0, 4, 23, 7, 21, 
    8, 6, 0, 8, 0, 0, 0, 0, 0, 0, 13, 5, 0, 18, 0, 
    2, 0, 0, 11, 1, 0, 0, 0, 0, 0, 16, 12, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 15, 3, 0, 1, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 11, 5, 1, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 2, 3, 0, 0, 19, 7, 1, 0, 0, 4, 7, 
    14, 0, 0, 0, 0, 14, 0, 0, 8, 2, 0, 5, 1, 7, 5, 
    12, 0, 0, 0, 6, 6, 1, 4, 6, 7, 2, 11, 0, 8, 8, 
    10, 9, 8, 11, 10, 11, 10, 6, 11, 0, 8, 7, 7, 11, 11, 
    12, 14, 12, 12, 9, 8, 9, 8, 27, 0, 11, 8, 11, 13, 4, 
    
    -- channel=96
    37, 30, 17, 32, 37, 34, 33, 35, 34, 35, 35, 34, 41, 40, 39, 
    31, 28, 29, 42, 65, 63, 54, 62, 61, 60, 55, 60, 49, 40, 40, 
    32, 24, 29, 49, 53, 57, 58, 65, 55, 53, 58, 58, 51, 36, 41, 
    29, 27, 26, 66, 53, 51, 50, 61, 55, 52, 59, 57, 59, 36, 35, 
    28, 27, 25, 17, 26, 24, 27, 30, 25, 24, 31, 42, 38, 33, 33, 
    35, 19, 16, 40, 29, 32, 35, 34, 31, 31, 34, 33, 35, 36, 37, 
    41, 22, 8, 11, 40, 43, 38, 37, 37, 33, 35, 33, 33, 33, 35, 
    44, 35, 35, 19, 0, 32, 50, 43, 36, 35, 36, 34, 34, 33, 32, 
    46, 42, 39, 38, 0, 20, 23, 26, 37, 39, 44, 36, 33, 33, 34, 
    50, 43, 42, 24, 0, 8, 21, 24, 18, 4, 16, 23, 38, 43, 39, 
    49, 41, 40, 31, 41, 7, 26, 60, 37, 21, 36, 23, 56, 43, 38, 
    26, 18, 15, 14, 14, 8, 14, 26, 13, 13, 16, 17, 16, 15, 17, 
    18, 18, 12, 11, 10, 11, 12, 13, 6, 8, 7, 8, 9, 7, 7, 
    9, 14, 11, 14, 11, 12, 12, 14, 12, 9, 11, 10, 9, 9, 23, 
    7, 10, 10, 11, 12, 20, 14, 19, 15, 14, 10, 10, 18, 12, 0, 
    
    -- channel=97
    43, 47, 40, 34, 34, 37, 38, 39, 38, 38, 39, 40, 44, 51, 51, 
    42, 46, 48, 9, 9, 10, 10, 6, 11, 15, 13, 16, 42, 47, 47, 
    40, 45, 47, 12, 25, 23, 15, 20, 28, 33, 31, 28, 37, 49, 47, 
    41, 44, 37, 0, 15, 14, 17, 8, 7, 7, 10, 16, 20, 45, 46, 
    44, 43, 49, 41, 30, 29, 31, 33, 34, 34, 32, 44, 42, 49, 46, 
    51, 52, 40, 43, 54, 50, 51, 51, 50, 53, 53, 44, 46, 46, 48, 
    51, 38, 24, 18, 19, 34, 44, 47, 48, 48, 46, 47, 46, 45, 44, 
    53, 51, 67, 48, 20, 14, 27, 41, 45, 45, 46, 46, 47, 47, 46, 
    54, 53, 53, 59, 30, 6, 0, 11, 22, 30, 36, 45, 46, 46, 45, 
    52, 51, 51, 51, 16, 2, 5, 7, 1, 0, 0, 11, 24, 35, 42, 
    50, 46, 50, 47, 49, 32, 15, 38, 51, 40, 33, 28, 40, 40, 41, 
    34, 26, 25, 22, 19, 31, 30, 17, 22, 22, 27, 29, 22, 18, 21, 
    22, 19, 23, 24, 23, 21, 19, 14, 11, 9, 7, 5, 5, 2, 0, 
    0, 0, 0, 0, 3, 1, 1, 3, 9, 7, 7, 8, 6, 8, 30, 
    7, 6, 7, 8, 8, 8, 11, 12, 14, 14, 14, 14, 14, 45, 29, 
    
    -- channel=98
    0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 1, 2, 0, 12, 9, 4, 0, 0, 0, 0, 
    0, 0, 5, 16, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 12, 6, 6, 10, 7, 4, 0, 0, 0, 0, 
    0, 29, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 107, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 105, 139, 69, 41, 91, 97, 94, 84, 10, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    1, 0, 0, 0, 0, 7, 12, 8, 14, 15, 5, 0, 8, 9, 0, 
    
    -- channel=99
    49, 51, 24, 36, 45, 41, 36, 36, 33, 37, 37, 36, 38, 43, 42, 
    51, 53, 41, 34, 55, 64, 56, 60, 61, 61, 61, 58, 55, 49, 46, 
    51, 48, 52, 33, 41, 36, 37, 42, 40, 40, 38, 40, 67, 47, 47, 
    45, 49, 47, 20, 34, 35, 25, 42, 36, 37, 43, 45, 40, 48, 48, 
    41, 48, 41, 39, 43, 43, 40, 44, 44, 40, 44, 51, 45, 47, 47, 
    46, 41, 49, 51, 30, 31, 36, 36, 32, 33, 36, 44, 48, 46, 45, 
    50, 25, 3, 52, 83, 65, 50, 48, 45, 42, 47, 46, 48, 50, 50, 
    56, 46, 24, 0, 0, 77, 86, 57, 46, 45, 45, 44, 45, 44, 46, 
    58, 49, 46, 38, 0, 24, 50, 75, 80, 68, 60, 45, 45, 46, 46, 
    59, 49, 47, 39, 0, 16, 20, 16, 25, 41, 72, 82, 81, 67, 52, 
    60, 50, 48, 36, 0, 0, 0, 6, 0, 0, 0, 0, 25, 34, 46, 
    73, 71, 70, 71, 75, 51, 51, 73, 64, 47, 59, 48, 62, 63, 62, 
    18, 24, 17, 18, 17, 15, 21, 36, 35, 39, 42, 46, 48, 49, 47, 
    10, 28, 23, 18, 12, 12, 13, 13, 7, 3, 4, 4, 5, 3, 0, 
    0, 4, 4, 4, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 22, 
    
    -- channel=100
    19, 30, 35, 23, 26, 28, 27, 27, 26, 27, 26, 27, 23, 18, 19, 
    26, 33, 31, 15, 6, 1, 5, 1, 2, 3, 6, 6, 21, 23, 23, 
    26, 33, 26, 7, 4, 3, 0, 1, 5, 4, 5, 6, 12, 24, 22, 
    27, 34, 24, 20, 16, 20, 16, 16, 22, 19, 15, 14, 25, 25, 28, 
    26, 32, 31, 31, 31, 31, 32, 28, 30, 29, 27, 24, 27, 26, 30, 
    21, 28, 27, 24, 27, 24, 23, 24, 25, 23, 22, 24, 29, 29, 29, 
    19, 36, 39, 34, 21, 22, 28, 29, 27, 26, 25, 26, 27, 27, 29, 
    18, 25, 21, 12, 26, 19, 12, 21, 28, 28, 26, 26, 27, 28, 31, 
    14, 18, 21, 21, 33, 12, 17, 24, 12, 13, 22, 28, 29, 28, 30, 
    12, 19, 22, 22, 38, 20, 11, 7, 15, 35, 36, 22, 9, 13, 25, 
    13, 23, 22, 27, 23, 20, 27, 13, 7, 23, 11, 25, 12, 18, 28, 
    11, 22, 21, 21, 22, 24, 11, 16, 38, 33, 30, 32, 34, 46, 44, 
    14, 21, 20, 13, 8, 10, 11, 15, 20, 19, 19, 20, 20, 21, 24, 
    22, 25, 23, 19, 17, 19, 18, 15, 13, 12, 11, 9, 11, 12, 12, 
    10, 11, 13, 11, 10, 9, 11, 7, 9, 9, 8, 6, 8, 8, 9, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 1, 6, 17, 20, 14, 5, 0, 0, 0, 
    0, 0, 0, 8, 0, 1, 9, 3, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 28, 27, 23, 25, 22, 21, 4, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 86, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 106, 128, 76, 103, 118, 101, 119, 88, 76, 29, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 
    0, 0, 0, 0, 0, 9, 11, 11, 11, 14, 5, 0, 18, 51, 0, 
    
    -- channel=103
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 7, 0, 0, 
    5, 0, 0, 0, 1, 0, 0, 0, 0, 0, 6, 3, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    4, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 25, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 17, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 5, 10, 0, 4, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 7, 1, 0, 0, 5, 2, 11, 5, 0, 
    13, 0, 0, 0, 1, 0, 7, 48, 0, 0, 4, 0, 35, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 25, 
    0, 0, 0, 0, 0, 7, 0, 3, 0, 0, 0, 0, 22, 0, 0, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 36, 35, 28, 30, 33, 33, 23, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 70, 83, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 81, 57, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 51, 107, 93, 42, 6, 0, 0, 0, 0, 
    0, 0, 0, 5, 13, 24, 12, 0, 13, 62, 117, 127, 88, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    84, 92, 101, 107, 112, 88, 60, 64, 74, 49, 50, 37, 42, 56, 56, 
    0, 0, 0, 0, 0, 0, 3, 22, 35, 43, 47, 54, 58, 59, 64, 
    27, 33, 30, 22, 18, 17, 14, 11, 6, 3, 2, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 1, 1, 2, 4, 4, 4, 4, 3, 2, 0, 
    0, 0, 2, 4, 3, 1, 3, 3, 3, 3, 5, 7, 1, 8, 10, 
    
    -- channel=108
    137, 168, 173, 149, 147, 163, 163, 158, 163, 163, 164, 163, 165, 176, 184, 
    142, 169, 179, 153, 116, 124, 130, 126, 133, 131, 137, 140, 167, 181, 187, 
    140, 169, 168, 129, 123, 111, 117, 110, 125, 129, 127, 132, 159, 185, 188, 
    145, 167, 160, 125, 127, 136, 130, 126, 135, 136, 127, 133, 143, 180, 183, 
    160, 165, 170, 162, 140, 139, 143, 144, 147, 147, 143, 149, 176, 180, 184, 
    170, 171, 154, 164, 175, 171, 172, 177, 177, 174, 173, 174, 179, 182, 185, 
    172, 187, 149, 90, 104, 161, 180, 186, 187, 185, 179, 181, 180, 180, 181, 
    173, 192, 193, 176, 94, 69, 127, 180, 186, 182, 179, 181, 181, 181, 181, 
    174, 193, 195, 195, 158, 46, 53, 73, 108, 145, 165, 184, 182, 180, 181, 
    173, 190, 193, 187, 142, 25, 34, 49, 55, 54, 41, 77, 112, 151, 176, 
    167, 187, 189, 194, 162, 139, 77, 87, 147, 132, 108, 108, 99, 154, 166, 
    115, 128, 123, 117, 112, 117, 100, 104, 127, 120, 123, 125, 128, 127, 131, 
    86, 87, 86, 80, 74, 73, 67, 67, 73, 64, 63, 60, 62, 62, 58, 
    54, 43, 43, 41, 43, 37, 35, 36, 39, 36, 32, 32, 32, 34, 58, 
    47, 34, 34, 33, 35, 38, 43, 42, 49, 45, 40, 36, 42, 70, 79, 
    
    -- channel=109
    56, 65, 57, 40, 46, 48, 45, 46, 45, 46, 45, 45, 47, 48, 51, 
    64, 72, 59, 0, 0, 0, 0, 0, 0, 0, 2, 10, 44, 51, 51, 
    61, 72, 59, 1, 5, 3, 0, 0, 12, 11, 10, 13, 40, 54, 54, 
    60, 70, 44, 0, 6, 11, 8, 2, 6, 0, 0, 8, 21, 53, 59, 
    60, 70, 66, 56, 50, 51, 51, 50, 51, 49, 46, 55, 52, 60, 61, 
    56, 63, 62, 57, 59, 57, 57, 56, 55, 57, 55, 59, 60, 57, 59, 
    54, 57, 38, 41, 45, 55, 58, 58, 57, 56, 56, 57, 58, 57, 58, 
    56, 62, 48, 22, 30, 40, 46, 52, 54, 52, 53, 55, 57, 58, 62, 
    53, 54, 52, 46, 17, 11, 22, 32, 36, 43, 52, 55, 57, 58, 60, 
    48, 48, 50, 44, 14, 9, 5, 3, 13, 25, 36, 33, 38, 47, 55, 
    50, 51, 53, 42, 21, 18, 21, 21, 22, 22, 19, 22, 32, 43, 51, 
    45, 43, 42, 42, 44, 38, 39, 47, 53, 49, 54, 51, 59, 61, 57, 
    29, 30, 31, 28, 26, 25, 28, 34, 33, 33, 33, 35, 36, 33, 31, 
    11, 11, 11, 8, 4, 7, 7, 6, 5, 4, 5, 5, 6, 10, 25, 
    3, 7, 6, 5, 3, 5, 4, 3, 4, 3, 3, 1, 14, 31, 29, 
    
    -- channel=110
    10, 4, 0, 0, 1, 0, 0, 2, 0, 1, 1, 1, 9, 8, 10, 
    6, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 10, 10, 
    5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 12, 
    2, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 9, 
    1, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 13, 3, 7, 7, 
    8, 1, 0, 9, 1, 2, 4, 4, 1, 2, 5, 2, 6, 7, 9, 
    13, 0, 0, 0, 10, 8, 7, 7, 7, 4, 6, 6, 6, 6, 8, 
    16, 10, 12, 0, 0, 2, 14, 10, 6, 6, 7, 6, 6, 5, 6, 
    17, 14, 11, 12, 0, 0, 0, 0, 8, 6, 10, 5, 5, 5, 7, 
    18, 13, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 10, 9, 8, 
    19, 9, 11, 0, 0, 0, 0, 5, 0, 0, 0, 0, 5, 0, 5, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=111
    31, 34, 29, 27, 27, 24, 24, 22, 21, 23, 24, 24, 20, 23, 25, 
    38, 47, 36, 8, 16, 25, 22, 22, 22, 23, 24, 20, 27, 30, 29, 
    39, 46, 45, 2, 0, 0, 0, 0, 0, 0, 0, 0, 25, 32, 31, 
    38, 44, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 35, 37, 
    35, 44, 38, 33, 32, 35, 33, 31, 35, 30, 28, 29, 24, 37, 37, 
    32, 49, 53, 27, 24, 23, 22, 22, 22, 24, 23, 31, 36, 32, 34, 
    30, 23, 27, 69, 58, 35, 34, 34, 32, 34, 35, 36, 37, 38, 38, 
    32, 35, 15, 0, 33, 61, 44, 31, 34, 32, 31, 33, 34, 34, 37, 
    32, 32, 31, 20, 14, 17, 43, 69, 56, 42, 32, 32, 35, 37, 38, 
    28, 30, 30, 42, 23, 23, 13, 6, 20, 51, 76, 74, 54, 37, 33, 
    30, 29, 32, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 32, 
    60, 64, 66, 68, 69, 56, 46, 50, 60, 50, 51, 44, 51, 60, 57, 
    22, 22, 23, 21, 22, 22, 25, 36, 42, 46, 48, 52, 54, 54, 54, 
    27, 30, 30, 23, 20, 20, 19, 18, 15, 12, 12, 12, 12, 6, 0, 
    7, 10, 10, 9, 7, 2, 4, 1, 2, 2, 7, 7, 0, 16, 40, 
    
    -- channel=112
    163, 185, 170, 156, 168, 170, 167, 164, 166, 167, 170, 170, 175, 191, 198, 
    166, 193, 188, 144, 150, 177, 174, 172, 178, 182, 178, 177, 201, 203, 205, 
    164, 187, 193, 158, 140, 127, 126, 134, 140, 142, 147, 162, 194, 204, 206, 
    162, 182, 172, 122, 134, 137, 131, 132, 144, 138, 135, 140, 159, 198, 204, 
    170, 182, 185, 171, 158, 159, 159, 164, 168, 162, 158, 176, 188, 199, 201, 
    181, 187, 189, 182, 175, 174, 179, 183, 179, 177, 179, 190, 197, 195, 199, 
    187, 165, 124, 136, 179, 198, 199, 202, 201, 198, 198, 199, 199, 201, 203, 
    194, 203, 182, 118, 88, 144, 196, 206, 202, 196, 194, 195, 196, 195, 197, 
    197, 209, 210, 193, 100, 57, 96, 148, 185, 197, 197, 198, 198, 198, 199, 
    195, 205, 209, 205, 100, 34, 44, 53, 66, 80, 118, 164, 188, 198, 199, 
    193, 204, 208, 174, 101, 52, 28, 63, 94, 60, 54, 48, 95, 155, 181, 
    180, 193, 190, 187, 187, 163, 150, 168, 175, 162, 165, 161, 167, 172, 174, 
    94, 97, 94, 89, 88, 84, 84, 99, 103, 102, 103, 106, 112, 111, 105, 
    57, 57, 54, 49, 42, 36, 36, 37, 36, 29, 26, 28, 27, 25, 38, 
    34, 30, 27, 27, 25, 25, 27, 29, 29, 26, 25, 25, 27, 54, 76, 
    
    -- channel=113
    62, 75, 61, 55, 63, 66, 64, 64, 64, 65, 65, 63, 68, 73, 73, 
    63, 73, 69, 44, 37, 34, 31, 38, 35, 36, 41, 50, 70, 71, 74, 
    60, 71, 58, 52, 47, 53, 44, 54, 61, 59, 53, 58, 67, 73, 75, 
    61, 71, 61, 55, 56, 54, 55, 57, 56, 52, 55, 57, 66, 69, 74, 
    66, 72, 71, 61, 55, 54, 55, 59, 57, 53, 54, 67, 74, 73, 74, 
    67, 62, 49, 71, 76, 76, 78, 78, 76, 73, 73, 76, 73, 74, 77, 
    70, 71, 48, 11, 34, 67, 77, 78, 77, 73, 72, 71, 71, 70, 72, 
    72, 77, 72, 65, 16, 15, 50, 72, 72, 71, 71, 72, 73, 73, 75, 
    70, 76, 74, 69, 19, 4, 1, 3, 24, 48, 68, 76, 73, 71, 74, 
    68, 72, 74, 56, 0, 0, 0, 5, 3, 0, 0, 0, 25, 54, 73, 
    69, 73, 73, 69, 74, 57, 43, 62, 72, 46, 63, 47, 67, 70, 69, 
    24, 22, 16, 13, 12, 9, 18, 32, 30, 37, 35, 42, 44, 43, 42, 
    24, 29, 24, 19, 15, 13, 15, 15, 11, 7, 6, 5, 5, 4, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 0, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 63, 9, 0, 0, 0, 33, 29, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 
    24, 26, 26, 23, 20, 20, 14, 11, 9, 9, 5, 1, 4, 12, 0, 
    4, 2, 3, 0, 5, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    
    -- channel=115
    11, 7, 13, 11, 16, 12, 14, 15, 16, 16, 15, 16, 17, 13, 14, 
    6, 6, 5, 0, 0, 2, 4, 2, 3, 5, 5, 7, 13, 9, 11, 
    6, 5, 0, 16, 10, 10, 9, 16, 17, 9, 16, 16, 9, 7, 8, 
    6, 5, 0, 2, 0, 0, 6, 0, 0, 0, 0, 0, 4, 5, 9, 
    6, 4, 8, 4, 8, 9, 11, 9, 6, 10, 9, 11, 7, 9, 8, 
    8, 0, 1, 14, 10, 10, 9, 7, 7, 9, 10, 6, 9, 10, 10, 
    11, 18, 14, 0, 0, 10, 7, 6, 7, 6, 6, 6, 6, 6, 7, 
    10, 9, 15, 26, 0, 0, 5, 10, 7, 7, 7, 7, 7, 8, 7, 
    10, 10, 11, 12, 10, 7, 3, 0, 0, 3, 11, 9, 7, 7, 7, 
    10, 10, 11, 0, 12, 5, 8, 12, 12, 1, 0, 0, 0, 9, 9, 
    9, 10, 10, 17, 30, 27, 24, 24, 24, 26, 28, 27, 15, 12, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 5, 3, 4, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 4, 5, 11, 11, 10, 8, 9, 10, 11, 11, 11, 13, 18, 26, 
    15, 12, 12, 13, 15, 17, 15, 19, 19, 18, 15, 14, 23, 14, 10, 
    
    -- channel=116
    57, 80, 89, 70, 70, 74, 73, 71, 74, 73, 74, 75, 76, 85, 88, 
    59, 85, 90, 82, 60, 73, 73, 70, 77, 76, 75, 73, 85, 91, 92, 
    61, 80, 93, 92, 71, 67, 71, 70, 76, 76, 81, 89, 74, 91, 92, 
    65, 78, 79, 77, 59, 66, 71, 62, 69, 65, 52, 56, 71, 85, 91, 
    69, 77, 87, 87, 72, 72, 71, 76, 78, 75, 69, 73, 91, 89, 91, 
    68, 89, 89, 71, 85, 83, 85, 88, 87, 84, 84, 87, 89, 89, 89, 
    68, 76, 64, 61, 58, 77, 89, 92, 92, 93, 90, 92, 90, 91, 92, 
    69, 89, 84, 65, 61, 47, 63, 86, 94, 90, 88, 88, 89, 89, 90, 
    70, 88, 93, 86, 88, 13, 28, 50, 64, 77, 81, 91, 91, 89, 90, 
    68, 89, 93, 103, 74, 10, 8, 12, 19, 26, 38, 58, 65, 75, 87, 
    65, 91, 90, 73, 53, 42, 6, 15, 42, 44, 17, 25, 24, 68, 79, 
    65, 90, 85, 82, 81, 76, 69, 71, 84, 82, 80, 81, 83, 86, 87, 
    34, 44, 46, 39, 35, 34, 36, 41, 43, 40, 39, 38, 41, 40, 37, 
    18, 15, 13, 10, 8, 5, 6, 4, 5, 2, 0, 1, 1, 0, 0, 
    10, 5, 3, 3, 1, 0, 4, 0, 2, 2, 4, 0, 0, 15, 22, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 38, 35, 33, 34, 33, 31, 28, 21, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 6, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 7, 5, 0, 8, 9, 12, 13, 7, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 35, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 36, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 50, 37, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 3, 0, 0, 29, 56, 54, 31, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 27, 31, 33, 36, 27, 5, 8, 22, 8, 6, 1, 1, 15, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 11, 13, 17, 20, 21, 22, 
    10, 17, 16, 10, 6, 5, 4, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=118
    79, 93, 78, 79, 85, 89, 85, 84, 82, 84, 86, 85, 87, 92, 97, 
    78, 91, 91, 90, 101, 113, 109, 114, 114, 114, 114, 111, 105, 104, 103, 
    77, 87, 95, 114, 96, 94, 95, 102, 101, 96, 96, 98, 107, 98, 105, 
    73, 87, 88, 100, 95, 91, 92, 97, 99, 101, 99, 103, 95, 99, 102, 
    77, 86, 89, 86, 86, 86, 84, 87, 89, 87, 85, 93, 98, 95, 98, 
    85, 81, 92, 99, 74, 79, 82, 87, 84, 79, 80, 88, 98, 97, 96, 
    90, 82, 48, 65, 118, 111, 101, 101, 99, 96, 97, 98, 98, 100, 103, 
    93, 99, 85, 42, 17, 84, 122, 110, 102, 100, 97, 97, 96, 95, 96, 
    94, 103, 101, 96, 35, 27, 49, 92, 119, 114, 109, 99, 97, 97, 98, 
    96, 103, 104, 95, 60, 17, 27, 30, 31, 48, 80, 108, 119, 113, 103, 
    98, 104, 103, 96, 46, 0, 1, 22, 25, 3, 8, 0, 33, 65, 90, 
    100, 111, 110, 111, 113, 101, 80, 95, 105, 98, 90, 93, 91, 103, 103, 
    44, 51, 43, 40, 36, 36, 37, 47, 57, 56, 59, 61, 66, 68, 65, 
    31, 39, 36, 29, 22, 20, 20, 19, 15, 9, 8, 9, 8, 8, 0, 
    13, 11, 10, 7, 8, 9, 4, 5, 3, 0, 0, 0, 5, 0, 6, 
    
    -- channel=119
    16, 32, 24, 13, 13, 17, 14, 13, 13, 13, 13, 12, 12, 17, 18, 
    23, 33, 32, 3, 0, 0, 0, 0, 0, 0, 0, 0, 15, 20, 18, 
    22, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 21, 20, 
    23, 33, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 23, 
    24, 32, 31, 27, 16, 17, 15, 15, 16, 16, 13, 17, 23, 27, 26, 
    25, 28, 28, 29, 32, 30, 30, 30, 29, 30, 28, 28, 27, 25, 25, 
    20, 30, 8, 0, 7, 27, 26, 27, 26, 26, 25, 25, 26, 24, 23, 
    20, 28, 26, 22, 0, 0, 16, 22, 21, 22, 22, 24, 26, 26, 27, 
    18, 22, 22, 23, 4, 0, 0, 0, 1, 15, 23, 24, 25, 25, 26, 
    15, 18, 19, 9, 4, 0, 0, 0, 0, 0, 0, 0, 5, 20, 24, 
    14, 20, 20, 30, 9, 17, 3, 0, 20, 8, 14, 6, 4, 17, 16, 
    6, 9, 4, 2, 2, 5, 13, 15, 12, 13, 19, 19, 25, 19, 17, 
    1, 7, 7, 7, 4, 4, 8, 9, 8, 6, 7, 5, 6, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    
    -- channel=120
    130, 136, 126, 122, 126, 132, 133, 131, 133, 133, 135, 132, 139, 147, 148, 
    130, 141, 140, 87, 98, 95, 92, 98, 99, 103, 100, 104, 144, 144, 146, 
    128, 138, 137, 84, 98, 101, 91, 99, 108, 113, 116, 119, 133, 146, 148, 
    129, 137, 119, 87, 94, 97, 96, 98, 98, 93, 94, 109, 117, 142, 144, 
    136, 137, 135, 119, 115, 114, 118, 120, 117, 113, 117, 132, 139, 145, 144, 
    145, 132, 112, 139, 140, 139, 140, 140, 137, 138, 140, 141, 144, 146, 150, 
    149, 135, 113, 72, 97, 133, 145, 147, 146, 143, 141, 141, 141, 141, 142, 
    154, 153, 147, 127, 62, 78, 118, 144, 144, 140, 141, 141, 143, 141, 143, 
    157, 156, 153, 145, 69, 54, 60, 72, 92, 116, 134, 143, 142, 142, 142, 
    156, 151, 152, 140, 45, 28, 43, 52, 55, 45, 49, 70, 96, 124, 140, 
    151, 147, 150, 136, 130, 99, 84, 116, 129, 93, 112, 94, 129, 134, 136, 
    96, 88, 84, 81, 78, 71, 73, 87, 87, 90, 89, 93, 93, 93, 96, 
    75, 72, 69, 64, 64, 59, 56, 57, 54, 51, 49, 49, 50, 48, 43, 
    44, 42, 42, 43, 41, 39, 39, 41, 42, 37, 37, 38, 37, 40, 79, 
    38, 38, 39, 41, 39, 49, 48, 52, 52, 50, 44, 40, 52, 90, 60, 
    
    -- channel=121
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 6, 0, 3, 1, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 12, 19, 17, 19, 15, 15, 19, 15, 0, 0, 0, 
    0, 0, 0, 20, 5, 0, 8, 5, 3, 3, 3, 4, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 19, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 7, 8, 12, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 38, 20, 15, 26, 20, 27, 23, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 5, 8, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 5, 8, 5, 6, 8, 11, 12, 12, 14, 13, 12, 15, 
    14, 15, 13, 15, 15, 15, 19, 19, 18, 20, 19, 18, 12, 17, 0, 
    
    -- channel=123
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=124
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 32, 12, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 5, 0, 0, 3, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 29, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 78, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 151, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 42, 72, 0, 0, 14, 31, 3, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 2, 0, 1, 0, 3, 0, 2, 0, 0, 0, 8, 
    
    -- channel=125
    17, 13, 7, 17, 17, 18, 18, 18, 17, 19, 18, 19, 20, 18, 19, 
    17, 11, 11, 19, 43, 44, 43, 42, 41, 42, 40, 34, 26, 22, 23, 
    17, 10, 14, 16, 19, 19, 21, 22, 14, 15, 19, 16, 30, 18, 21, 
    14, 12, 7, 21, 26, 24, 15, 25, 27, 27, 34, 31, 30, 22, 18, 
    13, 10, 8, 6, 15, 13, 16, 13, 16, 15, 18, 18, 16, 15, 17, 
    20, 8, 13, 19, 4, 4, 6, 7, 6, 7, 8, 9, 16, 17, 17, 
    24, 12, 3, 23, 37, 24, 17, 16, 16, 14, 16, 16, 17, 18, 19, 
    26, 17, 15, 0, 0, 31, 36, 25, 18, 18, 18, 17, 15, 15, 15, 
    28, 22, 21, 24, 0, 12, 25, 39, 39, 29, 25, 17, 17, 17, 16, 
    30, 24, 23, 18, 10, 10, 15, 14, 16, 25, 35, 40, 38, 29, 19, 
    29, 22, 23, 23, 2, 0, 0, 7, 0, 0, 0, 0, 6, 10, 19, 
    31, 27, 31, 31, 32, 27, 13, 18, 25, 12, 15, 11, 12, 17, 20, 
    9, 6, 3, 4, 4, 3, 1, 6, 9, 10, 11, 13, 14, 14, 16, 
    18, 19, 19, 18, 17, 15, 13, 14, 13, 11, 10, 10, 9, 9, 9, 
    9, 8, 9, 9, 10, 9, 6, 9, 9, 7, 6, 8, 10, 0, 10, 
    
    -- channel=126
    41, 57, 62, 54, 45, 56, 58, 54, 54, 54, 56, 56, 53, 57, 65, 
    44, 58, 67, 56, 52, 61, 65, 61, 64, 64, 64, 56, 60, 69, 67, 
    44, 60, 75, 62, 46, 36, 41, 34, 40, 44, 46, 45, 54, 66, 70, 
    43, 58, 58, 38, 41, 42, 43, 37, 42, 51, 42, 47, 38, 67, 67, 
    54, 58, 65, 63, 53, 53, 55, 54, 56, 61, 53, 50, 59, 65, 66, 
    62, 66, 67, 68, 52, 52, 51, 56, 57, 54, 53, 52, 67, 67, 66, 
    61, 69, 53, 46, 65, 66, 66, 68, 69, 69, 66, 68, 67, 68, 67, 
    60, 72, 77, 53, 14, 39, 63, 72, 70, 70, 66, 68, 66, 65, 64, 
    61, 74, 73, 79, 79, 11, 17, 57, 75, 73, 63, 66, 67, 68, 67, 
    61, 71, 73, 84, 100, 5, 12, 14, 11, 33, 43, 73, 75, 69, 66, 
    60, 70, 73, 80, 48, 11, 0, 0, 15, 17, 0, 0, 0, 30, 56, 
    63, 76, 79, 80, 78, 90, 53, 41, 68, 62, 52, 56, 44, 58, 59, 
    28, 32, 30, 29, 29, 29, 24, 26, 45, 43, 44, 45, 50, 52, 46, 
    30, 27, 31, 23, 22, 18, 16, 16, 19, 14, 11, 11, 8, 4, 10, 
    19, 10, 8, 6, 10, 7, 6, 5, 8, 6, 6, 8, 1, 14, 22, 
    
    -- channel=127
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 23, 12, 7, 13, 7, 10, 3, 6, 0, 0, 0, 
    5, 0, 0, 0, 0, 10, 7, 10, 0, 3, 8, 9, 4, 0, 0, 
    1, 0, 0, 7, 7, 5, 0, 13, 7, 1, 12, 9, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 20, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 2, 37, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 22, 37, 33, 20, 5, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 18, 23, 18, 22, 22, 37, 28, 21, 5, 0, 
    10, 0, 0, 0, 0, 0, 3, 21, 0, 0, 0, 0, 24, 6, 0, 
    20, 5, 8, 9, 12, 0, 6, 17, 0, 0, 1, 0, 0, 0, 0, 
    8, 0, 0, 2, 6, 4, 6, 12, 4, 9, 9, 12, 11, 9, 9, 
    14, 18, 15, 19, 17, 18, 18, 19, 17, 17, 20, 19, 18, 16, 26, 
    10, 17, 16, 19, 17, 19, 13, 19, 14, 14, 15, 17, 21, 23, 13, 
    
    -- channel=128
    10, 0, 9, 0, 0, 20, 2, 11, 7, 13, 0, 38, 0, 19, 11, 
    13, 2, 0, 1, 0, 8, 2, 16, 5, 10, 0, 47, 0, 22, 3, 
    0, 13, 5, 0, 0, 21, 11, 0, 16, 0, 24, 45, 11, 13, 11, 
    0, 36, 0, 3, 7, 21, 0, 0, 23, 9, 26, 31, 20, 19, 0, 
    0, 41, 0, 0, 33, 21, 0, 27, 14, 20, 13, 29, 21, 16, 0, 
    0, 37, 20, 0, 24, 36, 24, 40, 21, 28, 20, 40, 10, 17, 0, 
    0, 26, 25, 20, 28, 45, 48, 39, 37, 43, 49, 44, 21, 18, 0, 
    0, 24, 21, 18, 53, 18, 56, 50, 54, 54, 41, 58, 30, 21, 0, 
    20, 18, 6, 13, 36, 45, 48, 52, 50, 52, 45, 46, 27, 12, 0, 
    9, 4, 0, 18, 18, 35, 54, 54, 52, 46, 46, 40, 19, 8, 25, 
    0, 31, 0, 24, 10, 20, 64, 51, 46, 39, 49, 45, 27, 23, 10, 
    41, 46, 8, 14, 6, 27, 53, 57, 49, 35, 56, 43, 34, 23, 6, 
    10, 51, 37, 15, 7, 24, 37, 19, 54, 53, 48, 41, 20, 17, 0, 
    0, 5, 52, 48, 15, 13, 18, 22, 36, 50, 53, 29, 0, 18, 32, 
    0, 4, 22, 51, 46, 27, 12, 22, 14, 37, 29, 32, 12, 20, 47, 
    
    -- channel=129
    32, 23, 31, 33, 25, 16, 32, 26, 42, 34, 38, 29, 48, 15, 24, 
    39, 34, 42, 35, 21, 11, 18, 22, 43, 37, 41, 27, 58, 41, 42, 
    25, 14, 31, 27, 11, 21, 45, 43, 28, 25, 33, 39, 64, 47, 58, 
    32, 36, 42, 14, 16, 53, 55, 16, 25, 23, 53, 48, 62, 52, 46, 
    34, 48, 50, 36, 23, 55, 40, 28, 62, 54, 60, 53, 62, 52, 41, 
    24, 40, 62, 42, 53, 35, 36, 47, 54, 47, 48, 46, 62, 51, 42, 
    30, 40, 48, 60, 41, 25, 23, 28, 25, 25, 25, 29, 51, 58, 49, 
    29, 39, 39, 56, 29, 26, 17, 37, 31, 31, 27, 32, 32, 48, 25, 
    43, 52, 45, 47, 43, 17, 33, 31, 25, 24, 37, 24, 40, 31, 26, 
    47, 33, 27, 33, 28, 45, 20, 29, 39, 33, 25, 33, 19, 23, 47, 
    35, 32, 44, 47, 50, 21, 42, 40, 30, 34, 20, 27, 32, 39, 57, 
    52, 73, 70, 52, 48, 51, 32, 35, 33, 33, 29, 31, 33, 34, 61, 
    35, 50, 72, 79, 55, 52, 45, 24, 14, 28, 40, 24, 27, 25, 59, 
    32, 15, 40, 72, 85, 64, 56, 43, 37, 26, 26, 30, 11, 24, 45, 
    46, 19, 31, 54, 75, 83, 82, 62, 42, 26, 20, 17, 35, 47, 63, 
    
    -- channel=130
    13, 30, 4, 0, 27, 0, 5, 0, 0, 0, 7, 0, 41, 0, 10, 
    11, 26, 3, 0, 32, 0, 0, 0, 6, 0, 10, 0, 68, 9, 13, 
    0, 0, 0, 0, 29, 11, 21, 0, 0, 0, 0, 0, 27, 5, 8, 
    19, 2, 9, 16, 25, 0, 0, 4, 0, 45, 0, 0, 0, 0, 4, 
    20, 0, 54, 0, 0, 0, 39, 14, 9, 7, 0, 0, 0, 0, 34, 
    15, 0, 0, 90, 0, 0, 9, 0, 9, 0, 0, 0, 0, 0, 60, 
    42, 0, 0, 5, 0, 0, 14, 0, 0, 0, 2, 0, 0, 0, 56, 
    10, 0, 0, 0, 27, 0, 0, 0, 13, 26, 0, 0, 26, 0, 24, 
    11, 0, 0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 50, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 14, 7, 0, 
    3, 0, 19, 0, 0, 24, 0, 0, 0, 0, 0, 0, 3, 4, 0, 
    45, 45, 61, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 17, 28, 19, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    6, 0, 0, 0, 36, 11, 0, 37, 0, 0, 0, 0, 0, 0, 11, 
    12, 29, 0, 0, 0, 40, 27, 1, 0, 0, 0, 0, 59, 30, 0, 
    
    -- channel=131
    0, 0, 0, 0, 0, 1, 0, 0, 3, 6, 0, 13, 0, 18, 0, 
    0, 0, 0, 0, 0, 10, 4, 0, 0, 0, 0, 24, 0, 0, 0, 
    2, 6, 0, 0, 0, 0, 0, 0, 15, 0, 14, 21, 0, 0, 0, 
    0, 13, 0, 0, 0, 1, 0, 0, 3, 0, 15, 1, 17, 2, 0, 
    0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 5, 8, 0, 
    0, 49, 12, 0, 4, 11, 0, 18, 0, 5, 0, 0, 0, 20, 0, 
    0, 24, 24, 2, 0, 15, 0, 13, 8, 16, 10, 6, 1, 5, 0, 
    0, 17, 1, 13, 22, 0, 30, 10, 14, 2, 0, 38, 0, 9, 0, 
    0, 0, 7, 16, 33, 0, 24, 23, 19, 26, 11, 18, 16, 10, 0, 
    0, 8, 0, 14, 23, 48, 16, 25, 21, 24, 13, 14, 5, 0, 0, 
    0, 12, 0, 18, 0, 0, 50, 29, 25, 22, 25, 18, 0, 0, 7, 
    0, 0, 0, 0, 4, 11, 39, 37, 27, 8, 28, 16, 1, 6, 0, 
    30, 61, 0, 0, 0, 17, 32, 25, 52, 23, 36, 7, 1, 0, 0, 
    0, 21, 66, 9, 0, 0, 0, 0, 4, 39, 26, 5, 0, 0, 7, 
    0, 0, 27, 55, 12, 0, 0, 0, 0, 33, 42, 13, 0, 0, 24, 
    
    -- channel=132
    2, 7, 0, 7, 14, 0, 0, 0, 0, 0, 3, 0, 3, 0, 7, 
    2, 4, 3, 7, 15, 0, 7, 0, 0, 0, 1, 0, 4, 0, 0, 
    8, 1, 6, 13, 14, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    12, 0, 6, 5, 7, 0, 0, 9, 0, 0, 0, 0, 0, 0, 11, 
    7, 0, 4, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 3, 22, 
    11, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 12, 
    9, 0, 2, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 2, 21, 
    0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 4, 
    1, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 4, 
    11, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 
    
    -- channel=133
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=134
    18, 23, 30, 6, 0, 17, 7, 0, 0, 0, 0, 8, 0, 0, 10, 
    14, 31, 2, 3, 0, 0, 0, 11, 8, 9, 0, 12, 19, 63, 15, 
    0, 0, 0, 0, 0, 42, 60, 2, 0, 0, 0, 23, 9, 12, 15, 
    0, 42, 17, 0, 25, 39, 0, 0, 11, 15, 40, 16, 0, 7, 0, 
    5, 8, 21, 0, 25, 7, 0, 55, 34, 44, 0, 0, 0, 0, 0, 
    0, 0, 0, 58, 33, 0, 13, 32, 7, 0, 0, 25, 0, 0, 0, 
    24, 9, 0, 0, 0, 0, 15, 0, 0, 0, 6, 3, 0, 3, 2, 
    0, 0, 2, 0, 22, 0, 0, 2, 14, 37, 10, 0, 11, 0, 0, 
    23, 22, 0, 0, 0, 23, 3, 0, 0, 0, 0, 0, 0, 0, 4, 
    1, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 7, 11, 15, 0, 0, 0, 0, 0, 0, 0, 0, 13, 22, 
    63, 99, 56, 21, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 3, 35, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 18, 0, 22, 33, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 37, 25, 1, 0, 0, 0, 0, 46, 43, 36, 
    
    -- channel=135
    3, 0, 3, 0, 0, 30, 0, 10, 0, 5, 0, 37, 0, 25, 1, 
    3, 0, 0, 0, 0, 12, 11, 7, 0, 0, 0, 39, 0, 15, 0, 
    0, 0, 0, 0, 0, 34, 6, 0, 21, 0, 35, 36, 0, 0, 0, 
    0, 44, 0, 0, 8, 13, 0, 0, 14, 0, 28, 0, 0, 0, 0, 
    0, 48, 0, 0, 20, 0, 0, 24, 10, 0, 0, 18, 0, 0, 0, 
    0, 43, 12, 0, 4, 0, 0, 9, 0, 0, 0, 6, 0, 10, 0, 
    0, 22, 16, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 21, 0, 0, 4, 0, 10, 0, 1, 0, 0, 21, 0, 0, 0, 
    9, 0, 0, 3, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 27, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 21, 0, 32, 0, 0, 40, 0, 0, 0, 0, 0, 0, 12, 0, 
    27, 2, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 42, 0, 0, 0, 11, 0, 0, 28, 0, 0, 0, 0, 11, 0, 
    0, 0, 51, 13, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 14, 40, 10, 0, 0, 0, 0, 0, 0, 8, 0, 24, 24, 
    
    -- channel=136
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=137
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 15, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 24, 0, 5, 0, 0, 0, 0, 11, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 16, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 
    2, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 10, 
    0, 0, 17, 13, 24, 0, 0, 0, 0, 0, 0, 0, 26, 32, 0, 
    0, 23, 7, 13, 8, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    56, 67, 0, 0, 0, 2, 7, 51, 49, 0, 0, 0, 0, 28, 7, 
    0, 78, 74, 0, 0, 0, 0, 0, 0, 6, 0, 2, 31, 7, 0, 
    0, 0, 49, 56, 0, 0, 0, 0, 10, 32, 58, 12, 0, 0, 0, 
    
    -- channel=139
    16, 2, 24, 11, 11, 16, 18, 8, 23, 11, 16, 4, 26, 16, 5, 
    3, 1, 15, 11, 2, 20, 13, 7, 16, 14, 18, 8, 16, 19, 17, 
    12, 3, 5, 6, 0, 15, 23, 23, 6, 11, 20, 7, 20, 11, 16, 
    11, 20, 14, 5, 0, 36, 30, 1, 21, 0, 38, 17, 22, 8, 22, 
    4, 23, 7, 11, 9, 16, 11, 10, 28, 23, 29, 6, 20, 7, 13, 
    0, 24, 5, 0, 33, 11, 0, 17, 14, 14, 14, 11, 15, 10, 12, 
    0, 21, 5, 5, 7, 9, 6, 13, 5, 6, 0, 4, 9, 11, 2, 
    0, 13, 3, 6, 7, 0, 7, 7, 4, 6, 4, 1, 3, 10, 0, 
    4, 10, 3, 4, 6, 0, 6, 0, 5, 3, 2, 4, 1, 3, 0, 
    9, 1, 4, 15, 9, 13, 0, 1, 0, 4, 0, 6, 7, 7, 3, 
    6, 16, 8, 16, 8, 0, 13, 0, 0, 2, 0, 5, 10, 0, 24, 
    0, 29, 21, 19, 11, 6, 10, 7, 0, 0, 8, 7, 9, 14, 8, 
    16, 11, 13, 25, 17, 18, 9, 11, 0, 0, 8, 0, 13, 1, 21, 
    20, 18, 20, 16, 24, 27, 24, 10, 6, 9, 0, 3, 5, 18, 3, 
    22, 17, 30, 25, 15, 15, 26, 30, 13, 11, 9, 0, 1, 19, 39, 
    
    -- channel=140
    58, 45, 40, 55, 46, 3, 52, 42, 67, 67, 79, 49, 110, 19, 55, 
    84, 74, 72, 62, 48, 0, 32, 39, 73, 65, 76, 47, 131, 52, 85, 
    62, 53, 66, 60, 39, 19, 60, 66, 57, 62, 46, 66, 148, 100, 104, 
    59, 43, 84, 58, 35, 62, 90, 52, 30, 69, 65, 90, 141, 117, 107, 
    73, 65, 124, 59, 49, 104, 97, 35, 89, 86, 110, 97, 134, 120, 105, 
    74, 53, 127, 124, 76, 89, 88, 92, 119, 108, 105, 85, 140, 112, 106, 
    81, 63, 102, 131, 111, 85, 91, 94, 91, 83, 94, 114, 122, 113, 117, 
    84, 71, 103, 117, 110, 90, 82, 103, 109, 110, 106, 98, 138, 108, 94, 
    89, 105, 104, 104, 95, 123, 94, 111, 115, 113, 115, 110, 113, 96, 83, 
    103, 99, 80, 69, 82, 75, 116, 120, 127, 129, 114, 113, 101, 66, 78, 
    104, 60, 94, 75, 99, 92, 88, 143, 131, 121, 106, 107, 104, 93, 105, 
    115, 142, 145, 96, 105, 93, 109, 127, 130, 125, 111, 108, 102, 89, 122, 
    88, 107, 173, 156, 121, 89, 111, 99, 76, 121, 116, 118, 91, 71, 106, 
    77, 29, 77, 158, 170, 125, 104, 105, 79, 106, 113, 113, 77, 41, 103, 
    81, 35, 22, 92, 165, 181, 152, 128, 93, 79, 80, 92, 94, 85, 87, 
    
    -- channel=141
    10, 7, 13, 25, 15, 7, 10, 13, 11, 12, 12, 16, 0, 7, 8, 
    21, 12, 20, 25, 10, 5, 11, 10, 13, 16, 11, 17, 0, 16, 19, 
    15, 4, 19, 22, 6, 6, 17, 18, 19, 13, 6, 24, 11, 23, 17, 
    15, 16, 18, 6, 7, 13, 11, 6, 14, 5, 13, 22, 19, 22, 19, 
    18, 29, 20, 12, 2, 12, 4, 6, 16, 17, 11, 15, 17, 30, 15, 
    10, 27, 32, 17, 16, 0, 0, 4, 5, 0, 0, 9, 15, 34, 6, 
    10, 24, 32, 21, 0, 0, 0, 0, 0, 0, 0, 0, 4, 29, 12, 
    15, 25, 26, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 14, 
    18, 25, 29, 27, 18, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 
    27, 22, 17, 16, 17, 17, 0, 0, 0, 0, 0, 0, 0, 9, 21, 
    19, 8, 14, 24, 25, 11, 8, 0, 0, 0, 0, 0, 0, 17, 31, 
    15, 7, 5, 28, 23, 22, 2, 0, 0, 0, 0, 0, 0, 10, 34, 
    23, 15, 0, 8, 16, 25, 10, 0, 0, 0, 0, 0, 0, 10, 30, 
    8, 10, 8, 3, 5, 14, 15, 9, 14, 0, 0, 0, 0, 7, 20, 
    10, 0, 9, 12, 6, 8, 12, 14, 2, 0, 0, 0, 1, 16, 17, 
    
    -- channel=142
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 4, 0, 0, 
    0, 6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 4, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 17, 3, 0, 0, 0, 0, 0, 0, 0, 
    8, 2, 0, 0, 0, 6, 1, 4, 2, 0, 0, 0, 0, 0, 2, 
    0, 31, 15, 3, 0, 4, 2, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 26, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 31, 28, 12, 4, 2, 0, 0, 0, 0, 0, 0, 13, 
    
    -- channel=143
    5, 0, 9, 20, 22, 6, 13, 10, 23, 18, 19, 7, 12, 13, 5, 
    7, 4, 16, 22, 17, 19, 16, 10, 8, 14, 15, 8, 0, 0, 12, 
    36, 18, 18, 26, 12, 0, 0, 27, 17, 33, 5, 7, 4, 13, 17, 
    15, 0, 18, 9, 0, 6, 28, 15, 18, 0, 3, 16, 17, 15, 34, 
    18, 16, 6, 20, 0, 9, 8, 0, 1, 2, 16, 14, 14, 22, 28, 
    18, 28, 16, 0, 11, 7, 0, 0, 5, 10, 5, 4, 16, 24, 16, 
    3, 18, 27, 17, 3, 0, 0, 0, 3, 0, 0, 0, 8, 22, 7, 
    16, 16, 19, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 25, 
    4, 15, 31, 24, 23, 0, 0, 0, 0, 0, 0, 0, 14, 17, 3, 
    26, 25, 27, 27, 15, 28, 0, 0, 0, 0, 0, 0, 0, 12, 4, 
    27, 10, 12, 8, 19, 4, 3, 0, 0, 3, 0, 0, 0, 2, 22, 
    0, 0, 0, 21, 21, 14, 3, 0, 0, 0, 0, 0, 0, 11, 26, 
    47, 26, 0, 0, 10, 24, 9, 19, 10, 0, 0, 0, 0, 12, 38, 
    21, 49, 25, 0, 0, 5, 14, 0, 3, 2, 0, 2, 9, 22, 0, 
    20, 0, 34, 21, 0, 0, 3, 8, 24, 11, 19, 0, 0, 0, 12, 
    
    -- channel=144
    33, 9, 23, 35, 5, 6, 32, 35, 59, 65, 50, 63, 52, 23, 33, 
    59, 43, 44, 44, 5, 7, 21, 33, 50, 52, 45, 71, 59, 38, 61, 
    70, 57, 50, 45, 4, 1, 31, 49, 54, 41, 38, 85, 103, 78, 79, 
    22, 34, 53, 36, 8, 49, 65, 18, 39, 33, 52, 101, 119, 100, 79, 
    40, 86, 77, 34, 51, 79, 40, 19, 58, 70, 88, 100, 115, 110, 50, 
    45, 85, 113, 53, 59, 83, 69, 91, 93, 89, 77, 95, 116, 109, 40, 
    40, 66, 108, 119, 95, 87, 73, 87, 89, 93, 91, 103, 101, 108, 51, 
    60, 73, 100, 118, 96, 74, 90, 101, 97, 87, 97, 120, 108, 107, 47, 
    67, 88, 100, 101, 122, 105, 101, 111, 114, 117, 109, 119, 116, 96, 47, 
    98, 91, 69, 81, 86, 103, 120, 125, 127, 129, 111, 110, 76, 48, 59, 
    78, 66, 61, 62, 81, 84, 113, 145, 136, 121, 114, 102, 85, 73, 97, 
    77, 102, 80, 83, 87, 90, 125, 139, 137, 116, 111, 109, 88, 93, 100, 
    119, 151, 140, 107, 89, 102, 124, 116, 117, 122, 125, 104, 78, 68, 95, 
    50, 65, 128, 137, 112, 92, 94, 67, 82, 121, 124, 108, 59, 52, 72, 
    48, 6, 52, 136, 151, 127, 105, 95, 94, 105, 114, 83, 38, 36, 99, 
    
    -- channel=145
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 10, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 16, 19, 7, 3, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 15, 16, 0, 
    0, 18, 16, 0, 0, 0, 0, 1, 1, 7, 0, 0, 12, 17, 0, 
    0, 5, 19, 14, 6, 4, 1, 16, 4, 0, 0, 13, 5, 15, 0, 
    0, 7, 13, 14, 0, 6, 14, 11, 2, 9, 16, 15, 9, 13, 0, 
    0, 8, 16, 13, 37, 0, 14, 15, 23, 28, 17, 31, 21, 11, 0, 
    12, 13, 0, 3, 5, 33, 19, 24, 25, 22, 17, 22, 0, 0, 0, 
    7, 0, 0, 0, 10, 1, 28, 39, 27, 29, 20, 16, 10, 0, 5, 
    0, 5, 0, 7, 0, 14, 31, 35, 37, 16, 19, 18, 9, 10, 17, 
    30, 46, 14, 7, 6, 6, 27, 29, 30, 21, 28, 16, 0, 11, 1, 
    0, 4, 21, 10, 4, 14, 11, 0, 6, 31, 26, 15, 1, 0, 0, 
    0, 0, 0, 21, 10, 5, 2, 14, 14, 22, 28, 6, 0, 0, 7, 
    0, 0, 0, 0, 23, 21, 7, 5, 0, 0, 0, 3, 7, 7, 22, 
    
    -- channel=146
    0, 8, 0, 0, 23, 0, 0, 0, 0, 10, 4, 0, 0, 12, 0, 
    0, 0, 0, 0, 28, 0, 28, 0, 0, 0, 10, 0, 17, 0, 0, 
    0, 26, 5, 0, 37, 0, 0, 0, 21, 5, 15, 0, 0, 0, 0, 
    26, 0, 0, 10, 19, 0, 0, 73, 0, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 3, 0, 0, 33, 
    17, 0, 0, 6, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 16, 3, 0, 7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 7, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 11, 0, 
    0, 0, 21, 0, 0, 0, 0, 5, 0, 0, 0, 0, 35, 0, 46, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 0, 0, 
    
    -- channel=147
    18, 25, 19, 23, 12, 25, 20, 26, 21, 33, 22, 37, 14, 24, 29, 
    27, 31, 22, 22, 16, 15, 22, 28, 24, 25, 21, 35, 28, 23, 22, 
    13, 31, 27, 16, 22, 33, 28, 15, 32, 15, 30, 35, 24, 32, 20, 
    21, 33, 12, 24, 36, 28, 26, 33, 21, 36, 27, 37, 23, 27, 5, 
    23, 26, 30, 8, 36, 32, 32, 38, 28, 34, 26, 45, 29, 25, 5, 
    22, 18, 31, 41, 28, 31, 22, 29, 39, 36, 35, 49, 29, 26, 10, 
    27, 20, 26, 29, 21, 28, 30, 22, 22, 22, 28, 30, 32, 31, 20, 
    29, 26, 30, 22, 31, 21, 28, 20, 30, 31, 22, 23, 23, 30, 19, 
    32, 26, 22, 27, 13, 36, 15, 23, 26, 26, 23, 20, 9, 17, 37, 
    19, 27, 25, 22, 30, 0, 30, 24, 19, 21, 26, 21, 21, 23, 32, 
    20, 31, 27, 26, 23, 40, 16, 20, 23, 11, 24, 22, 22, 30, 21, 
    43, 35, 42, 31, 26, 24, 20, 20, 21, 20, 23, 18, 24, 30, 34, 
    16, 30, 49, 45, 37, 19, 17, 4, 18, 26, 12, 24, 16, 35, 28, 
    19, 16, 40, 49, 49, 44, 33, 37, 24, 14, 26, 15, 17, 26, 57, 
    15, 31, 16, 39, 44, 54, 51, 41, 17, 10, 6, 34, 34, 34, 27, 
    
    -- channel=148
    0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 4, 0, 15, 0, 0, 
    7, 18, 0, 0, 6, 0, 0, 0, 0, 5, 0, 0, 6, 0, 8, 
    23, 0, 0, 12, 3, 0, 0, 11, 0, 18, 0, 4, 25, 14, 15, 
    0, 0, 17, 2, 0, 0, 7, 0, 0, 0, 0, 10, 21, 22, 25, 
    14, 0, 18, 17, 0, 9, 5, 0, 0, 2, 15, 12, 20, 30, 21, 
    24, 0, 19, 21, 0, 12, 29, 11, 26, 13, 10, 16, 30, 16, 20, 
    16, 0, 20, 37, 34, 20, 14, 20, 25, 26, 29, 33, 22, 23, 24, 
    17, 0, 28, 30, 16, 50, 15, 33, 25, 24, 40, 29, 49, 21, 28, 
    10, 21, 32, 20, 44, 37, 37, 36, 40, 35, 37, 43, 52, 32, 8, 
    35, 26, 21, 9, 2, 28, 43, 42, 51, 47, 44, 38, 21, 8, 0, 
    26, 0, 14, 0, 30, 18, 16, 53, 50, 50, 37, 29, 26, 13, 18, 
    10, 16, 17, 10, 15, 20, 30, 42, 49, 51, 31, 41, 30, 13, 19, 
    37, 19, 30, 24, 13, 13, 40, 52, 24, 40, 42, 43, 27, 13, 19, 
    6, 13, 0, 19, 27, 8, 8, 2, 27, 36, 39, 51, 24, 1, 0, 
    12, 0, 0, 0, 27, 32, 19, 4, 26, 29, 38, 17, 10, 0, 0, 
    
    -- channel=149
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 9, 6, 0, 17, 1, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 4, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 11, 5, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 3, 0, 0, 3, 3, 0, 0, 
    5, 21, 0, 0, 0, 0, 0, 18, 28, 0, 3, 1, 0, 0, 0, 
    0, 17, 23, 0, 0, 0, 0, 0, 0, 8, 2, 6, 4, 0, 0, 
    0, 0, 6, 8, 0, 0, 0, 0, 0, 13, 18, 4, 0, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 6, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 
    9, 20, 0, 0, 0, 0, 0, 0, 9, 0, 6, 8, 24, 0, 1, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 9, 0, 4, 42, 17, 11, 
    0, 12, 12, 0, 3, 0, 0, 0, 0, 0, 0, 14, 26, 26, 3, 
    0, 16, 29, 0, 0, 22, 24, 14, 3, 11, 13, 4, 20, 31, 0, 
    0, 0, 25, 27, 25, 43, 39, 27, 40, 48, 47, 30, 32, 10, 5, 
    5, 10, 16, 32, 61, 18, 55, 50, 53, 38, 36, 73, 39, 25, 4, 
    7, 0, 19, 25, 44, 67, 44, 65, 55, 68, 60, 54, 58, 32, 6, 
    10, 24, 9, 15, 37, 49, 69, 65, 66, 67, 60, 54, 45, 6, 0, 
    14, 16, 0, 4, 0, 28, 56, 71, 76, 64, 67, 59, 36, 14, 2, 
    17, 2, 0, 0, 19, 11, 57, 78, 75, 60, 59, 56, 38, 25, 7, 
    30, 76, 42, 0, 0, 26, 47, 61, 83, 73, 65, 58, 34, 12, 0, 
    0, 0, 62, 45, 0, 0, 12, 24, 8, 69, 74, 51, 34, 0, 11, 
    0, 0, 0, 50, 54, 5, 0, 2, 20, 57, 66, 59, 0, 0, 0, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 3, 
    0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    
    -- channel=152
    65, 38, 65, 63, 27, 48, 57, 55, 73, 71, 68, 86, 66, 48, 64, 
    76, 67, 66, 69, 21, 33, 41, 63, 72, 75, 63, 96, 85, 82, 80, 
    60, 61, 70, 51, 20, 55, 82, 67, 67, 44, 76, 103, 113, 99, 102, 
    48, 93, 71, 54, 39, 99, 89, 26, 77, 59, 95, 122, 119, 108, 74, 
    57, 110, 99, 44, 81, 100, 57, 77, 90, 106, 110, 96, 117, 108, 48, 
    39, 97, 115, 88, 107, 96, 66, 106, 108, 102, 85, 122, 110, 108, 48, 
    61, 90, 102, 119, 83, 78, 87, 88, 83, 81, 88, 104, 96, 116, 60, 
    68, 92, 108, 110, 111, 57, 93, 97, 93, 102, 95, 103, 106, 105, 38, 
    90, 103, 83, 91, 92, 111, 86, 94, 105, 105, 94, 100, 77, 64, 66, 
    99, 74, 71, 89, 86, 73, 103, 116, 105, 108, 97, 95, 72, 73, 86, 
    67, 92, 73, 86, 92, 97, 114, 118, 114, 93, 93, 93, 82, 83, 113, 
    115, 149, 114, 106, 93, 95, 114, 114, 107, 94, 109, 91, 79, 91, 107, 
    88, 117, 146, 132, 106, 105, 99, 64, 80, 105, 98, 88, 72, 62, 104, 
    68, 47, 114, 152, 136, 119, 107, 97, 99, 99, 107, 80, 33, 85, 105, 
    60, 52, 58, 123, 151, 151, 136, 126, 84, 75, 66, 70, 79, 87, 137, 
    
    -- channel=153
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=154
    19, 19, 25, 11, 13, 19, 19, 12, 18, 9, 16, 7, 32, 10, 18, 
    10, 23, 13, 10, 14, 18, 8, 18, 16, 17, 16, 8, 29, 24, 20, 
    12, 10, 10, 8, 14, 25, 27, 20, 1, 14, 15, 6, 24, 14, 16, 
    13, 19, 17, 19, 18, 30, 20, 4, 20, 16, 29, 18, 9, 10, 15, 
    14, 7, 19, 16, 23, 16, 21, 26, 22, 24, 24, 1, 14, 7, 13, 
    14, 3, 2, 23, 28, 14, 26, 25, 24, 18, 19, 23, 18, 0, 22, 
    21, 11, 0, 9, 21, 24, 31, 26, 23, 22, 23, 27, 17, 11, 14, 
    13, 8, 11, 5, 24, 24, 22, 26, 27, 32, 29, 13, 32, 14, 7, 
    13, 14, 1, 0, 2, 29, 21, 19, 28, 20, 21, 21, 13, 8, 21, 
    12, 3, 11, 12, 6, 0, 20, 22, 18, 23, 21, 23, 24, 20, 8, 
    8, 19, 19, 7, 16, 16, 9, 18, 19, 15, 20, 23, 29, 10, 19, 
    13, 38, 38, 18, 7, 6, 15, 18, 13, 19, 24, 26, 28, 18, 4, 
    2, 0, 24, 30, 22, 8, 8, 17, 0, 19, 17, 24, 32, 11, 10, 
    21, 6, 0, 16, 33, 24, 18, 21, 17, 16, 20, 24, 21, 23, 3, 
    19, 30, 13, 1, 16, 29, 31, 17, 16, 13, 9, 12, 29, 20, 24, 
    
    -- channel=155
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=156
    0, 24, 0, 0, 59, 0, 0, 0, 0, 0, 30, 0, 93, 0, 0, 
    0, 14, 5, 0, 68, 0, 0, 0, 6, 0, 31, 0, 90, 0, 7, 
    0, 0, 0, 4, 60, 0, 0, 1, 0, 34, 0, 0, 41, 0, 0, 
    38, 0, 9, 23, 6, 0, 8, 48, 0, 49, 0, 0, 21, 0, 54, 
    32, 0, 63, 15, 0, 0, 70, 0, 0, 0, 0, 0, 0, 0, 109, 
    52, 0, 0, 75, 0, 0, 19, 0, 2, 0, 13, 0, 15, 0, 126, 
    50, 0, 0, 8, 14, 0, 8, 0, 0, 0, 0, 0, 17, 0, 101, 
    26, 0, 0, 0, 15, 15, 0, 0, 7, 0, 0, 0, 28, 0, 97, 
    0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 6, 0, 13, 0, 67, 
    0, 8, 20, 0, 2, 0, 0, 0, 0, 3, 0, 4, 49, 3, 0, 
    52, 0, 29, 0, 0, 14, 0, 0, 9, 3, 0, 6, 18, 0, 0, 
    0, 0, 50, 0, 27, 0, 0, 0, 0, 23, 0, 2, 19, 0, 0, 
    0, 0, 25, 19, 17, 0, 0, 16, 0, 3, 0, 23, 31, 0, 0, 
    35, 0, 0, 0, 27, 3, 0, 30, 0, 0, 0, 19, 73, 0, 0, 
    50, 16, 0, 0, 0, 15, 14, 0, 8, 0, 0, 19, 35, 0, 0, 
    
    -- channel=157
    11, 2, 4, 6, 0, 12, 5, 12, 18, 25, 12, 23, 9, 22, 11, 
    12, 2, 11, 7, 0, 13, 16, 12, 12, 12, 13, 24, 17, 2, 8, 
    11, 25, 13, 7, 0, 12, 3, 3, 23, 4, 30, 20, 23, 14, 15, 
    8, 17, 3, 9, 4, 16, 16, 18, 14, 11, 21, 18, 32, 18, 11, 
    0, 28, 6, 4, 19, 24, 13, 8, 17, 10, 26, 37, 29, 18, 6, 
    4, 31, 25, 0, 16, 22, 20, 22, 22, 30, 33, 19, 26, 24, 0, 
    1, 19, 28, 19, 27, 30, 30, 29, 35, 27, 29, 33, 33, 19, 5, 
    12, 20, 15, 22, 24, 17, 39, 32, 32, 27, 24, 34, 24, 29, 5, 
    15, 13, 18, 26, 25, 22, 25, 34, 31, 40, 36, 27, 36, 32, 4, 
    10, 23, 10, 22, 21, 33, 30, 27, 35, 31, 33, 30, 24, 14, 23, 
    15, 24, 9, 22, 12, 10, 36, 33, 28, 34, 35, 36, 28, 19, 11, 
    20, 15, 13, 12, 16, 23, 31, 41, 36, 27, 33, 31, 37, 24, 25, 
    26, 60, 43, 21, 15, 19, 25, 32, 48, 34, 33, 33, 24, 35, 16, 
    13, 29, 64, 47, 27, 19, 23, 21, 10, 35, 35, 27, 23, 21, 37, 
    9, 9, 32, 56, 48, 30, 24, 28, 18, 33, 34, 38, 11, 21, 24, 
    
    -- channel=158
    18, 10, 0, 13, 28, 0, 16, 4, 21, 24, 43, 0, 67, 0, 17, 
    21, 15, 22, 15, 27, 0, 13, 0, 26, 12, 41, 0, 73, 0, 26, 
    35, 31, 27, 18, 23, 0, 6, 21, 16, 22, 25, 0, 68, 27, 46, 
    26, 0, 25, 27, 2, 0, 42, 32, 0, 37, 0, 16, 73, 39, 59, 
    26, 0, 55, 19, 4, 26, 41, 0, 18, 20, 44, 25, 58, 44, 75, 
    34, 1, 55, 46, 0, 34, 41, 10, 31, 31, 38, 5, 65, 46, 73, 
    31, 0, 27, 55, 42, 28, 33, 22, 41, 32, 28, 22, 49, 31, 74, 
    38, 15, 28, 52, 40, 19, 26, 42, 35, 27, 34, 32, 52, 37, 55, 
    24, 21, 38, 42, 37, 63, 16, 39, 33, 44, 51, 35, 70, 42, 49, 
    34, 43, 40, 30, 33, 29, 49, 35, 48, 48, 43, 47, 47, 20, 19, 
    52, 20, 40, 13, 27, 37, 23, 55, 50, 55, 44, 47, 47, 28, 23, 
    36, 15, 52, 23, 45, 26, 33, 56, 53, 55, 38, 42, 49, 25, 50, 
    39, 60, 74, 56, 53, 32, 43, 57, 43, 52, 39, 50, 39, 17, 47, 
    37, 4, 46, 69, 61, 45, 49, 56, 4, 42, 48, 54, 51, 16, 36, 
    49, 16, 0, 44, 76, 56, 50, 46, 47, 46, 42, 51, 35, 6, 0, 
    
    -- channel=159
    17, 8, 28, 19, 0, 45, 20, 28, 32, 29, 7, 49, 0, 42, 19, 
    14, 10, 16, 17, 0, 42, 20, 36, 16, 29, 7, 59, 0, 33, 14, 
    21, 25, 16, 12, 0, 36, 28, 22, 28, 5, 33, 54, 0, 20, 13, 
    4, 43, 11, 10, 13, 45, 24, 5, 49, 1, 38, 50, 6, 15, 0, 
    4, 52, 0, 11, 42, 27, 0, 34, 26, 32, 31, 42, 15, 13, 0, 
    0, 57, 12, 0, 41, 26, 6, 33, 16, 23, 12, 42, 12, 18, 0, 
    0, 41, 30, 11, 14, 27, 21, 29, 22, 24, 21, 29, 6, 24, 0, 
    6, 34, 25, 17, 13, 13, 36, 23, 18, 21, 23, 25, 5, 18, 0, 
    15, 25, 15, 19, 38, 1, 28, 19, 23, 25, 15, 29, 9, 21, 0, 
    19, 12, 11, 33, 18, 39, 21, 19, 19, 13, 18, 15, 0, 15, 29, 
    0, 33, 5, 28, 27, 14, 46, 17, 9, 15, 22, 17, 10, 14, 21, 
    14, 20, 0, 32, 6, 32, 36, 22, 16, 5, 24, 17, 20, 24, 17, 
    35, 50, 12, 10, 15, 29, 29, 17, 43, 13, 20, 10, 9, 32, 22, 
    6, 55, 63, 25, 6, 22, 29, 10, 41, 27, 19, 11, 0, 46, 25, 
    1, 21, 70, 64, 23, 11, 13, 27, 22, 33, 30, 14, 3, 22, 60, 
    
    -- channel=160
    53, 62, 63, 70, 68, 67, 63, 60, 31, 33, 41, 37, 42, 46, 32, 
    63, 61, 69, 71, 75, 74, 69, 75, 50, 22, 43, 44, 54, 44, 44, 
    42, 69, 70, 75, 76, 75, 72, 74, 75, 48, 59, 45, 49, 52, 49, 
    49, 63, 69, 77, 74, 82, 74, 68, 73, 76, 64, 39, 46, 52, 51, 
    51, 68, 71, 75, 77, 70, 64, 68, 48, 76, 66, 24, 47, 45, 50, 
    83, 62, 76, 70, 64, 82, 34, 36, 45, 64, 43, 16, 38, 41, 50, 
    58, 81, 62, 60, 70, 59, 55, 51, 58, 52, 25, 15, 30, 42, 42, 
    43, 85, 59, 59, 76, 66, 68, 70, 57, 57, 22, 10, 37, 59, 19, 
    60, 84, 62, 35, 65, 72, 42, 56, 55, 34, 9, 14, 43, 69, 4, 
    59, 83, 58, 0, 63, 62, 42, 87, 29, 21, 25, 22, 44, 84, 0, 
    59, 75, 47, 6, 25, 18, 37, 54, 24, 13, 13, 35, 40, 79, 19, 
    64, 66, 59, 53, 41, 54, 52, 24, 4, 6, 0, 9, 44, 44, 62, 
    72, 73, 53, 64, 41, 50, 71, 45, 27, 20, 11, 20, 26, 35, 42, 
    54, 74, 54, 57, 42, 61, 71, 57, 56, 46, 50, 56, 48, 49, 41, 
    71, 72, 67, 69, 63, 68, 62, 62, 58, 59, 67, 71, 61, 52, 59, 
    
    -- channel=161
    23, 22, 10, 6, 9, 5, 2, 1, 7, 0, 0, 0, 0, 0, 0, 
    18, 21, 8, 13, 12, 13, 6, 0, 1, 0, 0, 0, 0, 0, 0, 
    23, 21, 13, 13, 15, 12, 9, 9, 10, 10, 11, 0, 0, 0, 0, 
    18, 25, 15, 14, 17, 7, 10, 4, 7, 8, 5, 3, 0, 0, 0, 
    9, 17, 18, 13, 19, 13, 10, 13, 7, 0, 5, 12, 0, 0, 0, 
    0, 14, 23, 22, 15, 31, 34, 25, 4, 5, 2, 1, 0, 0, 0, 
    7, 9, 31, 20, 20, 32, 20, 18, 33, 27, 11, 0, 0, 0, 0, 
    1, 9, 24, 25, 28, 41, 24, 31, 36, 32, 24, 1, 0, 10, 8, 
    3, 8, 30, 15, 18, 11, 20, 7, 6, 4, 0, 0, 0, 11, 8, 
    0, 9, 33, 7, 21, 12, 12, 20, 11, 0, 0, 0, 0, 18, 29, 
    2, 1, 22, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 34, 
    0, 0, 15, 23, 14, 3, 7, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 2, 2, 19, 21, 0, 0, 4, 2, 0, 0, 0, 0, 0, 1, 
    0, 0, 7, 0, 4, 1, 2, 0, 2, 4, 4, 10, 8, 5, 7, 
    0, 0, 0, 4, 5, 7, 0, 0, 0, 0, 0, 2, 3, 2, 0, 
    
    -- channel=162
    42, 16, 0, 0, 0, 0, 0, 0, 5, 0, 0, 7, 5, 0, 9, 
    0, 0, 0, 0, 0, 3, 5, 0, 20, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 3, 53, 13, 13, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 16, 2, 0, 0, 13, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 17, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 56, 31, 13, 17, 15, 0, 0, 0, 
    5, 0, 0, 0, 0, 7, 6, 0, 0, 0, 36, 6, 0, 9, 14, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 
    7, 0, 0, 29, 0, 0, 2, 1, 16, 0, 21, 13, 0, 0, 71, 
    0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 
    0, 0, 0, 58, 27, 35, 19, 6, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 0, 2, 31, 40, 37, 32, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 10, 13, 20, 29, 24, 36, 8, 0, 
    0, 0, 3, 0, 18, 0, 0, 0, 0, 0, 0, 0, 4, 8, 0, 
    
    -- channel=163
    0, 0, 10, 13, 9, 10, 4, 7, 0, 4, 12, 1, 1, 14, 0, 
    6, 9, 4, 13, 15, 5, 0, 12, 0, 0, 20, 14, 20, 9, 4, 
    4, 23, 8, 15, 13, 12, 4, 7, 4, 0, 5, 0, 17, 16, 9, 
    0, 26, 15, 17, 14, 14, 12, 5, 20, 16, 0, 0, 13, 11, 14, 
    22, 18, 14, 13, 14, 10, 12, 8, 0, 30, 9, 0, 15, 16, 19, 
    43, 13, 15, 12, 12, 14, 5, 28, 15, 26, 11, 0, 21, 10, 19, 
    36, 37, 21, 17, 4, 27, 15, 0, 6, 5, 0, 0, 8, 8, 15, 
    4, 54, 19, 20, 28, 14, 3, 31, 25, 25, 0, 0, 14, 18, 0, 
    5, 45, 17, 0, 60, 32, 6, 42, 42, 36, 17, 0, 17, 38, 0, 
    13, 45, 27, 0, 84, 38, 7, 39, 0, 0, 0, 0, 22, 50, 0, 
    12, 39, 34, 0, 7, 33, 34, 54, 6, 0, 10, 20, 7, 64, 0, 
    20, 23, 31, 0, 0, 0, 0, 5, 0, 0, 0, 10, 25, 29, 44, 
    17, 28, 11, 41, 0, 18, 21, 0, 0, 0, 0, 0, 13, 4, 29, 
    19, 37, 14, 14, 16, 15, 34, 8, 1, 0, 0, 0, 0, 0, 19, 
    22, 23, 14, 14, 4, 23, 18, 23, 18, 10, 18, 20, 8, 6, 4, 
    
    -- channel=164
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 0, 0, 7, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 8, 5, 0, 0, 0, 8, 
    0, 0, 0, 13, 1, 16, 1, 0, 7, 4, 5, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 15, 13, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=165
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=166
    21, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 
    0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 44, 42, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 9, 0, 0, 39, 65, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 7, 11, 0, 0, 0, 8, 0, 0, 28, 4, 
    4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 12, 18, 0, 8, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 53, 31, 53, 44, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 4, 25, 37, 36, 29, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 15, 25, 36, 51, 45, 32, 0, 
    0, 13, 0, 11, 18, 6, 0, 0, 0, 0, 2, 2, 3, 0, 13, 
    
    -- channel=167
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 2, 4, 0, 2, 
    0, 9, 0, 0, 0, 0, 0, 0, 1, 0, 3, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 5, 0, 1, 
    61, 0, 3, 0, 0, 27, 0, 0, 0, 11, 0, 0, 11, 0, 3, 
    6, 21, 0, 0, 5, 0, 0, 0, 9, 0, 0, 0, 5, 0, 0, 
    0, 39, 0, 0, 6, 0, 0, 6, 0, 0, 0, 0, 18, 20, 0, 
    0, 26, 0, 0, 1, 11, 0, 0, 0, 0, 0, 0, 21, 26, 0, 
    0, 30, 0, 0, 72, 0, 0, 35, 0, 0, 1, 0, 19, 49, 0, 
    0, 11, 0, 0, 0, 0, 4, 3, 0, 0, 0, 23, 0, 43, 0, 
    0, 0, 16, 0, 0, 3, 0, 0, 0, 1, 0, 0, 27, 0, 34, 
    0, 7, 0, 23, 0, 0, 14, 0, 0, 0, 0, 10, 0, 3, 0, 
    0, 14, 0, 0, 0, 3, 7, 0, 2, 0, 0, 3, 0, 0, 7, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 3, 
    
    -- channel=168
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=169
    0, 10, 23, 28, 26, 33, 27, 25, 11, 12, 12, 14, 12, 15, 5, 
    11, 11, 23, 24, 27, 28, 34, 33, 24, 21, 14, 15, 13, 16, 13, 
    10, 8, 24, 26, 27, 28, 33, 40, 22, 0, 8, 18, 28, 19, 15, 
    0, 9, 20, 23, 25, 33, 35, 35, 33, 23, 28, 25, 21, 26, 20, 
    2, 11, 17, 27, 23, 31, 20, 18, 29, 37, 28, 12, 15, 17, 16, 
    10, 13, 19, 20, 26, 0, 0, 8, 0, 17, 25, 13, 11, 16, 19, 
    29, 5, 3, 5, 4, 5, 0, 0, 0, 0, 1, 4, 7, 14, 20, 
    20, 15, 0, 2, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 15, 
    20, 12, 0, 12, 0, 5, 17, 24, 10, 19, 5, 7, 11, 2, 0, 
    29, 20, 0, 8, 0, 8, 1, 0, 27, 13, 0, 7, 10, 0, 0, 
    26, 24, 0, 0, 33, 32, 20, 54, 17, 18, 12, 0, 18, 12, 0, 
    20, 30, 0, 0, 2, 0, 12, 22, 16, 5, 0, 15, 11, 33, 0, 
    29, 22, 28, 0, 4, 17, 21, 10, 0, 0, 0, 0, 13, 15, 36, 
    34, 27, 17, 29, 2, 18, 25, 23, 11, 4, 0, 1, 1, 13, 0, 
    18, 28, 21, 21, 10, 22, 33, 24, 27, 27, 26, 23, 22, 20, 17, 
    
    -- channel=170
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 3, 0, 
    17, 0, 0, 0, 4, 0, 0, 42, 14, 0, 3, 12, 7, 0, 0, 
    0, 13, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 6, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 19, 13, 7, 52, 47, 73, 70, 15, 0, 0, 0, 
    0, 0, 0, 0, 81, 19, 11, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 11, 18, 0, 0, 71, 48, 56, 53, 14, 29, 8, 0, 25, 0, 
    2, 0, 5, 0, 0, 0, 0, 0, 5, 8, 7, 21, 12, 34, 14, 
    0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    1, 12, 0, 1, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=171
    2, 26, 17, 19, 20, 22, 18, 15, 14, 7, 7, 7, 6, 10, 2, 
    12, 17, 12, 20, 23, 20, 20, 22, 19, 8, 9, 8, 10, 10, 5, 
    17, 19, 16, 17, 19, 19, 21, 18, 18, 10, 20, 8, 11, 7, 7, 
    0, 20, 17, 18, 19, 16, 18, 13, 17, 14, 11, 12, 10, 9, 8, 
    5, 15, 16, 16, 19, 19, 7, 11, 11, 14, 7, 13, 10, 10, 9, 
    0, 10, 19, 16, 14, 8, 9, 15, 1, 11, 10, 0, 14, 9, 10, 
    25, 0, 12, 12, 1, 21, 0, 5, 15, 8, 2, 0, 7, 12, 11, 
    8, 14, 8, 5, 8, 6, 6, 13, 4, 5, 7, 1, 0, 14, 7, 
    8, 9, 6, 0, 26, 0, 11, 14, 10, 9, 0, 1, 5, 13, 1, 
    6, 10, 3, 7, 20, 5, 0, 19, 13, 0, 0, 14, 10, 13, 9, 
    8, 5, 9, 0, 11, 6, 0, 18, 0, 1, 7, 8, 8, 13, 10, 
    0, 11, 4, 3, 12, 7, 11, 14, 1, 5, 8, 9, 3, 8, 10, 
    5, 7, 5, 7, 1, 9, 5, 7, 5, 6, 9, 10, 17, 0, 18, 
    9, 0, 6, 0, 7, 10, 13, 5, 5, 8, 6, 16, 9, 14, 15, 
    6, 13, 1, 7, 1, 16, 12, 8, 8, 3, 9, 11, 7, 11, 4, 
    
    -- channel=172
    98, 63, 62, 58, 65, 55, 52, 47, 54, 20, 25, 31, 28, 28, 42, 
    89, 89, 70, 71, 68, 68, 62, 51, 58, 23, 13, 26, 35, 42, 34, 
    97, 75, 77, 76, 79, 78, 73, 54, 70, 72, 40, 43, 30, 34, 40, 
    101, 80, 80, 78, 86, 78, 75, 65, 59, 72, 69, 57, 27, 26, 38, 
    69, 77, 85, 85, 84, 81, 79, 82, 69, 47, 70, 73, 22, 32, 36, 
    10, 95, 87, 94, 87, 96, 118, 75, 70, 50, 66, 52, 11, 26, 30, 
    9, 77, 115, 103, 94, 111, 109, 103, 83, 94, 83, 38, 12, 24, 26, 
    55, 43, 113, 97, 109, 132, 112, 115, 125, 122, 105, 41, 13, 44, 50, 
    61, 61, 116, 98, 89, 99, 108, 74, 74, 69, 54, 10, 0, 51, 81, 
    65, 57, 122, 105, 12, 85, 96, 63, 83, 27, 17, 14, 0, 56, 119, 
    74, 61, 105, 89, 1, 5, 11, 20, 38, 11, 0, 1, 11, 38, 123, 
    66, 66, 79, 97, 60, 37, 37, 37, 4, 0, 0, 0, 0, 20, 69, 
    57, 72, 76, 70, 85, 53, 45, 60, 39, 19, 10, 0, 0, 12, 28, 
    58, 48, 78, 56, 61, 50, 48, 67, 50, 50, 44, 43, 49, 36, 41, 
    58, 58, 68, 64, 71, 66, 56, 52, 51, 45, 45, 56, 64, 57, 42, 
    
    -- channel=173
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=174
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 8, 3, 0, 6, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 2, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=175
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 27, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 5, 10, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=176
    51, 55, 62, 61, 58, 53, 45, 48, 38, 24, 24, 21, 19, 38, 32, 
    94, 84, 64, 68, 66, 62, 53, 50, 30, 12, 23, 33, 42, 40, 31, 
    85, 77, 76, 77, 79, 74, 61, 58, 56, 35, 35, 36, 39, 40, 41, 
    86, 84, 81, 84, 89, 83, 74, 65, 68, 68, 58, 40, 26, 31, 43, 
    79, 83, 86, 85, 85, 83, 72, 68, 61, 67, 75, 51, 31, 40, 42, 
    52, 82, 84, 92, 84, 93, 105, 100, 71, 61, 64, 27, 21, 29, 38, 
    54, 104, 114, 100, 88, 123, 109, 67, 63, 83, 61, 18, 14, 23, 32, 
    46, 87, 113, 102, 121, 121, 106, 122, 129, 118, 75, 28, 21, 38, 30, 
    55, 93, 113, 96, 121, 119, 110, 105, 109, 105, 55, 0, 16, 71, 42, 
    57, 91, 130, 71, 73, 116, 81, 71, 57, 22, 0, 0, 20, 83, 58, 
    72, 93, 121, 37, 10, 39, 39, 63, 40, 7, 8, 5, 19, 90, 85, 
    71, 78, 89, 57, 32, 19, 31, 22, 0, 0, 0, 0, 12, 58, 78, 
    69, 74, 83, 95, 73, 57, 46, 31, 8, 0, 0, 0, 8, 14, 49, 
    68, 76, 78, 73, 61, 46, 68, 58, 40, 35, 24, 29, 26, 34, 36, 
    56, 73, 67, 66, 66, 67, 69, 62, 58, 48, 51, 60, 59, 47, 43, 
    
    -- channel=177
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 2, 0, 0, 0, 0, 4, 6, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 2, 1, 1, 3, 6, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 12, 6, 0, 25, 20, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 9, 12, 11, 15, 16, 6, 29, 31, 21, 0, 0, 0, 0, 0, 
    0, 15, 14, 7, 29, 23, 16, 27, 23, 27, 7, 0, 0, 12, 0, 
    3, 23, 23, 0, 13, 14, 2, 0, 0, 0, 0, 0, 0, 14, 0, 
    3, 21, 28, 0, 0, 8, 0, 26, 0, 0, 0, 0, 0, 25, 4, 
    5, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 6, 
    1, 11, 11, 15, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 5, 
    8, 10, 4, 3, 0, 0, 8, 1, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 0, 0, 0, 3, 8, 3, 2, 2, 0, 7, 2, 0, 0, 
    9, 17, 7, 11, 11, 8, 0, 0, 0, 0, 2, 5, 4, 0, 3, 
    
    -- channel=178
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 61, 41, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 0, 0, 31, 7, 0, 0, 0, 0, 
    0, 0, 0, 57, 0, 32, 39, 0, 43, 9, 11, 15, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 31, 22, 17, 7, 11, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=179
    34, 26, 24, 24, 26, 24, 25, 25, 18, 16, 15, 19, 19, 13, 15, 
    29, 28, 31, 27, 27, 28, 26, 26, 26, 17, 13, 10, 15, 16, 16, 
    21, 28, 31, 29, 30, 30, 31, 27, 28, 32, 20, 17, 10, 15, 18, 
    32, 24, 29, 30, 27, 32, 23, 28, 24, 26, 31, 19, 16, 16, 15, 
    25, 27, 30, 33, 30, 27, 25, 27, 19, 20, 26, 16, 15, 13, 16, 
    35, 32, 27, 26, 30, 37, 20, 2, 23, 21, 13, 15, 11, 15, 14, 
    11, 32, 24, 29, 38, 17, 29, 35, 23, 21, 16, 15, 15, 16, 12, 
    17, 22, 23, 24, 31, 26, 27, 21, 20, 25, 15, 10, 19, 22, 10, 
    14, 25, 22, 19, 17, 35, 11, 11, 14, 3, 6, 16, 19, 21, 14, 
    19, 20, 23, 9, 0, 16, 15, 23, 11, 21, 17, 7, 16, 23, 13, 
    13, 19, 16, 15, 20, 7, 13, 0, 7, 10, 4, 10, 14, 14, 14, 
    18, 16, 23, 28, 15, 21, 17, 14, 18, 12, 10, 7, 14, 7, 19, 
    18, 16, 19, 20, 21, 15, 19, 15, 18, 20, 15, 19, 11, 25, 6, 
    11, 17, 12, 25, 18, 21, 13, 17, 20, 15, 22, 19, 23, 16, 12, 
    19, 16, 19, 17, 24, 13, 15, 13, 15, 16, 16, 18, 18, 18, 20, 
    
    -- channel=180
    16, 9, 15, 14, 9, 9, 5, 5, 9, 3, 0, 0, 0, 7, 12, 
    32, 22, 16, 13, 10, 13, 13, 3, 0, 5, 0, 7, 6, 11, 6, 
    32, 8, 22, 17, 19, 17, 13, 15, 7, 4, 0, 16, 12, 7, 10, 
    36, 20, 20, 20, 25, 23, 23, 20, 18, 13, 18, 16, 0, 4, 10, 
    22, 20, 23, 21, 20, 24, 24, 18, 30, 15, 26, 23, 0, 8, 7, 
    0, 23, 19, 28, 30, 12, 48, 45, 23, 10, 28, 15, 0, 2, 5, 
    10, 23, 41, 30, 27, 39, 35, 12, 12, 31, 33, 10, 0, 0, 5, 
    17, 9, 41, 35, 32, 44, 46, 32, 48, 36, 42, 19, 0, 0, 24, 
    21, 16, 42, 55, 18, 35, 59, 31, 30, 43, 22, 0, 0, 2, 34, 
    20, 16, 46, 53, 0, 43, 40, 0, 38, 7, 0, 0, 0, 0, 35, 
    32, 27, 39, 19, 0, 7, 3, 13, 19, 3, 0, 0, 0, 8, 28, 
    27, 29, 17, 23, 11, 0, 11, 8, 0, 0, 0, 0, 0, 23, 0, 
    26, 21, 35, 22, 47, 20, 8, 14, 0, 0, 0, 0, 0, 0, 12, 
    29, 23, 35, 29, 14, 7, 17, 23, 9, 12, 1, 0, 4, 8, 0, 
    8, 25, 26, 24, 24, 21, 25, 21, 17, 17, 13, 14, 22, 15, 10, 
    
    -- channel=181
    3, 0, 13, 16, 16, 18, 19, 14, 9, 5, 9, 4, 7, 7, 6, 
    10, 12, 16, 15, 17, 15, 16, 17, 10, 2, 14, 16, 11, 8, 11, 
    7, 16, 12, 19, 16, 21, 16, 23, 18, 0, 0, 1, 16, 18, 8, 
    14, 10, 18, 17, 21, 23, 26, 18, 24, 22, 12, 9, 14, 14, 15, 
    14, 13, 15, 17, 20, 13, 12, 5, 12, 29, 20, 6, 14, 14, 14, 
    32, 6, 13, 13, 18, 5, 0, 23, 15, 10, 15, 16, 10, 12, 14, 
    1, 26, 11, 8, 6, 9, 19, 0, 0, 0, 2, 2, 3, 8, 12, 
    6, 19, 12, 15, 2, 4, 3, 9, 5, 0, 0, 0, 4, 0, 0, 
    16, 7, 6, 10, 19, 27, 20, 40, 34, 37, 38, 13, 6, 8, 0, 
    18, 20, 5, 2, 42, 14, 26, 2, 3, 14, 0, 0, 4, 8, 0, 
    17, 25, 17, 13, 0, 39, 37, 45, 37, 9, 13, 13, 1, 24, 0, 
    27, 16, 15, 0, 0, 0, 0, 3, 6, 4, 0, 5, 18, 25, 24, 
    18, 24, 15, 25, 0, 8, 18, 3, 0, 0, 0, 0, 0, 9, 23, 
    20, 33, 23, 16, 19, 11, 19, 18, 8, 0, 0, 0, 0, 0, 7, 
    25, 9, 21, 13, 5, 14, 21, 27, 19, 21, 16, 16, 12, 10, 9, 
    
    -- channel=182
    41, 15, 50, 54, 51, 46, 47, 38, 26, 23, 32, 23, 22, 29, 32, 
    59, 56, 54, 52, 57, 52, 48, 53, 35, 7, 30, 36, 42, 38, 33, 
    51, 58, 53, 62, 61, 61, 56, 50, 56, 23, 20, 29, 40, 47, 39, 
    56, 49, 61, 64, 63, 70, 66, 56, 61, 64, 47, 35, 40, 36, 43, 
    59, 57, 60, 60, 64, 65, 65, 57, 44, 69, 62, 38, 36, 40, 45, 
    64, 55, 57, 62, 60, 66, 49, 58, 64, 55, 51, 32, 24, 33, 40, 
    11, 84, 68, 67, 58, 58, 75, 48, 26, 35, 41, 22, 13, 25, 33, 
    33, 62, 74, 65, 71, 71, 60, 74, 69, 69, 38, 18, 21, 34, 15, 
    54, 62, 70, 49, 80, 88, 70, 76, 83, 73, 63, 18, 13, 50, 25, 
    64, 64, 79, 39, 67, 72, 75, 66, 29, 32, 11, 2, 18, 58, 26, 
    65, 69, 74, 46, 0, 39, 64, 64, 66, 16, 15, 29, 16, 63, 55, 
    76, 61, 68, 36, 17, 19, 15, 24, 3, 0, 0, 0, 30, 39, 76, 
    67, 74, 50, 76, 43, 55, 62, 32, 4, 0, 0, 0, 0, 28, 29, 
    63, 77, 67, 54, 62, 44, 60, 63, 40, 27, 20, 16, 14, 16, 39, 
    68, 57, 70, 57, 53, 56, 61, 70, 56, 55, 53, 57, 52, 45, 41, 
    
    -- channel=183
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=184
    62, 82, 58, 65, 62, 57, 50, 52, 40, 27, 33, 37, 39, 44, 33, 
    87, 78, 64, 71, 71, 68, 56, 58, 45, 24, 32, 32, 44, 41, 37, 
    75, 85, 76, 74, 78, 72, 68, 58, 62, 62, 59, 38, 35, 37, 45, 
    70, 79, 76, 80, 80, 72, 64, 59, 61, 65, 58, 44, 32, 41, 43, 
    61, 85, 82, 81, 82, 72, 70, 81, 56, 58, 64, 42, 38, 36, 43, 
    61, 79, 96, 84, 70, 104, 92, 62, 50, 63, 53, 19, 30, 33, 41, 
    68, 84, 95, 90, 92, 105, 82, 89, 97, 92, 50, 23, 30, 38, 34, 
    43, 84, 92, 79, 115, 108, 90, 107, 103, 103, 71, 24, 30, 65, 30, 
    51, 87, 99, 65, 107, 92, 78, 62, 69, 46, 11, 9, 36, 78, 40, 
    49, 87, 109, 46, 48, 81, 51, 89, 43, 17, 25, 21, 33, 91, 63, 
    58, 70, 89, 23, 35, 19, 23, 36, 8, 7, 9, 17, 34, 75, 74, 
    46, 69, 75, 82, 38, 48, 46, 21, 8, 6, 1, 5, 26, 37, 69, 
    60, 61, 69, 69, 63, 44, 55, 44, 32, 25, 21, 26, 27, 24, 49, 
    52, 56, 55, 57, 51, 57, 61, 49, 51, 47, 45, 57, 50, 50, 36, 
    57, 71, 57, 61, 64, 63, 52, 44, 46, 42, 51, 58, 55, 47, 51, 
    
    -- channel=185
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=186
    43, 55, 46, 50, 50, 51, 50, 44, 40, 28, 31, 35, 32, 33, 33, 
    43, 45, 46, 49, 52, 54, 57, 53, 55, 34, 28, 30, 35, 38, 32, 
    40, 39, 48, 48, 50, 52, 56, 51, 53, 52, 47, 43, 37, 34, 37, 
    29, 38, 44, 48, 48, 53, 50, 52, 45, 46, 48, 46, 35, 37, 34, 
    27, 40, 46, 48, 50, 51, 38, 46, 45, 40, 43, 41, 31, 33, 33, 
    14, 40, 46, 45, 44, 36, 35, 21, 29, 34, 37, 26, 27, 33, 32, 
    35, 25, 36, 39, 38, 35, 26, 39, 41, 35, 33, 27, 27, 35, 32, 
    39, 28, 34, 29, 32, 32, 45, 29, 25, 26, 40, 28, 20, 36, 36, 
    44, 33, 32, 34, 26, 18, 40, 24, 22, 16, 11, 21, 22, 28, 38, 
    42, 31, 23, 44, 0, 24, 27, 42, 48, 25, 27, 37, 25, 26, 39, 
    43, 30, 21, 29, 34, 10, 15, 24, 22, 26, 18, 21, 33, 18, 29, 
    32, 43, 24, 45, 43, 45, 46, 40, 25, 20, 20, 18, 18, 25, 20, 
    42, 37, 39, 21, 43, 37, 37, 47, 40, 35, 33, 30, 31, 26, 29, 
    41, 27, 38, 36, 30, 38, 37, 45, 40, 41, 42, 46, 46, 44, 31, 
    37, 47, 40, 43, 42, 43, 44, 36, 39, 38, 43, 41, 42, 43, 38, 
    
    -- channel=187
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=188
    50, 0, 6, 0, 6, 0, 14, 0, 32, 0, 0, 6, 0, 0, 25, 
    0, 14, 1, 0, 0, 2, 12, 1, 39, 12, 0, 0, 0, 9, 0, 
    29, 0, 0, 0, 0, 6, 16, 0, 9, 42, 0, 17, 0, 0, 0, 
    22, 0, 0, 0, 0, 4, 7, 7, 0, 2, 8, 34, 7, 0, 0, 
    4, 0, 0, 0, 0, 2, 6, 0, 17, 0, 0, 59, 0, 0, 0, 
    0, 9, 0, 0, 7, 0, 28, 0, 30, 0, 10, 49, 0, 0, 0, 
    0, 0, 1, 10, 0, 0, 29, 41, 0, 0, 50, 40, 0, 0, 0, 
    13, 0, 12, 0, 0, 16, 6, 0, 0, 8, 63, 37, 0, 0, 30, 
    12, 0, 1, 21, 0, 0, 35, 0, 0, 1, 65, 22, 0, 0, 86, 
    24, 0, 0, 109, 0, 0, 63, 0, 42, 26, 12, 10, 0, 0, 111, 
    18, 0, 0, 123, 0, 0, 3, 0, 55, 15, 0, 0, 0, 0, 86, 
    17, 0, 0, 37, 37, 8, 0, 31, 22, 3, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 33, 15, 0, 35, 32, 17, 17, 0, 0, 0, 0, 
    5, 0, 24, 0, 38, 0, 0, 33, 5, 16, 13, 0, 14, 0, 19, 
    0, 0, 15, 0, 9, 0, 0, 7, 4, 5, 0, 0, 7, 19, 0, 
    
    -- channel=189
    41, 23, 38, 43, 46, 44, 43, 38, 28, 18, 25, 22, 24, 21, 21, 
    40, 45, 44, 46, 48, 46, 43, 45, 38, 15, 25, 26, 29, 26, 27, 
    35, 49, 43, 50, 49, 51, 48, 48, 50, 24, 21, 19, 28, 34, 26, 
    43, 43, 47, 49, 51, 52, 51, 46, 48, 51, 41, 26, 29, 28, 30, 
    38, 42, 47, 51, 51, 45, 41, 39, 31, 48, 46, 27, 28, 29, 30, 
    50, 42, 47, 46, 49, 50, 19, 33, 38, 35, 32, 29, 22, 26, 29, 
    17, 54, 45, 43, 43, 41, 46, 25, 20, 23, 21, 14, 17, 24, 25, 
    26, 45, 43, 44, 43, 42, 37, 46, 38, 37, 16, 10, 21, 26, 12, 
    33, 42, 39, 29, 50, 54, 34, 55, 49, 41, 40, 21, 19, 36, 10, 
    39, 45, 39, 13, 53, 38, 41, 42, 22, 25, 11, 9, 19, 43, 10, 
    35, 46, 42, 28, 10, 32, 34, 45, 37, 15, 15, 24, 16, 45, 31, 
    43, 36, 45, 25, 19, 17, 14, 21, 12, 9, 3, 7, 27, 27, 53, 
    35, 46, 35, 47, 20, 27, 37, 25, 10, 4, 2, 5, 7, 21, 32, 
    33, 45, 39, 34, 36, 33, 36, 36, 30, 20, 22, 19, 18, 17, 29, 
    45, 29, 39, 35, 31, 36, 37, 41, 36, 34, 35, 39, 34, 32, 28, 
    
    -- channel=190
    45, 0, 24, 21, 29, 20, 25, 12, 31, 4, 7, 5, 6, 0, 22, 
    38, 42, 29, 27, 25, 28, 26, 17, 27, 4, 2, 9, 8, 14, 13, 
    40, 36, 27, 29, 30, 32, 31, 19, 32, 27, 0, 10, 8, 15, 10, 
    54, 25, 34, 29, 38, 33, 35, 25, 21, 31, 21, 29, 11, 4, 13, 
    24, 29, 34, 32, 38, 31, 31, 25, 25, 19, 28, 45, 10, 11, 13, 
    1, 28, 29, 35, 33, 34, 41, 40, 47, 11, 25, 38, 0, 10, 9, 
    0, 35, 47, 44, 30, 36, 62, 38, 7, 21, 39, 19, 0, 6, 7, 
    16, 0, 50, 38, 32, 54, 35, 44, 50, 48, 53, 23, 0, 3, 14, 
    27, 0, 45, 40, 45, 46, 59, 48, 51, 45, 63, 18, 0, 8, 48, 
    28, 0, 52, 67, 6, 27, 67, 12, 27, 18, 5, 0, 0, 1, 67, 
    33, 12, 51, 73, 0, 14, 27, 12, 52, 9, 5, 6, 0, 0, 80, 
    34, 17, 31, 45, 11, 0, 0, 9, 4, 0, 0, 0, 0, 0, 46, 
    17, 28, 22, 31, 43, 23, 17, 22, 6, 0, 0, 0, 0, 3, 5, 
    25, 18, 40, 13, 36, 16, 9, 32, 16, 9, 8, 0, 5, 0, 15, 
    29, 8, 31, 17, 22, 20, 22, 29, 20, 21, 12, 15, 20, 20, 8, 
    
    -- channel=191
    13, 40, 34, 41, 36, 41, 33, 39, 15, 29, 30, 25, 28, 34, 15, 
    33, 32, 38, 39, 40, 39, 38, 42, 19, 23, 38, 31, 33, 24, 27, 
    19, 42, 39, 41, 41, 40, 35, 47, 37, 13, 32, 23, 34, 32, 29, 
    20, 40, 38, 43, 42, 40, 37, 38, 45, 37, 31, 20, 30, 36, 32, 
    31, 38, 38, 42, 40, 37, 31, 32, 28, 49, 37, 8, 38, 32, 32, 
    69, 27, 40, 38, 36, 43, 9, 27, 21, 41, 26, 8, 38, 33, 36, 
    67, 47, 27, 26, 34, 39, 16, 2, 26, 28, 4, 8, 32, 34, 32, 
    21, 63, 22, 29, 40, 18, 27, 31, 20, 16, 0, 8, 35, 33, 12, 
    23, 54, 22, 18, 46, 37, 13, 43, 34, 29, 6, 17, 49, 46, 0, 
    21, 57, 20, 0, 63, 44, 5, 37, 9, 15, 17, 20, 44, 57, 0, 
    22, 49, 23, 0, 40, 38, 32, 55, 11, 24, 29, 30, 38, 67, 0, 
    25, 35, 28, 9, 15, 21, 26, 14, 17, 22, 17, 38, 45, 50, 27, 
    34, 31, 32, 33, 15, 28, 34, 12, 9, 14, 14, 23, 38, 29, 49, 
    26, 45, 19, 37, 14, 32, 41, 17, 24, 18, 20, 28, 20, 32, 20, 
    29, 35, 23, 31, 24, 30, 32, 31, 31, 28, 36, 36, 26, 22, 34, 
    
    -- channel=192
    142, 134, 140, 136, 127, 116, 116, 103, 99, 71, 77, 66, 9, 37, 58, 
    131, 118, 113, 110, 103, 94, 94, 87, 83, 77, 80, 32, 12, 49, 68, 
    88, 86, 90, 87, 87, 86, 86, 84, 82, 85, 42, 14, 34, 64, 64, 
    78, 83, 84, 83, 88, 89, 93, 89, 86, 73, 0, 29, 64, 70, 70, 
    81, 86, 86, 85, 91, 85, 81, 87, 94, 52, 3, 19, 55, 65, 69, 
    86, 86, 84, 83, 87, 86, 58, 35, 25, 24, 51, 0, 26, 46, 59, 
    87, 86, 78, 82, 59, 30, 2, 0, 8, 62, 56, 0, 0, 14, 38, 
    87, 83, 80, 44, 17, 28, 12, 45, 63, 55, 35, 0, 1, 14, 49, 
    83, 84, 18, 18, 0, 8, 46, 65, 36, 42, 18, 0, 49, 47, 38, 
    91, 97, 0, 7, 0, 8, 56, 36, 30, 0, 40, 30, 30, 20, 1, 
    85, 16, 0, 0, 0, 28, 49, 30, 0, 0, 0, 58, 5, 0, 0, 
    59, 10, 12, 0, 11, 18, 58, 26, 0, 8, 0, 26, 29, 0, 9, 
    44, 14, 16, 0, 36, 29, 40, 26, 0, 24, 0, 0, 24, 0, 12, 
    41, 17, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 2, 
    37, 12, 3, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 5, 
    
    -- channel=193
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 16, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 44, 48, 37, 36, 52, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 37, 0, 0, 0, 
    0, 0, 0, 0, 5, 1, 9, 10, 55, 65, 63, 58, 0, 0, 14, 
    0, 0, 0, 5, 10, 0, 14, 67, 59, 53, 39, 2, 0, 22, 50, 
    0, 19, 28, 0, 0, 0, 0, 53, 50, 49, 43, 43, 49, 42, 29, 
    0, 26, 15, 1, 0, 0, 20, 50, 38, 0, 0, 15, 35, 30, 0, 
    0, 0, 32, 10, 0, 16, 25, 57, 46, 0, 6, 0, 21, 20, 0, 
    0, 2, 29, 6, 20, 41, 45, 44, 38, 10, 15, 0, 12, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 4, 10, 4, 4, 2, 0, 0, 3, 0, 0, 0, 0, 0, 
    
    -- channel=194
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 8, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 23, 3, 0, 
    0, 0, 0, 0, 0, 0, 3, 8, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 45, 68, 60, 20, 8, 0, 0, 
    0, 0, 0, 0, 0, 17, 19, 0, 0, 0, 61, 88, 0, 21, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 156, 23, 0, 0, 
    0, 0, 3, 12, 0, 0, 15, 106, 122, 36, 0, 0, 48, 6, 54, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 30, 53, 0, 
    0, 21, 80, 0, 14, 0, 0, 0, 0, 0, 0, 99, 34, 0, 0, 
    0, 0, 33, 2, 12, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 32, 16, 0, 0, 0, 57, 6, 15, 0, 0, 18, 12, 
    0, 0, 0, 65, 30, 59, 0, 0, 83, 0, 52, 0, 0, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 2, 0, 
    0, 10, 32, 51, 25, 28, 22, 18, 15, 0, 0, 14, 6, 6, 3, 
    
    -- channel=195
    13, 10, 23, 15, 14, 12, 19, 6, 16, 24, 11, 3, 0, 22, 6, 
    16, 7, 16, 17, 18, 15, 19, 10, 12, 8, 9, 0, 0, 16, 7, 
    24, 25, 19, 16, 16, 14, 15, 11, 9, 10, 7, 0, 0, 17, 8, 
    16, 15, 14, 11, 14, 15, 14, 7, 6, 4, 0, 15, 17, 12, 9, 
    17, 16, 15, 15, 19, 14, 23, 21, 5, 0, 0, 0, 10, 9, 9, 
    16, 15, 14, 14, 21, 12, 4, 17, 52, 61, 24, 0, 22, 10, 9, 
    15, 16, 13, 19, 11, 49, 42, 17, 27, 33, 81, 0, 0, 35, 14, 
    17, 14, 11, 0, 4, 9, 5, 0, 0, 12, 46, 8, 0, 0, 9, 
    17, 18, 0, 24, 11, 20, 16, 70, 58, 58, 46, 0, 15, 0, 40, 
    19, 19, 0, 15, 0, 8, 48, 70, 43, 46, 84, 0, 13, 30, 24, 
    21, 87, 0, 1, 0, 5, 34, 52, 35, 4, 36, 115, 38, 29, 16, 
    27, 0, 38, 0, 0, 35, 56, 39, 0, 6, 0, 48, 49, 0, 0, 
    14, 16, 48, 0, 8, 6, 50, 36, 0, 22, 0, 0, 75, 0, 8, 
    9, 19, 41, 12, 60, 78, 80, 78, 23, 41, 14, 0, 30, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 25, 14, 0, 0, 0, 0, 
    
    -- channel=196
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 24, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 28, 6, 0, 0, 
    0, 0, 0, 0, 0, 6, 36, 43, 28, 17, 12, 38, 24, 9, 0, 
    0, 0, 0, 0, 18, 4, 15, 15, 10, 0, 20, 37, 12, 14, 0, 
    0, 0, 20, 28, 24, 21, 18, 0, 12, 24, 28, 50, 11, 10, 0, 
    0, 0, 36, 24, 28, 13, 3, 23, 30, 29, 11, 12, 13, 23, 23, 
    0, 19, 38, 24, 23, 15, 13, 26, 36, 50, 34, 21, 33, 32, 34, 
    0, 27, 22, 30, 16, 15, 13, 24, 47, 19, 25, 13, 26, 40, 13, 
    5, 22, 23, 38, 18, 23, 18, 35, 50, 14, 25, 21, 14, 38, 7, 
    0, 12, 19, 24, 21, 32, 36, 38, 40, 11, 33, 29, 20, 24, 10, 
    0, 21, 33, 26, 23, 23, 21, 21, 19, 15, 18, 22, 13, 12, 10, 
    
    -- channel=197
    0, 0, 7, 16, 15, 11, 7, 6, 0, 0, 0, 0, 0, 0, 0, 
    13, 7, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=198
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 21, 0, 
    0, 0, 0, 0, 0, 0, 6, 9, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 47, 71, 54, 38, 2, 0, 0, 
    0, 0, 0, 0, 0, 39, 85, 36, 0, 0, 84, 35, 0, 3, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 5, 18, 47, 19, 0, 0, 
    0, 0, 16, 30, 0, 7, 0, 107, 201, 156, 9, 0, 0, 8, 82, 
    0, 0, 0, 0, 0, 0, 13, 63, 0, 0, 0, 0, 49, 121, 48, 
    0, 106, 27, 0, 0, 0, 4, 0, 0, 0, 0, 80, 87, 11, 0, 
    0, 0, 0, 0, 0, 43, 53, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 15, 14, 2, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 23, 81, 96, 40, 0, 0, 19, 37, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 22, 53, 30, 33, 26, 14, 8, 0, 0, 0, 5, 6, 11, 
    
    -- channel=199
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 18, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 8, 0, 
    0, 0, 0, 0, 1, 0, 0, 1, 0, 5, 0, 0, 1, 1, 0, 
    2, 1, 0, 0, 0, 1, 6, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 6, 14, 27, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 39, 15, 0, 0, 14, 30, 0, 31, 0, 0, 
    0, 0, 0, 12, 1, 0, 0, 0, 3, 76, 41, 0, 0, 19, 0, 
    0, 0, 29, 0, 0, 7, 4, 45, 54, 0, 0, 0, 0, 19, 32, 
    0, 21, 0, 21, 0, 10, 62, 31, 0, 0, 0, 0, 46, 15, 14, 
    26, 49, 0, 4, 0, 12, 54, 11, 0, 0, 37, 0, 0, 0, 0, 
    16, 15, 0, 0, 0, 44, 40, 1, 0, 0, 0, 88, 0, 0, 0, 
    10, 0, 24, 0, 20, 22, 50, 0, 0, 3, 0, 23, 21, 0, 0, 
    12, 12, 31, 0, 48, 19, 13, 0, 0, 35, 0, 0, 36, 0, 5, 
    3, 8, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 8, 0, 4, 
    4, 0, 16, 0, 3, 5, 0, 0, 0, 19, 0, 0, 3, 3, 11, 
    
    -- channel=200
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 11, 
    0, 0, 0, 0, 1, 0, 1, 3, 9, 0, 0, 4, 18, 17, 8, 
    
    -- channel=201
    112, 127, 135, 142, 136, 129, 123, 114, 108, 84, 75, 59, 41, 16, 49, 
    137, 123, 126, 130, 120, 108, 104, 96, 88, 78, 67, 52, 0, 19, 63, 
    102, 103, 102, 101, 93, 87, 87, 81, 77, 71, 44, 0, 7, 34, 59, 
    80, 83, 83, 83, 83, 83, 81, 79, 70, 65, 17, 0, 34, 67, 69, 
    76, 85, 86, 85, 84, 77, 60, 62, 48, 39, 0, 0, 51, 68, 67, 
    83, 86, 85, 84, 76, 43, 0, 0, 0, 0, 0, 0, 2, 31, 61, 
    86, 85, 86, 72, 52, 19, 0, 3, 1, 0, 0, 0, 2, 0, 35, 
    85, 85, 56, 40, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 67, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    71, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    18, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=202
    0, 0, 4, 12, 15, 15, 15, 9, 13, 34, 3, 0, 26, 16, 0, 
    8, 0, 10, 16, 16, 11, 9, 6, 1, 0, 0, 0, 0, 0, 0, 
    32, 32, 17, 9, 3, 0, 0, 0, 0, 0, 7, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 7, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 66, 79, 0, 0, 38, 0, 0, 
    0, 0, 0, 0, 0, 56, 68, 72, 46, 0, 0, 0, 0, 40, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 
    0, 0, 7, 30, 25, 29, 0, 0, 9, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 10, 18, 5, 5, 0, 77, 87, 0, 0, 0, 22, 
    13, 113, 4, 0, 5, 0, 0, 0, 40, 63, 68, 104, 27, 43, 74, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 15, 19, 0, 
    10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 62, 27, 10, 
    0, 16, 55, 59, 102, 149, 161, 163, 90, 14, 15, 3, 46, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 34, 7, 0, 0, 0, 
    
    -- channel=203
    47, 42, 44, 40, 38, 33, 34, 29, 25, 20, 23, 16, 12, 0, 16, 
    32, 28, 27, 25, 23, 20, 23, 21, 19, 20, 16, 14, 3, 9, 16, 
    20, 15, 14, 17, 18, 16, 19, 21, 22, 16, 20, 0, 5, 22, 19, 
    15, 14, 14, 15, 17, 18, 18, 19, 21, 17, 12, 0, 13, 18, 18, 
    15, 14, 13, 14, 15, 20, 17, 11, 0, 9, 0, 0, 13, 15, 16, 
    15, 13, 14, 16, 12, 2, 7, 0, 0, 0, 0, 0, 0, 9, 11, 
    14, 13, 16, 10, 14, 0, 0, 0, 1, 0, 6, 0, 0, 10, 4, 
    12, 13, 6, 5, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 3, 
    12, 5, 2, 0, 3, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    1, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    14, 0, 9, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 7, 
    8, 5, 9, 0, 2, 0, 0, 0, 0, 3, 0, 0, 15, 0, 6, 
    6, 0, 0, 1, 0, 0, 1, 1, 3, 9, 0, 0, 8, 7, 6, 
    
    -- channel=204
    21, 19, 13, 15, 15, 6, 3, 6, 0, 11, 6, 0, 4, 0, 0, 
    12, 18, 6, 0, 0, 0, 0, 0, 0, 0, 0, 18, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 33, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 12, 16, 37, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 4, 15, 29, 54, 86, 67, 7, 3, 0, 0, 
    0, 0, 0, 0, 0, 37, 77, 96, 94, 109, 143, 109, 0, 18, 0, 
    0, 0, 0, 0, 15, 42, 60, 30, 7, 24, 147, 187, 19, 0, 0, 
    0, 0, 4, 36, 52, 29, 57, 67, 106, 142, 199, 169, 51, 0, 30, 
    0, 1, 31, 34, 46, 8, 39, 137, 195, 205, 200, 124, 33, 69, 111, 
    0, 68, 127, 21, 25, 0, 29, 160, 179, 158, 130, 170, 134, 140, 120, 
    0, 77, 107, 28, 0, 6, 55, 165, 156, 72, 13, 49, 156, 120, 67, 
    0, 38, 68, 46, 0, 29, 89, 181, 165, 14, 22, 3, 99, 97, 0, 
    0, 31, 63, 66, 45, 112, 127, 174, 156, 25, 61, 9, 28, 55, 0, 
    0, 15, 35, 25, 13, 34, 43, 49, 52, 10, 46, 12, 0, 0, 0, 
    6, 23, 29, 27, 7, 10, 9, 3, 0, 0, 15, 2, 0, 0, 0, 
    
    -- channel=205
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 15, 25, 30, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 15, 0, 26, 63, 12, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 13, 22, 49, 66, 39, 0, 1, 0, 
    0, 0, 0, 14, 18, 15, 28, 49, 57, 57, 46, 0, 0, 11, 35, 
    0, 0, 21, 23, 7, 11, 41, 64, 63, 57, 48, 29, 46, 48, 33, 
    0, 37, 27, 18, 0, 17, 55, 63, 51, 21, 29, 52, 55, 43, 14, 
    0, 15, 37, 16, 9, 38, 56, 63, 33, 11, 9, 34, 43, 28, 0, 
    0, 17, 43, 23, 35, 48, 63, 62, 28, 23, 16, 13, 36, 11, 0, 
    0, 2, 32, 24, 40, 42, 42, 42, 17, 22, 21, 5, 14, 0, 0, 
    0, 0, 20, 17, 18, 18, 14, 10, 4, 17, 11, 0, 0, 0, 1, 
    
    -- channel=206
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 24, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 22, 13, 20, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 2, 12, 12, 0, 24, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 6, 0, 0, 0, 25, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=207
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 23, 0, 11, 4, 0, 0, 
    0, 0, 0, 0, 0, 12, 43, 49, 28, 0, 35, 0, 16, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 57, 1, 0, 0, 
    0, 0, 0, 16, 29, 23, 2, 17, 39, 35, 43, 10, 0, 0, 7, 
    0, 0, 7, 24, 21, 21, 18, 43, 41, 81, 43, 0, 0, 26, 46, 
    0, 55, 28, 28, 11, 0, 23, 40, 77, 40, 64, 63, 51, 59, 42, 
    0, 17, 27, 19, 0, 29, 26, 37, 38, 12, 13, 42, 35, 43, 2, 
    0, 16, 30, 5, 0, 0, 33, 40, 29, 7, 6, 24, 52, 29, 5, 
    0, 16, 54, 49, 74, 91, 95, 95, 49, 26, 26, 21, 36, 16, 6, 
    0, 0, 3, 5, 8, 6, 9, 10, 8, 29, 30, 9, 6, 5, 3, 
    
    -- channel=208
    34, 32, 31, 29, 23, 17, 16, 10, 13, 21, 5, 5, 4, 0, 0, 
    22, 20, 16, 9, 6, 3, 3, 1, 0, 0, 0, 0, 0, 0, 0, 
    22, 15, 4, 0, 0, 0, 0, 0, 0, 1, 36, 17, 0, 6, 3, 
    0, 0, 0, 0, 0, 3, 6, 7, 8, 18, 17, 8, 16, 10, 0, 
    0, 0, 1, 2, 4, 15, 29, 28, 28, 28, 9, 8, 2, 0, 0, 
    0, 0, 1, 0, 7, 26, 75, 114, 153, 143, 119, 39, 13, 8, 0, 
    0, 3, 1, 0, 34, 77, 82, 44, 22, 53, 175, 88, 0, 10, 0, 
    4, 3, 9, 27, 33, 35, 33, 6, 27, 139, 209, 149, 29, 0, 14, 
    4, 7, 28, 44, 36, 21, 53, 174, 225, 225, 201, 62, 10, 44, 116, 
    0, 69, 59, 29, 5, 7, 93, 187, 198, 204, 195, 132, 117, 141, 136, 
    39, 136, 84, 21, 0, 0, 92, 180, 172, 66, 60, 148, 173, 140, 62, 
    14, 41, 64, 10, 0, 48, 136, 191, 98, 10, 0, 62, 124, 65, 0, 
    0, 37, 69, 17, 27, 75, 146, 182, 85, 27, 22, 15, 82, 28, 0, 
    0, 34, 69, 53, 83, 118, 132, 134, 64, 43, 36, 0, 0, 0, 0, 
    5, 6, 0, 0, 0, 0, 0, 0, 0, 10, 29, 0, 0, 0, 0, 
    
    -- channel=209
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 31, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 40, 24, 8, 8, 72, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 32, 76, 40, 0, 0, 0, 
    0, 0, 0, 8, 0, 2, 5, 49, 83, 103, 80, 9, 0, 0, 28, 
    0, 0, 0, 0, 0, 0, 20, 84, 69, 73, 62, 0, 27, 50, 50, 
    2, 65, 7, 0, 0, 0, 38, 65, 67, 24, 33, 72, 69, 50, 19, 
    5, 0, 8, 0, 0, 12, 54, 65, 24, 0, 0, 31, 41, 11, 0, 
    0, 4, 21, 0, 0, 19, 60, 69, 1, 0, 0, 0, 37, 0, 0, 
    0, 4, 23, 5, 43, 65, 74, 66, 8, 13, 6, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=210
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 47, 79, 58, 18, 0, 22, 0, 18, 4, 
    0, 0, 0, 0, 8, 0, 12, 21, 0, 0, 0, 0, 30, 17, 0, 
    0, 0, 0, 23, 15, 29, 7, 0, 0, 0, 0, 92, 2, 0, 0, 
    0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    0, 0, 56, 0, 42, 6, 0, 0, 0, 130, 7, 11, 0, 0, 88, 
    0, 7, 0, 22, 9, 0, 0, 0, 43, 7, 11, 0, 7, 29, 32, 
    0, 0, 0, 34, 0, 0, 0, 0, 33, 0, 0, 0, 0, 76, 10, 
    0, 0, 0, 24, 2, 45, 54, 63, 108, 0, 42, 21, 25, 52, 9, 
    0, 11, 29, 0, 1, 1, 0, 8, 14, 0, 7, 48, 12, 11, 6, 
    
    -- channel=211
    31, 33, 33, 36, 34, 30, 28, 27, 21, 14, 17, 17, 2, 10, 15, 
    32, 28, 24, 23, 19, 19, 18, 20, 17, 17, 26, 8, 12, 14, 13, 
    17, 16, 16, 14, 16, 16, 17, 19, 19, 20, 7, 13, 14, 14, 14, 
    14, 14, 15, 16, 15, 15, 16, 20, 19, 20, 1, 13, 16, 17, 13, 
    12, 13, 13, 13, 14, 13, 15, 20, 34, 18, 11, 10, 7, 8, 13, 
    13, 13, 13, 12, 18, 26, 8, 0, 0, 2, 29, 7, 10, 9, 9, 
    13, 11, 10, 16, 4, 4, 2, 2, 5, 33, 0, 26, 5, 1, 5, 
    12, 13, 19, 5, 5, 8, 12, 48, 38, 15, 10, 0, 19, 21, 24, 
    11, 23, 6, 7, 0, 15, 26, 3, 4, 12, 5, 15, 14, 17, 4, 
    23, 20, 3, 3, 6, 3, 25, 1, 10, 0, 3, 31, 6, 5, 0, 
    13, 0, 11, 0, 13, 25, 16, 7, 0, 17, 0, 0, 1, 0, 1, 
    5, 16, 0, 3, 17, 0, 20, 7, 0, 12, 5, 1, 10, 0, 15, 
    6, 7, 0, 19, 22, 18, 7, 12, 2, 12, 8, 4, 0, 7, 6, 
    6, 0, 0, 1, 0, 0, 0, 0, 0, 9, 5, 4, 0, 11, 9, 
    5, 12, 15, 7, 9, 9, 7, 7, 7, 0, 0, 13, 8, 10, 12, 
    
    -- channel=212
    0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    1, 3, 7, 2, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    7, 5, 2, 0, 0, 0, 0, 0, 0, 0, 8, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 3, 1, 0, 18, 10, 9, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 35, 74, 81, 59, 21, 79, 0, 10, 0, 
    0, 2, 1, 0, 15, 30, 23, 21, 0, 0, 49, 75, 20, 0, 0, 
    2, 2, 0, 25, 17, 8, 3, 0, 0, 56, 91, 99, 24, 0, 0, 
    4, 0, 24, 12, 18, 0, 8, 48, 102, 93, 90, 63, 0, 23, 41, 
    0, 10, 68, 8, 15, 0, 16, 66, 88, 117, 66, 74, 62, 67, 74, 
    18, 48, 38, 14, 0, 0, 25, 70, 92, 39, 21, 11, 86, 74, 38, 
    0, 19, 0, 22, 0, 0, 34, 87, 73, 0, 0, 13, 32, 52, 0, 
    0, 4, 2, 25, 0, 21, 49, 80, 76, 0, 19, 16, 0, 34, 0, 
    0, 2, 19, 27, 23, 38, 46, 50, 23, 0, 9, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    
    -- channel=213
    49, 59, 70, 73, 70, 65, 64, 58, 56, 55, 46, 26, 8, 26, 26, 
    68, 59, 62, 65, 62, 55, 53, 48, 44, 40, 22, 18, 8, 5, 28, 
    56, 62, 57, 53, 49, 44, 43, 41, 36, 32, 5, 2, 3, 10, 27, 
    44, 43, 41, 40, 41, 40, 37, 31, 31, 22, 12, 18, 25, 33, 38, 
    38, 42, 44, 43, 41, 34, 27, 26, 4, 0, 0, 0, 18, 36, 33, 
    40, 42, 41, 42, 32, 10, 0, 0, 6, 19, 0, 0, 16, 10, 31, 
    42, 43, 41, 33, 17, 26, 30, 35, 26, 0, 0, 0, 0, 12, 21, 
    44, 40, 20, 0, 7, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    43, 26, 8, 16, 0, 2, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 13, 25, 0, 0, 0, 1, 
    35, 34, 0, 0, 0, 0, 0, 0, 1, 29, 24, 45, 0, 9, 24, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 1, 0, 2, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 3, 1, 
    14, 5, 7, 11, 25, 52, 58, 61, 35, 0, 2, 0, 12, 4, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 0, 0, 0, 
    
    -- channel=214
    73, 83, 93, 93, 91, 84, 83, 76, 73, 62, 55, 44, 23, 32, 34, 
    98, 87, 86, 89, 85, 76, 72, 66, 60, 52, 47, 26, 7, 8, 39, 
    82, 85, 79, 73, 66, 63, 61, 56, 52, 52, 40, 31, 9, 23, 44, 
    59, 59, 59, 57, 59, 61, 63, 56, 54, 50, 20, 14, 36, 46, 50, 
    54, 60, 62, 62, 65, 62, 61, 68, 62, 31, 1, 0, 40, 48, 45, 
    60, 63, 61, 61, 65, 58, 44, 57, 80, 102, 59, 0, 26, 36, 41, 
    63, 64, 61, 61, 50, 64, 62, 38, 35, 41, 72, 45, 0, 27, 33, 
    65, 65, 58, 38, 29, 26, 22, 3, 0, 13, 88, 67, 26, 0, 11, 
    66, 67, 26, 43, 15, 14, 29, 64, 100, 118, 99, 48, 26, 5, 41, 
    71, 58, 7, 11, 0, 0, 46, 85, 95, 84, 129, 72, 36, 57, 57, 
    67, 82, 57, 0, 0, 0, 17, 81, 68, 60, 21, 112, 85, 61, 47, 
    54, 24, 30, 0, 0, 6, 62, 79, 39, 7, 0, 16, 77, 23, 6, 
    38, 21, 31, 0, 0, 13, 43, 85, 31, 13, 0, 0, 48, 21, 0, 
    23, 22, 25, 28, 37, 75, 88, 93, 68, 24, 28, 0, 0, 0, 0, 
    26, 11, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 
    
    -- channel=215
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 7, 20, 32, 27, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 25, 26, 23, 25, 0, 0, 0, 24, 
    0, 0, 5, 0, 0, 0, 0, 29, 21, 14, 22, 19, 24, 22, 0, 
    0, 12, 7, 0, 0, 0, 4, 31, 13, 0, 0, 6, 24, 4, 2, 
    0, 0, 20, 4, 0, 8, 10, 31, 30, 0, 0, 0, 10, 17, 0, 
    0, 0, 24, 5, 10, 29, 26, 22, 15, 6, 0, 0, 2, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=216
    38, 28, 28, 23, 17, 12, 14, 9, 8, 8, 11, 4, 0, 11, 5, 
    19, 22, 7, 1, 0, 0, 3, 2, 2, 6, 18, 7, 9, 20, 3, 
    8, 0, 0, 0, 0, 4, 3, 9, 10, 10, 37, 19, 18, 29, 8, 
    0, 0, 2, 2, 5, 6, 14, 20, 25, 23, 10, 21, 23, 7, 1, 
    1, 0, 0, 1, 5, 17, 30, 32, 61, 72, 46, 26, 10, 1, 3, 
    1, 0, 1, 1, 10, 53, 93, 81, 73, 63, 146, 27, 14, 21, 0, 
    1, 1, 0, 5, 36, 33, 44, 10, 17, 71, 158, 94, 9, 11, 0, 
    2, 1, 18, 32, 33, 41, 40, 91, 137, 178, 160, 70, 30, 13, 78, 
    0, 13, 27, 38, 22, 26, 63, 168, 152, 156, 144, 31, 44, 93, 106, 
    4, 120, 44, 33, 2, 15, 83, 143, 144, 99, 98, 123, 121, 113, 87, 
    24, 47, 63, 26, 0, 45, 107, 138, 104, 14, 32, 95, 105, 81, 2, 
    7, 43, 77, 11, 23, 65, 127, 142, 53, 34, 21, 38, 99, 29, 11, 
    3, 41, 74, 32, 83, 116, 142, 141, 59, 48, 45, 17, 61, 0, 2, 
    11, 28, 35, 14, 25, 27, 31, 30, 7, 48, 30, 4, 2, 0, 0, 
    15, 20, 33, 34, 18, 23, 20, 14, 7, 15, 16, 0, 0, 1, 10, 
    
    -- channel=217
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=218
    107, 103, 102, 101, 96, 89, 86, 83, 75, 50, 60, 58, 35, 17, 54, 
    93, 89, 86, 83, 79, 73, 73, 71, 66, 65, 57, 51, 24, 34, 59, 
    65, 62, 66, 68, 66, 65, 68, 68, 67, 64, 46, 15, 34, 51, 60, 
    58, 63, 64, 66, 66, 67, 68, 71, 68, 63, 22, 10, 48, 58, 58, 
    60, 65, 64, 66, 64, 66, 53, 53, 53, 60, 25, 24, 48, 54, 56, 
    64, 65, 65, 64, 57, 48, 38, 25, 6, 0, 9, 36, 7, 40, 51, 
    65, 64, 65, 55, 50, 9, 0, 0, 3, 0, 0, 28, 23, 10, 31, 
    62, 64, 52, 45, 18, 16, 12, 21, 35, 27, 0, 0, 20, 16, 28, 
    63, 55, 32, 0, 5, 3, 0, 3, 0, 0, 0, 5, 19, 29, 5, 
    55, 47, 19, 3, 10, 8, 0, 0, 0, 0, 0, 12, 13, 0, 1, 
    49, 0, 0, 12, 13, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 7, 0, 12, 14, 2, 0, 0, 2, 11, 13, 0, 0, 2, 17, 
    34, 5, 0, 8, 7, 7, 0, 0, 10, 2, 19, 15, 0, 1, 18, 
    34, 14, 0, 0, 0, 0, 0, 0, 0, 2, 0, 17, 2, 11, 19, 
    30, 20, 8, 20, 12, 13, 14, 15, 18, 2, 6, 14, 19, 19, 18, 
    
    -- channel=219
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=220
    0, 9, 0, 2, 9, 5, 0, 15, 0, 0, 9, 6, 13, 0, 12, 
    0, 7, 11, 6, 4, 6, 0, 7, 2, 9, 0, 13, 32, 0, 9, 
    0, 10, 7, 7, 1, 3, 3, 2, 4, 0, 0, 40, 10, 0, 14, 
    1, 0, 1, 6, 0, 1, 0, 0, 0, 0, 37, 0, 6, 4, 13, 
    0, 1, 1, 4, 0, 0, 0, 0, 0, 11, 43, 0, 4, 7, 3, 
    1, 3, 4, 3, 0, 0, 0, 0, 0, 11, 0, 121, 0, 17, 3, 
    0, 4, 10, 0, 0, 0, 7, 28, 2, 0, 0, 195, 22, 0, 5, 
    1, 8, 0, 0, 1, 0, 23, 0, 0, 0, 0, 131, 81, 0, 0, 
    4, 0, 0, 0, 41, 0, 0, 0, 0, 0, 41, 154, 0, 0, 0, 
    0, 0, 117, 0, 59, 0, 0, 0, 0, 10, 0, 65, 0, 0, 12, 
    0, 0, 94, 17, 34, 0, 0, 0, 45, 83, 0, 0, 27, 17, 93, 
    0, 0, 0, 66, 0, 0, 0, 0, 169, 0, 18, 0, 0, 107, 20, 
    0, 0, 0, 68, 0, 0, 0, 0, 168, 0, 37, 0, 0, 113, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 90, 0, 36, 46, 0, 31, 0, 
    0, 7, 3, 16, 0, 0, 2, 6, 8, 0, 17, 42, 0, 0, 0, 
    
    -- channel=221
    75, 81, 91, 93, 89, 80, 79, 71, 63, 67, 56, 36, 15, 25, 31, 
    86, 76, 72, 71, 67, 61, 59, 56, 51, 48, 42, 26, 17, 12, 34, 
    61, 61, 55, 54, 52, 48, 48, 50, 46, 44, 24, 15, 15, 20, 35, 
    45, 45, 45, 45, 46, 47, 48, 48, 46, 36, 26, 17, 29, 41, 43, 
    39, 44, 45, 46, 46, 45, 45, 48, 43, 21, 3, 0, 24, 39, 38, 
    42, 44, 44, 46, 43, 42, 10, 4, 17, 37, 12, 0, 19, 19, 33, 
    45, 44, 43, 42, 26, 32, 31, 20, 23, 24, 24, 0, 0, 11, 19, 
    45, 43, 38, 12, 24, 9, 12, 4, 0, 0, 14, 3, 0, 3, 1, 
    42, 42, 16, 21, 4, 11, 17, 10, 19, 32, 19, 12, 14, 0, 6, 
    43, 25, 0, 1, 0, 2, 9, 24, 18, 8, 41, 0, 0, 5, 8, 
    37, 39, 9, 0, 0, 3, 0, 17, 3, 24, 11, 49, 11, 11, 19, 
    38, 4, 11, 0, 0, 0, 16, 10, 0, 0, 0, 10, 22, 0, 5, 
    28, 8, 12, 0, 0, 0, 4, 16, 0, 4, 0, 0, 26, 0, 5, 
    19, 12, 8, 3, 14, 31, 35, 36, 24, 9, 9, 0, 12, 2, 0, 
    15, 9, 0, 0, 0, 0, 0, 0, 0, 7, 1, 2, 0, 0, 0, 
    
    -- channel=222
    4, 13, 12, 13, 15, 10, 8, 12, 2, 18, 13, 0, 0, 3, 0, 
    9, 13, 7, 5, 5, 3, 0, 3, 0, 0, 0, 2, 16, 0, 0, 
    8, 12, 4, 1, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 26, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 12, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 23, 39, 69, 47, 29, 0, 8, 0, 
    0, 0, 0, 0, 0, 14, 47, 43, 25, 0, 24, 103, 0, 1, 0, 
    0, 0, 0, 0, 27, 4, 16, 0, 0, 0, 66, 111, 44, 0, 0, 
    0, 0, 0, 24, 23, 0, 0, 10, 64, 87, 86, 89, 0, 0, 9, 
    0, 0, 51, 0, 20, 0, 0, 52, 72, 79, 84, 66, 10, 42, 59, 
    0, 30, 88, 8, 6, 0, 0, 56, 88, 78, 2, 33, 75, 73, 66, 
    0, 13, 30, 20, 0, 0, 5, 60, 107, 0, 8, 0, 54, 60, 8, 
    0, 2, 15, 18, 0, 2, 0, 66, 100, 0, 16, 0, 15, 58, 0, 
    0, 0, 21, 32, 14, 51, 61, 70, 88, 0, 28, 8, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 13, 0, 0, 0, 
    
    -- channel=223
    73, 74, 83, 81, 73, 70, 72, 62, 65, 51, 50, 37, 23, 43, 36, 
    76, 66, 66, 64, 62, 57, 59, 53, 53, 48, 46, 28, 12, 43, 41, 
    60, 53, 54, 52, 54, 50, 49, 51, 47, 47, 36, 10, 27, 42, 37, 
    48, 49, 49, 47, 50, 48, 51, 47, 48, 41, 9, 40, 35, 42, 42, 
    47, 48, 49, 47, 50, 47, 51, 43, 40, 13, 0, 24, 40, 44, 45, 
    47, 47, 47, 48, 47, 42, 27, 21, 28, 4, 0, 0, 39, 29, 42, 
    49, 47, 42, 44, 44, 36, 10, 7, 19, 50, 28, 0, 5, 26, 36, 
    48, 42, 41, 28, 19, 25, 5, 5, 11, 24, 0, 0, 0, 18, 26, 
    44, 39, 26, 19, 0, 26, 37, 31, 2, 0, 0, 0, 16, 21, 13, 
    39, 49, 0, 19, 0, 32, 56, 10, 0, 0, 10, 0, 2, 0, 0, 
    58, 30, 0, 4, 5, 29, 51, 0, 0, 0, 37, 51, 0, 0, 0, 
    42, 11, 5, 0, 20, 34, 40, 0, 0, 14, 4, 58, 6, 0, 13, 
    38, 15, 13, 0, 25, 0, 23, 0, 0, 23, 0, 19, 41, 0, 30, 
    33, 22, 17, 6, 36, 27, 25, 20, 0, 36, 0, 0, 33, 7, 25, 
    26, 12, 6, 0, 10, 11, 11, 12, 13, 40, 8, 4, 20, 21, 25, 
    
    -- channel=224
    11, 8, 18, 11, 16, 22, 10, 12, 7, 6, 5, 2, 3, 8, 6, 
    10, 8, 14, 11, 14, 21, 20, 18, 12, 14, 17, 19, 20, 21, 17, 
    8, 10, 2, 13, 11, 19, 22, 31, 33, 26, 23, 25, 22, 17, 15, 
    11, 15, 10, 5, 15, 21, 26, 31, 31, 30, 26, 22, 25, 19, 24, 
    35, 37, 9, 2, 13, 32, 27, 19, 30, 30, 32, 32, 38, 38, 38, 
    37, 32, 9, 0, 20, 34, 14, 18, 29, 28, 26, 33, 43, 46, 35, 
    28, 29, 29, 0, 13, 27, 18, 26, 28, 20, 22, 31, 30, 35, 18, 
    33, 38, 28, 34, 15, 32, 23, 31, 30, 16, 19, 22, 26, 28, 29, 
    43, 56, 58, 23, 44, 20, 40, 21, 26, 17, 19, 17, 27, 25, 24, 
    62, 58, 31, 15, 33, 19, 34, 21, 24, 22, 22, 14, 22, 20, 31, 
    53, 36, 0, 16, 15, 15, 25, 25, 27, 24, 23, 20, 25, 37, 29, 
    13, 15, 15, 16, 0, 16, 32, 3, 19, 26, 26, 23, 25, 46, 29, 
    14, 16, 22, 25, 19, 15, 25, 18, 18, 33, 20, 16, 28, 39, 44, 
    22, 24, 21, 22, 32, 34, 26, 25, 24, 21, 20, 18, 22, 39, 41, 
    17, 23, 32, 31, 41, 40, 30, 34, 35, 31, 31, 30, 30, 38, 38, 
    
    -- channel=225
    24, 22, 19, 21, 26, 29, 26, 18, 17, 16, 12, 9, 6, 2, 3, 
    23, 22, 19, 17, 32, 36, 35, 29, 15, 14, 14, 15, 18, 17, 15, 
    21, 21, 18, 9, 31, 35, 37, 38, 32, 30, 28, 24, 18, 13, 7, 
    20, 20, 14, 18, 33, 37, 39, 44, 32, 32, 32, 25, 11, 13, 11, 
    36, 48, 50, 18, 37, 43, 51, 46, 45, 40, 41, 37, 20, 16, 17, 
    43, 43, 48, 20, 32, 45, 51, 46, 46, 46, 44, 42, 25, 14, 14, 
    35, 33, 42, 14, 27, 33, 45, 48, 49, 46, 46, 44, 30, 13, 9, 
    36, 39, 43, 46, 31, 31, 42, 46, 53, 53, 49, 43, 38, 19, 13, 
    43, 43, 60, 59, 54, 37, 38, 45, 52, 54, 52, 51, 45, 28, 1, 
    73, 73, 67, 56, 56, 54, 41, 42, 53, 54, 55, 55, 42, 13, 0, 
    66, 64, 23, 36, 37, 39, 33, 34, 49, 51, 43, 46, 37, 16, 3, 
    37, 24, 27, 38, 32, 35, 42, 17, 30, 42, 47, 47, 26, 13, 4, 
    24, 20, 20, 24, 34, 31, 29, 32, 40, 48, 56, 53, 27, 6, 12, 
    19, 23, 22, 8, 0, 14, 15, 28, 26, 27, 38, 42, 37, 3, 2, 
    13, 0, 0, 0, 0, 9, 12, 5, 1, 7, 11, 14, 9, 0, 0, 
    
    -- channel=226
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 24, 26, 23, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 9, 4, 0, 0, 0, 
    0, 1, 42, 0, 0, 3, 4, 0, 0, 0, 0, 0, 0, 3, 6, 
    35, 36, 38, 24, 0, 0, 11, 11, 0, 0, 0, 0, 0, 11, 11, 
    0, 0, 28, 24, 19, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 79, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 83, 18, 17, 0, 0, 7, 4, 0, 0, 0, 6, 
    0, 11, 56, 49, 25, 34, 2, 5, 0, 0, 8, 3, 0, 0, 0, 
    35, 4, 0, 7, 0, 2, 0, 10, 0, 0, 1, 6, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 13, 10, 
    0, 0, 0, 1, 15, 0, 0, 15, 0, 0, 0, 10, 1, 0, 25, 
    0, 0, 0, 0, 12, 15, 0, 7, 0, 0, 2, 0, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=227
    5, 3, 12, 11, 7, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 12, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 6, 2, 5, 0, 0, 0, 0, 0, 0, 0, 1, 2, 7, 5, 
    3, 5, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 4, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    22, 24, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 4, 
    29, 26, 17, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 17, 8, 
    20, 19, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    22, 25, 7, 0, 12, 0, 9, 0, 0, 0, 0, 0, 0, 0, 10, 
    16, 33, 43, 16, 31, 14, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    51, 45, 0, 25, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    63, 52, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 
    17, 23, 16, 8, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 10, 
    8, 7, 12, 15, 12, 4, 0, 0, 0, 1, 12, 0, 0, 0, 9, 
    11, 15, 7, 0, 5, 13, 0, 0, 0, 0, 0, 3, 0, 0, 4, 
    
    -- channel=228
    9, 9, 7, 8, 0, 0, 0, 3, 8, 7, 8, 10, 9, 9, 11, 
    9, 9, 6, 7, 0, 0, 0, 0, 0, 5, 3, 2, 0, 0, 1, 
    9, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 
    7, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 9, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 12, 29, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 27, 17, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=229
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 12, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 13, 15, 16, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 4, 3, 15, 22, 17, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 15, 18, 22, 26, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 6, 10, 5, 11, 19, 20, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 6, 5, 17, 23, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 8, 5, 14, 21, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 7, 4, 8, 19, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 9, 8, 8, 8, 15, 8, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 2, 8, 3, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 2, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=230
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 30, 39, 38, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 31, 20, 11, 0, 0, 0, 
    0, 0, 21, 4, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 2, 
    60, 74, 43, 0, 0, 3, 22, 6, 0, 0, 0, 0, 6, 13, 17, 
    11, 0, 0, 4, 15, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 
    0, 6, 0, 8, 57, 47, 12, 0, 1, 0, 0, 0, 0, 0, 4, 
    9, 24, 72, 67, 28, 24, 5, 3, 0, 0, 3, 0, 0, 0, 0, 
    86, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 6, 3, 0, 0, 3, 
    0, 0, 0, 0, 7, 16, 0, 0, 4, 7, 11, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=231
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 10, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 2, 1, 0, 1, 0, 9, 0, 0, 0, 0, 0, 
    13, 7, 0, 0, 0, 21, 0, 0, 0, 0, 1, 1, 2, 0, 0, 
    0, 0, 0, 0, 5, 17, 0, 0, 0, 0, 0, 9, 2, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 5, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 9, 0, 3, 0, 0, 4, 0, 0, 0, 4, 3, 0, 
    2, 12, 13, 0, 0, 0, 10, 0, 3, 0, 0, 0, 8, 0, 0, 
    2, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 2, 20, 0, 10, 9, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 1, 14, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=232
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=233
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 13, 20, 
    0, 1, 6, 11, 17, 5, 1, 9, 17, 9, 9, 5, 7, 22, 25, 
    
    -- channel=234
    0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 13, 15, 4, 0, 3, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 5, 0, 0, 12, 33, 5, 0, 0, 0, 0, 0, 0, 12, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 25, 5, 24, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 35, 49, 39, 45, 19, 23, 0, 0, 2, 0, 0, 0, 0, 
    94, 80, 11, 0, 0, 9, 0, 0, 15, 0, 0, 0, 0, 0, 0, 
    29, 22, 5, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 30, 19, 0, 0, 0, 5, 25, 37, 1, 0, 0, 8, 
    19, 30, 11, 0, 0, 0, 0, 0, 0, 0, 7, 17, 6, 1, 4, 
    
    -- channel=235
    2, 1, 1, 3, 11, 15, 13, 6, 4, 7, 5, 5, 5, 5, 4, 
    2, 3, 7, 0, 23, 29, 27, 25, 11, 6, 7, 7, 7, 7, 6, 
    3, 4, 8, 9, 26, 36, 41, 38, 23, 14, 9, 10, 5, 4, 4, 
    5, 4, 3, 19, 30, 37, 37, 42, 40, 30, 20, 15, 6, 4, 8, 
    0, 2, 19, 3, 30, 33, 34, 35, 45, 45, 43, 30, 16, 8, 12, 
    0, 0, 4, 0, 22, 36, 32, 32, 40, 40, 47, 38, 22, 10, 8, 
    0, 0, 0, 0, 21, 24, 32, 37, 38, 33, 44, 39, 28, 15, 5, 
    0, 0, 3, 0, 6, 14, 26, 35, 38, 33, 39, 43, 37, 19, 8, 
    0, 0, 0, 0, 12, 16, 21, 28, 36, 32, 37, 43, 38, 22, 14, 
    0, 0, 0, 0, 13, 25, 23, 24, 38, 33, 37, 41, 35, 17, 11, 
    0, 0, 0, 15, 21, 30, 29, 21, 36, 34, 34, 35, 30, 20, 14, 
    0, 0, 0, 7, 16, 29, 27, 16, 31, 30, 31, 31, 24, 21, 11, 
    0, 0, 0, 3, 8, 14, 29, 23, 31, 28, 32, 30, 26, 23, 18, 
    2, 8, 13, 11, 7, 16, 14, 27, 24, 27, 27, 25, 29, 19, 18, 
    10, 9, 10, 13, 13, 19, 17, 14, 18, 22, 22, 22, 17, 18, 17, 
    
    -- channel=236
    67, 64, 59, 64, 65, 69, 65, 54, 50, 43, 36, 28, 19, 14, 17, 
    65, 63, 54, 54, 59, 54, 65, 56, 45, 42, 42, 41, 41, 43, 43, 
    58, 57, 48, 32, 47, 45, 47, 51, 54, 68, 67, 66, 58, 52, 42, 
    54, 56, 60, 29, 38, 47, 48, 50, 56, 57, 68, 69, 55, 51, 41, 
    88, 107, 114, 58, 38, 51, 76, 70, 58, 57, 57, 64, 61, 62, 57, 
    125, 133, 136, 62, 51, 57, 85, 73, 64, 63, 61, 54, 57, 66, 64, 
    119, 121, 124, 103, 38, 51, 78, 68, 70, 72, 64, 52, 58, 52, 54, 
    114, 122, 125, 112, 111, 57, 80, 65, 81, 88, 70, 56, 54, 50, 51, 
    128, 146, 176, 164, 141, 119, 82, 85, 79, 88, 77, 66, 55, 52, 38, 
    191, 206, 200, 190, 127, 128, 80, 94, 79, 86, 85, 77, 55, 43, 14, 
    225, 219, 173, 104, 78, 80, 63, 63, 77, 79, 78, 72, 52, 43, 28, 
    167, 141, 113, 96, 79, 42, 54, 60, 42, 60, 75, 79, 51, 34, 49, 
    89, 81, 80, 76, 79, 61, 49, 63, 52, 66, 97, 83, 59, 32, 39, 
    65, 65, 63, 49, 37, 43, 47, 50, 47, 46, 64, 73, 53, 30, 26, 
    49, 36, 28, 21, 15, 37, 45, 34, 24, 26, 29, 35, 33, 12, 15, 
    
    -- channel=237
    17, 16, 14, 14, 3, 0, 6, 8, 9, 7, 7, 6, 3, 2, 1, 
    17, 15, 12, 7, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 
    15, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 22, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 21, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 18, 14, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 19, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 34, 38, 12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 40, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 33, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 15, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=238
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    2, 9, 13, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    22, 22, 14, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=239
    16, 17, 14, 19, 12, 1, 11, 13, 12, 13, 14, 13, 11, 6, 2, 
    16, 15, 16, 11, 6, 6, 0, 0, 9, 3, 0, 0, 0, 0, 0, 
    18, 16, 22, 9, 1, 0, 0, 0, 0, 0, 0, 0, 2, 5, 5, 
    13, 9, 0, 4, 0, 0, 0, 0, 0, 4, 2, 1, 0, 1, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 16, 8, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 19, 8, 0, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    12, 7, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 37, 16, 16, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 34, 31, 31, 25, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 51, 19, 5, 3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    31, 24, 15, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 7, 11, 10, 0, 0, 0, 0, 0, 10, 13, 0, 0, 0, 0, 
    12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=240
    60, 56, 60, 65, 63, 58, 53, 48, 39, 33, 27, 18, 8, 3, 0, 
    58, 52, 54, 47, 49, 53, 51, 41, 35, 28, 20, 17, 18, 23, 24, 
    54, 51, 43, 37, 30, 24, 27, 29, 40, 54, 54, 54, 51, 48, 38, 
    45, 45, 22, 9, 16, 13, 15, 26, 40, 58, 68, 59, 48, 42, 30, 
    61, 80, 80, 24, 18, 36, 46, 34, 28, 33, 47, 52, 52, 49, 44, 
    126, 136, 100, 27, 19, 42, 59, 43, 32, 28, 27, 39, 55, 64, 58, 
    130, 127, 112, 49, 33, 59, 56, 42, 46, 39, 27, 37, 52, 59, 52, 
    114, 119, 125, 100, 48, 29, 43, 43, 60, 54, 33, 29, 37, 38, 37, 
    125, 136, 135, 124, 121, 89, 68, 53, 60, 57, 40, 28, 34, 44, 40, 
    174, 211, 229, 181, 136, 104, 79, 61, 56, 60, 53, 38, 34, 24, 5, 
    242, 234, 153, 100, 90, 75, 59, 49, 56, 61, 53, 34, 28, 24, 11, 
    216, 169, 110, 79, 37, 18, 37, 32, 29, 40, 49, 44, 28, 38, 26, 
    99, 92, 81, 76, 58, 39, 46, 35, 32, 52, 69, 59, 34, 28, 35, 
    60, 65, 70, 58, 41, 35, 29, 33, 32, 49, 63, 50, 35, 20, 30, 
    56, 43, 26, 14, 18, 37, 37, 23, 13, 14, 23, 32, 22, 11, 13, 
    
    -- channel=241
    2, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 1, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 39, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    36, 33, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 25, 26, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 34, 26, 18, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 55, 72, 36, 34, 14, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 84, 51, 30, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    80, 64, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 8, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 3, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=242
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 9, 7, 9, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 13, 0, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 3, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 3, 
    0, 0, 42, 40, 0, 29, 0, 12, 0, 0, 0, 6, 0, 0, 0, 
    0, 53, 9, 0, 13, 15, 0, 0, 15, 4, 0, 0, 0, 0, 0, 
    8, 3, 8, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 23, 0, 0, 0, 0, 0, 17, 11, 0, 0, 0, 
    0, 18, 20, 1, 0, 0, 0, 5, 0, 0, 0, 3, 15, 0, 0, 
    
    -- channel=243
    15, 15, 15, 12, 22, 29, 17, 16, 16, 14, 13, 13, 13, 14, 16, 
    16, 16, 13, 22, 24, 27, 33, 27, 18, 19, 21, 21, 20, 17, 15, 
    15, 15, 7, 26, 32, 39, 41, 43, 34, 22, 20, 18, 15, 11, 12, 
    18, 20, 23, 22, 43, 46, 47, 43, 39, 26, 27, 22, 18, 17, 19, 
    28, 25, 9, 34, 36, 41, 44, 45, 46, 44, 40, 34, 22, 21, 21, 
    19, 18, 16, 28, 42, 39, 39, 48, 47, 49, 49, 44, 25, 22, 18, 
    15, 17, 20, 33, 16, 33, 42, 48, 44, 44, 45, 46, 31, 16, 13, 
    22, 21, 15, 22, 33, 33, 38, 45, 43, 43, 48, 46, 36, 25, 19, 
    25, 32, 37, 27, 30, 22, 32, 42, 43, 44, 48, 47, 40, 24, 14, 
    26, 19, 5, 22, 22, 19, 27, 46, 46, 45, 47, 49, 42, 27, 17, 
    17, 9, 24, 20, 28, 31, 35, 39, 43, 41, 43, 49, 39, 28, 14, 
    3, 13, 22, 23, 35, 42, 38, 34, 39, 44, 42, 42, 32, 22, 24, 
    15, 16, 19, 18, 21, 30, 29, 33, 37, 44, 38, 38, 36, 22, 22, 
    19, 17, 15, 16, 22, 22, 31, 27, 38, 35, 35, 45, 33, 24, 20, 
    12, 17, 22, 21, 19, 20, 24, 25, 25, 26, 27, 28, 30, 22, 17, 
    
    -- channel=244
    15, 16, 12, 19, 12, 0, 6, 5, 8, 3, 0, 0, 0, 0, 0, 
    14, 12, 8, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    11, 8, 15, 0, 0, 0, 0, 0, 0, 7, 10, 10, 15, 14, 9, 
    5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 7, 10, 1, 
    10, 22, 33, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 
    44, 51, 33, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 18, 
    47, 47, 35, 36, 4, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 
    34, 39, 48, 32, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    39, 40, 44, 78, 28, 35, 1, 5, 0, 0, 0, 0, 0, 0, 7, 
    70, 91, 110, 73, 36, 19, 10, 6, 0, 0, 0, 0, 0, 0, 0, 
    102, 106, 94, 20, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    92, 65, 50, 23, 12, 0, 0, 8, 0, 0, 0, 0, 0, 0, 4, 
    34, 25, 20, 21, 16, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 15, 18, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 6, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=245
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 8, 25, 8, 12, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    25, 32, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    9, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 
    0, 0, 2, 14, 16, 1, 0, 0, 0, 0, 5, 0, 0, 10, 12, 
    4, 16, 15, 6, 10, 7, 1, 8, 7, 4, 5, 9, 7, 10, 13, 
    
    -- channel=246
    15, 13, 21, 23, 14, 14, 8, 13, 6, 3, 2, 0, 0, 0, 0, 
    15, 11, 16, 10, 0, 0, 5, 0, 5, 4, 0, 0, 0, 0, 0, 
    12, 13, 7, 9, 0, 0, 0, 0, 3, 5, 12, 15, 18, 21, 19, 
    8, 10, 2, 0, 0, 0, 0, 0, 0, 16, 17, 17, 26, 16, 12, 
    10, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 23, 18, 
    48, 56, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 39, 33, 
    60, 60, 52, 6, 0, 8, 0, 0, 0, 0, 0, 0, 10, 38, 34, 
    47, 50, 47, 50, 6, 0, 0, 0, 0, 0, 0, 0, 0, 12, 18, 
    50, 62, 56, 14, 50, 21, 26, 0, 0, 0, 0, 0, 0, 3, 28, 
    62, 83, 98, 90, 48, 49, 17, 0, 0, 0, 0, 0, 0, 5, 19, 
    116, 111, 70, 44, 24, 21, 4, 9, 0, 0, 0, 0, 0, 14, 9, 
    114, 102, 61, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 20, 
    47, 41, 38, 29, 17, 0, 0, 0, 0, 0, 0, 0, 4, 15, 31, 
    25, 21, 23, 31, 31, 20, 0, 0, 0, 0, 11, 0, 0, 19, 21, 
    22, 28, 23, 13, 19, 23, 12, 16, 9, 2, 0, 6, 10, 15, 22, 
    
    -- channel=247
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=248
    64, 60, 63, 59, 66, 73, 61, 55, 49, 45, 38, 31, 26, 27, 26, 
    62, 60, 60, 48, 64, 65, 69, 62, 47, 47, 49, 51, 51, 51, 47, 
    58, 57, 42, 46, 55, 61, 64, 70, 71, 75, 67, 66, 55, 47, 38, 
    57, 61, 54, 38, 58, 68, 70, 69, 68, 70, 75, 63, 56, 50, 45, 
    96, 109, 94, 39, 56, 78, 88, 73, 74, 73, 76, 75, 67, 62, 59, 
    113, 113, 92, 41, 65, 88, 82, 79, 81, 74, 74, 76, 71, 65, 58, 
    101, 100, 100, 69, 52, 66, 79, 80, 86, 78, 71, 75, 69, 58, 43, 
    105, 111, 108, 86, 77, 77, 79, 79, 95, 87, 74, 73, 71, 57, 55, 
    119, 137, 157, 126, 129, 101, 91, 76, 91, 90, 84, 75, 74, 60, 31, 
    175, 178, 144, 130, 106, 95, 81, 81, 93, 94, 92, 79, 72, 43, 22, 
    178, 163, 83, 86, 81, 68, 77, 64, 85, 86, 78, 78, 66, 54, 27, 
    109, 93, 88, 76, 60, 59, 77, 53, 65, 79, 87, 82, 52, 51, 42, 
    75, 70, 71, 75, 65, 59, 59, 64, 68, 89, 100, 81, 63, 44, 48, 
    65, 68, 60, 43, 39, 53, 51, 59, 57, 63, 73, 79, 61, 36, 38, 
    45, 33, 34, 29, 31, 49, 51, 35, 31, 38, 43, 45, 37, 26, 24, 
    
    -- channel=249
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=250
    9, 10, 9, 9, 18, 20, 19, 14, 15, 15, 14, 15, 16, 17, 19, 
    9, 11, 12, 12, 28, 25, 28, 28, 17, 18, 21, 25, 26, 25, 25, 
    10, 10, 13, 20, 31, 37, 37, 38, 30, 26, 23, 24, 19, 17, 18, 
    13, 13, 23, 32, 35, 38, 43, 45, 39, 24, 24, 23, 19, 22, 26, 
    20, 22, 31, 32, 36, 31, 40, 45, 46, 43, 38, 30, 23, 32, 34, 
    10, 7, 12, 28, 35, 34, 32, 39, 41, 47, 48, 33, 25, 30, 29, 
    1, 3, 6, 36, 28, 21, 34, 38, 36, 42, 46, 38, 31, 22, 19, 
    7, 9, 14, 11, 40, 35, 42, 42, 34, 37, 44, 44, 31, 22, 25, 
    10, 9, 17, 33, 26, 38, 32, 45, 30, 32, 42, 44, 32, 26, 26, 
    16, 11, 0, 14, 7, 23, 25, 42, 34, 31, 38, 44, 34, 27, 33, 
    0, 0, 1, 5, 18, 18, 27, 26, 35, 32, 34, 41, 35, 33, 38, 
    0, 0, 7, 18, 30, 31, 27, 35, 30, 28, 34, 38, 35, 30, 40, 
    2, 3, 8, 17, 27, 36, 26, 31, 36, 28, 31, 32, 39, 38, 32, 
    13, 19, 20, 19, 21, 31, 35, 32, 36, 27, 18, 29, 32, 35, 35, 
    19, 20, 27, 35, 34, 33, 36, 35, 41, 38, 34, 31, 34, 38, 38, 
    
    -- channel=251
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=252
    0, 0, 0, 0, 0, 0, 5, 5, 5, 0, 4, 9, 7, 0, 7, 
    0, 4, 0, 0, 0, 0, 8, 4, 8, 2, 2, 1, 0, 0, 4, 
    0, 0, 6, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 
    0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 10, 1, 8, 8, 
    0, 0, 33, 42, 0, 0, 0, 12, 0, 0, 0, 0, 0, 6, 2, 
    0, 0, 64, 39, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 9, 83, 0, 0, 14, 0, 0, 6, 5, 0, 0, 0, 13, 
    0, 0, 0, 21, 73, 0, 6, 0, 0, 14, 10, 0, 0, 0, 6, 
    0, 0, 0, 11, 12, 35, 0, 9, 0, 6, 7, 6, 0, 0, 18, 
    0, 0, 0, 79, 0, 52, 0, 30, 0, 0, 0, 15, 0, 22, 9, 
    0, 8, 94, 2, 0, 11, 0, 0, 0, 0, 4, 10, 0, 7, 16, 
    14, 19, 42, 20, 29, 0, 0, 24, 0, 0, 0, 7, 14, 0, 34, 
    6, 0, 0, 0, 27, 7, 0, 18, 0, 0, 0, 5, 27, 0, 0, 
    0, 0, 0, 11, 2, 0, 0, 0, 0, 0, 0, 6, 7, 5, 0, 
    4, 8, 5, 8, 0, 0, 3, 14, 3, 0, 0, 0, 11, 0, 0, 
    
    -- channel=253
    10, 9, 12, 12, 22, 23, 13, 13, 8, 9, 8, 6, 5, 5, 3, 
    10, 9, 12, 16, 22, 31, 29, 20, 12, 13, 10, 8, 4, 3, 4, 
    11, 12, 10, 18, 29, 31, 37, 38, 22, 10, 12, 15, 13, 14, 16, 
    11, 12, 8, 13, 30, 31, 33, 37, 38, 34, 26, 22, 18, 14, 15, 
    9, 7, 2, 15, 24, 33, 28, 30, 41, 39, 40, 31, 23, 22, 20, 
    19, 23, 22, 7, 25, 29, 32, 33, 37, 39, 40, 39, 28, 30, 24, 
    24, 25, 25, 0, 21, 38, 37, 37, 33, 30, 39, 37, 26, 28, 21, 
    22, 22, 20, 25, 7, 16, 28, 37, 36, 30, 35, 34, 33, 24, 19, 
    23, 28, 24, 4, 27, 13, 35, 32, 38, 33, 33, 33, 33, 20, 24, 
    15, 19, 27, 32, 41, 34, 36, 36, 36, 33, 35, 34, 30, 20, 21, 
    33, 31, 27, 49, 35, 47, 33, 41, 40, 35, 38, 38, 28, 22, 15, 
    38, 45, 22, 22, 22, 33, 29, 14, 39, 35, 30, 32, 25, 32, 20, 
    24, 22, 23, 19, 19, 14, 30, 26, 27, 31, 27, 29, 24, 27, 33, 
    21, 18, 22, 28, 33, 27, 25, 30, 33, 31, 43, 34, 27, 30, 32, 
    19, 29, 31, 23, 26, 32, 26, 29, 31, 29, 33, 35, 32, 26, 29, 
    
    -- channel=254
    22, 22, 18, 24, 27, 31, 30, 25, 15, 14, 14, 10, 5, 0, 0, 
    22, 22, 17, 21, 24, 26, 39, 29, 20, 11, 8, 5, 1, 0, 4, 
    21, 21, 22, 12, 25, 20, 20, 28, 24, 15, 16, 20, 17, 19, 19, 
    17, 15, 22, 0, 14, 13, 12, 15, 24, 37, 34, 35, 23, 19, 13, 
    10, 14, 40, 20, 6, 13, 20, 23, 25, 27, 30, 36, 23, 19, 14, 
    35, 46, 70, 13, 11, 2, 34, 35, 21, 19, 23, 23, 24, 25, 23, 
    48, 50, 54, 38, 3, 16, 40, 28, 23, 26, 28, 17, 30, 26, 29, 
    41, 41, 48, 52, 31, 0, 20, 17, 28, 37, 28, 21, 28, 20, 22, 
    36, 37, 47, 41, 58, 46, 32, 25, 30, 38, 30, 27, 20, 22, 22, 
    41, 54, 79, 111, 55, 77, 28, 44, 29, 34, 33, 33, 20, 25, 8, 
    86, 98, 95, 72, 49, 62, 34, 29, 28, 33, 32, 32, 19, 16, 6, 
    98, 96, 70, 33, 27, 13, 20, 14, 14, 24, 24, 28, 20, 9, 24, 
    52, 38, 40, 31, 34, 9, 7, 37, 11, 14, 34, 37, 32, 9, 19, 
    28, 24, 29, 32, 23, 19, 7, 17, 12, 13, 35, 33, 27, 16, 6, 
    23, 24, 18, 9, 0, 11, 18, 17, 5, 7, 2, 12, 16, 3, 6, 
    
    -- channel=255
    14, 13, 20, 13, 24, 25, 18, 16, 14, 16, 16, 14, 16, 19, 14, 
    14, 12, 20, 19, 27, 42, 30, 30, 20, 18, 18, 17, 17, 17, 14, 
    16, 15, 15, 27, 34, 44, 49, 49, 35, 21, 19, 20, 18, 17, 18, 
    17, 18, 3, 28, 43, 44, 46, 51, 51, 41, 31, 24, 19, 15, 20, 
    15, 12, 0, 11, 43, 47, 37, 38, 51, 51, 51, 38, 29, 21, 23, 
    15, 11, 0, 7, 31, 50, 35, 36, 46, 47, 48, 53, 41, 28, 22, 
    13, 11, 3, 0, 33, 47, 32, 43, 42, 37, 43, 56, 41, 33, 18, 
    15, 13, 10, 5, 0, 34, 28, 45, 44, 30, 40, 49, 42, 34, 20, 
    16, 14, 0, 0, 11, 5, 27, 33, 45, 33, 37, 41, 48, 36, 23, 
    5, 6, 0, 0, 29, 0, 40, 27, 43, 38, 37, 37, 48, 26, 25, 
    0, 0, 0, 21, 35, 33, 44, 37, 44, 41, 37, 38, 42, 27, 24, 
    2, 3, 0, 9, 13, 44, 42, 19, 45, 45, 37, 35, 33, 42, 17, 
    10, 16, 15, 18, 8, 22, 40, 24, 41, 49, 29, 33, 32, 40, 32, 
    20, 22, 25, 25, 28, 25, 32, 33, 37, 45, 38, 33, 36, 36, 40, 
    23, 26, 29, 28, 40, 35, 30, 30, 34, 34, 42, 37, 30, 36, 35, 
    
    -- channel=256
    0, 53, 73, 52, 45, 60, 58, 59, 48, 1, 71, 66, 69, 69, 68, 
    1, 27, 74, 59, 45, 32, 51, 60, 50, 16, 81, 59, 61, 65, 65, 
    3, 8, 80, 55, 59, 13, 26, 40, 35, 52, 54, 58, 55, 58, 56, 
    11, 51, 62, 30, 63, 39, 31, 24, 36, 58, 46, 71, 53, 35, 59, 
    42, 56, 47, 23, 60, 46, 34, 15, 35, 49, 55, 71, 54, 30, 53, 
    47, 48, 45, 39, 53, 39, 28, 28, 37, 47, 48, 73, 53, 34, 41, 
    47, 52, 34, 62, 38, 45, 23, 47, 30, 43, 48, 72, 58, 51, 39, 
    38, 52, 34, 82, 36, 39, 36, 26, 54, 39, 37, 47, 74, 43, 55, 
    31, 46, 58, 58, 52, 51, 36, 21, 51, 41, 48, 35, 51, 43, 69, 
    41, 44, 52, 49, 46, 41, 50, 42, 31, 54, 33, 54, 54, 42, 48, 
    47, 30, 60, 52, 52, 30, 55, 48, 41, 27, 49, 51, 49, 37, 37, 
    46, 31, 61, 51, 46, 43, 56, 51, 41, 26, 55, 42, 52, 38, 37, 
    41, 35, 58, 48, 29, 50, 59, 48, 37, 31, 50, 40, 35, 45, 40, 
    39, 32, 55, 53, 38, 55, 41, 44, 34, 35, 44, 40, 30, 48, 47, 
    34, 38, 41, 57, 41, 36, 29, 43, 25, 43, 39, 42, 38, 41, 43, 
    
    -- channel=257
    0, 0, 26, 29, 29, 30, 32, 36, 36, 16, 11, 46, 39, 40, 37, 
    0, 0, 20, 21, 41, 38, 35, 39, 40, 26, 30, 51, 47, 43, 40, 
    0, 0, 17, 21, 38, 35, 14, 18, 18, 23, 49, 50, 54, 57, 56, 
    25, 23, 58, 38, 30, 47, 36, 26, 21, 24, 49, 55, 63, 59, 52, 
    64, 50, 58, 36, 30, 40, 42, 25, 19, 20, 50, 60, 64, 63, 52, 
    57, 53, 56, 38, 42, 40, 30, 21, 29, 25, 38, 62, 71, 69, 61, 
    59, 50, 42, 33, 30, 30, 39, 27, 45, 32, 41, 60, 71, 77, 70, 
    61, 45, 24, 39, 54, 35, 42, 26, 30, 43, 36, 45, 51, 68, 61, 
    60, 40, 39, 41, 50, 56, 45, 41, 29, 23, 43, 13, 26, 39, 51, 
    71, 55, 49, 41, 46, 44, 43, 50, 31, 34, 36, 26, 26, 38, 23, 
    66, 53, 47, 51, 53, 44, 37, 37, 49, 36, 21, 35, 31, 29, 28, 
    63, 58, 48, 52, 50, 39, 45, 41, 42, 30, 28, 31, 34, 32, 24, 
    62, 64, 50, 48, 38, 1, 39, 36, 33, 23, 25, 25, 27, 22, 25, 
    60, 58, 46, 53, 56, 26, 38, 24, 24, 16, 25, 21, 21, 18, 30, 
    48, 53, 43, 46, 48, 44, 27, 20, 17, 12, 21, 24, 23, 25, 23, 
    
    -- channel=258
    3, 0, 0, 0, 0, 0, 0, 0, 40, 35, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 14, 0, 0, 0, 0, 47, 0, 1, 0, 0, 0, 
    1, 0, 0, 0, 0, 34, 0, 0, 0, 2, 0, 0, 0, 0, 7, 
    110, 56, 0, 0, 0, 25, 55, 22, 0, 0, 0, 0, 0, 0, 0, 
    38, 7, 0, 23, 0, 0, 0, 11, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 19, 0, 0, 0, 9, 6, 0, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 2, 0, 0, 0, 0, 11, 22, 
    0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 18, 0, 0, 19, 21, 29, 0, 0, 0, 23, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 29, 47, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    
    -- channel=259
    0, 42, 44, 14, 16, 24, 15, 16, 3, 0, 42, 31, 19, 19, 18, 
    0, 17, 73, 23, 24, 7, 32, 31, 26, 0, 46, 27, 21, 21, 21, 
    0, 5, 76, 13, 52, 0, 26, 45, 39, 21, 42, 39, 29, 27, 21, 
    0, 0, 32, 5, 71, 18, 0, 4, 20, 41, 46, 45, 32, 32, 43, 
    0, 15, 24, 0, 55, 42, 24, 6, 25, 37, 48, 53, 34, 4, 32, 
    21, 25, 29, 0, 44, 38, 26, 5, 21, 27, 41, 62, 35, 0, 11, 
    19, 22, 17, 36, 25, 27, 15, 28, 23, 37, 31, 61, 37, 20, 0, 
    12, 28, 0, 72, 17, 34, 24, 12, 49, 19, 33, 65, 68, 38, 24, 
    5, 24, 25, 41, 31, 29, 10, 13, 36, 9, 35, 0, 60, 48, 55, 
    10, 8, 37, 33, 41, 49, 45, 16, 0, 26, 28, 28, 9, 21, 41, 
    24, 6, 47, 27, 27, 17, 52, 39, 28, 23, 21, 25, 31, 17, 19, 
    27, 10, 48, 40, 37, 26, 34, 30, 28, 2, 29, 25, 38, 11, 11, 
    21, 13, 40, 40, 32, 24, 51, 34, 27, 9, 34, 21, 35, 30, 18, 
    18, 7, 30, 45, 17, 5, 33, 29, 17, 11, 29, 18, 10, 29, 23, 
    19, 14, 14, 60, 26, 22, 17, 30, 10, 14, 21, 21, 8, 20, 30, 
    
    -- channel=260
    15, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    14, 1, 0, 0, 4, 2, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    13, 9, 0, 0, 4, 16, 10, 3, 3, 2, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 11, 4, 7, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 10, 7, 12, 7, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 12, 16, 6, 4, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 16, 15, 4, 6, 2, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 4, 14, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 1, 12, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 8, 6, 8, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 5, 3, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 2, 1, 1, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 4, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    
    -- channel=261
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=262
    0, 0, 0, 0, 0, 0, 0, 2, 26, 8, 3, 20, 8, 4, 0, 
    0, 0, 0, 0, 19, 1, 0, 0, 0, 0, 50, 8, 2, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 22, 0, 0, 6, 13, 
    112, 111, 85, 0, 0, 10, 51, 12, 0, 0, 0, 5, 9, 0, 0, 
    39, 54, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 19, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 9, 0, 0, 0, 0, 4, 15, 
    0, 0, 0, 0, 4, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 7, 0, 34, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 19, 36, 3, 0, 0, 17, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=263
    2, 39, 13, 0, 0, 3, 0, 0, 0, 0, 55, 0, 0, 0, 0, 
    1, 8, 38, 10, 2, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 
    0, 0, 73, 0, 20, 0, 0, 0, 0, 25, 2, 0, 0, 0, 0, 
    0, 46, 15, 0, 31, 0, 0, 0, 5, 19, 0, 17, 0, 0, 3, 
    0, 0, 0, 0, 24, 0, 0, 0, 2, 10, 18, 8, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 3, 0, 22, 0, 0, 0, 
    0, 0, 0, 8, 0, 5, 0, 13, 0, 2, 0, 16, 0, 0, 0, 
    0, 0, 0, 54, 0, 0, 0, 0, 22, 0, 0, 0, 19, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 9, 0, 0, 0, 11, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 4, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 9, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 8, 0, 2, 0, 0, 
    0, 0, 7, 0, 0, 0, 7, 0, 0, 0, 5, 0, 0, 2, 0, 
    0, 0, 6, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 6, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    
    -- channel=264
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=265
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=266
    0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 23, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 8, 0, 0, 0, 19, 46, 44, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 7, 82, 29, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 56, 55, 27, 
    0, 0, 0, 0, 0, 24, 1, 0, 0, 0, 7, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 0, 8, 7, 0, 3, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 23, 6, 7, 12, 2, 2, 1, 22, 11, 0, 
    0, 0, 6, 0, 0, 0, 4, 11, 12, 7, 0, 0, 0, 0, 0, 
    17, 0, 9, 7, 0, 0, 20, 14, 7, 0, 0, 0, 0, 0, 6, 
    
    -- channel=267
    3, 0, 16, 4, 1, 7, 8, 6, 1, 0, 0, 10, 8, 9, 9, 
    3, 0, 27, 0, 0, 0, 0, 3, 5, 0, 7, 0, 2, 3, 4, 
    3, 1, 23, 0, 0, 0, 0, 3, 0, 0, 12, 0, 0, 0, 0, 
    6, 0, 28, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    1, 6, 4, 0, 3, 0, 0, 0, 0, 0, 0, 3, 0, 0, 7, 
    2, 1, 4, 0, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 11, 
    4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    3, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 5, 0, 3, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 12, 1, 2, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 7, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 3, 0, 0, 3, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 2, 0, 0, 
    2, 8, 2, 0, 0, 0, 4, 0, 0, 0, 6, 0, 4, 0, 1, 
    2, 10, 1, 0, 0, 0, 2, 0, 0, 0, 8, 0, 0, 1, 2, 
    1, 14, 0, 0, 0, 0, 0, 3, 3, 0, 2, 3, 0, 6, 1, 
    
    -- channel=268
    0, 0, 94, 115, 107, 103, 115, 115, 128, 92, 49, 132, 138, 136, 134, 
    0, 0, 57, 105, 135, 126, 112, 131, 140, 124, 75, 164, 159, 151, 147, 
    0, 0, 28, 107, 137, 158, 89, 83, 100, 102, 133, 162, 176, 174, 174, 
    89, 47, 96, 134, 120, 168, 139, 105, 80, 90, 156, 162, 200, 190, 169, 
    163, 137, 162, 143, 107, 155, 154, 122, 81, 93, 144, 177, 207, 196, 151, 
    167, 160, 165, 147, 129, 150, 146, 110, 103, 105, 138, 171, 216, 208, 160, 
    172, 160, 149, 130, 142, 132, 142, 106, 139, 120, 139, 173, 212, 220, 196, 
    173, 149, 143, 111, 168, 149, 143, 126, 118, 130, 141, 120, 175, 208, 190, 
    180, 133, 140, 138, 174, 179, 170, 149, 92, 129, 128, 115, 90, 142, 148, 
    190, 158, 156, 162, 160, 163, 167, 174, 146, 115, 127, 104, 112, 123, 112, 
    189, 173, 152, 176, 175, 170, 132, 156, 163, 134, 100, 111, 122, 122, 101, 
    183, 178, 143, 180, 179, 155, 147, 157, 154, 131, 92, 119, 121, 125, 109, 
    181, 169, 145, 176, 164, 103, 132, 144, 136, 108, 93, 108, 104, 103, 105, 
    176, 160, 133, 171, 173, 129, 137, 117, 107, 87, 88, 98, 94, 80, 105, 
    151, 145, 122, 152, 173, 153, 116, 92, 90, 66, 87, 93, 96, 87, 97, 
    
    -- channel=269
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 1, 0, 0, 14, 4, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 2, 0, 0, 25, 14, 4, 0, 0, 0, 21, 13, 9, 8, 4, 
    0, 2, 9, 0, 25, 18, 7, 3, 3, 14, 18, 20, 24, 22, 17, 
    0, 7, 10, 0, 23, 25, 15, 6, 7, 16, 18, 22, 21, 9, 11, 
    8, 13, 7, 0, 19, 24, 13, 8, 12, 18, 19, 24, 24, 7, 5, 
    5, 4, 0, 0, 17, 22, 17, 15, 20, 23, 21, 22, 23, 18, 11, 
    7, 5, 0, 3, 20, 22, 22, 15, 7, 15, 11, 11, 14, 21, 16, 
    5, 8, 0, 14, 22, 26, 27, 13, 5, 0, 0, 0, 7, 3, 9, 
    10, 13, 18, 13, 25, 28, 26, 22, 3, 0, 0, 0, 0, 0, 0, 
    16, 14, 20, 16, 16, 14, 18, 20, 12, 0, 0, 0, 1, 0, 0, 
    17, 9, 24, 24, 17, 4, 9, 11, 9, 0, 0, 1, 2, 0, 0, 
    14, 6, 19, 27, 10, 0, 2, 3, 0, 0, 0, 0, 2, 0, 0, 
    10, 0, 12, 26, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 10, 28, 19, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=270
    0, 0, 5, 0, 0, 4, 0, 6, 0, 0, 8, 6, 7, 8, 6, 
    0, 0, 4, 5, 0, 0, 4, 7, 1, 0, 15, 12, 11, 11, 9, 
    0, 0, 7, 0, 14, 0, 0, 0, 0, 1, 8, 20, 17, 18, 15, 
    0, 0, 4, 0, 15, 0, 0, 0, 0, 7, 8, 30, 18, 5, 23, 
    7, 5, 11, 0, 10, 6, 0, 0, 0, 0, 17, 29, 21, 6, 19, 
    13, 13, 10, 0, 8, 2, 0, 0, 0, 0, 6, 36, 27, 10, 13, 
    14, 14, 0, 8, 0, 4, 0, 0, 0, 0, 9, 31, 31, 27, 14, 
    12, 14, 0, 23, 4, 0, 1, 0, 4, 3, 0, 19, 36, 20, 27, 
    3, 8, 5, 10, 15, 8, 0, 0, 3, 0, 0, 0, 10, 14, 33, 
    17, 11, 12, 4, 11, 12, 13, 3, 0, 4, 0, 0, 0, 0, 0, 
    21, 3, 20, 13, 13, 0, 10, 9, 4, 0, 0, 0, 0, 0, 0, 
    20, 4, 22, 16, 8, 1, 8, 7, 0, 0, 0, 0, 1, 0, 0, 
    15, 11, 21, 13, 0, 0, 9, 4, 0, 0, 0, 0, 0, 0, 0, 
    12, 6, 21, 19, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 6, 11, 19, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=271
    9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 13, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 13, 0, 0, 11, 9, 15, 21, 13, 0, 7, 7, 0, 0, 0, 
    0, 0, 0, 4, 17, 0, 0, 0, 1, 8, 13, 2, 5, 19, 8, 
    0, 0, 2, 0, 14, 16, 11, 8, 7, 9, 8, 4, 8, 6, 12, 
    1, 6, 7, 0, 9, 19, 13, 2, 2, 6, 13, 11, 10, 0, 3, 
    1, 1, 12, 0, 9, 11, 14, 2, 7, 10, 12, 9, 13, 0, 0, 
    8, 4, 0, 0, 9, 14, 10, 17, 4, 14, 18, 39, 10, 21, 5, 
    4, 5, 0, 2, 3, 0, 7, 4, 9, 0, 1, 0, 31, 25, 13, 
    0, 0, 5, 3, 20, 32, 15, 0, 0, 0, 6, 0, 0, 0, 14, 
    6, 12, 7, 3, 3, 11, 17, 19, 4, 11, 0, 0, 0, 0, 4, 
    11, 6, 12, 12, 14, 3, 0, 4, 10, 0, 0, 3, 1, 0, 0, 
    10, 7, 10, 16, 19, 4, 6, 8, 8, 0, 0, 2, 15, 0, 0, 
    10, 5, 9, 14, 0, 0, 4, 4, 5, 0, 0, 0, 1, 0, 0, 
    13, 0, 14, 19, 9, 11, 8, 0, 1, 0, 0, 0, 0, 0, 1, 
    
    -- channel=272
    0, 43, 111, 111, 107, 107, 109, 112, 95, 58, 82, 132, 132, 134, 130, 
    0, 23, 96, 115, 129, 119, 127, 138, 143, 82, 113, 162, 153, 149, 145, 
    0, 3, 67, 112, 161, 134, 100, 117, 121, 100, 146, 174, 174, 171, 166, 
    10, 11, 106, 130, 161, 152, 107, 84, 78, 123, 168, 187, 206, 200, 190, 
    127, 136, 158, 115, 138, 170, 153, 109, 91, 120, 160, 200, 211, 175, 170, 
    165, 166, 167, 130, 149, 168, 144, 98, 98, 120, 155, 201, 217, 176, 152, 
    166, 160, 148, 140, 137, 137, 131, 120, 131, 134, 152, 201, 222, 202, 167, 
    168, 162, 123, 143, 163, 160, 139, 134, 137, 142, 157, 181, 216, 216, 197, 
    160, 141, 130, 157, 176, 169, 156, 121, 118, 131, 130, 100, 137, 168, 187, 
    168, 153, 168, 167, 177, 192, 188, 155, 120, 125, 127, 109, 108, 120, 139, 
    185, 165, 168, 175, 176, 157, 161, 178, 161, 133, 107, 116, 131, 117, 109, 
    186, 161, 170, 192, 189, 158, 160, 164, 160, 110, 107, 126, 134, 122, 98, 
    178, 158, 169, 188, 164, 124, 158, 159, 142, 106, 109, 115, 121, 113, 102, 
    172, 145, 153, 183, 157, 131, 142, 129, 111, 88, 97, 102, 90, 95, 110, 
    154, 133, 138, 180, 173, 153, 121, 106, 84, 77, 92, 98, 87, 95, 108, 
    
    -- channel=273
    0, 0, 18, 22, 15, 16, 18, 23, 33, 2, 25, 36, 32, 29, 26, 
    0, 0, 8, 28, 46, 23, 23, 32, 32, 13, 48, 46, 40, 35, 32, 
    0, 0, 11, 33, 58, 34, 9, 5, 6, 32, 49, 44, 51, 53, 51, 
    21, 32, 48, 19, 49, 53, 42, 23, 19, 36, 43, 63, 66, 46, 47, 
    38, 50, 39, 20, 47, 50, 41, 19, 21, 33, 42, 66, 62, 31, 32, 
    40, 39, 33, 30, 48, 43, 30, 23, 35, 40, 40, 61, 59, 39, 26, 
    35, 35, 13, 41, 40, 45, 34, 40, 37, 44, 41, 59, 60, 58, 41, 
    29, 33, 22, 51, 46, 45, 43, 32, 34, 30, 27, 10, 47, 48, 49, 
    30, 31, 48, 48, 60, 70, 59, 34, 20, 25, 32, 18, 9, 12, 35, 
    39, 41, 49, 51, 47, 43, 55, 55, 40, 37, 14, 20, 31, 23, 15, 
    45, 34, 51, 53, 56, 37, 42, 47, 42, 17, 17, 30, 34, 21, 15, 
    41, 33, 51, 58, 49, 38, 46, 47, 37, 12, 27, 25, 34, 23, 17, 
    37, 23, 43, 56, 34, 20, 38, 32, 22, 11, 19, 20, 13, 16, 20, 
    30, 15, 31, 55, 45, 50, 22, 19, 9, 4, 16, 17, 8, 16, 24, 
    16, 16, 20, 50, 48, 31, 7, 11, 0, 8, 11, 16, 15, 17, 15, 
    
    -- channel=274
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=275
    7, 17, 24, 25, 24, 26, 28, 30, 31, 15, 30, 23, 28, 30, 30, 
    7, 15, 15, 24, 23, 17, 20, 26, 17, 20, 27, 28, 28, 28, 27, 
    7, 10, 22, 20, 14, 16, 13, 9, 14, 31, 19, 28, 28, 28, 29, 
    28, 35, 18, 16, 12, 18, 24, 15, 14, 17, 18, 27, 21, 17, 30, 
    29, 29, 26, 26, 13, 14, 12, 13, 13, 17, 20, 27, 26, 28, 29, 
    29, 26, 25, 31, 13, 11, 14, 20, 14, 19, 21, 26, 31, 37, 34, 
    31, 30, 19, 31, 21, 22, 9, 17, 11, 17, 21, 26, 31, 36, 41, 
    29, 26, 21, 17, 14, 17, 14, 8, 22, 15, 17, 7, 34, 23, 40, 
    32, 27, 20, 11, 23, 22, 18, 12, 13, 27, 14, 35, 13, 22, 33, 
    34, 29, 18, 21, 18, 9, 18, 26, 26, 20, 12, 22, 28, 17, 22, 
    33, 26, 24, 23, 23, 17, 16, 16, 19, 8, 28, 19, 18, 20, 14, 
    30, 29, 22, 18, 15, 19, 22, 19, 16, 22, 21, 17, 17, 19, 23, 
    31, 29, 27, 20, 9, 22, 16, 18, 16, 20, 19, 19, 9, 21, 20, 
    31, 34, 32, 20, 19, 20, 11, 20, 16, 23, 17, 20, 16, 20, 19, 
    30, 35, 27, 19, 23, 14, 15, 18, 16, 23, 19, 18, 23, 15, 19, 
    
    -- channel=276
    0, 3, 20, 38, 47, 32, 37, 35, 30, 47, 6, 43, 47, 45, 45, 
    0, 6, 0, 33, 49, 64, 45, 44, 52, 43, 18, 60, 59, 55, 54, 
    0, 0, 0, 37, 52, 75, 44, 40, 42, 26, 45, 60, 68, 67, 66, 
    9, 0, 24, 60, 41, 66, 58, 38, 23, 40, 56, 57, 88, 85, 61, 
    47, 46, 55, 53, 35, 68, 69, 55, 29, 42, 51, 57, 82, 74, 52, 
    56, 59, 57, 57, 47, 73, 64, 44, 33, 45, 59, 54, 83, 71, 46, 
    57, 57, 66, 31, 51, 51, 63, 45, 54, 43, 60, 56, 82, 76, 70, 
    64, 57, 65, 21, 76, 64, 56, 72, 33, 63, 63, 66, 58, 82, 67, 
    59, 45, 47, 63, 65, 65, 76, 56, 44, 56, 37, 42, 37, 52, 50, 
    58, 59, 63, 63, 67, 78, 70, 68, 67, 40, 52, 30, 40, 45, 47, 
    63, 69, 49, 73, 69, 71, 50, 72, 65, 60, 32, 39, 47, 48, 43, 
    66, 57, 49, 79, 82, 70, 57, 64, 68, 52, 28, 48, 42, 53, 37, 
    64, 52, 46, 72, 71, 63, 48, 62, 57, 45, 29, 43, 46, 35, 35, 
    64, 49, 39, 63, 67, 66, 58, 46, 44, 32, 26, 36, 35, 26, 35, 
    54, 34, 43, 54, 72, 68, 55, 32, 33, 20, 29, 30, 30, 32, 33, 
    
    -- channel=277
    0, 9, 12, 0, 0, 7, 1, 0, 0, 0, 5, 0, 0, 1, 3, 
    0, 1, 24, 8, 0, 0, 5, 0, 0, 0, 0, 0, 0, 1, 3, 
    0, 0, 13, 1, 0, 0, 9, 25, 22, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 7, 0, 0, 32, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 30, 29, 11, 
    0, 0, 0, 0, 0, 11, 1, 0, 0, 0, 4, 7, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 7, 6, 0, 1, 7, 0, 0, 4, 4, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 2, 0, 2, 1, 0, 0, 
    0, 0, 0, 0, 4, 27, 10, 8, 9, 4, 4, 4, 12, 10, 0, 
    0, 0, 0, 0, 0, 0, 6, 11, 12, 7, 2, 2, 3, 4, 0, 
    3, 0, 0, 1, 0, 0, 11, 10, 7, 3, 3, 1, 0, 0, 6, 
    
    -- channel=278
    0, 19, 72, 65, 56, 67, 62, 62, 57, 12, 55, 63, 74, 72, 73, 
    0, 5, 68, 75, 64, 46, 72, 71, 72, 49, 44, 78, 79, 79, 80, 
    0, 0, 49, 60, 89, 62, 54, 69, 81, 71, 50, 86, 86, 84, 80, 
    0, 0, 15, 56, 96, 83, 42, 36, 42, 59, 81, 91, 94, 87, 95, 
    51, 42, 63, 55, 70, 90, 79, 57, 51, 63, 78, 90, 98, 70, 69, 
    73, 70, 74, 61, 71, 83, 78, 57, 45, 57, 72, 96, 95, 68, 51, 
    69, 72, 65, 83, 65, 74, 62, 70, 55, 66, 69, 91, 97, 86, 53, 
    64, 79, 73, 88, 71, 77, 78, 52, 86, 56, 72, 89, 119, 95, 89, 
    61, 66, 86, 69, 94, 77, 66, 62, 53, 70, 68, 46, 65, 94, 90, 
    66, 58, 83, 88, 82, 98, 107, 77, 42, 66, 62, 67, 55, 54, 65, 
    78, 64, 88, 80, 83, 71, 84, 93, 88, 59, 69, 57, 69, 66, 55, 
    76, 68, 80, 97, 92, 91, 74, 83, 77, 62, 52, 66, 75, 61, 54, 
    71, 61, 75, 94, 87, 85, 87, 84, 78, 60, 59, 63, 63, 72, 54, 
    68, 52, 64, 91, 80, 68, 70, 74, 63, 53, 51, 55, 49, 52, 60, 
    68, 53, 49, 94, 85, 72, 68, 66, 49, 43, 49, 52, 47, 44, 60, 
    
    -- channel=279
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 12, 2, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=280
    9, 44, 106, 95, 95, 97, 101, 106, 104, 57, 89, 123, 119, 120, 116, 
    9, 29, 93, 91, 120, 98, 102, 119, 115, 67, 128, 140, 133, 128, 121, 
    9, 17, 84, 100, 134, 102, 71, 82, 78, 95, 142, 145, 147, 148, 144, 
    71, 80, 136, 96, 125, 125, 107, 81, 77, 104, 135, 158, 157, 144, 147, 
    127, 138, 140, 90, 122, 127, 116, 78, 81, 96, 132, 171, 169, 138, 140, 
    139, 136, 137, 111, 124, 119, 102, 80, 100, 106, 126, 170, 175, 155, 138, 
    142, 136, 105, 129, 115, 117, 105, 97, 107, 113, 128, 169, 177, 175, 149, 
    137, 129, 94, 129, 127, 122, 109, 104, 110, 106, 117, 105, 159, 164, 163, 
    138, 118, 116, 124, 144, 150, 132, 102, 90, 99, 117, 93, 100, 116, 148, 
    150, 133, 136, 135, 135, 132, 137, 129, 117, 117, 90, 95, 104, 103, 103, 
    155, 133, 142, 144, 146, 119, 127, 129, 123, 95, 88, 104, 110, 91, 88, 
    152, 136, 143, 147, 140, 109, 133, 129, 122, 82, 102, 98, 112, 98, 84, 
    148, 132, 139, 146, 119, 75, 127, 116, 100, 81, 95, 90, 86, 86, 90, 
    141, 127, 130, 151, 123, 116, 101, 97, 82, 67, 88, 86, 74, 84, 98, 
    118, 126, 111, 144, 135, 118, 80, 80, 65, 77, 78, 87, 80, 86, 86, 
    
    -- channel=281
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=282
    15, 8, 31, 25, 25, 26, 32, 30, 29, 33, 6, 29, 34, 34, 34, 
    16, 12, 22, 13, 13, 19, 15, 19, 19, 23, 20, 20, 24, 27, 28, 
    17, 16, 15, 21, 0, 15, 10, 8, 6, 9, 17, 5, 11, 14, 19, 
    47, 28, 35, 19, 0, 7, 25, 22, 15, 6, 7, 4, 9, 11, 3, 
    23, 25, 16, 19, 2, 0, 9, 14, 11, 3, 4, 7, 8, 17, 11, 
    15, 12, 14, 19, 6, 1, 6, 8, 15, 8, 6, 1, 6, 20, 20, 
    16, 12, 15, 17, 9, 1, 11, 2, 12, 5, 6, 5, 6, 12, 19, 
    16, 9, 25, 10, 9, 5, 0, 16, 4, 7, 10, 0, 0, 7, 8, 
    20, 8, 14, 15, 2, 9, 9, 13, 9, 13, 18, 30, 3, 0, 2, 
    15, 14, 7, 11, 2, 0, 0, 7, 30, 18, 15, 19, 23, 23, 13, 
    10, 14, 0, 9, 10, 10, 1, 2, 6, 19, 13, 19, 16, 16, 20, 
    9, 15, 1, 1, 7, 6, 15, 10, 12, 18, 20, 14, 13, 20, 19, 
    12, 15, 3, 1, 9, 4, 13, 10, 12, 19, 16, 14, 11, 10, 20, 
    14, 20, 5, 0, 8, 28, 16, 15, 17, 14, 18, 17, 18, 16, 18, 
    10, 20, 9, 0, 5, 14, 14, 16, 21, 20, 16, 19, 20, 22, 14, 
    
    -- channel=283
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=284
    2, 0, 0, 3, 0, 0, 0, 0, 28, 49, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 90, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 0, 0, 17, 0, 34, 31, 23, 0, 0, 0, 0, 0, 12, 0, 
    33, 0, 0, 62, 0, 0, 20, 51, 0, 0, 0, 0, 0, 43, 0, 
    0, 0, 0, 29, 0, 0, 29, 23, 0, 0, 0, 0, 0, 46, 0, 
    0, 0, 23, 0, 0, 0, 25, 0, 2, 0, 0, 0, 0, 14, 19, 
    7, 0, 62, 0, 8, 0, 15, 0, 0, 0, 0, 0, 0, 1, 0, 
    35, 0, 13, 0, 0, 0, 9, 54, 0, 13, 0, 29, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 25, 27, 0, 16, 0, 0, 0, 0, 
    0, 19, 0, 0, 0, 32, 0, 0, 26, 19, 0, 0, 0, 18, 0, 
    0, 35, 0, 0, 0, 29, 0, 0, 5, 55, 0, 0, 0, 13, 16, 
    0, 15, 0, 0, 41, 0, 0, 0, 19, 28, 0, 0, 0, 0, 3, 
    8, 17, 0, 0, 37, 0, 0, 1, 14, 9, 0, 0, 16, 0, 0, 
    8, 8, 0, 0, 11, 11, 30, 0, 27, 0, 0, 0, 9, 0, 0, 
    
    -- channel=285
    0, 18, 48, 34, 32, 42, 39, 39, 28, 3, 34, 36, 42, 43, 43, 
    0, 6, 53, 37, 24, 18, 35, 39, 33, 19, 25, 36, 39, 43, 43, 
    0, 1, 48, 28, 32, 12, 24, 38, 39, 33, 25, 41, 36, 35, 34, 
    0, 6, 12, 23, 39, 23, 7, 13, 21, 26, 38, 37, 30, 31, 44, 
    26, 17, 34, 23, 30, 30, 24, 16, 21, 24, 40, 40, 39, 36, 41, 
    36, 35, 38, 25, 27, 25, 27, 21, 16, 19, 33, 49, 43, 36, 37, 
    39, 39, 36, 41, 27, 28, 18, 20, 19, 21, 29, 47, 44, 40, 31, 
    37, 36, 25, 51, 21, 24, 25, 7, 42, 23, 31, 48, 61, 43, 43, 
    34, 32, 30, 32, 31, 22, 13, 19, 31, 28, 34, 23, 49, 56, 54, 
    38, 23, 29, 33, 32, 35, 34, 24, 8, 30, 32, 38, 27, 29, 41, 
    40, 26, 39, 32, 31, 25, 38, 33, 32, 26, 37, 28, 29, 31, 27, 
    40, 33, 35, 32, 33, 32, 32, 32, 29, 29, 29, 29, 34, 26, 28, 
    39, 40, 36, 33, 29, 35, 44, 36, 35, 27, 34, 29, 31, 37, 27, 
    39, 39, 38, 36, 27, 13, 37, 36, 33, 30, 30, 28, 25, 30, 30, 
    41, 42, 30, 40, 30, 28, 30, 35, 27, 26, 29, 28, 26, 23, 33, 
    
    -- channel=286
    0, 0, 39, 43, 36, 37, 41, 39, 48, 30, 0, 36, 49, 49, 52, 
    0, 0, 22, 40, 40, 37, 44, 45, 57, 68, 0, 58, 59, 56, 56, 
    0, 0, 0, 32, 46, 69, 32, 39, 59, 41, 19, 61, 65, 62, 62, 
    6, 0, 0, 58, 41, 74, 42, 31, 23, 11, 62, 55, 73, 80, 70, 
    68, 19, 60, 65, 23, 62, 68, 56, 28, 20, 50, 56, 85, 93, 58, 
    70, 59, 70, 66, 37, 58, 69, 48, 29, 22, 40, 59, 86, 92, 61, 
    69, 62, 67, 56, 49, 49, 61, 30, 49, 36, 46, 56, 85, 90, 65, 
    75, 62, 72, 25, 65, 53, 64, 43, 54, 42, 61, 53, 81, 93, 82, 
    81, 50, 61, 27, 74, 55, 53, 67, 16, 55, 55, 40, 25, 84, 57, 
    82, 53, 59, 62, 59, 75, 79, 66, 41, 42, 54, 45, 32, 41, 34, 
    77, 73, 58, 62, 64, 72, 49, 64, 78, 56, 48, 33, 42, 54, 41, 
    74, 85, 45, 71, 74, 69, 47, 60, 65, 67, 22, 46, 48, 53, 45, 
    74, 80, 51, 72, 81, 43, 53, 63, 67, 53, 32, 45, 45, 50, 39, 
    75, 73, 45, 68, 79, 38, 54, 55, 55, 39, 29, 39, 43, 23, 41, 
    72, 67, 41, 60, 72, 68, 60, 42, 45, 23, 32, 37, 38, 24, 38, 
    
    -- channel=287
    16, 70, 42, 19, 23, 32, 27, 28, 6, 0, 51, 27, 25, 27, 25, 
    17, 50, 59, 25, 5, 12, 24, 26, 15, 0, 61, 16, 18, 22, 22, 
    17, 28, 70, 30, 18, 0, 16, 33, 19, 14, 33, 20, 9, 12, 11, 
    0, 27, 46, 10, 31, 0, 0, 1, 17, 40, 12, 27, 2, 1, 20, 
    0, 27, 15, 0, 36, 6, 0, 0, 18, 30, 22, 30, 5, 0, 34, 
    12, 18, 14, 2, 23, 6, 0, 0, 12, 23, 21, 35, 6, 0, 22, 
    16, 18, 9, 19, 10, 11, 0, 14, 1, 16, 19, 35, 11, 0, 2, 
    12, 22, 0, 42, 0, 7, 0, 7, 18, 16, 14, 40, 32, 6, 14, 
    1, 22, 3, 31, 1, 0, 0, 0, 39, 9, 14, 9, 52, 21, 41, 
    3, 14, 15, 8, 15, 11, 2, 0, 0, 22, 10, 22, 21, 16, 37, 
    10, 3, 21, 9, 6, 0, 26, 11, 0, 7, 19, 23, 19, 8, 19, 
    15, 0, 31, 5, 5, 0, 19, 10, 6, 0, 34, 16, 19, 8, 10, 
    12, 10, 32, 6, 0, 17, 25, 14, 7, 7, 31, 16, 21, 18, 15, 
    10, 12, 37, 12, 0, 12, 17, 17, 12, 17, 27, 19, 11, 31, 19, 
    15, 17, 34, 22, 0, 5, 7, 22, 10, 31, 23, 21, 13, 26, 23, 
    
    -- channel=288
    50, 50, 46, 25, 44, 47, 49, 54, 54, 48, 45, 55, 45, 43, 41, 
    52, 52, 39, 0, 13, 20, 16, 15, 29, 42, 47, 57, 52, 34, 59, 
    51, 52, 38, 0, 24, 15, 14, 4, 3, 11, 58, 58, 40, 32, 56, 
    52, 45, 41, 0, 42, 40, 3, 8, 12, 18, 16, 61, 51, 36, 39, 
    54, 44, 7, 0, 25, 8, 1, 8, 12, 13, 12, 53, 60, 46, 55, 
    62, 35, 28, 0, 16, 14, 0, 0, 1, 9, 6, 31, 68, 52, 52, 
    54, 24, 31, 13, 11, 1, 0, 0, 7, 3, 6, 27, 42, 49, 61, 
    45, 2, 63, 10, 0, 9, 7, 0, 0, 3, 0, 0, 26, 23, 75, 
    38, 0, 46, 0, 27, 16, 22, 16, 34, 39, 21, 29, 35, 15, 69, 
    39, 0, 29, 0, 9, 0, 7, 26, 11, 13, 4, 11, 16, 0, 67, 
    44, 0, 14, 4, 0, 18, 32, 0, 41, 5, 13, 41, 0, 31, 49, 
    30, 0, 34, 22, 0, 0, 8, 0, 29, 22, 23, 14, 0, 7, 65, 
    30, 11, 14, 15, 0, 0, 1, 6, 16, 73, 32, 0, 0, 23, 55, 
    31, 17, 3, 10, 7, 0, 5, 9, 17, 24, 29, 0, 0, 24, 51, 
    18, 17, 5, 0, 7, 0, 6, 9, 11, 14, 19, 3, 0, 22, 63, 
    
    -- channel=289
    63, 59, 57, 44, 43, 48, 63, 69, 68, 68, 62, 61, 64, 70, 59, 
    65, 65, 68, 32, 17, 11, 10, 18, 28, 39, 53, 55, 58, 61, 61, 
    61, 61, 60, 18, 7, 17, 14, 14, 11, 11, 40, 62, 55, 48, 54, 
    61, 59, 46, 32, 22, 40, 26, 16, 20, 33, 26, 42, 54, 66, 41, 
    59, 62, 32, 7, 12, 5, 9, 12, 17, 13, 26, 47, 57, 63, 62, 
    47, 57, 27, 13, 0, 0, 6, 0, 0, 0, 13, 9, 45, 61, 61, 
    36, 33, 14, 15, 15, 10, 5, 3, 10, 17, 4, 8, 22, 37, 53, 
    31, 7, 13, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 
    44, 20, 13, 5, 0, 22, 14, 19, 34, 41, 44, 40, 34, 26, 31, 
    41, 13, 8, 0, 0, 0, 0, 0, 1, 0, 0, 0, 11, 0, 5, 
    39, 24, 8, 0, 0, 0, 2, 1, 0, 1, 0, 1, 11, 6, 11, 
    31, 2, 5, 19, 6, 0, 0, 0, 5, 10, 21, 25, 0, 0, 0, 
    23, 24, 21, 19, 3, 3, 0, 0, 0, 39, 54, 40, 0, 0, 1, 
    27, 26, 13, 19, 5, 1, 0, 0, 1, 2, 3, 21, 0, 0, 0, 
    21, 19, 22, 10, 2, 1, 0, 0, 0, 0, 0, 14, 0, 0, 4, 
    
    -- channel=290
    4, 3, 1, 0, 0, 0, 10, 16, 0, 0, 0, 0, 26, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 66, 0, 20, 32, 44, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 45, 0, 0, 3, 0, 0, 5, 0, 0, 0, 18, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 2, 0, 0, 36, 51, 
    0, 0, 26, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 43, 0, 0, 0, 0, 4, 69, 93, 79, 113, 107, 41, 0, 0, 
    4, 38, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 68, 2, 11, 0, 0, 21, 10, 0, 7, 0, 11, 0, 6, 0, 
    0, 39, 0, 35, 44, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 
    0, 113, 28, 0, 41, 27, 0, 0, 0, 0, 28, 53, 8, 0, 0, 
    0, 0, 17, 0, 0, 38, 11, 1, 0, 0, 0, 15, 19, 0, 0, 
    0, 0, 19, 0, 0, 14, 13, 7, 0, 0, 0, 0, 26, 0, 0, 
    
    -- channel=291
    29, 29, 33, 12, 32, 29, 25, 20, 40, 39, 33, 43, 13, 19, 5, 
    43, 43, 37, 0, 57, 69, 60, 73, 84, 71, 41, 51, 45, 22, 38, 
    49, 49, 40, 0, 50, 38, 28, 21, 35, 45, 68, 51, 32, 20, 47, 
    49, 49, 34, 0, 73, 66, 32, 56, 50, 41, 46, 77, 35, 8, 25, 
    52, 44, 31, 8, 77, 57, 48, 58, 59, 52, 49, 71, 55, 24, 4, 
    65, 46, 7, 0, 63, 51, 39, 53, 58, 57, 65, 70, 78, 48, 50, 
    59, 39, 40, 0, 20, 43, 46, 34, 43, 56, 31, 58, 90, 79, 67, 
    54, 8, 51, 18, 40, 33, 28, 25, 45, 47, 27, 49, 74, 64, 108, 
    22, 0, 58, 5, 42, 29, 30, 5, 0, 0, 0, 0, 9, 30, 102, 
    32, 0, 69, 0, 50, 21, 44, 49, 58, 55, 53, 56, 68, 20, 83, 
    42, 0, 15, 8, 5, 32, 26, 0, 68, 17, 29, 44, 2, 33, 60, 
    49, 0, 52, 10, 0, 12, 52, 8, 55, 37, 38, 54, 0, 62, 63, 
    55, 0, 4, 47, 0, 0, 4, 11, 13, 61, 23, 5, 0, 22, 63, 
    48, 48, 15, 45, 23, 0, 0, 4, 20, 80, 63, 21, 0, 30, 65, 
    50, 42, 23, 16, 27, 4, 0, 8, 16, 29, 51, 33, 0, 29, 65, 
    
    -- channel=292
    6, 4, 9, 15, 5, 7, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    8, 8, 11, 32, 38, 42, 45, 44, 30, 13, 2, 1, 2, 1, 0, 
    12, 12, 17, 49, 51, 54, 58, 59, 63, 55, 12, 0, 7, 4, 0, 
    12, 13, 22, 55, 35, 31, 48, 64, 58, 51, 36, 8, 8, 2, 0, 
    11, 15, 35, 63, 45, 55, 66, 62, 57, 56, 51, 19, 3, 11, 5, 
    11, 17, 25, 55, 48, 59, 65, 58, 59, 56, 49, 32, 14, 12, 12, 
    14, 26, 25, 36, 44, 57, 57, 56, 48, 42, 43, 34, 30, 23, 8, 
    8, 35, 10, 25, 54, 61, 63, 52, 39, 40, 43, 30, 37, 48, 17, 
    14, 29, 3, 50, 32, 23, 22, 30, 18, 11, 14, 14, 15, 30, 11, 
    19, 42, 18, 37, 28, 46, 45, 37, 46, 57, 57, 54, 47, 55, 19, 
    21, 41, 23, 31, 35, 30, 29, 44, 31, 48, 47, 34, 52, 28, 18, 
    35, 55, 20, 25, 35, 26, 30, 40, 12, 22, 21, 22, 42, 35, 23, 
    39, 44, 27, 31, 39, 30, 20, 21, 24, 0, 3, 24, 31, 23, 19, 
    39, 42, 43, 33, 34, 34, 19, 19, 15, 26, 45, 50, 31, 20, 26, 
    47, 47, 47, 42, 32, 31, 24, 25, 27, 31, 33, 39, 29, 23, 24, 
    
    -- channel=293
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=294
    11, 11, 3, 0, 0, 18, 41, 63, 24, 0, 0, 0, 20, 22, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 35, 39, 39, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 11, 0, 0, 3, 29, 0, 0, 0, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 75, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 4, 0, 0, 0, 0, 15, 58, 141, 147, 132, 150, 118, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 41, 0, 0, 0, 0, 21, 0, 19, 0, 
    0, 0, 0, 52, 17, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 63, 66, 0, 4, 14, 0, 0, 0, 72, 67, 29, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 14, 15, 10, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 11, 9, 0, 0, 0, 0, 5, 0, 20, 
    
    -- channel=295
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 34, 5, 0, 0, 0, 0, 42, 0, 0, 0, 13, 
    0, 0, 0, 0, 35, 18, 0, 0, 0, 8, 0, 27, 0, 0, 0, 
    0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 
    5, 0, 0, 0, 22, 6, 0, 0, 0, 0, 0, 3, 28, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 14, 3, 
    0, 0, 41, 0, 0, 0, 0, 0, 0, 5, 0, 0, 26, 2, 57, 
    0, 0, 0, 0, 21, 0, 4, 4, 10, 7, 0, 5, 4, 0, 45, 
    0, 0, 21, 0, 15, 0, 0, 14, 0, 0, 0, 0, 2, 0, 53, 
    0, 0, 0, 0, 0, 26, 30, 0, 56, 0, 0, 34, 0, 15, 23, 
    0, 0, 49, 0, 0, 0, 0, 0, 20, 3, 4, 0, 0, 10, 53, 
    0, 0, 0, 0, 0, 0, 0, 6, 16, 72, 0, 0, 0, 26, 40, 
    0, 0, 0, 0, 0, 0, 2, 5, 5, 12, 14, 0, 0, 22, 42, 
    0, 0, 0, 0, 0, 0, 0, 1, 3, 3, 4, 3, 0, 21, 52, 
    
    -- channel=296
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=297
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=298
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 52, 60, 77, 97, 89, 61, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 18, 0, 0, 9, 22, 
    0, 0, 0, 0, 1, 0, 0, 8, 0, 0, 0, 33, 0, 0, 2, 
    0, 0, 40, 20, 8, 29, 27, 8, 11, 11, 0, 1, 0, 0, 0, 
    13, 7, 0, 0, 38, 5, 3, 26, 30, 17, 40, 29, 4, 0, 0, 
    6, 27, 25, 0, 0, 1, 7, 0, 5, 24, 22, 44, 77, 71, 3, 
    13, 40, 0, 0, 22, 0, 0, 14, 54, 49, 34, 65, 61, 39, 27, 
    0, 0, 2, 55, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 46, 0, 36, 13, 37, 49, 35, 44, 53, 47, 49, 29, 24, 
    0, 0, 0, 0, 3, 15, 0, 0, 16, 0, 0, 0, 1, 0, 9, 
    7, 16, 20, 0, 0, 11, 75, 36, 46, 25, 0, 39, 29, 56, 27, 
    2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 7, 0, 8, 0, 0, 0, 0, 0, 57, 53, 12, 0, 0, 6, 
    9, 0, 0, 13, 4, 0, 0, 0, 0, 4, 27, 14, 0, 0, 0, 
    
    -- channel=299
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=300
    204, 198, 197, 173, 145, 154, 167, 182, 198, 206, 201, 197, 207, 188, 187, 
    219, 219, 217, 165, 108, 101, 108, 120, 129, 153, 176, 186, 199, 195, 174, 
    220, 219, 215, 171, 80, 112, 113, 120, 107, 104, 124, 192, 197, 175, 149, 
    220, 217, 199, 172, 83, 147, 163, 130, 133, 133, 142, 148, 197, 187, 147, 
    215, 219, 175, 132, 81, 108, 126, 113, 121, 129, 145, 139, 196, 218, 191, 
    186, 208, 170, 128, 50, 88, 97, 85, 87, 92, 101, 114, 163, 222, 219, 
    165, 169, 125, 123, 86, 94, 94, 79, 74, 89, 89, 79, 118, 155, 204, 
    153, 124, 86, 131, 80, 78, 63, 53, 26, 26, 32, 19, 37, 82, 141, 
    167, 130, 82, 96, 57, 76, 96, 103, 94, 105, 129, 101, 98, 109, 121, 
    182, 133, 51, 62, 32, 55, 39, 49, 113, 89, 99, 90, 92, 94, 75, 
    174, 148, 60, 50, 27, 21, 58, 70, 41, 87, 70, 80, 87, 72, 88, 
    165, 127, 30, 83, 63, 9, 11, 43, 8, 86, 92, 88, 82, 33, 48, 
    146, 153, 83, 93, 73, 34, 1, 3, 14, 66, 157, 140, 44, 19, 52, 
    142, 147, 120, 84, 63, 53, 10, 12, 22, 54, 94, 124, 27, 12, 61, 
    139, 131, 126, 77, 50, 44, 27, 27, 30, 40, 52, 81, 36, 16, 64, 
    
    -- channel=301
    32, 32, 32, 23, 22, 24, 26, 30, 36, 34, 30, 31, 25, 25, 20, 
    42, 42, 39, 34, 45, 49, 50, 49, 45, 32, 26, 30, 30, 18, 23, 
    44, 45, 40, 32, 64, 74, 73, 72, 73, 58, 35, 34, 25, 9, 19, 
    44, 43, 41, 46, 66, 64, 74, 86, 82, 81, 58, 31, 27, 15, 10, 
    42, 42, 47, 53, 72, 78, 75, 84, 81, 82, 73, 49, 38, 30, 24, 
    36, 37, 33, 53, 60, 67, 72, 74, 73, 73, 75, 62, 48, 45, 44, 
    31, 26, 24, 34, 64, 74, 72, 65, 66, 66, 44, 43, 44, 42, 41, 
    16, 15, 16, 23, 62, 48, 48, 40, 39, 39, 37, 39, 50, 57, 50, 
    24, 17, 20, 26, 43, 39, 45, 36, 26, 34, 29, 26, 47, 53, 53, 
    30, 23, 21, 13, 42, 34, 41, 44, 50, 55, 54, 52, 51, 44, 53, 
    34, 21, 22, 21, 21, 28, 39, 35, 40, 43, 41, 42, 43, 38, 55, 
    48, 23, 22, 31, 19, 18, 32, 15, 32, 28, 38, 41, 18, 37, 44, 
    58, 31, 37, 39, 24, 14, 11, 14, 22, 33, 41, 30, 18, 21, 54, 
    55, 54, 43, 35, 35, 15, 10, 15, 20, 46, 47, 32, 9, 28, 57, 
    62, 59, 47, 35, 32, 19, 16, 18, 24, 31, 40, 31, 13, 25, 57, 
    
    -- channel=302
    20, 15, 12, 0, 8, 8, 13, 17, 21, 22, 17, 25, 15, 15, 12, 
    23, 24, 17, 0, 0, 0, 0, 0, 7, 13, 22, 23, 21, 9, 28, 
    23, 24, 13, 0, 0, 0, 0, 0, 0, 0, 19, 23, 10, 4, 27, 
    23, 17, 12, 0, 0, 0, 0, 0, 0, 0, 0, 27, 18, 6, 1, 
    24, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 23, 12, 15, 
    25, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 24, 24, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 24, 28, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=303
    9, 8, 14, 19, 11, 3, 0, 0, 11, 16, 18, 15, 0, 8, 1, 
    18, 17, 24, 38, 47, 53, 57, 64, 60, 36, 22, 18, 19, 17, 9, 
    24, 25, 23, 22, 32, 32, 30, 31, 42, 50, 18, 14, 21, 17, 17, 
    24, 28, 24, 36, 44, 32, 51, 60, 48, 41, 45, 30, 5, 3, 14, 
    23, 25, 51, 44, 50, 68, 57, 60, 60, 57, 46, 25, 13, 0, 0, 
    25, 33, 12, 44, 53, 48, 57, 64, 62, 61, 68, 48, 30, 24, 24, 
    25, 31, 30, 13, 30, 52, 54, 45, 48, 53, 39, 46, 55, 47, 23, 
    21, 31, 3, 23, 52, 36, 44, 52, 58, 50, 54, 60, 51, 53, 31, 
    6, 7, 20, 36, 30, 36, 17, 0, 0, 0, 0, 0, 0, 37, 35, 
    13, 30, 30, 15, 43, 32, 47, 50, 44, 58, 57, 53, 55, 42, 36, 
    20, 12, 16, 17, 25, 26, 6, 42, 26, 35, 33, 13, 44, 20, 30, 
    33, 36, 17, 6, 13, 28, 60, 26, 45, 21, 21, 54, 25, 51, 31, 
    37, 0, 13, 33, 13, 15, 15, 16, 15, 2, 6, 17, 24, 12, 28, 
    36, 40, 33, 33, 29, 13, 7, 11, 17, 51, 48, 39, 14, 21, 32, 
    44, 37, 30, 32, 30, 17, 10, 13, 19, 28, 42, 29, 13, 19, 26, 
    
    -- channel=304
    198, 198, 196, 166, 154, 153, 161, 178, 207, 214, 210, 209, 188, 182, 167, 
    230, 229, 219, 163, 141, 148, 156, 172, 190, 196, 192, 205, 213, 192, 190, 
    237, 237, 216, 124, 94, 112, 116, 110, 108, 124, 164, 206, 202, 172, 176, 
    235, 232, 208, 134, 134, 177, 173, 159, 151, 149, 166, 193, 195, 164, 157, 
    236, 227, 194, 120, 125, 158, 149, 146, 157, 165, 159, 178, 217, 194, 164, 
    224, 221, 163, 103, 94, 114, 116, 124, 125, 133, 152, 172, 212, 237, 236, 
    197, 180, 150, 103, 97, 122, 120, 97, 108, 126, 105, 123, 178, 211, 235, 
    178, 128, 119, 128, 100, 78, 62, 66, 68, 65, 62, 76, 102, 137, 206, 
    166, 103, 122, 92, 83, 106, 111, 69, 49, 72, 69, 41, 87, 132, 194, 
    182, 104, 89, 50, 64, 64, 70, 111, 136, 127, 131, 123, 132, 101, 153, 
    186, 98, 59, 43, 28, 42, 62, 65, 78, 84, 75, 86, 82, 91, 145, 
    184, 94, 56, 68, 33, 25, 71, 43, 75, 110, 103, 134, 78, 68, 125, 
    173, 96, 73, 101, 52, 9, 1, 7, 24, 107, 151, 108, 35, 30, 114, 
    165, 161, 118, 92, 71, 27, 0, 11, 42, 109, 139, 99, 14, 38, 122, 
    161, 146, 114, 74, 62, 35, 17, 21, 34, 57, 91, 74, 17, 33, 122, 
    
    -- channel=305
    70, 72, 69, 39, 49, 53, 61, 72, 72, 65, 59, 64, 65, 54, 48, 
    79, 79, 67, 27, 30, 36, 27, 22, 32, 35, 44, 63, 62, 39, 56, 
    80, 79, 68, 39, 61, 75, 80, 74, 61, 38, 55, 70, 52, 27, 35, 
    80, 76, 67, 44, 66, 77, 72, 71, 79, 78, 47, 55, 61, 47, 27, 
    78, 73, 45, 35, 63, 56, 58, 67, 65, 69, 70, 66, 78, 76, 82, 
    71, 61, 64, 32, 31, 58, 53, 46, 45, 53, 48, 51, 78, 80, 80, 
    60, 40, 35, 42, 64, 55, 53, 43, 49, 43, 25, 31, 35, 49, 76, 
    49, 9, 45, 46, 40, 37, 32, 16, 1, 6, 1, 0, 22, 45, 75, 
    60, 24, 37, 0, 36, 31, 46, 49, 66, 71, 68, 63, 76, 54, 62, 
    64, 13, 13, 6, 13, 15, 14, 30, 34, 38, 30, 32, 40, 20, 60, 
    64, 24, 14, 12, 0, 11, 51, 13, 35, 38, 35, 62, 22, 50, 56, 
    64, 2, 20, 42, 4, 0, 0, 0, 7, 22, 42, 25, 0, 1, 50, 
    68, 63, 47, 36, 20, 0, 0, 0, 4, 68, 69, 40, 0, 11, 61, 
    69, 56, 40, 30, 22, 0, 0, 0, 13, 17, 36, 16, 0, 17, 59, 
    61, 61, 46, 13, 16, 4, 3, 7, 11, 18, 25, 15, 0, 15, 72, 
    
    -- channel=306
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 2, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 21, 0, 0, 11, 41, 15, 0, 14, 37, 4, 5, 29, 0, 0, 
    0, 0, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 23, 11, 0, 23, 6, 27, 26, 0, 39, 0, 
    0, 17, 0, 10, 1, 15, 0, 0, 38, 0, 12, 0, 0, 0, 0, 
    0, 36, 10, 0, 0, 0, 0, 80, 0, 12, 0, 0, 65, 12, 0, 
    0, 5, 0, 0, 17, 0, 6, 5, 2, 0, 0, 0, 7, 8, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 22, 27, 29, 0, 0, 
    0, 0, 0, 8, 0, 14, 0, 0, 0, 0, 0, 32, 5, 0, 0, 
    
    -- channel=307
    24, 27, 17, 16, 14, 13, 19, 23, 21, 22, 22, 24, 31, 25, 34, 
    19, 20, 11, 6, 0, 0, 0, 0, 0, 16, 24, 21, 22, 26, 29, 
    17, 17, 13, 6, 0, 0, 0, 0, 0, 0, 21, 18, 15, 27, 29, 
    18, 14, 18, 0, 0, 0, 0, 0, 0, 0, 5, 14, 27, 18, 25, 
    19, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 21, 28, 30, 
    16, 6, 16, 0, 0, 0, 0, 0, 0, 0, 0, 10, 15, 18, 17, 
    8, 5, 4, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 
    1, 5, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    9, 9, 1, 0, 0, 0, 1, 11, 15, 14, 13, 17, 2, 0, 5, 
    13, 2, 0, 13, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    8, 8, 1, 3, 0, 0, 9, 0, 6, 0, 0, 11, 0, 3, 7, 
    0, 0, 0, 3, 1, 0, 0, 6, 0, 5, 0, 0, 14, 0, 18, 
    0, 20, 0, 0, 7, 0, 2, 3, 6, 4, 2, 0, 0, 7, 5, 
    0, 0, 0, 0, 0, 4, 6, 3, 0, 0, 1, 0, 8, 0, 4, 
    0, 0, 0, 0, 0, 3, 5, 3, 1, 0, 0, 0, 5, 2, 7, 
    
    -- channel=308
    84, 81, 81, 87, 58, 68, 65, 74, 82, 86, 87, 78, 81, 74, 66, 
    99, 98, 100, 109, 68, 71, 86, 86, 80, 74, 68, 76, 82, 81, 53, 
    102, 102, 99, 96, 36, 58, 70, 72, 68, 77, 46, 75, 92, 73, 50, 
    101, 99, 99, 95, 54, 88, 106, 88, 82, 87, 103, 57, 79, 78, 66, 
    99, 100, 113, 82, 48, 93, 82, 82, 89, 93, 86, 77, 86, 83, 72, 
    86, 102, 83, 89, 38, 57, 76, 70, 66, 66, 71, 73, 70, 102, 101, 
    84, 88, 71, 54, 68, 80, 73, 66, 66, 73, 70, 61, 75, 88, 88, 
    77, 85, 34, 70, 53, 44, 39, 45, 31, 23, 37, 32, 31, 68, 58, 
    87, 83, 43, 66, 32, 60, 54, 43, 27, 45, 41, 25, 39, 80, 73, 
    86, 94, 20, 47, 21, 38, 34, 54, 68, 65, 70, 59, 56, 68, 53, 
    87, 85, 33, 22, 23, 9, 20, 64, 2, 47, 33, 17, 67, 33, 70, 
    95, 95, 0, 33, 43, 13, 27, 23, 28, 47, 42, 69, 64, 17, 43, 
    83, 70, 54, 38, 39, 21, 0, 0, 7, 10, 74, 64, 38, 3, 42, 
    86, 84, 74, 38, 38, 30, 0, 3, 15, 35, 57, 60, 19, 5, 44, 
    86, 80, 70, 51, 28, 23, 10, 9, 14, 24, 38, 32, 26, 1, 37, 
    
    -- channel=309
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 14, 23, 33, 29, 17, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 1, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    0, 0, 2, 4, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 12, 0, 0, 2, 5, 3, 13, 5, 6, 0, 0, 
    8, 15, 17, 0, 0, 0, 0, 0, 0, 0, 0, 6, 26, 30, 1, 
    8, 17, 12, 0, 6, 0, 4, 10, 20, 18, 15, 21, 19, 14, 16, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 18, 0, 6, 1, 11, 21, 6, 19, 20, 18, 16, 11, 10, 
    0, 0, 0, 0, 0, 6, 0, 0, 15, 0, 0, 0, 1, 0, 0, 
    0, 0, 9, 0, 0, 0, 29, 15, 11, 4, 0, 5, 7, 21, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 14, 25, 3, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 9, 7, 0, 0, 0, 
    
    -- channel=310
    89, 86, 93, 74, 83, 74, 66, 61, 79, 96, 90, 101, 82, 61, 67, 
    108, 107, 101, 79, 85, 97, 96, 107, 117, 109, 95, 99, 104, 80, 88, 
    116, 116, 110, 61, 70, 61, 65, 58, 59, 59, 94, 97, 91, 79, 77, 
    116, 114, 108, 78, 74, 100, 85, 96, 89, 78, 61, 113, 102, 64, 60, 
    118, 111, 100, 90, 77, 86, 104, 86, 88, 94, 92, 87, 108, 97, 68, 
    123, 111, 97, 47, 64, 81, 68, 78, 82, 82, 90, 97, 115, 116, 116, 
    105, 106, 92, 74, 44, 66, 81, 58, 64, 72, 58, 68, 102, 129, 127, 
    103, 77, 91, 65, 77, 59, 44, 41, 51, 57, 39, 52, 82, 89, 124, 
    88, 53, 62, 67, 57, 54, 68, 41, 7, 10, 19, 0, 19, 59, 104, 
    101, 47, 68, 34, 43, 48, 48, 76, 89, 84, 90, 87, 92, 68, 92, 
    104, 56, 21, 34, 15, 38, 44, 15, 75, 46, 52, 62, 33, 63, 69, 
    106, 52, 58, 32, 5, 11, 44, 54, 31, 78, 59, 59, 62, 46, 87, 
    106, 60, 13, 61, 37, 0, 1, 7, 15, 57, 60, 46, 13, 28, 59, 
    90, 95, 69, 58, 45, 15, 0, 2, 21, 59, 100, 62, 16, 23, 73, 
    96, 88, 64, 42, 39, 24, 6, 11, 19, 35, 59, 61, 2, 24, 70, 
    
    -- channel=311
    6, 5, 5, 0, 0, 5, 15, 11, 13, 9, 0, 3, 3, 0, 0, 
    13, 12, 10, 3, 12, 12, 5, 7, 6, 3, 0, 0, 2, 0, 0, 
    13, 12, 18, 6, 35, 45, 44, 44, 38, 12, 6, 8, 0, 0, 0, 
    13, 13, 7, 27, 34, 55, 47, 52, 56, 53, 24, 0, 4, 0, 0, 
    11, 12, 13, 22, 44, 32, 41, 52, 46, 44, 45, 21, 13, 16, 2, 
    3, 11, 11, 28, 27, 38, 38, 39, 41, 33, 36, 23, 6, 13, 13, 
    0, 5, 0, 11, 38, 42, 48, 38, 35, 45, 22, 11, 8, 6, 11, 
    4, 0, 0, 12, 30, 27, 20, 13, 14, 17, 3, 6, 14, 13, 17, 
    1, 0, 0, 0, 15, 13, 30, 41, 16, 20, 42, 24, 23, 30, 25, 
    9, 0, 5, 0, 15, 6, 7, 0, 25, 9, 15, 14, 20, 11, 7, 
    7, 10, 0, 3, 0, 8, 24, 9, 17, 15, 13, 22, 13, 11, 18, 
    19, 1, 9, 12, 7, 0, 0, 0, 0, 10, 23, 6, 0, 11, 0, 
    29, 22, 16, 21, 11, 0, 0, 0, 0, 14, 36, 29, 1, 2, 13, 
    24, 31, 17, 23, 13, 4, 0, 0, 1, 12, 5, 16, 0, 0, 18, 
    32, 31, 25, 17, 10, 5, 0, 1, 3, 6, 10, 20, 0, 2, 12, 
    
    -- channel=312
    166, 164, 160, 117, 123, 124, 138, 162, 171, 166, 161, 163, 161, 155, 145, 
    174, 174, 162, 84, 78, 85, 79, 82, 104, 127, 144, 164, 161, 146, 161, 
    174, 174, 152, 78, 80, 93, 91, 90, 81, 89, 132, 165, 150, 129, 141, 
    173, 169, 145, 73, 103, 112, 100, 94, 99, 102, 113, 147, 151, 143, 120, 
    172, 166, 104, 58, 85, 87, 78, 83, 92, 96, 109, 133, 166, 163, 162, 
    159, 150, 115, 54, 47, 73, 66, 61, 61, 78, 77, 102, 167, 174, 174, 
    138, 105, 89, 75, 74, 64, 63, 51, 61, 66, 56, 77, 106, 126, 172, 
    117, 55, 98, 85, 56, 53, 49, 36, 18, 19, 24, 20, 47, 81, 157, 
    122, 62, 96, 15, 70, 62, 70, 64, 99, 102, 98, 96, 108, 85, 125, 
    131, 52, 56, 32, 36, 38, 39, 64, 70, 73, 65, 68, 80, 44, 114, 
    133, 55, 53, 38, 20, 28, 68, 37, 61, 64, 63, 95, 40, 84, 97, 
    119, 32, 49, 78, 25, 19, 27, 13, 47, 60, 80, 80, 23, 32, 93, 
    110, 97, 76, 77, 46, 18, 11, 16, 27, 126, 121, 85, 12, 34, 94, 
    115, 96, 76, 63, 50, 23, 19, 26, 41, 59, 82, 62, 13, 39, 88, 
    97, 96, 82, 34, 44, 29, 29, 32, 35, 44, 54, 47, 15, 39, 109, 
    
    -- channel=313
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=314
    3, 4, 3, 4, 0, 4, 5, 12, 4, 0, 3, 0, 8, 13, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 7, 8, 0, 0, 0, 0, 0, 24, 19, 23, 27, 12, 0, 0, 
    0, 8, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 10, 1, 3, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 8, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 12, 0, 3, 16, 10, 7, 0, 1, 5, 13, 6, 0, 0, 
    0, 0, 0, 0, 0, 11, 13, 10, 6, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 5, 9, 7, 2, 0, 0, 0, 12, 0, 0, 
    
    -- channel=315
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=316
    0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 18, 
    0, 0, 7, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 
    0, 0, 25, 122, 0, 0, 0, 11, 0, 0, 0, 0, 1, 28, 0, 
    0, 0, 6, 129, 0, 0, 26, 0, 0, 0, 0, 0, 7, 23, 0, 
    0, 3, 41, 85, 0, 0, 17, 0, 0, 0, 10, 0, 0, 35, 0, 
    0, 17, 49, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 40, 0, 59, 0, 0, 20, 1, 0, 0, 7, 0, 0, 0, 0, 
    3, 60, 0, 48, 4, 20, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    15, 85, 0, 73, 0, 0, 1, 51, 0, 0, 51, 6, 0, 0, 0, 
    22, 110, 0, 55, 0, 14, 0, 0, 6, 0, 0, 0, 0, 31, 0, 
    0, 138, 0, 24, 4, 0, 0, 35, 0, 19, 0, 0, 33, 0, 0, 
    0, 139, 0, 0, 58, 0, 0, 70, 0, 5, 0, 0, 89, 0, 0, 
    0, 101, 0, 0, 53, 33, 0, 0, 0, 0, 5, 81, 43, 0, 0, 
    0, 13, 45, 11, 3, 61, 0, 0, 0, 0, 0, 81, 43, 0, 0, 
    0, 6, 34, 31, 0, 31, 1, 0, 0, 0, 0, 46, 37, 0, 0, 
    
    -- channel=317
    28, 25, 27, 22, 23, 23, 20, 14, 23, 33, 31, 37, 28, 26, 28, 
    30, 30, 27, 6, 15, 17, 20, 31, 36, 46, 41, 37, 38, 37, 38, 
    32, 32, 29, 0, 0, 0, 0, 0, 0, 7, 37, 34, 32, 38, 47, 
    32, 30, 27, 0, 0, 3, 0, 0, 0, 0, 4, 46, 37, 23, 29, 
    34, 30, 11, 0, 0, 0, 0, 0, 0, 0, 0, 21, 32, 27, 15, 
    42, 29, 9, 0, 5, 0, 0, 0, 0, 0, 4, 18, 39, 32, 33, 
    34, 30, 25, 6, 0, 0, 0, 0, 0, 0, 0, 10, 35, 43, 42, 
    28, 18, 30, 0, 0, 0, 0, 0, 1, 5, 0, 4, 15, 10, 47, 
    15, 0, 17, 15, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 
    23, 0, 24, 0, 3, 0, 4, 7, 15, 11, 14, 15, 14, 5, 23, 
    25, 0, 0, 0, 0, 5, 0, 0, 23, 0, 2, 8, 0, 0, 7, 
    16, 0, 17, 0, 0, 0, 11, 11, 4, 16, 3, 4, 2, 16, 19, 
    13, 0, 0, 8, 0, 0, 0, 0, 0, 11, 0, 0, 0, 3, 2, 
    4, 10, 0, 5, 0, 0, 0, 0, 0, 20, 26, 10, 0, 0, 6, 
    6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 0, 1, 6, 
    
    -- channel=318
    73, 64, 77, 70, 61, 51, 46, 42, 54, 80, 78, 79, 79, 58, 72, 
    81, 79, 91, 78, 44, 41, 43, 59, 67, 69, 81, 70, 81, 86, 71, 
    86, 86, 92, 86, 19, 20, 17, 20, 16, 15, 35, 68, 79, 83, 53, 
    85, 88, 83, 96, 11, 43, 56, 49, 45, 36, 22, 64, 83, 75, 46, 
    84, 92, 73, 86, 14, 31, 65, 36, 40, 42, 52, 25, 64, 82, 50, 
    74, 95, 83, 59, 11, 29, 33, 36, 37, 37, 49, 37, 55, 87, 85, 
    59, 86, 58, 73, 0, 22, 41, 21, 18, 28, 28, 13, 39, 72, 86, 
    63, 68, 35, 47, 40, 29, 19, 32, 28, 24, 30, 26, 16, 20, 41, 
    64, 57, 12, 70, 18, 28, 36, 18, 0, 0, 12, 0, 0, 25, 13, 
    76, 69, 23, 34, 1, 24, 4, 18, 47, 35, 49, 41, 42, 49, 0, 
    70, 81, 10, 21, 3, 5, 0, 15, 17, 31, 27, 15, 28, 28, 0, 
    63, 78, 12, 18, 15, 0, 9, 56, 0, 50, 27, 27, 64, 14, 0, 
    58, 63, 0, 38, 30, 5, 0, 0, 0, 0, 38, 63, 17, 0, 0, 
    45, 64, 58, 36, 24, 25, 0, 0, 0, 0, 47, 80, 16, 0, 0, 
    55, 48, 50, 32, 19, 18, 0, 0, 0, 5, 15, 56, 5, 0, 0, 
    
    -- channel=319
    0, 3, 0, 0, 4, 4, 1, 5, 10, 1, 4, 7, 0, 9, 0, 
    0, 0, 0, 0, 0, 4, 6, 6, 12, 17, 12, 14, 4, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 29, 9, 0, 0, 35, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 1, 26, 0, 0, 19, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 21, 7, 0, 0, 
    11, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 9, 24, 0, 0, 
    13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 17, 27, 14, 7, 
    1, 0, 24, 0, 0, 0, 0, 0, 4, 3, 0, 14, 21, 8, 33, 
    0, 0, 33, 0, 6, 2, 0, 0, 0, 0, 0, 0, 7, 0, 40, 
    0, 0, 22, 0, 14, 0, 12, 18, 0, 0, 0, 0, 0, 0, 45, 
    0, 0, 9, 0, 5, 14, 3, 0, 22, 0, 0, 4, 0, 0, 32, 
    0, 0, 18, 0, 0, 17, 33, 0, 50, 0, 0, 14, 0, 20, 45, 
    0, 0, 0, 0, 0, 0, 13, 16, 20, 38, 0, 0, 0, 16, 44, 
    0, 0, 0, 0, 0, 0, 12, 15, 18, 35, 7, 0, 0, 28, 33, 
    0, 0, 0, 0, 1, 0, 7, 8, 10, 11, 14, 0, 0, 23, 39, 
    
    
    others => 0);
end gold_package;
