library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -2193, 2019, -1031, 1628, 448, -1727, 1097, -480, -829, 207,

    -- weights
    -- filter=0 channel=0
    0, 0, 0, -1, -1, 0, 1, 0, -1, 1, 0, -1, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 1, 2, 0, -1, 1, -1, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, -2, 1, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 1, 0, 0, -2, -1, 0, 0, 0, 1, 0, 1, -1, -1, 0, -2, 1, 0, 1, 0, -1, 0, 1, 0, -3, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, -1, 2, 0, 0, 0, 0, 1, 0, -1, 0, -1, -2, 1, -1, 0, -2, -2, 0, 0, 0, -2, 0, -1, -1, -1, 0, 0, -2, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -2, -2, -2, 1, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, 0, 1, 1, 1, -1, 1, 0, 0, -1, 0, -1, 0, -1, 0, -2, -1, 0, -1, -1, -1, 0, -1, -1, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, 0, 1, -2, -2, -1, -1, 0, 0, -1, 1, -2, 0, -2, 0, 0, -1, 1, 1, -1, 2, 1, 0, -1, 0, 0, 0, 0, 1, 0, 2, -1, 0, 0, 1, 0, -2, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, -1, -1, 1, -1, -1, -1, -1, 1, -1, -1, 2, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 2, 0, -1, 0, -1, 1, -2, 0, -3, 0, -1, 0, -1, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, -2, -1, 1, -2, 0, 0, 1, 0, -1, -2, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -2, 1, 0, -2, 0, -1, 0, -1, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, 0, 1, 0, 1, -1, 1, 1, 0, 1, -1, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, -1, 2, 0, 1, 1, 0, 0, -1, -1, -2, -1, 0, 0, 0, -1, -1, 1, 0, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 1, 2, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, -1, -1, -1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 2, -1, -1, 0, 1, 1, -1, 0, 1, 0, -1, -2, -2, 0, -1, 0, 0, 2, 0, 0, 0, 2, 1, 0, 0, -1, 0, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, -3, -3, -1, -2, 0, 0, -1, 0, -1, 0, -1, 0, -1, 0, -1, 1, 0, -2, -1, -2, -1, 0, -2, 0, 0, -1, -1, 0, -1, 0, -2, -2, 0, -2, -1, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, 1, -1, -2, -2, -3, -2, 1, -1, -1, 0, 0, -2, 0, 0, 0, -1, 0, -1, 1, 1, 1, 0, 0, 0, -1, 0, -2, -2, 1, -3, -2, 0, 0, -2, -1, -1, 0, -2, 0, 0, -1, -1, 1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, -1, -2, 0, -2, -2, -1, -1, 1, 0, 0, 1, 1, 0, -1, 0, 1, 0, 0, -1, 0, 2, 0, -2, -1, 1, 0, -1, 0, 1, 1, 0, -1, -1, 0, -2, -3, -2, 0, -2, -2, 0, 0, -2, -1, 0, -1, 0, 1, 2, 0, 0, 1, 0, -1, 0, -1, -1, 1, 2, 0, 1, -1, -2, 1, 0, -2, -2, -1, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, -2, -1, 0, 1, 0, 0, -1, -2, -1, 0, 0, -2, 0, -1, -2, -2, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 0, 1, 0, -2, -1, -1, -1, -2, -1, -1, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 1, -1, 2, 0, 0, 0, 0, 1, -2, 0, 0, 0, 0, -3, -1, 0, 0, 0, -1, 0, 0, -1, 1, 1, -1, 0, 0, 0, 1, 0, 0, 1, 1, -1, 2, -1, 0, 0, -2, -1, -2, 1, -2, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, -2, -1, 1, 0, -1, 0, 0, 0, 1, -1, 0, -2, 0, 0, 1, 0, 0, 0, 1, -1, 2, -1, 0, 0, -1, 1, 0, 0, 1, 0, -1, -1, 0, 1, 1, -2, 0, 0, 1, 1, -1, 0, -1, 0, 1, 1, 1, 2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -2, 1, 0, -1, 0, 0, 1, 0, 1, 1, -1, -2, 0, 0, -1, 0, 0, 1, 1, 1, 3, 0, 3, 2, 0, 0, 1, 4, 3, 1, 4, 1, 1, 0, 1, 0, 0, 1, 0, -2, -3, -5, -3, -6, -7, -5, 1, 0, 1, 0, 1, 0, 1, 0, 0, -2, 0, 1, 1, 2, 0, 3, 0, 1, 3, 0, 1, 1, 3, 2, 0, -3, -4, -4, -3, -3, -2, 0, 0, -1, 0, 0, -1, 0, 0, -3, -2, 0, 0, -1, 0, 2, 0, 2, 3, 0, 4, 2, 1, 2, 0, 1, -1, -3, -3, -2, 0, -1, -1, 0, 0, 0, 1, -2, -4, -2, -3, -4, -2, 0, 0, 0, 2, 2, 2, 4, 2, 3, 1, 2, 0, 2, 0, -2, -1, 0, 1, 2, 0, 0, 2, 2, 0, 0, -2, -4, -1, -5, -1, -2, -2, -2, 0, 0, 2, 1, 2, 3, 4, 3, 0, 0, 0, -2, 0, -1, 0, 1, 1, 2, 0, 2, 1, 2, 0, -1, -2, -1, -4, -4, 0, -1, -1, 1, 0, 1, 5, 3, 3, 1, 0, 2, 0, 1, 1, 0, 0, 0, 2, 3, 0, 4, 2, 0, 0, -1, -1, -1, 0, -3, -2, -3, 0, 2, 1, 3, 4, 2, 3, 3, 4, 4, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 3, 2, 3, 0, 2, 0, -2, -3, 0, -2, 1, 2, 0, 2, 2, 4, 3, 2, 2, 0, 1, 1, 0, 0, -1, 1, 0, 1, 1, 0, 1, 1, 2, 1, 3, 0, -4, -2, -2, 0, 1, -1, 0, 0, 1, 1, 5, 5, 5, 4, 3, 2, 0, -1, 2, 1, 2, 4, 4, 3, 3, 1, 0, 1, 0, -1, -1, 0, -2, -1, 1, -2, 1, 1, 0, 0, 2, 4, 5, 4, 3, 0, 0, 0, 1, 1, 2, 3, 0, 5, 0, 4, 0, 1, 0, -1, 0, -4, 0, -1, 0, 0, 0, 1, 3, 3, 1, 2, 4, 5, 1, 3, 2, 2, 0, 0, 1, 1, 5, 3, 2, 2, 2, 1, 2, 1, -2, 0, -2, 0, 0, 0, 0, 0, 2, 1, 3, 3, 1, 2, 2, 2, 2, -1, 3, 3, 3, 1, 3, 3, 4, 2, 1, 0, 2, 0, 1, -3, -1, -3, -3, -3, 0, 0, 0, 0, 0, 1, 4, 2, 3, 1, 4, 2, 2, 2, 0, 2, 2, 5, 4, 5, 5, 4, 2, 1, 0, 0, -2, -1, -3, -4, -3, 0, 2, 0, 4, 2, 2, 1, 1, 3, 1, 1, 2, 0, 0, 2, 2, 4, 1, 2, 4, 3, 1, 2, -1, -2, -2, -3, -4, -1, -2, -1, 1, 4, 2, 5, 4, 3, 4, 0, 1, -1, 2, 0, 1, 4, 3, 3, 3, 5, 4, 1, 0, 1, 0, -4, -3, -3, -3, -3, -6, -1, 0, 0, 3, 3, 5, 2, 0, 4, 4, -1, 2, 0, 4, 1, 1, 3, 5, 5, 1, 4, 0, -1, 0, 0, -3, -6, -5, -5, -2, -4, 0, 0, 3, 3, 3, 3, 4, 4, 4, -1, 0, 1, 3, 2, 0, 3, 1, 2, 2, 1, 0, -2, 0, 0, -1, -1, -1, -5, -3, -2, 0, 2, 0, 0, 2, 1, 1, 4, 2, 0, 0, 1, 0, 3, 0, 2, 4, 3, 1, 1, 2, 1, -1, 0, -1, 0, -1, -3, 0, -2, -1, 1, 3, 2, 2, 1, 4, 2, 0, 0, 1, 0, 1, 1, 1, 1, 3, 5, 3, 4, 3, -1, 1, 0, 0, 1, -2, -1, 0, 0, 2, 2, 2, 3, 4, 2, 1, 0, 2, -1, 0, 1, 1, 4, 4, 2, 3, 2, 0, 3, 0, 0, 0, -1, 0, 1, -1, 3, 1, 2, 1, 3, 2, 1, 0, 1, 1, -1, 1, -1, 0, 1, 4, 4, 1, 3, 0, 0, 2, 4, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 3, 3, 0, 0, 0, 1, -2, 0, 1, 0, 1, 3, 2, 3, 0, 3, 1, 2, 0, -1, -2, -2, 0, 2, 0, 1, 4, 0, 3, 4, 4, 4, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 2, 1, 1, 2, 2, 0, 1, 0, 0, 0, 0, 0, 1, 2, 2, 4, 3, 2, 3, 1, 3, 0, 2, 0, 0, -1, 0, 0, 0, 0, 3, 0, 1, 0, 1, -2, 0, -2, -3, -1, -2, 1, 1, 0, 4, 3, 5, 3, 4, 3, 2, 1, 3, -1, 0, 1, 0, 2, 2, 1, 0, 0, 1, -1, 1, -3, -2, -5, -3, -4, -1, 0, 0, 1, 2, 5, 1, 4, 1, 3, 3, 3, 1, 0, -2, 1, 0, 0, 2, 3, 2, 0, 1, -1, -3, -2, -5, -5, -4, -1, -2, 0, 1, 2, 2, 5, 3, 4, 3, 1, 0, -1, 0, -2, -1, -1, 2, 0, 1, 2, 2, 2, 1, 0, 0, -4, -1, -2, -1, -1, -3, 1, 0, 5, 4, 5, 2, 5, 0, 3, 0, 0, 0, -4, -3, 0, -2, 2, 1, 0, 0, 0, 1, -1, -1, 0, -3, 0, -2, -4, 0, 1, 3, 3, 2, 2, 1, 1, 3, 2, 1, -2, -3, -3, -5, 0, 0, -1, -1, 1, 1, 0, 2, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 3, 0, 3, 0, 1, 0, 0, 0, -3, -4, -3, -4, 2, 4, 0, 3, 2, 3, 0, 0, 2, 2, 0, 2, 0, 2, 2, 0, 1, 0, 1, 1, 0, 2, 0, 0, 0, -2, -3, -1, -3, -4, 3, 0, 0, 1, 0, 3, 0, 2, 1, 2, 0, 0, -1, 0, 2, 3, 0, 3, 0, 2, 0, 1, 2, 1, -1, -1, -1, -1, 0, -1, 3, 2, 2, 3, 0, 0, 0, 0, 0, 0, -1, 1, -2, -1, 0, 0, 2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 3, 1, 1, 0, 0, -2, 0, -1, 0, -1, 0, -1, 1, 0, 1, 0, 1, 0, 4, 1, 1, 1, 2, 0, -1, 0, 1, 1, 3, 2, 3, 0, 0, 2, -1, -3, 0, 0, -2, 0, 0, 0, -1, 0, 0, 3, 1, 4, 4, 0, 0, 0, 0, 1, -1, -1, 1, 3, 2, 1, 4, 0, 2, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 0, 1, 1, 1, 3, 2, 4, 1, 3, 1, 2, 0, 0, 2, 1, 2, 4, 3, 3, 0, 0, 1, 1, 0, 2, 1, 0, 0, -1, 1, -1, 2, 1, 1, 3, 1, 3, 2, 0, 2, 0, 0, 0, 3, 0, 2, 2, 1, 1, 0, 0, 2, 2, 2, 0, -1, 1, 1, 0, -1, 0, 2, 0, 3, 4, 4, 0, 0, 2, 0, 0, 2, 1, 0, 1, 1, 2, 4, 4, 3, 3, 2, 2, 1, 2, 2, 0, -1, -2, -1, 0, 1, 0, 1, 1, 1, 1, 2, 2, 3, 1, 2, -1, 1, 2, 1, 3, 2, 1, 1, 4, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 3, 3, 2, 3, 0, 0, 1, 0, 2, 0, 3, 0, 2, 1, 2, 1, 0, 2, 0, 0, 0, -1, 0, -1, 0, 1, -1, 0, -1, 2, 0, 1, 3, 2, 1, 2, 0, 2, 3, 2, 1, 1, 3, 2, 1, 3, 3, 3, 2, 0, 0, 0, 1, 0, 1, 2, 0, 2, 1, 3, 3, 1, 2, 1, 4, 3, 0, 0, 2, 3, 3, 1, 2, 2, 2, 2, 4, 3, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 2, 0, 2, 2, 1, 1, 1, 3, 1, 1, 0, 1, 3, 1, 2, 4, 2, 1, 1, 2, 1, 2, -1, 1, 0, -2, 0, -2, 1, 1, 0, 2, 1, 3, 4, 4, 1, 0, 0, 2, 4, 2, 1, 4, 1, 4, 2, 2, 1, 1, 2, 0, 0, 1, 0, -1, -2, 0, 0, 2, 0, 3, 0, 1, 3, 4, 3, 3, 0, 1, 0, 0, 3, 2, 3, 2, 2, 3, 2, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, -1, 0, 2, 3, 0, 3, 0, 0, 2, 0, 3, 2, 1, 3, 0, 0, 1, 2, 1, 2, 1, 3, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, 3, 1, 3, 3, 1, 3, 2, 3, 0, 2, 3, 0, 0, 1, 2, 0, 4, 0, 2, 1, 1, 1, -1, -3, -2, -2, -1, 0, 2, 0, 0, 3, 0, 3, 3, 3, 3, 0, 0, 3, 0, 1, 0, 3, 3, 3, 3, 2, 1, 1, 0, 0, 0, -2, 0, 0, 0, 1, 1, 0, 1, 2, 3, 1, 3, 4, 2, 2, 2, 1, 0, 1, 3, 3, 4, 3, 1, 1, 1, 2, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 2, 3, 3, 1, 3, 3, 3, 1, 1, 0, 2, 1, 1, 1, 2, 1, 2, 0, 3, 2, 2, 0, 0, 0, 1, 1, 3, 3, 2, 1, 1, 2, 2, 4, 4, 1, 0, 1, 0, 1, 0, 0, 1, 2, 0, 3, 1, 3, 0, 1, 0, 1, 1, 1, 0, 0, 2, 0, 1, 4, 1, 3, 3, 1, 1, 3, 0, 1, 0, 2, 0, 2, 3, 0, 0, 3, 2, 2, 0, 0, 1, -1, 0, 0, 0, 2, 3, 0, 1, 4, 3, 1, 2, 1, 3, 3, 0, 1, 1, 1, 3, 3, 0, 2, 3, 1, 1, 0, 0, 2, 0, 0, 1, -1, 0, 0, 0, 3, 3, 2, 2, 4, 3, 0, 1, 3, 0, 2, 3, 2, 2, 3, 0, 1, 0, 1, 0, 2, 0, 0, 0, -2, 0, 0, 0, 1, 1, 2, 2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 3, 0, 2, 2, 0, 2, 3, 2, 2, 0, -1, 0, -2, -2, 0, 0, 1, 1, 0, 3, 3, 3, 3, 2, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 3, 2, 2, -1, 1, 0, -1, 0, 0, -1, 1, -1, 0, 2, 3, 2, 3, 0, 0, 0, -1, -1, 0, -1, 3, 3, 3, 0, 1, 2, 2, 2, 0, 2, 0, -2, -2, -2, 0, 0, 2, 0, 2, 2, 1, 3, 2, 0, 2, 1, 1, 2, 0, -2, 0, 0, 0, 0, 1, 3, 0, 1, 3, 2, 2, 0, 0, 0, 0, 1, 2, 1, 0, 2, 0, 2, 0, 2, 0, 0, 0, 0, -2, -3, 2, 0, 2, 2, 2, 2, 1, 0, 2, 1, 1, 2, 0, 1, -1, 0, 3, 0, 2, 3, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, -1, 0, -1, 1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, 0, 1, 0, 0, 2, 2, 0, 0, 0, 0, 1, -2, 2, 1, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, 1, 0, -1, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 1, 1, 0, 0, 0, -1, 1, 1, 0, 1, 2, 1, 2, -1, 0, 1, -1, 0, 1, 2, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, -2, -1, 0, 2, 0, 1, 1, 0, -1, 0, 2, 0, 0, -2, 1, 1, 1, 1, 0, 1, -1, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, 1, -1, 0, 0, 2, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, -1, 1, 0, -1, 0, 1, 1, 0, -1, 0, 1, 1, 1, -2, -1, 1, -1, 1, 1, 0, 1, 0, 0, 0, 1, -1, 1, 1, 2, -1, -1, 0, -1, -1, -1, 0, 0, -1, 0, 1, -1, -1, 0, -1, 1, -2, 0, 0, -2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, 1, -1, 0, -1, 0, 1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 1, -1, 1, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, -1, 1, -1, 0, 1, 0, 0, 2, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, -1, 0, 1, 0, 0, 1, 0, 0, 1, -1, -1, -1, -1, 1, 1, 1, 0, -1, 1, 1, 0, -1, -1, -1, -1, 0, 0, 1, 0, -1, -1, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 1, -1, 0, 0, -2, 0, -1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, -1, 0, 0, -1, 1, -1, -2, 0, 2, -1, 0, -1, 1, 0, 1, 1, 0, 1, -1, 0, 1, 2, 0, 0, -1, 0, 0, 0, 0, 2, 0, 1, -1, 2, -1, 0, -1, 1, 0, 0, 2, -1, -2, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 1, -1, -1, -2, -1, 0, 0, 0, -1, -1, 0, -1, 1, -2, 1, 0, -1, 0, 1, -1, 1, 1, 0, 1, 1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, 1, 0, 1, 0, 2, 0, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, -1, 1, -1, 0, -1, 1, 0, -1, -1, 1, -1, -1, 0, 0, -1, 0, 0, -2, 1, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, -1, 0, -1, 0, 1, 0, 1, 0, 1, -1, -1, 0, 0, 0, -1, 1, -1, -1, -1, 0, 1, 1, 1, 2, -1, 1, 0, 0, 2, -1, -1, 0, 1, -1, -1, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 1, 0, 0, -1, -1, 1, -1, 1, 0, 0, -2, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, 1, -2, 0, -1, 0, -1, 1, 0, 0, 0, 0, -1, 1, 1, 0, 1, 1, 0, 1, 0, -1, 1, 0, -1, 0, 1, 1, 0, 0, -1, -1, 1, 0, -1, 1, 0, 0, 1, 1, -1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, 2, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, -1, 1, 0, 1, 1, 1, 1, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 2, -1, 0, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 2, 1, 2, 0, -1, -1, 1, -1, -1, 1, -1, 1, 1, 1, 1, 0, 0, 1, 1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, -1, -1, 0, 1, 0, -1, 0, -1, 0, 1, 1, 1, 0, 1, -1, 1, 1, 1, 0, -1, -1, -1, 1, 0, -1, 0, 1, 0, 1, 0, -1, 1, 0, 0, 1, -1, 0, 0, 2, 1, 2, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, -2, 0, 0, 0, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -3, -3, -1, -1, -4, -4, 0, 0, -1, 0, -1, 1, -1, -2, 1, 0, -1, -2, -1, -1, 0, -3, -3, -2, -2, -2, -3, -1, -2, -4, -4, -3, -3, -3, -4, -2, -1, -1, -1, -2, -2, 1, 1, 0, 0, -2, 1, -1, -1, 0, -2, -2, -2, 0, -4, -3, -3, -1, -3, 0, -5, -4, -4, -4, -2, -2, -3, -3, 0, -1, -3, -1, 0, 0, 1, 0, 0, 0, -2, 0, 2, 0, 1, -1, 0, 0, 0, -1, 0, -3, -2, -2, -4, -3, -3, -2, -1, -3, -2, -4, -4, -1, 0, 2, 0, -1, 0, 1, 0, 1, 1, 0, 0, 0, 0, -3, -2, -1, 0, 0, -4, -3, -6, -5, -2, -1, -2, -4, -4, -2, -3, -1, -1, 0, -2, 0, 0, -1, 0, 0, -2, 0, 0, 1, -3, -3, -3, -1, -3, -2, -1, -3, -2, -5, -1, -1, -1, -2, 0, -1, -1, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -2, -2, -1, -3, 0, -3, -5, -3, -3, -3, -4, -1, -1, 0, -1, 0, -1, -1, -3, 0, 0, 0, -1, 1, 1, -1, 1, -1, -2, 0, 0, -2, 0, 0, 0, 0, -4, -3, -3, -4, -1, -2, -2, 0, -3, 0, -1, -1, -3, -1, -3, 0, -3, 0, -2, -1, -1, 1, -1, 0, 0, 1, 0, 0, 0, 0, -3, -4, -5, 0, -3, 0, -2, 0, -2, 1, -1, 0, 0, -2, -2, -1, -2, -1, -1, 0, 0, -1, -3, -2, 0, -1, 1, -1, 0, -1, -4, -4, -1, -3, 0, -2, -3, -2, 0, 0, 0, 0, -1, -1, -3, -2, -2, -1, -3, -4, -2, -2, -3, -1, 0, -1, -2, -1, -2, 0, -4, -5, -1, -4, 0, -1, -1, -3, -1, -3, 0, -3, -1, -1, -1, -1, -1, -1, -2, 0, -1, -1, -2, -1, -1, -1, 1, -2, -2, -2, -4, -2, -3, -2, -2, -2, 0, 0, 0, -3, -2, -2, -4, -1, -4, -2, -1, 0, 0, -1, -1, -1, -3, -1, -3, -1, -2, -2, 0, -1, -1, -2, -5, -2, -4, 0, -3, -2, -3, 0, -1, -2, -2, -2, -3, 0, -3, -3, -4, 0, -4, 0, 0, 0, -1, -2, -2, 0, 1, 2, -5, -3, -5, -4, -4, 0, 0, -1, -1, 0, -2, -2, -4, -3, 0, -2, -3, -2, -3, -5, -4, 0, -2, -1, -3, -1, -2, -1, 2, 1, -4, -5, -2, -3, -1, -1, -2, -2, -2, -2, -1, -2, -3, -1, -2, -2, -3, -2, -5, -3, -4, 0, 0, 0, -2, -3, 0, -1, 0, 0, -5, -2, -1, -2, -3, -3, -3, -2, -1, -2, 0, 0, 0, -2, -2, -4, -5, -3, -3, -4, -3, -3, -2, -2, -3, -4, -1, 0, 1, 1, -6, -5, -4, -3, -2, 0, -1, -1, -4, -2, 0, -1, -1, 0, -1, -3, -4, -5, -5, -4, -3, -5, -3, -3, -2, -4, -2, -1, 0, 0, -4, -3, -2, -3, 0, -3, -2, -2, -1, -1, -1, -2, -3, 0, 0, -3, -1, -4, -7, -6, -4, -4, -5, -3, -2, -2, 0, -2, 0, 0, -3, -3, -4, -4, -4, -1, -2, 0, -2, -3, 0, -2, -1, 0, -1, -1, 0, -1, -2, -2, -3, -3, -1, -3, 0, -3, -2, -1, 0, 1, -2, -3, -4, -3, 0, 0, -2, -3, -2, -1, -2, 0, -2, 0, -1, 0, -2, -2, -1, -4, -4, -1, 0, -3, -2, -1, -1, 0, -1, 0, -6, -4, -2, 0, -1, -1, -3, 0, 0, -1, 0, 0, -2, -2, 1, -1, -2, -2, -2, -2, -1, -1, -1, 0, 0, -2, 0, -1, -2, 0, -3, -1, -3, -1, 0, 0, 0, -1, -1, 0, 0, 1, 0, -3, -1, 1, 0, -1, -2, -2, -1, -3, -4, -3, -1, -2, 0, -3, -1, 0, -2, -4, -2, 0, -2, -3, -3, -1, 0, -1, 1, 0, 0, -2, 0, -1, -1, 0, -1, -1, -4, -2, -1, -1, -1, -1, -1, 0, -3, -1, -3, -1, 0, -1, -3, -4, -1, -1, -1, -2, 0, 1, 0, 1, -1, -2, -3, -1, -3, -3, -2, -4, 0, -3, -1, -1, 0, -1, -1, -1, -4, -2, -2, -1, -1, -2, 0, -2, -3, 0, 0, -1, 0, 0, 0, 0, -3, 0, -3, -2, -3, 0, 0, -3, -2, 0, -3, 0, -1, -1, -1, -3, -3, -2, 0, 0, -2, 0, -2, -2, -2, -1, -3, 0, -1, -1, 0, -3, -3, 0, -2, -3, 1, 0, 0, -1, -1, 0, -1, -1, -5, -2, -3, -3, 0, -2, 0, -2, -2, -3, -4, -1, 0, 0, -3, 0, -2, 0, -1, 0, 0, -1, 1, -1, -1, -1, -1, 0, 0, 0, -5, -2, -3, 0, 0, -3, -1, -4, -3, -5, -1, 0, -1, -4, -3, -1, 0, 1, 0, -1, 0, 2, 0, 0, 0, 1, 0, -2, 0, 0, -2, -3, -3, -5, -2, -4, -3, -2, -4, -3, -2, -4, -4, -2, -1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, 0, -3, -3, -2, -3, 0, -1, -3, -3, -3, -3, -1, -1, -1, -1, 0, -1, 0, 0, 1, -1, 0, 0, -2, -1, 0, 0, -1, -2, -1, -1, 0, -1, 1, -1, 0, 0, 0, 0, -1, 1, 1, -1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, -1, 1, 0, 1, 0, 0, 1, 1, 2, 1, 1, 0, 1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, 0, -1, -2, 1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 1, -1, 0, -1, 1, 0, -1, -2, 0, -1, 1, 1, -1, 1, 0, 1, -2, 1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, 0, 0, -2, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, 0, -1, 1, 1, 1, 0, 1, 0, 0, -1, 1, 0, -2, 0, -2, 1, 0, 0, -1, 0, 1, 1, 1, -1, 1, 0, 1, 1, 0, 0, -1, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 1, -2, 0, 1, 0, -1, 1, 1, 0, -2, 1, 0, 0, 0, -1, 0, 2, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, -1, 1, -2, 0, 0, -1, 0, -1, 0, 0, -1, 1, -1, -1, 1, -1, 0, 0, 0, -1, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -2, 0, 0, -1, -1, -1, 0, 0, 0, 1, 1, 1, 2, 0, 0, -1, 0, 0, -1, -2, -1, 0, 0, 0, -1, 1, -1, -1, 1, 1, 1, 1, 1, 2, 0, 0, 0, 1, 1, 0, -1, -1, 2, 0, 1, 0, 0, 0, 0, 1, 0, -2, 0, 0, -1, 1, -1, -1, 1, -1, 0, 1, 0, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, -2, -2, -2, 1, 0, 1, 1, 0, 1, -2, 0, -1, -2, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 1, 1, -2, 0, 0, 0, 1, 1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -2, -1, 0, -1, 0, -1, -1, -1, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 0, -1, 1, 1, 2, 0, 2, 2, 0, 0, -1, 1, -1, 0, 0, 0, -1, -2, 0, 0, 1, -2, -1, -1, 0, -2, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, -1, 0, 1, 0, -1, 1, -2, -1, 0, 0, 1, -2, 0, 0, -1, 0, 1, -1, 0, 0, -1, -1, 1, 1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, 1, -1, 1, 0, -2, 0, 0, 0, -1, -2, 0, 1, -2, 0, 1, 0, 0, 0, 2, 2, -1, 0, 1, 1, 1, 1, -2, 0, 0, -2, -1, 0, 0, 0, -1, -1, 1, 0, -1, 0, -2, 0, 0, 0, 1, 1, 1, -1, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, -1, -1, 1, -1, -1, 0, 1, -1, 0, 2, 1, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, -2, -1, 0, -2, -1, -1, 0, 0, 1, 1, -2, 0, -2, 0, -1, -1, 1, -2, 1, -1, 0, 0, 0, 1, 0, 0, 2, -1, 1, -1, 1, 0, -1, 0, 0, -2, -2, -1, 0, 0, -1, -1, -2, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, -1, 0, 1, 0, 2, -1, 0, 0, 1, -2, 0, 1, 0, 0, -1, 1, 0, -2, 0, -1, -2, 0, -1, 0, 0, -1, 1, 1, 0, 2, 1, 0, 2, 0, -1, 1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 0, -2, 0, 0, -1, -1, 1, 1, 0, 0, 1, 1, 2, 0, 1, 2, 1, 1, -1, 2, -1, -2, 0, 0, -2, 0, 0, 1, 1, -1, 1, 1, 0, 1, -2, 0, 1, -1, -1, 0, -1, -1, 0, 0, 2, 1, 1, 1, -1, 1, -2, -2, 1, -1, 0, 1, 0, -2, 0, 0, -1, 1, 1, 0, 0, -1, 1, 1, 0, 1, 1, 1, 2, 0, 1, 2, 2, 2, -1, -1, -1, 1, -1, 0, -1, 0, -2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, -2, 0, 0, -1, 0, 1, 1, 0, 1, -1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 1, -1, -1, 0, 0, 1, 1, -2, -1, 1, -2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -2, -1, 1, -1, 0, -2, -2, 0, 0, 0, 0, 1, -1, 1, -1, 0, 1, 0, 0, 0, -1, 1, -2, 0, -1, 0, 1, -2, 1, 0, 0, 0, 0, 0, 1, 1, -2, -1, 0, 0, -1, 2, 0, 0, -2, 1, 0, 0, 0, 1, 0, 1, 0, -1, 0, 1, 1, 0, 0, -2, 1, 1, 0, 0, 1, 1, 0, -1, 0, -1, -1, 1, 0, 0, 1, 0, 0, 1, 0, 1, -1, 0, -1, -1, 1, 0, -1, -2, 0, 0, 1, 1, -1, 0, 1, -1, 0, -1, -1, -2, 1, 0, -2, -2, 0, 0, 1, 0, -1, 1, 0, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, -1, -2, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -2, 0, 0, 0, 1, -1, 0, 0, 1, 1, -1, 0, 0, -1, 1, -1, 0, 1, -1, 0, 0, -1, 0, -2, 0, 0, 0, 0, -1, -1, -1, -2, 1, 0, 0, 1, 1, -2, 0, 0, 0, 0, -1, 1, 0, -1, 1, 0, 1, 1, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 1, 0, -2, 0, -1, -1, -1, 1, 0, 0, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, -1, 0, -1, 1, 0, -1, 0, 1, -1, 1, 1, -1, 0, -1, -1, -1, 1, 0, 0, -2, 0, 0, 1, 0, -1, 1, 0, -2, -1, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, -1, 0, -2, 1, 0, 1, 1, -1, 1, -2, -1, 0, 1, -1, -1, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, -1, -1, 1, 0, 0, 2, 1, 2, 1, 0, 1, -1, 1, 0, -2, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 1, 1, -1, -1, -1, 1, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, -2, 1, -2, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, -1, 1, -1, -1, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, -1, 1, 0, 2, 1, 2, 2, -1, 1, -1, -2, -1, 1, -1, 0, 0, 1, 1, -1, 0, -1, 0, 1, 1, 1, -1, 0, 1, -1, 1, 0, 1, -1, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 1, 0, -1, -2, 0, 0, 1, 0, -1, 0, -1, 0, 1, -1, 0, 1, -1, 1, 0, -1, 2, -1, 2, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, -2, -1, -1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, -1, 1, 1, 2, 0, -1, 1, -1, 0, 0, 0, -2, 1, 1, 0, -1, -1, 1, 0, 0, -1, 0, 1, 0, 0, 1, 1, 1, 0, 2, 0, 1, 1, 0, 1, 0, 0, 1, 1, -1, 0, 0, -1, -1, -2, 0, -1, 0, 0, -1, 0, -1, -2, 1, -2, 0, 1, -2, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, -1, 0, -1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 1, -1, -1, 1, 0, 0, 0, 1, 0, 0, -1, 0, -1, 1, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, -2, 1, 0, 1, -1, 0, 2, -1, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, 1, -1, 1, 0, 1, 0, 1, 0, 0, -1, 1, 0, 1, -2, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 1, 0, -1, 1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 1, -1, 0, -1, 1, -1, -2, 0, 1, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, -1, 1, -2, -1, -1, -1, 0, 0, 1, 0, 0, -1, -2, -2, 0, 0, -2, 1, 1, 0, 0, -2, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, -2, 0, 0, 0, 0, 0, -2, 0, 1, 1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 1, 1, -2, -1, 1, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, 0, 0, 1, 0, -2, 0, -1, 1, -2, 0, -1, 1, 0, -2, 0, 0, 0, 0, 0, -2, 1, -1, 0, 1, -1, 0, 0, 0, -1, -2, 0, -2, -1, 0, 1, -1, 0, -1, 0, -2, -2, -1, 1, -2, -1, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, -2, -1, -1, 0, 0, -2, 1, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, 1, 0, -1, 0, 0, 1, 1, -1, -1, 0, 1, 1, -1, -2, -1, 0, 1, 0, 0, -2, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, -2, 0, -2, 0, 1, 0, 0, 0, -1, 1, 0, 1, 0, -2, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, 0, 1, 1, 1, 0, 1, 0, -1, -2, -1, -1, 0, -3, 0, -1, 0, -1, -3, -3, 0, 0, -2, -2, -3, 0, 0, -2, 0, -2, -2, 0, -2, -2, -3, 0, -2, -2, -3, -3, 0, 0, 0, -1, 0, -3, -2, -2, -2, 0, 0, -3, 0, 0, -1, -3, -1, 0, -1, 0, -2, 0, 0, -2, 0, 0, 0, -1, 0, -1, -1, -1, -1, -1, -3, -1, 0, 0, 0, -1, -1, -2, 0, -1, 0, -2, -1, -1, -2, -2, -1, -3, -1, -2, 0, -2, -2, -3, 0, -2, -3, -2, 0, -2, 0, 0, -3, -1, -1, -3, -1, -2, -3, 0, 0, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, -1, -2, 0, -3, 0, -1, -2, -3, 0, -1, -2, -2, 0, 0, -2, -1, -1, -2, 0, -2, -2, 0, 0, 0, 2, -1, -1, 0, 0, 0, -1, 1, -1, -2, -2, -2, -3, -2, 0, -1, -2, 0, -2, 0, -2, 0, -1, -1, 0, -2, 0, 0, 1, -1, 0, 0, 0, -2, -2, 0, -2, -1, 1, 0, -1, -1, -2, -2, 0, -1, -2, 0, -1, -2, 0, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, 0, -1, 0, -2, -2, -2, -1, 0, 0, -1, -1, 0, -3, -2, 0, -1, -2, -2, -2, 0, 0, 0, 0, 0, 0, 2, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, -3, 0, 0, -2, 0, -1, -2, 0, 0, -3, -1, 0, 0, -2, -1, 0, -1, 0, 0, -1, 1, -1, 0, 1, -1, 0, -1, -1, -2, -3, 0, -1, 0, -1, -2, -2, 0, 0, 0, -2, 0, -2, 0, -2, -1, -2, 0, 0, -1, 1, 0, 1, -1, 0, 0, 0, -2, -1, 0, -1, 0, -2, 0, 0, -2, -2, 0, 0, -2, -2, -1, -1, 0, -1, 0, 0, -1, -1, 1, 1, 1, 1, 0, 1, 0, 1, 0, -1, -1, -2, -2, -2, -2, 0, -1, -1, 0, -3, 0, -3, -2, 0, -2, 0, 0, 1, 0, 0, 2, 0, 1, -1, 1, 1, 0, 2, 0, -1, 0, 1, -3, -1, 0, -3, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, -1, 0, 0, -1, -2, -2, 0, 0, -2, -2, 0, -1, -3, -2, 0, -1, -2, -1, 0, 0, -2, 0, -1, 0, 0, 2, 0, 2, 0, 0, 0, 2, 0, 0, 0, 0, -1, 0, -2, -2, -1, -2, -3, -3, -3, -3, -2, -2, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 2, 1, 1, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, -2, -2, 0, 0, -1, 0, 0, -1, 0, -2, -2, -1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, -3, 0, -2, 0, -2, 0, -2, 0, 0, -2, 0, 0, 1, 0, 1, 1, 2, 2, 1, 0, 2, 0, 0, -1, 0, -2, -1, 0, -2, -3, -3, -1, -1, -1, -2, 0, -2, -1, 1, -1, 1, 0, 1, 2, 0, 2, 3, 3, 2, 0, 1, 0, 1, -1, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, -2, -3, 0, 0, -1, 0, 0, -1, 2, 0, 1, 0, 0, 2, 0, 0, -2, 0, -1, 0, 0, -1, -2, -2, -4, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 2, 0, 1, -1, 0, -1, -2, 0, 0, -1, -1, 0, 0, 0, -1, -3, 0, 0, -2, -2, 0, 1, -1, 1, 2, 0, 0, 0, -1, 0, -1, 1, 1, 1, -2, 0, 0, -2, -2, -2, -3, -2, -1, 0, -2, -2, -1, 0, 1, -2, 0, 1, -2, 0, 0, 0, -1, -1, 2, 1, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, -2, -2, 0, 0, -2, -1, 0, -1, 0, -2, -2, 0, 0, -1, -1, 0, -1, 0, 1, 2, 0, 1, 0, 0, 0, -2, 0, 0, 0, -2, -3, -4, 0, 0, 0, 0, 0, -3, -2, -2, 0, 0, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, -3, -3, -4, -2, -1, -2, 0, -1, -3, -2, -2, -1, 0, 0, 0, -2, -2, 0, 0, 0, 0, 1, -1, -1, 0, -2, 0, -2, 0, -2, -2, -3, -2, -1, -1, -2, -2, 0, 0, -2, 0, -2, 0, 0, -1, -3, -2, 2, -2, -1, -2, -2, -1, 0, 0, -2, 0, -3, -3, -2, -1, -4, 0, -3, 0, -1, 0, 0, 0, -3, 0, 0, 0, 0, 1, 0, -2, -1, 1, -2, -1, -1, -1, 0, 0, -1, 0, -1, -2, -4, -2, -2, -4, -1, -3, -3, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, 0, -2, 0, -3, -4, -2, -2, -2, -2, 0, -3, -2, -2, -2, -2, -1, 0, 0, -3, -2, 0, 1, 0, -2, 0, -1, 0, -1, 0, 0, -3, -1, 0, -3, -4, -1, -3, -2, -2, -2, 0, -6, -7, -8, -9, -8, -6, -6, -5, -3, -5, -4, -2, -4, -4, -3, -3, -6, -3, -2, -2, -1, 0, 0, -3, -2, -1, -1, 0, 0, 0, -10, -8, -9, -7, -9, -6, -7, -7, -6, -3, -1, -1, -1, -1, -2, -3, -4, -4, 0, -1, -3, -1, -2, -3, -4, -2, -2, 0, -1, 1, -10, -10, -10, -6, -7, -5, -4, -6, -5, -5, -1, 0, -2, 0, 0, -1, -3, -1, -3, 0, -3, 0, -3, -3, -1, -1, -2, -1, 0, 0, -7, -8, -10, -8, -6, -6, -6, -6, -6, -3, -1, 0, -2, 0, -1, -1, 0, -2, -1, -1, -2, -2, -1, -3, -2, -3, -3, -2, 0, 0, -7, -7, -10, -6, -5, -7, -4, -6, -7, -4, -2, -3, -2, 0, 0, 0, 1, 0, -2, -3, -2, -1, -2, -1, -1, -3, -3, -2, 0, 0, -10, -6, -8, -6, -6, -6, -4, -3, -6, -5, -4, -5, -3, -3, 0, -2, 0, -3, -1, -3, -3, -4, -3, -1, -2, -2, -3, -4, -3, 0, -8, -8, -8, -6, -5, -6, -6, -3, -5, -4, -4, -4, -3, -4, -2, 0, -3, -1, -1, -2, -2, -2, -4, -2, -4, -3, -5, -2, -2, -1, -9, -8, -9, -9, -6, -7, -4, -5, -4, -4, -5, -3, -2, -3, 0, 0, -2, -1, -3, -3, -5, -2, -3, -4, -5, -1, -3, -4, -3, -1, -7, -9, -8, -9, -8, -4, -4, -4, -2, -5, -4, -5, -5, -6, -3, -4, -4, -3, -4, -5, -2, -4, -6, -6, -2, -4, -2, -3, -1, -3, -7, -9, -8, -7, -8, -5, -8, -3, -4, -5, -1, -4, -4, -6, -2, -1, -1, -3, -6, -7, -4, -3, -5, -4, -5, -3, -3, -2, 0, 0, -9, -10, -7, -6, -6, -4, -4, -5, -7, -7, -6, -6, -7, -6, -4, 0, -2, -6, -3, -6, -4, -4, -2, -3, -4, -5, -5, -1, -1, -2, -9, -8, -6, -5, -5, -8, -6, -4, -7, -7, -6, -7, -4, -4, -2, -2, -3, -5, -5, -6, -6, -3, -5, -4, -5, -2, -3, -3, -2, -2, -6, -7, -9, -8, -6, -6, -5, -4, -7, -6, -6, -8, -4, -2, -3, 0, -1, -4, -3, -3, -5, -6, -3, -3, -4, -2, -1, -3, 0, 0, -8, -8, -9, -7, -7, -4, -7, -8, -5, -8, -5, -5, -5, -3, -3, -3, -2, -2, -4, -4, -6, -3, -7, -6, -3, -6, -4, -3, -2, 0, -10, -6, -9, -6, -8, -5, -7, -7, -7, -5, -6, -6, -4, -4, -4, -1, -3, -4, -4, -6, -3, -3, -5, -6, -4, -3, -5, -2, -1, 0, -8, -7, -6, -7, -5, -7, -8, -8, -5, -5, -8, -6, -4, -3, -1, -3, -3, -6, -6, -5, -5, -5, -3, -3, -5, -5, -2, 0, 1, -1, -8, -5, -5, -8, -5, -6, -6, -5, -8, -5, -3, -4, -4, -2, -3, -3, -4, -5, -6, -5, -6, -7, -6, -3, -4, -3, -2, -3, -2, -1, -9, -5, -7, -8, -4, -5, -8, -5, -6, -7, -2, -2, 0, -1, -3, -4, -4, -7, -7, -6, -7, -5, -6, -5, -5, -2, -4, -3, -2, 0, -11, -8, -8, -7, -6, -8, -4, -5, -7, -5, -4, -5, -4, -1, 0, -4, -3, -7, -8, -4, -8, -7, -3, -3, -4, -3, -4, 0, 0, 1, -10, -7, -6, -6, -6, -5, -6, -6, -6, -4, -3, -5, -5, -2, -1, -2, -3, -6, -5, -6, -7, -6, -2, -6, -3, -6, -4, -3, 0, -1, -9, -7, -4, -6, -5, -5, -7, -8, -4, -5, -5, -5, -1, -2, -1, -4, -5, -5, -7, -7, -8, -5, -6, -4, -5, -5, -1, -3, -2, 0, -7, -6, -6, -4, -7, -6, -6, -4, -3, -5, -5, -4, -2, -3, -3, -2, -2, -3, -6, -7, -7, -6, -3, -4, -6, -3, -1, -4, -1, 0, -6, -8, -6, -5, -6, -4, -8, -5, -3, -5, -1, -5, -3, -4, -1, -1, -3, -4, -7, -5, -6, -5, -4, -5, -2, -4, -2, -2, -2, -1, -10, -7, -6, -5, -5, -7, -5, -8, -4, -3, -3, -4, 0, -4, -4, -3, -3, -6, -3, -2, -3, -4, -5, -4, -2, -1, -3, -2, -1, 0, -7, -6, -7, -5, -5, -6, -4, -7, -6, -2, -5, -1, -3, -3, -2, -4, -2, -5, -2, -2, -4, -3, -3, -5, -2, -2, -2, -2, 1, 0, -6, -8, -7, -6, -6, -4, -5, -6, -4, -3, -1, -4, -2, -1, -2, -2, -3, -2, -5, -3, -1, -4, -5, -5, 0, -1, -1, -2, 0, 0, -7, -6, -7, -7, -4, -5, -4, -4, -6, -2, -1, -4, -3, 0, -3, -3, -4, -2, -4, -1, -2, -1, -2, 0, -2, 0, -2, 0, 0, 2, -5, -7, -6, -7, -8, -8, -7, -5, -7, -4, -4, -4, -5, -1, 0, -3, -3, -3, -2, -3, -1, -3, 0, 0, -2, 0, -1, 0, 2, 1, -7, -6, -6, -8, -6, -9, -8, -7, -10, -6, -8, -4, -5, -3, 0, -1, -1, -3, 0, 0, -2, -2, 0, 0, 0, 1, 0, -1, 2, 1, -7, -10, -10, -8, -6, -9, -8, -7, -9, -10, -7, -8, -7, -5, -3, -4, -2, -3, -2, -1, -1, 0, -1, 0, 1, -2, 1, 2, -1, 1, 1, 0, 0, 1, 1, 1, 2, 1, 0, 0, 1, 2, -1, 1, -1, 1, 0, 1, 0, 0, 1, -1, -1, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 2, 1, -1, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 2, -1, 0, 0, 0, 2, 0, -1, 0, 0, 1, 0, 0, -1, 1, -2, 0, -1, 1, 0, 1, -1, 0, -1, 0, 1, -1, 0, 0, -1, -1, 1, 0, 2, 1, 0, 1, 0, -1, 0, -1, 1, 0, -1, -1, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, 1, -1, -1, 0, 2, 0, 2, -1, 0, 2, -1, 0, 1, 0, 0, -1, 1, 0, 1, 0, -1, 1, 0, 0, -1, -1, -1, 0, -1, -1, 1, 1, 1, 0, 1, 1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 2, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 1, -1, 2, -1, -1, 0, 1, -1, -1, 2, 1, 0, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 2, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 2, 1, 2, -1, -1, 0, 1, 0, 1, 0, 0, -1, 2, 0, 1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 1, 0, 1, -1, -1, 1, 0, -1, 0, 1, 0, 0, 0, 1, -1, 2, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, 2, 0, 0, 1, 0, 0, 1, -1, 1, 2, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, 2, 0, 1, -1, -1, 2, 2, 0, 0, 1, 2, 0, 1, -1, 0, -1, 0, 2, 0, 1, 0, 1, -1, 1, 1, 1, 0, 0, -1, 1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 2, 2, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 1, 2, -1, 0, 0, 1, 1, 0, -1, 0, -1, 1, 1, 0, 0, -1, 0, 2, 0, 1, 0, 0, 2, 1, 0, 0, 1, 1, 0, 1, -1, 0, 0, 1, -1, -2, 0, -1, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, -1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 0, 1, -1, 1, 1, -1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 2, 0, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 1, -1, 0, 1, 1, 0, -1, 0, 0, 0, 1, -1, 1, -1, 0, -1, 2, 0, 1, 1, 0, 0, -1, 0, 0, 1, 2, -1, 0, 0, 1, 1, 1, -1, 0, 0, 2, 0, -1, -1, 0, -1, 1, 0, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 2, -1, 0, -1, 0, 1, 0, 2, 2, 1, -1, 0, 1, -1, 0, 1, 1, 0, 0, -1, 0, 0, 2, 2, 1, 0, 0, 0, 1, 0, -1, 0, 2, 0, 1, 1, 1, 1, 0, -1, 1, 0, 1, -1, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 2, 1, 0, 1, 1, 0, 1, -1, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 2, 0, 0, 0, 0, 0, 2, -1, 1, -1, 1, 0, -1, 1, 1, 0, 0, 0, 0, 1, 0, 1, 1, -1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, -1, 1, -1, 1, -1, 0, 0, -2, 0, 0, 0, -2, 0, 0, 0, -1, 1, 1, -1, 1, 0, 2, 2, 1, -1, 0, 1, 1, 1, -1, 0, -1, 1, 1, 0, 1, 0, 1, 1, 0, 1, -1, 0, 0, 0, 1, 1, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, -1, -1, 0, 2, 2, 1, 1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 2, 0, 0, -1, 0, 1, -1, 0, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 2, -1, 0, 0, 0, 1, 1, 0, -1, 1, 0, -1, -1, 0, 0, 0, 1, -1, 1, 2, 1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, -1, -1, -1, -1, -1, -1, 0, 1, 0, 0, -2, -2, 0, 0, -1, 0, 0, 1, 1, -1, 0, 0, 2, 0, 0, 1, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, -1, -1, -1, 1, 0, 0, 0, -1, 0, 0, 2, 1, -1, 0, -1, 1, -1, -1, 1, 0, -2, 1, 0, 0, -1, -1, 1, -2, 2, 0, -1, 1, 0, 0, 0, 0, 1, 1, 0, -2, 0, 1, 0, -1, -1, 1, 1, 1, 0, -1, 1, 0, 2, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 1, 0, 0, 2, 0, -1, 0, -1, 0, 1, 0, -1, 1, -1, 0, 0, 1, -1, 0, 0, -2, 0, 1, -2, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, 2, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 0, -1, 1, 0, 1, -1, 0, 0, -2, 1, 0, 0, -1, 0, -1, 1, 0, 0, -1, 0, -1, -2, -1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, -2, 0, 1, 1, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, -2, -1, 0, 1, 1, 0, -2, 0, -1, 0, 1, 2, 1, 0, -1, 0, 0, 1, 0, -1, 0, 0, -1, 1, -1, 0, 1, 0, -1, 2, -1, 0, 0, 0, 1, -1, 2, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 1, -1, 0, -1, -1, 0, 1, 1, 1, 0, 0, 1, 0, -1, 2, 1, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 1, -1, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 1, 0, 0, 2, 0, 0, -1, -1, -1, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, -1, -2, 0, -1, 0, 0, 1, 0, 0, -1, 1, 0, 1, -1, 1, -1, 0, 1, -1, 1, 1, 0, -1, -1, 1, 0, 2, -2, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, -1, -1, 0, 0, 1, -1, 2, 1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, 0, 1, -1, 1, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 2, 1, 0, 1, -1, -1, -1, -1, 0, -1, 2, -1, 0, 0, 1, 0, 0, 1, 1, 2, -1, 1, 1, 0, 0, 0, 0, 0, -1, 2, -2, 0, -1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, -1, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 1, 1, -1, 0, 1, 0, 1, -1, -2, 0, -1, 1, 0, 1, -1, 0, 0, -1, -1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 1, -2, 0, 0, 0, 1, 1, 1, -1, 1, -1, 2, 0, -2, 0, 0, -1, 1, -1, 0, 2, -2, -2, 0, 0, 1, 0, 0, -1, 1, 0, 1, 1, -1, 1, -1, 0, 0, -1, 1, 1, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, -1, 1, 0, 1, -1, 0, -1, -1, 0, 0, -1, 0, 1, -1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, -1, 0, -1, -1, 0, 0, 0, -1, -1, 1, -2, 1, 0, 1, 0, -1, 0, -2, 1, 1, 1, 0, 1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, -1, -1, 0, -2, 0, -1, -1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 2, 0, 1, 0, 1, 1, -1, 0, 1, 1, -1, 0, -1, -1, 0, 0, 0, 1, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, -1, -1, 1, -1, 0, 1, -1, 0, -1, -1, 0, -1, 1, 0, 1, -1, 1, 0, 0, 0, 0, 1, 0, 1, -1, 2, 0, 1, 0, 0, 0, 1, -1, 0, -1, 0, 1, 1, 0, -1, -1, -1, 1, 1, 0, -1, 0, 0, 1, 0, -1, -1, -1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 1, 1, 0, 0, 2, -2, -1, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, 0, 0, 2, 0, 0, -1, 1, -1, -1, 0, -2, 1, -1, 0, 0, -1, 0, -2, 0, 1, 0, 1, -1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 1, 0, 0, -2, 0, -2, 0, 0, -1, 1, 1, 0, 0, 0, 1, 1, 1, -1, -1, -1, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 2, 1, -1, 0, 0, 0, -1, 1, -2, 0, 0, -1, 0, 0, -4, -3, -3, 0, 0, 0, 1, -1, 0, 1, 1, 4, 4, 2, 3, 3, 2, 1, 2, 2, 0, -1, -2, -1, -2, -4, -6, -3, -5, -6, -2, -4, -4, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 2, 3, 3, 4, 1, 1, 3, 1, 2, 0, 0, -4, -3, -4, -2, -5, -5, -3, -3, -3, -3, 0, 0, -3, 0, -1, -3, -2, -2, 0, 1, 0, 3, 0, 2, 4, 3, 3, 3, 0, 2, 1, 0, -3, -2, -2, -3, -1, -5, -4, -3, -1, -3, -3, -5, -1, -1, -1, 0, 0, 1, 0, 1, 0, 1, 3, 5, 4, 4, 3, 0, 0, 0, 0, -2, -1, -3, -4, -3, -4, 0, 0, 0, -1, -2, -1, -3, 0, -3, -1, -1, 0, 1, 2, 3, 4, 3, 5, 5, 4, 3, 2, 0, 0, -2, -1, 0, -1, -1, -3, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, 0, 0, 0, 1, 5, 6, 4, 5, 5, 0, 1, 1, 2, 0, 2, 0, -1, -4, -4, -2, -1, 1, 0, 0, 0, 2, 3, 0, 0, 0, -2, -2, 1, 0, 3, 1, 1, 2, 5, 2, 3, 3, 4, 0, 1, 1, 0, -3, 0, 0, 1, 2, 0, 4, 1, 3, 4, 1, 2, 1, -2, -2, 0, 2, 3, 0, 0, 4, 1, 4, 3, 1, 4, 2, 3, 0, -1, -1, -4, 0, -1, 0, 2, 0, 1, 1, 3, 4, 1, -2, -1, -2, 1, 1, -2, 0, -1, 1, 0, 1, 4, 5, 2, 1, 3, 2, 0, -1, -3, -1, 1, 1, 1, 1, 2, 4, 3, 1, 2, 0, 0, 0, 3, 0, 1, -2, 0, 0, 3, 0, 2, 1, 3, 1, 4, 0, 0, -3, -2, 0, 0, 4, 3, 3, 1, 0, 3, 0, -1, -1, -2, 0, 3, 1, 0, 0, 0, 0, 3, 1, 0, 1, 1, 3, 3, 0, 3, 0, -1, 0, 1, 1, 4, 2, 2, 3, 1, -1, 0, 0, 0, 1, 0, 1, 0, -3, -1, -1, 0, 0, 0, 1, 0, 3, 4, 4, 3, -3, 1, 1, 0, 4, 3, 1, 2, 1, 0, 0, 2, 0, 0, -1, -2, -2, -1, -2, -3, 0, 2, 2, 0, 1, 1, 1, 3, 2, 3, -4, 0, 0, 1, 2, 1, 4, 1, 2, 3, 0, -1, 2, 0, 0, -3, -3, -4, -4, -4, -3, 1, 1, 3, 2, 0, 2, 2, 2, 4, 0, 0, 0, 0, 0, 2, 3, 0, 1, 2, 2, 0, 1, 0, -1, -1, -4, -7, -4, -4, -2, 0, 1, 3, 1, 2, 0, 2, 4, 6, -2, 0, 0, -1, 1, 1, 0, 4, 0, 3, 0, 2, 2, 1, -1, -2, -4, -7, -4, -4, -4, -3, 2, 1, 3, 0, 0, 3, 4, 5, -4, 0, 0, 1, -1, 0, 3, 2, 4, 1, 0, 1, 0, 0, 0, -4, -5, -6, -5, -4, -3, 0, 0, 1, 0, 1, 1, 4, 4, 4, -2, 0, -1, 0, 0, 1, 0, 4, 4, 2, 1, 4, 2, 0, 0, -1, -5, -5, -6, -3, -1, -1, 0, 1, 2, 2, 2, 3, 2, 4, -5, 0, 1, -1, 1, 2, 3, 3, 2, 2, 2, 1, 2, 2, 2, 2, -1, -1, -3, -2, 0, 0, 0, 2, 1, 2, 2, 4, 1, 0, -1, 0, -2, 1, 1, 1, 3, 0, 4, 3, 2, 3, 2, 1, 2, 1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 3, 0, 2, 0, -2, 0, 2, 4, 3, 2, 0, 0, 1, 1, 5, 3, 1, 1, 3, 1, 0, 1, 0, 1, 0, 0, 0, 3, 0, 1, 0, 1, 1, 1, -1, 0, 0, 2, 1, 0, 1, 0, 0, 5, 1, 1, 0, 4, 4, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 1, 0, -1, -2, 0, 2, 0, 3, 2, 1, 2, -1, 1, 3, 1, 0, 2, 0, 1, 1, 2, 2, 2, 0, 3, 0, 3, 2, 3, 1, 0, 0, -1, 0, 0, 2, 0, 2, -1, 1, 0, 1, 1, 4, 2, 0, 0, 1, -1, 0, -2, 0, 1, 1, 2, 2, 3, 1, 1, 3, 0, 0, -1, 0, -1, -2, 1, 0, 2, 0, 0, 0, -1, -1, 0, 0, -3, -2, 0, -3, -2, 0, 4, 4, 4, 4, 3, 4, 2, 0, 2, 2, 0, 0, -1, -2, -1, 1, 2, 0, 1, 0, 0, -1, -4, -3, -2, -2, 0, 0, 0, 3, 4, 3, 5, 6, 4, 4, 3, 3, 0, -1, -2, -3, -3, -1, -1, 1, 0, 0, 0, 0, 0, -1, -2, -3, -1, -1, -1, 2, 5, 4, 3, 3, 6, 6, 1, 3, 3, 0, 2, -1, 0, -3, -2, 0, 0, 0, 1, -1, -2, -2, 0, -3, -4, -1, -1, -3, -1, 3, 5, 3, 4, 4, 6, 4, 1, 1, 2, 0, -1, -2, -1, -2, -1, -4, 0, 0, -1, 0, 1, -2, -2, -4, -4, 0, 1, 0, 0, 3, 1, 2, 5, 5, 2, 2, 3, 1, 0, 1, -2, -1, -1, -5, -3, -3, -1, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 4, 2, 4, 1, 3, 2, 2, 0, -1, 0, 1, -2, -1, -2, -4, -6, 0, -1, 1, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 3, 2, 0, 2, 0, 0, 1, 1, 3, 0, 0, -2, -2, -2, -2, 0, -3, -1, -1, -1, 0, 2, 0, -1, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 2, 2, 0, 2, 3, 0, 0, -1, 1, 1, -1, 0, -2, 0, 0, 0, 0, 2, 2, 1, 1, 0, -1, 1, 0, -1, 0, 2, 1, 1, 2, 2, 1, 0, 2, 2, 0, 1, 0, 2, -1, 0, 1, 0, -1, 0, 1, 2, -1, -1, -1, -1, 0, 1, -1, 0, 0, 2, 2, 0, 2, 0, 1, 2, 2, 1, 2, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 4, 2, 1, 0, 2, 2, 0, 2, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 2, 0, 1, -1, 0, -1, -1, 0, 0, 2, 3, 2, 2, 4, 0, 2, 1, 1, 0, 2, 0, -1, -1, -1, 2, 0, 1, 0, 2, 1, 3, 2, 1, 0, 1, -1, 0, 1, -1, 0, 2, 0, 2, 0, 3, 1, 0, 2, 0, 0, 0, 0, -1, 0, 1, 3, 0, 1, 1, 2, 2, 2, 3, 2, 0, -2, -2, 0, 0, 1, -1, 0, 2, 3, 0, 0, 1, 2, 0, 0, 0, 1, 2, 1, 1, 2, 0, 0, 2, 0, 3, 1, 1, 0, 0, -3, 0, 0, -1, 0, 2, 2, 0, 2, 2, 1, 3, 2, 0, 2, 1, 2, -1, 0, 0, 1, 2, 2, 0, 1, 1, 0, 1, 0, -2, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 3, 0, 0, 2, 2, 2, -1, 1, 0, 0, -1, 0, -2, -1, -1, 0, 2, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 4, 0, 0, 3, 0, 0, 1, 2, -2, -2, 1, 0, -1, 1, 1, -1, 2, 0, 0, 1, 2, 3, 2, 1, 3, 1, 2, 1, 0, 0, 2, 1, 2, 3, 2, 1, 0, 0, 0, -1, 0, -2, 0, 0, -2, 0, 0, 2, 1, 1, 0, 1, 0, 3, 1, 0, 1, 2, 2, 1, 0, 0, 1, 4, 4, 1, 2, 2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 3, 4, 3, 0, 2, 0, 0, 0, 2, 1, 2, 3, 3, 1, 0, 1, 0, -1, 0, 0, -2, -1, 0, 0, -2, 1, 1, 2, 1, 3, 1, 3, 1, 4, -1, 0, 1, 1, 0, 0, 2, 2, 0, 1, 2, 2, 0, -1, 0, -2, -1, -2, 0, 0, 0, 0, 0, 1, 3, 3, 2, 3, 1, 0, -1, 0, 1, 0, 3, 1, 2, 2, 1, 0, 1, 1, 0, 1, 0, 0, 0, -2, 0, 0, -1, -1, 2, 1, 0, 0, 0, 2, 3, 0, 0, 0, 2, 2, 3, 0, 1, 3, 2, 0, 0, 1, 0, 1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 2, 0, 0, 3, 3, 1, 1, 0, 0, 0, 0, 2, 3, 1, 1, 1, 1, 2, 0, 1, 0, 1, -1, -1, -1, 0, 0, 2, 2, 3, 2, 3, 2, 0, 3, 1, 1, 0, 0, -1, 2, 0, 1, 2, 3, 0, 2, 3, 1, 1, 0, 1, 1, 1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 2, 3, 3, 1, 2, 1, 0, 0, 0, 2, 2, 1, 2, 0, 1, 3, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 3, 1, 2, 2, 0, 0, 0, 0, 2, 0, 3, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, -1, 0, -1, 0, 2, 2, 0, 2, 0, 0, 2, 2, 1, 0, 2, 1, 0, 1, 1, 0, 2, 1, 2, 2, 1, 2, 2, 0, 1, 1, 1, 1, -1, 2, 0, 0, 1, 0, 0, 1, 2, 0, 2, 1, 0, 1, 0, 1, 0, 0, 0, 3, 0, 0, 2, 0, 0, -1, 0, 0, 0, -1, 1, 0, 1, 0, 3, 2, 2, 1, 3, 2, 0, 0, 0, 0, 0, 0, 1, 1, 2, 0, 1, 0, 2, 2, 0, -1, 0, -1, -1, 0, 1, 0, 2, 3, 4, 1, 0, 2, 0, 0, 0, 2, 1, -1, -1, 2, 2, 1, 0, 0, 3, 1, 1, -1, -2, 0, 0, 0, 0, -1, 0, 3, 1, 2, 3, 2, 3, 2, 1, 0, 1, 2, -1, -1, 0, 0, 2, 0, 1, 0, 2, 2, 2, 0, 0, -2, -2, 0, -1, 1, 2, 0, 3, 3, 4, 1, 3, 0, 3, 1, -1, 0, 1, -2, 1, 2, 0, 2, 2, 2, 2, 0, -1, -2, 0, 0, -1, -1, 0, 2, 2, 1, 3, 0, 2, 3, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 3, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 3, 2, 2, 1, 0, 0, 2, 1, 2, 1, 0, 1, 0, 2, 0, -1, 2, -1, 2, 0, -1, 0, 0, -1, -3, 0, 2, 3, 3, 1, 0, 1, 2, 3, 6, 3, 6, 6, 5, 5, 4, 6, 4, 4, 4, 4, 0, 1, -3, -1, -4, -5, -2, -1, -2, 0, -1, 0, 2, 0, 0, -1, -1, 2, 0, 3, 4, 4, 5, 7, 6, 7, 7, 6, 5, 6, 2, 1, -1, -1, -2, -1, 0, -2, -1, -3, 0, 2, 1, -1, 0, -2, -4, 0, 0, 1, 1, 3, 3, 5, 3, 7, 8, 8, 5, 5, 5, 3, 0, 1, 1, 0, -1, -3, -2, 0, 0, 0, 2, 2, 0, -1, 0, -3, -2, 0, -1, 2, 0, 0, 2, 5, 8, 8, 8, 4, 6, 3, 0, 1, 1, -1, 2, -2, 0, 0, -1, 0, 1, 3, 0, 0, 0, 0, -1, -1, 0, -1, 0, 3, 4, 4, 8, 7, 6, 5, 2, 4, 3, 1, 3, 0, 2, -2, -2, 0, 0, 1, 3, 6, 3, 5, 2, 4, 0, 0, -2, 0, -1, 1, 2, 4, 6, 5, 5, 3, 4, 5, 5, 5, 5, 1, 0, -1, 0, 1, 1, 0, 2, 6, 5, 4, 3, 3, 3, -3, -4, -5, -3, 0, 2, 0, 3, 3, 4, 4, 4, 4, 5, 6, 7, 3, 1, -2, 0, 2, 2, 3, 6, 5, 6, 4, 5, 3, 5, 0, -5, -4, -3, 0, -2, -1, 0, 0, 3, 4, 7, 4, 6, 5, 7, 2, 2, 0, -2, 1, 3, 2, 5, 5, 3, 4, 5, 6, 2, -2, -3, -2, 1, 0, 0, 0, 0, 0, 0, 1, 5, 6, 8, 4, 7, 5, 3, -2, 1, 1, 2, 4, 5, 5, 5, 2, 5, 3, 1, -2, -3, -3, 0, 2, -2, 0, 0, -1, 1, 2, 2, 4, 7, 7, 6, 7, 3, -3, 1, 4, 3, 6, 8, 6, 4, 4, 5, 0, -1, 0, -1, -3, 0, -2, -3, -4, -3, -1, 2, 2, 3, 5, 3, 7, 7, 7, 8, 0, 0, 1, 3, 6, 6, 6, 4, 5, 2, 2, 0, 0, 0, 0, -4, -2, -7, -5, -2, 0, 1, 0, 0, 4, 5, 7, 6, 9, 8, -3, 0, 1, 1, 6, 5, 4, 5, 7, 3, 2, 0, 0, 0, 0, -4, -4, -9, -8, -7, -3, 1, 3, 2, 4, 2, 6, 8, 9, 8, 0, 0, 3, 2, 5, 2, 6, 7, 6, 5, 2, 3, 1, -2, -5, -6, -8, -11, -8, -6, -3, -2, 4, 5, 3, 2, 4, 7, 7, 10, -2, 1, 0, 3, 3, 2, 4, 5, 6, 3, 4, 1, 2, 0, -6, -8, -11, -10, -12, -10, -5, -1, 1, 1, 3, 2, 7, 9, 10, 9, -1, 1, 2, 2, 2, 3, 4, 6, 4, 5, 3, 1, 3, 1, -3, -6, -8, -10, -12, -8, -6, -6, 1, 3, 2, 3, 7, 10, 11, 11, -3, 0, 0, 3, 3, 3, 5, 5, 4, 7, 2, 2, 4, 1, 0, -6, -7, -9, -11, -10, -6, -2, 1, 1, 6, 6, 8, 9, 11, 6, -3, -1, 1, 0, 2, 4, 5, 4, 5, 4, 4, 6, 3, 1, 3, 0, -5, -5, -6, -5, -4, 0, -1, 3, 4, 4, 6, 7, 4, 6, -4, -1, 0, 4, 6, 4, 2, 3, 6, 4, 4, 6, 3, 1, 3, 0, -2, -2, 0, -3, 1, 0, 0, 1, 5, 6, 5, 6, 2, 2, -2, 2, 3, 2, 6, 4, 4, 4, 4, 4, 5, 5, 0, 1, 2, 2, 3, 0, 2, -1, 1, 2, 2, 3, 1, 4, 2, 2, 3, 2, 0, 1, 3, 5, 2, 5, 4, 3, 4, 6, 7, 4, 0, 2, 0, 4, 0, 1, 0, -1, 0, 0, 1, 2, 4, 3, 1, 3, 2, 0, 1, 2, 1, 2, 4, 2, 1, 3, 2, 4, 5, 4, 2, 1, -1, 0, 0, 0, 2, 3, 1, 2, 2, 4, 4, 2, 1, 3, 3, 0, 0, 3, 2, 4, 3, 2, 0, 1, 2, 2, 2, 2, 2, 1, -1, -4, 0, -1, 3, 1, 4, 5, 6, 5, 5, 4, 2, 5, 1, 1, 0, 0, 1, 2, 3, 3, 2, 3, 3, 3, 0, 0, -2, -3, 0, -2, -2, 0, 1, 2, 6, 6, 4, 6, 4, 5, 2, 2, 2, 2, -2, 0, 0, 0, 1, 0, 1, 1, 2, 0, 0, -2, -2, 0, -2, 0, 0, 4, 3, 4, 6, 7, 6, 7, 5, 6, 6, 0, 1, -1, -1, 1, 0, 2, 2, 4, 0, 0, 0, 0, -3, -1, -1, -2, 0, 0, 1, 5, 7, 8, 7, 10, 8, 8, 7, 6, 4, 3, -1, -3, -2, -2, 2, 1, 1, 3, 1, 0, -3, -4, -4, -3, -2, -2, 2, 2, 6, 5, 7, 10, 6, 9, 8, 8, 4, 4, 1, 0, 0, -1, -2, -4, -2, 0, 3, 0, 1, -1, 0, -3, -3, -1, -2, 0, 0, 3, 6, 8, 6, 7, 8, 7, 3, 4, 5, 3, 1, -1, -4, -2, -2, -4, -2, 0, 3, 0, 3, 1, 2, 0, 2, 4, 3, 2, 5, 5, 4, 4, 6, 5, 5, 5, 4, 2, 2, 0, 0, -3, -2, -3, -2, -2, 0, 0, 3, 5, 2, 2, 5, 5, 8, 7, 6, 5, 7, 5, 8, 8, 5, 4, 2, 0, 0, 1, -1, 0, -3, -5, -2, -7, 0, 1, 2, 1, 2, 0, 0, 1, 1, 3, 4, 0, 0, 3, 0, 3, 2, -1, -1, 1, 0, -1, -2, -2, -1, -1, -1, -4, -4, 0, 0, 1, 0, 2, 0, 0, 1, 2, 0, 2, 3, 3, 0, 1, 0, 2, 0, 0, 3, 1, -1, 1, 0, 0, -3, -1, 0, -4, -4, -1, 0, 0, 2, 3, 0, 0, 0, 0, 0, 2, 2, 2, 2, 1, 3, 2, 0, 0, 2, 0, 2, 1, 0, 1, 0, -1, -2, -1, -2, 0, 1, 1, 0, 3, 0, -1, -2, 0, -2, 0, 0, 1, 1, -1, 0, 3, 3, 1, 0, 2, 0, 0, 1, 0, 0, -2, -1, -1, -1, -2, 1, 0, 0, 2, 3, 1, -2, -1, -3, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 0, 0, 1, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 2, 0, 0, -1, 0, 0, -3, -1, -1, -2, 0, 0, 0, 1, 3, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 3, 4, 0, 0, 1, 0, -2, 0, 0, 0, 1, 1, 2, 3, 3, 3, 0, 1, 1, 2, 0, 0, 1, 0, 0, -2, 0, 0, 0, 1, 3, 3, 2, 1, 0, 1, 0, -2, -2, -2, 0, 0, 0, 1, 1, 0, 2, 1, 2, 0, 0, 2, 0, -2, 0, -2, 2, 0, 2, 0, 3, 0, 2, 0, 0, 0, 1, -1, 0, -3, 1, 0, 1, 0, 0, 1, 1, 3, 0, 1, 2, 3, 1, 1, 1, -2, 1, 2, 2, 1, 3, 2, 3, 0, 2, 0, 0, 0, 0, -2, 0, 1, -1, -2, 0, -1, 0, 3, 0, 1, 3, 0, 0, 0, 0, 0, -1, 2, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -3, -2, 0, 0, 0, -1, -2, 1, 0, 3, -1, 2, 0, 0, 3, 0, 0, -1, 1, 2, 0, 3, 3, 3, 0, 0, 2, 1, 0, -2, 0, -3, -3, -1, 0, 0, 1, 1, 0, 0, -1, 0, 1, 1, 2, 3, 1, 0, 2, 1, 2, 3, 3, 2, 3, 2, 0, -1, -1, -1, -1, -1, -4, -1, -1, 0, -1, 0, 1, 0, 0, 0, 2, 3, 3, 2, 1, 1, 2, 3, 3, 3, 1, 4, 1, 2, 3, 1, 0, -1, 0, -1, -3, -4, -1, -1, -2, 0, 1, 1, 3, 2, 0, 2, 2, 1, 0, -1, 1, 2, 2, 0, 0, 1, 2, 0, 2, 0, 0, -2, -2, -3, -4, -1, -4, -2, -1, 0, 3, 3, 0, 0, 0, 2, 4, 3, 3, 2, 1, 0, 1, 2, 1, 1, 2, 3, 1, 0, 0, 0, -2, -1, -2, -5, -3, -4, -4, 0, 1, 0, 4, 2, 0, 2, 2, 1, 0, 3, 0, 2, 0, 0, 0, 1, 1, 1, 0, 1, 0, -1, -1, -3, -2, -4, -4, -3, -3, 0, -2, 0, 3, 0, 2, 2, 3, 1, 1, 1, 0, 0, 1, 2, 3, 1, 2, 2, 2, 2, -1, 0, -2, 0, -3, -3, -4, -2, -2, -2, -3, 2, 3, 1, 1, 2, 1, 1, 0, 1, 2, 3, 1, 0, -1, -1, 1, 3, 0, -1, 0, 1, 0, 0, -3, -1, -4, -4, -1, -3, -3, 0, 0, 3, 0, 0, 1, 3, 2, 0, 0, 2, 2, 0, 2, 0, 0, 2, 1, 2, 1, -2, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, 2, 1, 2, 3, 0, 2, 0, 0, 0, 2, 0, 2, 0, 1, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 2, 1, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 2, -2, 0, -2, 0, 1, 0, 0, 1, 0, 1, -1, 2, 0, 2, -1, 2, 2, 1, 1, 0, 1, 0, 2, 1, 0, 1, 0, 2, 3, 0, 1, 0, 0, -1, 0, 1, -1, 1, 0, 0, -1, 0, 1, 0, 0, 1, 2, -1, 0, 0, 0, 3, 2, 0, -1, -1, 0, 0, 2, 2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 1, 0, 2, 0, 1, 1, 0, 0, 2, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, 2, 2, 0, 1, 1, 0, 0, 2, 1, 1, -1, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, -1, -1, 1, -2, -1, 1, -1, 0, 3, 0, 2, 1, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 2, 0, 0, 2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 1, 0, 0, 3, 3, 0, 2, 0, 2, 0, 1, -2, -2, -2, 1, 2, 1, 2, 1, -1, 0, 1, -2, -2, 0, 0, 0, 0, 1, 2, 0, 0, 3, 1, 2, 1, 2, 3, 0, 0, -1, 0, -2, -2, 2, 1, 2, 2, 0, -1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 3, 2, 0, 3, 1, 2, 1, 2, 2, 3, 0, -1, 0, -1, 0, -1, 1, 0, 3, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 2, 0, 3, 2, 0, 0, 0, 0, 1, 0, 0, -1, 0, -2, -1, -3, -1, 0, 1, -1, -1, -1, 2, -1, 0, 0, -1, 0, 1, 0, 0, 2, 1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 1, -1, 0, 0, 1, 1, 0, -1, 0, -1, 1, -1, 0, 1, -1, 0, 0, 2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, -1, 1, 0, 1, 0, -2, 0, 2, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, -1, 1, 1, -1, 1, 2, 0, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 1, 0, 2, 0, 0, 0, 2, -1, 0, 0, 1, 1, 1, 1, 0, 1, -1, 0, -1, 0, -2, 0, 1, 0, 0, 0, 1, 0, 0, -2, 0, 1, 0, 1, 0, 0, 1, -1, 0, 0, 1, 0, 0, -1, 1, 0, 1, 0, 1, -1, 0, 1, -1, 0, 0, 1, 1, 1, 1, -1, 0, 0, 0, -2, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, -1, 1, -1, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 2, 1, 0, 0, -2, 0, 0, 0, 2, 0, 0, 1, 1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, -1, 1, 0, -1, 0, 0, 1, -2, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 2, 1, 0, 0, -1, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 1, 0, 1, 1, 0, 0, 1, 0, 2, 1, -1, 0, 1, 1, 0, -1, 1, 0, -2, 1, -1, -1, 0, -1, 1, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -2, 0, 1, 1, 0, 1, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 1, -1, 0, -1, 0, -1, 2, -1, 1, -1, 0, 1, -2, 1, 0, 0, -2, -2, 1, -1, 0, 0, 0, -1, 0, 1, 0, -1, -2, -1, 0, 1, -1, 1, -1, 0, 0, 1, -1, -1, 1, 1, -1, 0, -1, 0, 0, 2, 1, -1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, 1, -1, 0, -1, 0, 0, -1, 0, 0, -2, -1, 1, 0, -1, -1, 0, 0, 2, -1, 0, 2, -1, 0, 0, -1, 0, 1, -1, -1, 0, 1, 0, 0, 1, -2, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, -1, 0, -2, 0, 0, 0, 0, -1, -1, 1, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 2, 1, -1, 0, -1, 2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, -1, 1, -1, 1, 1, 0, 0, -2, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 1, -1, 1, 0, -1, 0, 0, 0, -1, 1, 1, 0, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, 1, -1, -2, 0, 0, -1, 0, 2, 1, -1, 0, -1, 2, -1, 1, -1, 1, -1, 1, -1, 0, 1, 0, 1, 0, 1, -1, 1, 0, 0, 0, 1, 1, 1, 1, -1, 0, 1, -1, 0, 0, 1, 0, -1, -1, 1, 0, -1, -1, 0, 0, -1, 1, 1, -1, 1, -1, 0, 0, 1, 0, -1, 0, 0, 0, -2, 0, 1, -1, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 1, -2, 0, -1, -1, -2, 0, 1, 0, -2, 1, 1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 0, -1, 1, 0, 1, -1, -1, 0, 1, -1, 1, -1, 0, 2, 0, 0, -1, 1, 0, 2, 0, -1, 0, 1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, -2, 0, 0, -1, -1, -1, 0, -1, 0, 1, 0, -1, 0, 0, -1, -1, 0, 1, 2, 1, 0, 0, 0, -1, 0, 2, 0, -1, 0, -1, -2, 0, 0, -1, 0, -1, 0, -1, -1, 1, -1, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, 0, 0, -2, 0, -2, -1, 0, 0, 0, 1, 1, -1, 0, 0, 2, -1, 1, 1, 0, 1, 1, 0, -1, 1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 2, -1, 0, -1, -1, -1, -1, -1, -1, 2, 0, 0, -1, -2, 0, 1, 0, -1, 1, -1, 1, 1, -1, -1, -1, 0, 1, 0, -1, 1, 0, 1, -1, 1, 0, -1, 0, -1, 1, 2, 1, 1, 0, 0, 0, -1,
    -- filter=0 channel=1
    2, 1, 1, 3, 0, 0, 2, 0, 1, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 2, 3, 0, 3, 0, 2, 1, 0, 2, 2, 0, 4, 1, 1, 4, 3, 1, -1, 1, 3, 1, 1, 3, 1, 2, 0, 3, 1, -1, -1, 3, 1, 3, 3, 2, 1, 3, 4, 1, 2, 2, 3, 1, 2, 0, 2, 0, 4, 2, 1, 3, 3, 2, 2, 2, 3, 3, 1, 2, 0, 1, 1, 2, 1, 0, 2, 3, 3, 4, 2, 4, 1, 1, 2, 2, 3, 3, 3, 2, 4, 3, 2, 4, 5, 4, 2, 2, 0, 0, 2, 2, 1, 2, 2, 3, 3, 1, 0, 2, 0, 1, 2, 1, 3, 1, 4, 5, 1, 3, 2, 2, 2, 2, 3, 3, 3, 4, 0, 0, 1, 2, 0, 0, 0, 1, 3, 1, 3, 1, 3, 1, 2, 1, 4, 1, 1, 3, 1, 3, 1, 4, 3, 3, 1, 5, 3, 4, 1, 1, 0, 0, 0, 2, 0, 2, 2, 1, 1, 5, 2, 1, 1, 0, 3, 2, 3, 4, 4, 3, 1, 3, 1, 4, 2, 2, 4, 3, 2, 0, 0, 2, 2, 2, 0, 3, 3, 1, 2, 1, 2, 1, 1, 4, 2, 3, 2, 4, 2, 3, 2, 3, 4, 3, 4, 2, 3, 3, 1, 2, 1, 1, -1, -1, 1, 3, 3, 2, 4, 1, 5, 1, 1, 0, 3, 2, 5, 5, 2, 3, 3, 5, 3, 3, 1, 4, 3, 5, 3, 0, 0, -1, 0, 1, 2, 0, 0, 1, 5, 2, 4, 1, 1, 1, 3, 3, 2, 5, 2, 4, 1, 1, 1, 4, 4, 3, 2, 6, 1, 1, 0, 1, 0, 1, 1, 0, 3, 4, 5, 5, 5, 4, 2, 2, 5, 6, 4, 4, 3, 2, 2, 3, 3, 1, 3, 5, 4, 4, 5, 1, -1, 1, 0, 2, 0, 3, 1, 3, 4, 3, 2, 2, 4, 5, 2, 4, 4, 1, 1, 1, 3, 3, 1, 2, 5, 5, 5, 5, 2, 2, 0, 0, 0, 0, 2, 1, 3, 4, 4, 3, 3, 4, 4, 4, 1, 1, 4, 1, 3, 3, 2, 3, 4, 5, 5, 5, 4, 4, 5, 1, 0, 1, 3, 2, 0, 0, 1, 5, 6, 4, 4, 4, 2, 2, 1, 5, 4, 5, 3, 1, 4, 2, 2, 1, 3, 4, 8, 4, 5, 1, 0, 0, 0, 0, 0, 0, 4, 5, 6, 3, 5, 2, 4, 2, 1, 4, 4, 3, 1, 2, 4, 3, 1, 4, 5, 5, 4, 7, 5, 3, 0, -1, 1, 0, 0, 1, 3, 4, 3, 5, 4, 2, 5, 3, 3, 3, 3, 2, 1, 4, 1, 2, 3, 1, 5, 4, 6, 4, 3, 2, 2, 0, 0, 0, 0, 0, 1, 4, 1, 4, 4, 2, 3, 5, 3, 4, 5, 3, 2, 3, 1, 1, 2, 1, 4, 6, 5, 6, 5, 3, 3, 1, 0, 0, 0, 1, 3, 2, 4, 2, 1, 3, 2, 3, 4, 5, 4, 3, 3, 2, 4, 3, 3, 3, 5, 5, 5, 6, 3, 3, 0, 0, 0, 0, 1, 1, 3, 1, 3, 3, 3, 3, 3, 1, 2, 2, 4, 6, 1, 3, 2, 3, 1, 5, 5, 6, 5, 3, 5, 3, 1, 0, 1, 0, 1, 0, 2, 3, 2, 3, 5, 4, 3, 1, 1, 3, 2, 3, 3, 3, 3, 2, 3, 3, 3, 6, 4, 4, 4, 3, 0, 2, 0, 1, 0, 0, 1, 2, 4, 4, 1, 1, 1, 4, 5, 3, 4, 2, 4, 2, 2, 3, 5, 4, 3, 3, 3, 4, 3, 2, 2, 0, 2, 0, 2, 3, 1, 1, 4, 5, 1, 3, 0, 5, 4, 5, 2, 2, 2, 0, 5, 1, 5, 4, 3, 4, 3, 1, 1, 2, 0, 0, 0, 0, 1, 0, 2, 4, 1, 1, 3, 1, 1, 2, 4, 5, 2, 2, 0, 2, 5, 4, 2, 5, 4, 5, 5, 3, 4, 2, -1, 2, 1, 2, 2, 0, 2, 1, 0, 2, 0, 1, 2, 2, 3, 1, 4, 3, 5, 5, 5, 5, 3, 5, 3, 2, 3, 4, 1, 2, 0, 0, 1, 2, 0, 1, 1, 1, 2, 1, 0, 2, 2, 4, 2, 2, 4, 2, 4, 4, 1, 2, 4, 2, 5, 2, 4, 4, 0, 2, 1, 1, 0, 2, 2, 0, 1, 0, 2, 0, 0, 1, 2, 3, 4, 3, 4, 5, 3, 1, 4, 4, 2, 4, 4, 4, 4, 3, 0, 1, -1, 2, 1, 0, 1, 3, 1, 3, 0, 1, 3, 0, 1, 2, 4, 4, 5, 2, 5, 2, 4, 3, 3, 6, 4, 5, 2, 2, 0, 0, -1, 0, 0, 3, 3, 3, 2, 0, 0, 0, 2, 1, 0, 3, 3, 1, 1, 4, 4, 1, 1, 4, 2, 4, 3, 1, 2, 1, 0, 1, 0, 2, 0, 1, 1, 0, 3, 3, 3, 3, 1, 0, 0, 2, 2, 0, 3, 1, 2, 0, 2, 1, 3, 2, 0, 0, 1, -1, 0, -1, 0, 0, 4, 2, 1, 4, 0, 3, 3, 2, 3, 0, 1, 3, 3, 0, 0, 1, 1, 0, 0, -1, 0, 1, -1, 0, 0, -1, -2, 0, 0, -7, -5, -8, -5, -6, -4, -4, -2, -4, -5, -6, -4, -2, -1, -5, 0, -1, -1, 2, 0, 2, 7, 7, 7, 9, 9, 5, 9, 8, 6, -3, -3, -6, -4, -6, -2, -5, -1, -2, -3, -3, -3, 0, -1, -1, 0, -3, 1, 2, 0, 1, 4, 3, 3, 5, 6, 6, 4, 5, 6, -3, -6, -5, -4, -6, -5, -2, 0, 0, 1, 0, 0, 0, 0, 0, -4, -2, -2, 0, 1, -1, 0, 0, 0, 3, 2, 2, 4, 4, 7, -3, -6, -5, -4, -5, -4, -1, -1, -1, -2, 1, 0, -2, -1, -1, -3, -1, -2, 0, -1, 1, -1, 0, -3, -3, 0, -2, 0, 3, 3, -3, -4, -5, -2, -5, -3, -3, 0, 0, 0, 1, 0, 0, 1, 0, 1, -2, -2, -2, 0, 0, 0, -3, 0, -2, -1, -1, -2, 0, 3, -6, -4, -3, -5, -5, -3, -1, -2, -2, -1, 0, 1, 0, 0, 1, 2, 0, -1, -3, 0, -1, 0, 0, 0, -1, -3, -2, 0, 3, 1, -4, -5, -5, -2, -2, -3, -3, 0, -1, -1, 0, 2, 3, 2, 5, 4, 0, -1, -1, 1, 0, 1, 0, -2, -3, -2, -2, 0, 0, 1, -4, -1, -2, -2, -2, -3, 0, 0, -3, 0, 2, 1, 3, 4, 5, 2, 4, 1, -2, -1, 0, 1, 0, -1, -2, -1, -2, 2, 3, 1, -5, -2, 0, 1, 0, -2, -1, 0, -2, 1, 1, 1, 5, 3, 3, 3, 3, 0, -2, -1, -3, -1, 0, 0, -3, -1, -1, 0, -1, 3, -4, -1, 0, 1, 0, -1, -1, 1, 1, 0, 1, 5, 6, 4, 4, 3, 4, 1, -2, -2, -2, 0, -3, -2, -2, -3, -1, -2, 0, 0, -4, -2, -1, 1, 1, 0, 0, 1, 0, 3, 2, 3, 5, 5, 8, 4, 4, 1, 1, 0, -3, 0, -1, -1, -2, -1, -1, -1, -2, -1, -1, -1, 0, -1, 0, 0, 2, 1, 3, 5, 2, 5, 5, 8, 5, 4, 2, 2, -1, 0, -3, 0, -3, -3, -2, 0, -1, 0, 0, -1, -2, -2, 0, 0, 2, 2, 3, 3, 2, 5, 5, 9, 8, 7, 7, 3, 4, 3, 0, 0, -1, 0, 1, 0, -3, -1, -1, -5, -3, -1, -3, 0, -3, -2, 1, 2, 3, 4, 3, 6, 4, 8, 10, 7, 7, 8, 4, 0, 0, -1, -2, 0, -1, 2, -2, -1, -4, -2, -1, 0, -2, -1, -3, 0, 1, 3, 2, 5, 5, 3, 7, 7, 7, 8, 8, 5, 3, 0, 1, 0, -3, 0, -2, 0, 0, 0, -4, -1, -2, 0, -1, 0, 0, -1, 2, 2, 3, 4, 5, 3, 5, 9, 9, 9, 9, 7, 3, 0, 1, 0, -2, -3, -2, 0, 0, 0, -4, -2, -2, 0, -4, -3, -2, -1, 2, 1, 1, 5, 4, 3, 6, 9, 9, 9, 6, 6, 3, 1, 1, -1, -2, -2, 0, 2, 0, -1, -3, -4, 0, 0, -4, -2, 0, 0, 0, 1, 1, 1, 1, 5, 5, 5, 7, 10, 7, 6, 1, 2, -1, -1, 0, -1, 0, 0, 0, 0, -1, -4, -2, 1, -2, -3, -2, -1, 0, 3, 1, 1, 3, 4, 7, 5, 5, 9, 9, 5, 6, 3, 0, -1, 0, 1, 2, 1, 0, -2, -1, -3, 0, 1, -4, -4, -2, -1, 0, 0, 0, 0, 1, 2, 4, 3, 8, 5, 8, 6, 2, 2, 0, 0, 0, 0, 0, 0, -2, -3, -2, -2, 0, 0, -4, -4, -4, -1, 0, 2, 1, 3, 3, 4, 4, 4, 6, 7, 5, 6, 2, 0, 0, 0, -1, 0, 0, -3, -2, -4, -3, -2, 2, 3, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 4, 6, 4, 2, 2, 1, -1, 1, 0, -2, 1, -3, -1, -1, -3, 0, 0, 2, 1, -2, -3, -2, -1, 0, 0, 0, 0, -1, 0, 1, 3, 6, 2, 4, 0, 3, -1, 0, -1, 0, -2, -1, -2, -2, -1, 0, 1, 0, 4, -2, -4, -4, -1, -2, 0, -1, -1, -1, -1, 2, 1, 4, 1, 2, 3, 2, 0, 0, -1, 0, -3, 0, -1, -1, -2, 0, 0, 2, 3, -2, -2, -4, -2, -2, -3, -3, 0, -1, -1, 3, 4, 2, 3, 1, 2, 2, 1, -1, 1, 0, -3, -1, 0, -3, 0, -2, 0, 0, 5, -3, -2, -2, -3, -2, 0, -2, -4, 0, 1, 0, 2, 4, 5, 4, 1, 1, 0, 0, -1, -3, -2, -3, 0, 0, -3, -2, 0, 2, 5, -5, -1, -4, -2, -1, 0, -3, -5, -3, 0, 0, 2, 4, 2, 1, 2, 4, -1, 0, -2, -4, -1, -4, -2, -4, -4, -2, 0, 3, 4, -5, -2, -1, -4, -3, -1, -1, -4, -2, 0, 1, -1, -1, 1, 3, 2, 0, 0, 0, -2, 0, 0, -3, -1, -5, -4, 0, 0, 0, 2, -2, -4, -4, -4, -2, -3, -2, -3, -2, -3, 0, -1, -1, 0, 0, 1, 0, -2, -2, -1, -1, -1, 0, -2, -3, -2, 1, 3, 3, 3, -6, -4, -3, -3, -4, -4, -4, -4, -1, -3, -4, -2, -2, -3, 0, -3, -2, 1, 0, 0, 1, 0, 0, 1, 3, 2, 4, 6, 6, 7, -5, -4, -5, -5, -5, -2, -4, -5, -2, -4, -2, -1, -3, 0, 0, 0, -1, -2, 0, 0, 0, 0, 2, 2, 2, 3, 4, 4, 1, 1, -5, -4, -2, -1, -5, -2, -2, -1, 0, 0, -2, -2, 0, 0, -1, 0, 0, -1, 1, 1, 1, -1, 0, 0, 2, 4, 1, 2, 3, 0, -1, -3, -4, -1, -4, -2, -3, -1, 0, 0, 0, 1, 2, 0, 1, -2, -1, 1, 0, 0, 0, 0, 2, 0, 2, 2, 0, 0, 0, 2, -3, -3, -1, -2, -2, -2, -1, 0, 0, -1, 0, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 1, -2, 0, 0, -2, 0, 0, 1, 0, -4, -2, -4, -1, -4, -1, 0, 0, -1, 0, 1, -1, 2, 3, 0, 0, 1, 0, 1, 0, 2, 0, 0, -2, -2, 0, -1, -3, 0, -1, -5, -5, -3, -4, -4, -2, -3, 0, 1, 0, 1, 2, 1, 3, 3, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, -1, 0, 0, 0, 1, -3, -3, -1, -1, -1, 0, 0, 0, -1, 0, 1, 0, 2, 1, 3, 3, 0, 2, 2, 1, 0, -1, 1, 0, 0, 1, 0, 1, -1, 1, -4, -2, -2, -1, -3, 0, -1, -1, -1, 1, 2, 3, 3, 5, 3, 1, 2, 1, 0, 0, 0, 2, 2, 2, 1, -1, -1, 0, 0, -1, -2, -3, 0, -2, -1, -1, -1, 0, 0, 2, 2, 3, 6, 4, 2, 2, 2, 3, 2, 0, -1, 0, 2, 0, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 0, 0, -1, 1, 3, 4, 4, 4, 6, 5, 3, 2, 2, 0, 0, 0, 0, 2, 0, -1, 1, 0, 0, 0, 0, -2, -3, -4, -3, -1, -1, 0, 2, 0, 2, 4, 4, 4, 4, 4, 7, 6, 4, 3, 3, 1, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, -4, -1, 0, 0, 0, 1, 0, 1, 1, 6, 2, 5, 5, 5, 5, 4, 2, 3, 3, 3, 2, 0, 2, 0, -1, 1, 1, -1, 0, 0, -4, 0, -2, -1, -1, 2, 2, 1, 2, 6, 5, 4, 4, 6, 5, 3, 5, 4, 1, 0, 0, 0, 2, 0, 0, -2, -2, 0, -1, 0, -1, -2, -1, -3, 0, 0, 3, 2, 3, 5, 8, 5, 8, 6, 5, 6, 5, 5, 4, 4, 3, 0, 2, 2, 0, 0, 1, 0, 0, 0, -1, -1, -2, -1, 1, 0, 3, 3, 4, 5, 4, 5, 6, 5, 4, 6, 3, 3, 3, 4, 0, 2, 1, 0, 2, -1, 1, -2, 0, 1, -3, 0, 0, 0, 0, -1, 4, 2, 5, 4, 6, 4, 8, 7, 6, 4, 6, 1, 1, 3, 0, 0, 1, 0, 0, 0, -2, 0, -1, 0, -2, -1, 0, -1, 0, 2, 3, 1, 4, 4, 5, 6, 6, 9, 7, 4, 7, 3, 3, 0, 0, 2, 2, 3, 2, 1, 1, -2, 0, -1, -4, -4, 0, -2, 0, 0, 2, 4, 5, 6, 6, 5, 4, 6, 7, 7, 6, 1, 4, 2, 1, 0, 1, 1, 0, 0, 0, -2, 0, 0, -2, -2, -3, -3, 0, -1, 0, 1, 3, 5, 6, 5, 7, 7, 5, 4, 7, 3, 4, 1, 1, 1, 4, 3, 0, -1, -2, -1, 0, -2, -3, -4, -2, 0, -2, 0, 1, 2, 2, 2, 6, 3, 7, 7, 7, 5, 6, 2, 2, 1, 2, 1, 1, 3, 1, 0, -2, -1, -2, 0, -1, -1, -2, -2, -1, -1, 0, 2, 1, 3, 5, 4, 3, 6, 4, 2, 5, 2, 0, 3, 2, 0, 2, 0, -1, -2, -2, 0, 1, 2, -3, -3, -2, -4, -1, -1, 1, 0, 0, 3, 3, 5, 3, 5, 5, 1, 1, 1, 1, 0, 0, 2, 0, 1, 0, -1, -2, 0, 0, 0, -5, -2, -4, -2, -1, 0, 0, 1, 2, 1, 2, 2, 4, 4, 4, 1, 3, 3, 2, 1, 3, 0, 1, 2, -2, -1, 0, 1, 1, 0, -4, -3, -3, 0, 0, 0, -2, -2, 0, 1, 2, 3, 4, 2, 3, 3, 3, 3, 0, 1, 0, 1, 0, 1, -1, -1, 1, 1, 0, 0, -4, -1, -4, -1, 0, 0, 0, -2, 1, 2, 0, 0, 0, 4, 0, 0, 1, 2, 2, 2, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, -3, -2, -1, -1, 0, -2, 0, -3, -3, 0, -1, 0, 3, 4, 0, 3, 3, 0, 1, 0, 1, 0, 0, 0, 1, -2, -1, 0, 1, 1, -4, -1, -1, -3, -4, 0, -2, 0, 0, -2, -1, 0, 2, 1, 0, 2, 2, 0, 0, -1, 0, 0, -1, 0, -1, -3, -2, -1, -1, -1, -2, -4, -4, -1, -2, 0, -2, -1, -2, 0, 0, 0, -1, 0, -1, 1, 0, 1, 1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -1, -2, -3, -1, -3, -3, -2, -1, -2, -3, -2, 0, -2, 0, -2, 0, 0, -1, 0, 0, -1, -2, -3, -1, -2, -1, -2, -1, 0, 0, 0, -4, -1, -2, -2, -2, -2, -3, -3, -3, 0, -3, -3, -2, -1, -1, -1, 0, -1, -3, 0, -1, 0, -1, -1, 0, -1, 0, 0, 1, 0, -1, 0, 1, 1, -1, 0, -1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 1, 1, -1, -1, -1, 1, 1, 0, -1, 0, -1, 1, -1, 1, -1, 1, -1, 1, -1, 2, -1, 0, 1, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, -2, -1, 1, 0, -2, 0, 0, -1, 2, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 0, -1, -2, -2, 0, -1, 0, 1, -1, -1, 0, -1, 0, -1, -2, 0, 1, 1, -1, 0, 0, -1, 0, 0, -2, -1, -1, 1, 0, 0, 1, 1, 0, 0, 2, 0, 0, 1, 1, -1, 2, 0, -1, -1, -1, -1, 0, 0, 0, 1, 0, 0, 2, 0, -1, 0, -1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, -1, 0, -1, -1, 1, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, 0, -1, 1, -1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 2, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 1, -1, -1, -2, 1, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, 1, 0, 1, 0, 0, 1, 0, 2, 2, 0, 0, 0, -1, 1, 1, -1, 0, -1, 0, 1, 1, -1, -1, 1, 1, -1, 0, 1, 0, -1, 1, -1, 0, -1, 0, -1, 0, 1, 1, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, -1, 0, -1, -1, 1, 1, -2, 0, 1, 0, 0, 1, 0, 1, -1, 0, -1, 1, -1, -1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, -1, -1, -2, 0, -1, -2, -2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 2, 0, -2, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, -2, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 1, 0, -2, 0, 0, -1, 0, 1, 1, 1, -1, 1, 1, 2, 0, 0, 1, -1, -1, -1, 1, 1, 0, -1, 1, 0, 0, 0, -1, -1, 1, -1, 0, 1, 0, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, -1, 0, 1, -1, 0, 0, 0, 1, 1, 0, 0, -1, -2, 1, 0, -1, 1, -1, -1, -2, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, -2, 0, -1, -1, -1, 0, -2, 0, 1, 0, 1, -1, 0, -1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, 0, -1, 0, 1, 0, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, -1, 2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 1, 1, -1, 1, -1, 0, -1, 0, 0, 0, 1, -1, 0, -1, 1, -1, 0, 1, 0, 0, 0, 0, 0, 2, 0, -1, 1, -2, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 1, 0, -1, -1, 0, 1, 0, 1, -1, -1, 0, -1, 0, -1, 0, 0, -1, 1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 1, 1, 1, -2, -1, -1, 0, 1, 1, 1, 1, 1, -1, 0, 0, 0, 1, -2, 0, 1, 0, 1, 1, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 2, 1, -2, 0, -1, -1, -1, 0, 0, 0, -1, -2, 0, 1, 0, 1, 0, -1, 0, 0, 2, -1, -1, 0, -1, 0, -1, -1, 0, 0, -2, -1, -1, 0, 1, 0, -1, 2, -1, 0, -1, 0, 1, 1, 0, 0, 0, -2, 0, -1, 1, -1, -1, 0, 0, 0, 0, -1, 0, 2, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, 2, 0, -1, 0, 0, -1, 1, 0, 1, 2, 0, 0, -1, 0, 1, -1, -1, 1, 0, 0, -1, 0, 0, -1, -1, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 1, 1, 1, -1, -2, -1, 1, -1, -1, 0, 1, -1, 0, 1, 0, 1, 0, -1, -1, 1, -1, -1, 0, 0, 1, 1, 1, 0, -1, 0, 0, 0, 1, 0, -1, 2, 0, 0, 3, 1, 1, 3, 2, 2, 3, 4, 2, 1, 5, 3, 1, 5, 3, 4, 7, 8, 6, 7, 9, 8, 7, 7, 4, 3, 3, 3, 2, 0, 2, 2, 3, 2, 4, 3, 2, 0, 2, 3, 2, 0, 3, 1, 2, 3, 3, 4, 3, 5, 7, 7, 6, 5, 7, 4, 2, 2, 0, 0, 1, 2, 1, 4, 1, 2, 2, 2, 2, 2, 1, 0, 3, 3, 0, 0, 2, -1, 0, 0, 1, 2, 2, 2, 3, 0, 3, 0, 4, 0, 4, 5, 4, 2, 1, 0, 1, 0, 0, 2, 2, 0, 1, 1, 0, -2, -2, -2, -1, -3, 0, -2, 2, 2, 3, 1, 4, 0, 1, 2, 3, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, -2, -1, 0, -1, -2, 1, 3, 1, 4, 1, 2, 0, 1, 0, 2, 0, 0, 0, 1, 0, 0, 3, 3, 2, 2, -1, 1, 1, -1, -3, 0, -1, -1, 0, 0, 0, 0, 1, 1, 2, 1, 0, 3, 0, 2, 2, -1, 0, -2, 0, 2, 2, 5, 3, 1, 0, -1, 1, 0, 1, 0, -1, 0, 0, 0, 0, 2, 2, 2, 1, 2, 4, 0, 1, 0, 0, 0, 0, 1, 1, 1, 4, 2, 3, 1, 0, -1, -1, 1, -1, -2, 0, -2, 0, 0, 0, 1, 4, 5, 3, 4, 3, 3, 1, 1, 0, -2, -3, -3, -1, 0, 3, 3, 2, 4, 1, 0, 0, 0, 0, -3, -1, 0, -3, 0, 0, 1, 3, 2, 5, 5, 2, 4, 2, -1, 0, -3, -1, -2, -1, -1, 1, 3, 1, 3, -1, -2, 0, -2, 0, 0, -3, 0, 0, -1, -1, 1, 0, 4, 3, 5, 1, 4, 1, 1, 0, -1, -1, -2, 0, 0, 2, 1, 0, 3, 2, 2, 0, -2, 0, -4, -3, -3, -2, -3, 0, 0, 0, 3, 3, 2, 1, 4, 1, 1, -1, -3, -3, -1, 0, 0, 1, 0, 0, 0, 1, 3, 0, -1, -1, -2, -4, -1, -4, -4, -2, 0, -1, 3, 1, 1, 2, 1, 1, -1, -3, -3, -3, -3, -1, 0, 1, 2, 2, 2, 4, 3, 1, 0, 0, -2, 0, -3, -2, -4, -4, -2, 0, 2, 0, 0, 1, 0, 1, 0, -3, -5, -6, -3, -2, -2, 0, 0, 4, 0, 1, 2, -1, -1, 0, 1, -1, -3, -4, -6, -2, -1, 1, 2, 2, 2, 0, 0, 0, 1, 0, -4, -3, -4, -3, -2, 2, 4, 1, 0, 0, 0, 0, -2, 0, 0, -3, -1, -3, -6, -3, -3, 0, 5, 4, 3, 3, 0, 0, 0, -1, -4, -4, -2, -3, 0, 1, 4, 2, 3, 0, 0, 0, 0, -1, -3, -2, -3, -4, -4, -4, -1, -1, 3, 3, 3, 1, 2, 0, -2, -3, -4, -6, -6, -1, 0, 0, 4, 1, 0, 1, 2, -1, 0, 0, -1, 0, -1, -2, -2, -1, -1, 0, 0, 3, 3, 1, 4, 2, 0, -4, -5, -5, -3, -3, 0, 0, 2, 1, 1, 3, 0, 1, 0, -1, 0, 0, -2, -1, -2, -3, -1, 0, 0, 3, 4, 3, 4, 0, 0, 0, -3, -2, -1, 0, -1, 0, 3, 2, 1, 1, 2, 0, 0, -1, 0, -2, 0, -1, -3, -4, 0, 0, 1, 2, 3, 2, 2, 0, 1, 0, -2, 0, -2, -3, 1, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, -3, -3, -4, -4, -1, 0, 2, 2, 2, 3, 1, 4, 3, 0, -2, -3, -1, -2, -2, -1, 1, 4, 4, 0, 0, 1, 0, -2, 2, 0, -3, -2, -2, -1, 0, 0, 0, 2, 3, 1, 4, 4, 0, -1, -1, 0, -4, -3, -2, 1, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 3, 2, 2, 5, 3, 0, 0, -1, -3, -4, -3, 1, 1, 1, 1, 1, 1, 2, 0, 0, -2, -1, 0, -3, -5, -2, -1, -1, 0, 1, 4, 4, 1, 2, 4, 2, 0, 0, 1, -1, 0, 0, 2, 0, 1, 1, 0, 2, 1, 2, -3, -2, 0, -1, -2, -2, 1, 0, 2, 1, 3, 0, 3, 0, 1, 0, 1, -1, -1, 0, 0, 1, 2, 3, 2, 0, 1, 0, 0, 0, 0, 0, -1, -3, 0, 0, 1, 0, 1, 2, 2, 4, 4, 3, 0, 0, 0, 0, 0, 0, 3, 2, 1, 3, 3, 1, 2, -2, -1, -1, -1, 0, -1, -3, 0, -1, 0, 1, 3, 3, 4, 1, 4, 4, 3, 0, 0, 0, 2, 1, 1, 3, 4, 4, 3, 3, 0, 0, -1, -3, 0, -1, -3, -3, -3, -3, -3, -1, 2, 3, 2, 0, 1, 1, 1, 3, 3, 2, 1, 3, 3, 2, 3, 4, 2, 4, 1, 0, -2, -1, -1, 0, -2, -3, -3, 0, 0, 2, 0, 1, 1, 2, 1, 3, 2, 2, 0, 1, 3, 3, 3, 4, 2, 4, 3, 1, 3, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, 3, 5, 0, 4, 4, 2, 3, 4, 0, 2, 3, 4, 4, 4, 3, 4, 1, 4, 2, 3, 1, 2, 1, 0, 0, 3, 2, 0, 2, 4, 4, 3, 0, 1, 1, 2, 0, 0, 2, 0, 0, 0, 2, 0, 0, 2, 1, 0, 1, 2, 1, 1, 0, 0, 2, 3, 0, 2, 0, 0, -1, 0, 0, -1, -1, 0, 1, -1, 2, 0, 0, 1, -1, 0, 1, 0, 3, 3, 2, 3, 0, 1, 0, -1, 2, 1, 2, -1, 1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 1, 1, 1, 2, 3, 0, 0, 3, 0, 0, 0, 1, 0, 1, 2, 0, -1, -1, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 0, 0, 0, 1, 3, 0, 1, 1, -1, 1, 0, 1, 0, 1, 0, 0, -1, 0, 1, 1, -1, 1, 0, 2, 3, 1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 2, 0, 1, -1, 0, -2, 0, -2, 1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 1, 0, 1, 2, 0, 2, 0, 0, 0, -1, -1, 0, 0, -2, 0, 1, -1, 2, 0, -1, 2, -1, 2, 0, 2, 1, 0, 1, 2, 2, -1, 1, 1, 0, 0, 0, -1, 1, 2, 0, 0, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, -1, 2, 2, 0, 0, 0, 2, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 0, 3, 1, 1, -1, 2, -1, 0, 0, 2, -1, -1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 2, 2, -1, -1, 1, 1, -1, 2, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 1, 0, 0, 2, 1, 0, 2, 2, 0, 2, -1, 1, 0, -1, 1, 0, 2, 2, 1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 1, -2, 0, 1, 1, 1, 0, 0, 0, 0, 2, 1, 2, 0, -1, -1, 2, 0, 2, -1, 0, 2, 2, 1, 2, 0, 2, 0, 2, 0, 1, 0, 0, -1, 2, 0, 2, 0, 0, 0, 2, 2, 1, 0, 0, 2, 0, 1, 0, 2, 0, 1, 0, 0, 0, 2, 0, 1, 2, -1, 0, -1, 2, 0, 0, 0, -1, 2, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, 1, 1, 1, 2, 1, 0, 0, 0, 2, 0, 1, 0, -1, 0, -1, 2, 0, 1, 1, 1, 0, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 3, 2, 0, -1, 0, -1, 2, 1, -1, 2, 0, 0, 0, 0, 2, 0, 0, 0, 2, 2, 0, 2, -1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 1, 0, -1, 0, 0, -1, 2, 2, -1, -2, 0, -1, -1, 2, 0, 2, 2, 2, 0, 0, 0, 1, 0, 2, -1, 0, 0, 0, 0, -1, 2, -1, 2, 2, -1, 0, 0, 1, 1, -1, 0, 0, -1, 1, 1, 0, 2, 1, 2, 3, 0, 1, 2, 0, 0, 3, -1, 1, 0, -1, 2, -1, 0, 0, 0, 2, 0, 1, -1, 0, 1, 1, 0, 2, 0, 2, 3, 2, 2, 0, 2, 1, 0, 3, 2, 1, 0, -1, 0, -1, 0, 0, 1, 2, 2, 2, 0, 0, 2, 0, 0, 0, 1, -1, 0, 2, 0, 0, 0, 0, -1, 3, 0, 3, 3, 0, 1, 0, 0, 2, 0, 1, 1, -1, 0, 0, 1, 2, 2, 1, 0, 0, 0, 0, 0, 2, 0, 1, 3, 0, 1, 2, 0, 1, 2, 0, -1, 1, -1, 1, 1, 0, -1, 2, 0, 1, 2, 2, 1, 0, 0, 0, -1, 1, 2, 1, 0, 0, 0, 2, 2, 0, 0, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 2, 0, 1, 0, 2, 1, 2, 0, 3, 0, 0, 3, 1, 3, 0, 2, 1, 0, 0, -1, 2, 1, 1, 0, 2, 0, 1, 0, 0, 2, 0, 0, 1, 0, 1, 0, 0, 1, 2, 1, 0, 3, 2, 0, 2, 1, 0, 0, -2, 1, -1, 2, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 3, 0, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, -1, 1, 2, -1, -1, 1, 0, 1, 1, 0, 2, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 2, 2, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 1, 2, 0, 3, 0, 3, 1, 0, 0, 2, 1, 1, 2, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 2, 1, 2, 1, 0, 0, 1, 0, -1, 1, 0, 0, -2, 0, 0, 0, 1, 3, 0, 2, 1, 0, 0, 2, 2, 0, 1, 3, 3, 2, 1, 0, 2, 2, 3, 2, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, -1, 2, 0, 1, 0, 1, 3, 3, 3, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 2, 1, 0, 2, 0, 0, 2, 0, 1, 0, 0, 0, -1, 0, 1, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, -1, -1, 1, 3, 1, 1, 1, 3, 0, 2, 1, 0, 1, 0, 0, 2, -1, 0, 1, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, 2, 0, 0, -1, 2, 2, 0, 1, 0, 0, 2, 3, 0, 2, 0, 1, 2, 0, -1, 1, 1, 1, 0, 1, 2, 1, 2, 2, 2, 1, 0, 2, 0, 1, 2, 2, 3, 2, 1, 0, 1, 1, 0, -1, -1, 0, 1, 0, 1, -1, 1, 0, 2, 0, 2, 0, 0, 1, 0, -1, -1, 1, 0, 1, 0, 1, 0, 2, 2, 3, 0, 0, 0, 0, 0, 0, -1, 1, -2, 0, 2, 2, 1, 1, 1, 0, 1, 1, 1, 0, 0, 2, 2, 0, 3, 1, 1, 2, 2, 3, 0, 0, 3, 1, 1, 0, 0, 0, -2, 1, -1, -1, 0, 1, 2, 1, -1, 0, 0, 1, -1, 0, -1, -1, 3, 0, 0, 1, 3, 0, 1, 1, 1, -1, 1, 0, 0, -1, 0, 0, 0, 0, 2, 0, 2, 0, 3, 1, 0, 0, 0, 1, 1, 0, 0, 1, 2, 1, 0, 1, 3, 0, 0, -1, -1, -1, 0, 0, -1, 1, -1, 0, 0, 2, 2, 3, 1, 1, 0, 1, 0, 1, 1, 0, 2, 3, 2, 1, 0, 2, 1, 0, 1, -1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 3, 1, 0, 0, 2, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 1, 1, 0, 2, 0, 1, 0, 2, 1, 0, 2, 0, 1, 0, 2, 0, 0, 1, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 2, 0, 0, 2, 0, 0, 1, 0, 2, 0, 0, 0, 1, 1, -1, 1, 0, 1, 0, 1, 0, 0, 2, 0, 0, 0, 2, 0, 0, 1, 0, 2, 2, 1, 2, 0, 0, 0, 0, 0, 0, 2, 1, -1, 1, 0, 0, 0, 1, -1, 1, 0, 0, 2, 1, 2, 2, 2, 1, 2, 0, 1, 2, 0, 0, 2, 1, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 2, 0, -1, 0, 0, 2, 1, 0, 2, 0, 0, 2, 1, -1, 1, 1, 0, 0, -1, 0, -1, 0, -2, 0, 1, 1, 2, 0, 0, 1, 2, 2, 2, 0, 1, 0, 0, 0, 0, 2, 2, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, -2, 0, -2, 0, 1, 0, 2, 0, 0, 0, 2, 0, 0, 3, 3, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 1, -1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 3, 3, 1, 2, 1, 2, 0, 0, 0, 1, 1, 0, 0, -2, 0, -2, 0, 0, 0, 1, 2, 1, 2, 3, 2, 0, 2, 0, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 2, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 2, 2, 2, 2, 2, 1, 3, 0, 0, 0, 0, 3, 2, 1, 2, 0, 2, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 2, 2, 2, 3, 2, 0, 2, 0, 1, 0, -2, -1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 2, 2, 1, 0, 2, 0, 3, 0, 0, 2, 0, 2, 0, 0, 0, 1, 0, 0, 1, 1, -1, 2, 1, -1, 1, 2, 0, 0, 2, 1, 2, 2, 0, -1, 1, 2, 0, 2, 2, 2, 0, 2, 0, 1, 1, 1, -2, 0, -1, -1, 1, 0, 1, 0, 2, 1, 2, -1, 0, 0, 2, 0, -1, 1, 0, 0, 0, 0, 0, 2, 0, 1, 2, 0, -1, -2, -1, 0, 0, -1, 1, 2, -1, 1, 1, 1, 1, -1, -1, 1, 0, 1, 0, 1, 0, 2, 0, 3, 0, 0, 0, 0, 2, 2, 1, -1, -2, -2, -1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 2, 2, 2, 0, 0, 2, 0, 1, 2, 0, 1, 2, 0, 1, 0, 0, 1, 1, 0, -1, 0, 1, -1, 0, 0, 1, 0, 2, 0, 2, 2, -1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 1, 1, 0, 1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 0, 0, 3, 0, 0, 3, 1, 1, 0, 0, 1, 0, 2, 1, 0, 1, -1, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 1, -1, -2, 0, 0, 2, 2, 0, 0, 3, 0, 3, 0, 0, 1, 0, 0, 1, 3, 2, 1, 0, -2, 0, 1, 0, -2, 1, 0, 0, 0, 0, 0, 1, 2, 1, 3, 3, 2, 0, 3, 1, 1, 3, 3, 0, 2, 2, 1, 1, 2, -1, -2, 0, 1, 0, -2, -2, 0, 0, -1, -1, 0, -1, 1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, -1, 0, 1, 0, -1, 0, 0, -1, 0, 0, -2, -2, -2, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, -1, 1, -1, -2, -1, 0, -1, -3, -3, -3, -1, 0, 0, -2, 0, -1, -2, 1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, -3, -1, -1, -1, -3, -3, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -3, -3, -4, -3, -2, -4, -2, -3, -2, -1, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 2, -1, 0, -2, -1, -3, -3, -1, -1, -3, 0, -2, -1, 0, -1, 0, 0, 0, 1, 1, 2, 0, 1, 2, 1, 0, 0, -1, 0, -1, 1, 1, 0, 0, -1, -4, -4, -1, -4, -4, -4, 0, -3, 0, 0, 0, 2, 1, 0, -1, 0, 2, 1, 0, 0, 1, 0, -1, 1, -1, -1, -1, -3, -3, -3, -4, -5, -3, -4, -1, -1, -4, 0, 0, -1, 0, 0, -2, -1, 2, 1, 2, 3, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, -1, -4, -2, -3, -4, -5, -1, -5, -2, 0, 0, -1, 0, 0, 0, -1, 1, 2, 1, 1, 2, -1, 2, 1, -1, 0, -1, -1, 0, -1, -2, -2, -3, -5, -4, -4, -3, -3, -1, -1, 0, -1, -1, 0, 2, 0, 0, -1, 1, 0, 0, 2, 0, 1, 2, 1, 0, 0, -3, 0, -2, -3, -6, -1, -5, -3, -4, -2, -4, -3, 0, 0, -2, -2, -1, 0, 1, 0, 2, 2, 0, 0, -1, 0, 0, -1, 1, 1, 0, 0, -2, -3, -2, 0, -4, -2, -3, -3, -2, -1, 0, -2, -2, 0, 0, -1, 2, 0, 2, 0, 0, 2, 2, 1, 0, 0, -1, 0, 0, -3, -1, -3, -1, -3, -4, -3, -2, -3, -1, -3, 0, 0, -1, -1, 0, 0, 0, 0, 1, 3, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -2, -1, -2, -2, -2, -1, 0, 0, -3, -1, -1, 0, -1, 1, 0, -1, 0, 0, 3, 0, 1, 0, 0, 1, 1, 0, -2, -2, -1, -4, -3, -1, -6, -3, -5, -2, -3, -2, -2, 0, 0, -1, 0, 2, 1, -1, 0, 0, 0, 0, 1, -2, -1, 0, 1, 0, -1, -2, 0, -3, -5, -3, -5, -4, -4, -1, -1, 0, -3, 0, -1, 1, 0, 0, 2, 0, 0, 2, 2, 0, 0, 0, -1, 0, -1, 1, -1, 0, -1, -3, -6, -3, -1, -1, -3, 0, 0, -3, -1, -1, -1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 2, -1, 0, 0, 0, -1, -1, -2, -5, -1, -1, -2, -3, -1, 0, -1, -1, -2, -1, 0, 0, 1, 1, 0, 0, 0, 2, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -4, -5, -3, -3, -1, -1, 0, -1, -3, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, -1, 2, 0, 1, 1, 0, 1, 0, -2, 0, -2, -3, -3, -5, -4, -4, -3, -1, -3, -3, 0, -3, 0, 1, 0, -1, 1, 0, 2, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, -3, -3, -3, -4, -3, -4, -2, -1, -1, -1, -3, -3, 0, 0, 2, 1, 0, 0, 0, 0, 0, 2, 1, -1, 1, 0, -1, 1, 0, -2, -1, -2, -2, -6, -1, -2, -3, 0, -3, -2, -2, 0, -1, 0, 2, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, 1, -1, -1, 0, 0, -4, -2, -5, -5, -2, -1, -4, -1, -1, -3, -1, -2, 1, 0, 0, 1, 0, -1, 0, 0, 2, -1, 0, -2, 0, 0, 1, 0, -1, -2, -2, -4, -3, -3, -2, -2, -4, -2, -3, -1, -3, 0, 0, -2, -1, 2, 0, -1, -1, 0, 2, 1, 0, 0, -2, 1, -1, 0, -1, -2, -3, -1, -2, -5, -2, -4, -5, -5, -3, -4, -3, -2, -2, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -4, -2, -4, -5, -5, -4, -4, -1, -2, -2, 0, -2, 0, -2, 1, 1, 2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, -4, -3, -3, -5, -5, -1, -3, -4, -1, -1, -2, 0, -3, 1, 0, 1, 1, -1, -1, -1, -1, 0, 2, -1, 0, 1, 1, 0, 0, -3, -4, -1, -4, -3, -2, -1, -4, -1, 0, -2, -2, 0, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, -2, -2, -2, -4, -5, -4, -2, -2, -2, -1, 0, 1, -1, -1, 0, 1, 1, -1, -1, 0, -1, -2, 0, -2, 0, 0, -1, 0, 0, -3, -1, -2, -3, -2, -3, -3, 0, 0, 0, 0, 1, 3, 0, 3, 0, 3, 2, 0, 0, 0, -2, -1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -2, 0, -1, 0, 0, 1, 3, 1, 3, 2, 2, 2, 1, 1, 4, 4, 4, 7, 8, 6, 7, 7, 5, 4, 6, 7, 8, 6, 5, 7, 7, 4, 5, 6, 6, 6, 8, 8, 6, 4, 4, 7, 6, 4, 5, 9, 8, 6, 8, 9, 5, 7, 4, 7, 5, 6, 3, 1, 4, 1, 1, 3, 1, 1, 2, 3, 4, 1, 3, 6, 6, 5, 3, 6, 7, 6, 9, 9, 10, 8, 9, 7, 5, 3, 5, 4, 2, 1, 2, 0, 0, 0, 0, -1, -3, -1, -2, 0, -1, 0, 0, 5, 3, 3, 8, 8, 9, 9, 8, 6, 6, 4, 5, 4, 3, 0, 2, -1, 0, -1, 0, 0, -2, -4, -3, -4, -3, -1, -1, -3, 0, 1, 4, 5, 9, 6, 8, 6, 5, 8, 6, 3, 1, 0, 2, 0, 0, -1, -1, 1, -3, -4, -5, -2, -4, -6, -5, -4, -1, -2, -2, 0, 2, 0, 6, 5, 8, 4, 4, 3, 2, 0, 0, 0, 0, -3, -3, -3, 0, 0, -3, -1, -1, -2, -2, -5, -1, 0, -3, -3, 0, 0, 0, 1, 10, 6, 5, 3, 4, 4, 1, 3, 0, -3, -4, -4, 0, -1, -2, 0, -2, -2, -3, -4, -1, -3, -3, 0, -3, -1, 0, -1, 1, 2, 8, 10, 5, 5, 6, 5, 3, 0, 0, -6, -5, -5, -1, 0, 0, 0, -1, 0, 0, -2, 0, -3, -1, -2, 0, -2, -1, 0, 0, 0, 8, 9, 8, 7, 4, 4, 2, 0, -6, -7, -5, -9, -4, -5, -2, -4, -4, -4, 0, -2, -1, -1, -2, -1, 0, -1, -4, -2, 0, 0, 10, 10, 9, 7, 3, 0, -1, -4, -6, -8, -8, -11, -6, -7, -5, -5, -2, -1, 0, 0, -2, -1, -4, -2, -5, -2, -1, -1, -1, 0, 10, 8, 9, 5, 5, 0, -2, -3, -8, -10, -12, -13, -8, -5, -4, -3, 0, -1, -1, 1, 0, -2, 0, -2, -3, -4, -5, -4, 0, 0, 9, 10, 6, 6, 3, 1, -1, -8, -11, -11, -14, -14, -11, -8, -5, -2, -3, 0, -1, -2, -1, -2, -5, -3, -4, -6, -5, -4, -1, 0, 11, 6, 7, 4, 2, 2, -4, -7, -10, -12, -14, -14, -12, -10, -6, -7, -3, 1, 1, -1, 0, 0, -3, -5, -6, -6, -7, -4, -3, 2, 7, 7, 6, 4, 2, 0, -4, -11, -13, -15, -13, -16, -14, -7, -5, -6, -3, -3, -1, 0, -1, -1, -3, -2, -6, -7, -6, -3, -3, -2, 8, 8, 8, 6, 0, -3, -4, -10, -13, -16, -15, -14, -11, -7, -5, -3, -1, -1, -1, 0, -2, 0, -3, -2, -7, -7, -8, -4, -1, 0, 9, 7, 7, 5, 2, 0, -6, -9, -16, -14, -17, -16, -12, -7, -7, -5, -2, 0, 0, -1, 0, 0, -2, -4, -7, -7, -5, -4, -4, -1, 7, 8, 7, 5, 3, -1, -4, -10, -13, -17, -15, -17, -11, -7, -6, -3, -2, 0, 0, 1, 1, -2, -1, -2, -5, -6, -4, -6, -5, -3, 9, 7, 7, 7, 1, -2, -5, -9, -14, -16, -16, -13, -12, -7, -7, -4, -4, 0, -1, 2, 0, 0, 0, -5, -6, -7, -6, -4, -4, 0, 10, 8, 6, 5, 1, -1, -4, -10, -9, -11, -16, -14, -13, -8, -7, -5, -4, 0, 0, 1, 2, 0, 0, -5, -4, -7, -5, -4, -1, 0, 9, 10, 6, 8, 5, 2, -1, -4, -9, -10, -11, -13, -8, -6, -4, -3, -3, -2, 0, 0, 0, 0, -3, -2, -4, -6, -4, -2, -2, 0, 10, 10, 8, 6, 6, 1, -2, -6, -7, -11, -10, -11, -11, -7, -4, -1, 0, 0, 0, -1, 0, -2, -5, -2, -3, -2, -2, -1, 0, 0, 7, 9, 6, 6, 5, 2, -2, -2, -5, -10, -7, -9, -8, -3, -1, -3, -2, 0, 0, -3, -3, -1, -2, -3, -6, -4, -2, -2, -2, 0, 9, 6, 6, 9, 6, 1, 2, -1, -3, -4, -5, -8, -5, -5, -3, -3, 0, -2, -2, -3, -3, -1, -4, -3, -3, -3, -2, -3, -1, 1, 8, 9, 9, 6, 5, 4, 2, -1, 0, -3, -4, -5, -6, -5, -1, -1, -3, -3, -1, -3, -1, -5, -3, -2, -2, -2, 0, -2, -1, 0, 8, 8, 6, 7, 5, 4, 2, 0, 2, 0, -2, -4, -2, -2, -1, -3, -5, -5, -5, -3, -4, -5, -4, -3, -3, -1, 0, -1, 2, 1, 7, 7, 5, 5, 5, 4, 3, 3, 1, 0, 1, -2, 0, 1, 0, -2, -7, -5, -8, -3, -5, -2, -5, -4, -1, -2, 0, 1, 0, 2, 6, 8, 6, 7, 5, 4, 1, 2, 2, 1, 1, 0, 0, 0, -2, -1, -7, -8, -7, -5, -6, -3, -6, -5, -3, -4, -3, -1, 1, 3, 7, 8, 8, 4, 7, 6, 7, 6, 4, 2, 4, 3, 3, 3, 0, -3, -6, -6, -5, -6, -5, -4, -2, -5, -2, -1, -2, 0, 1, 5, 5, 5, 7, 8, 7, 7, 7, 7, 7, 4, 6, 4, 6, 5, 2, 1, -2, -2, -5, -2, -3, -4, -3, -4, 0, 0, 0, 2, 4, 5, 5, 6, 5, 5, 9, 8, 7, 7, 10, 10, 6, 8, 5, 8, 4, 4, 3, 0, 1, -1, 0, 1, 0, 0, 1, 0, 1, 1, 4, 1, 1, 0, -1, 1, 2, 0, 0, 0, 0, 0, -1, 2, 0, 2, 2, 0, 0, 1, 2, 0, 0, -1, 1, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 1, 1, -1, -1, 1, 0, 0, 0, -2, 0, 1, 0, -1, 0, 0, 0, 1, -1, 1, 2, -1, 1, 1, 0, 0, 0, 1, 2, -1, 0, 2, -1, 0, -2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 2, 0, 0, 0, -1, 0, 0, -1, 1, 0, 2, 0, 1, 1, -1, -2, 0, -2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, 0, -1, -1, 1, 2, 1, -2, -2, 1, 1, 1, 0, 0, 1, -1, 0, 0, 1, -1, -1, 0, -1, 1, 1, 1, -1, 0, 0, 0, 1, 0, 2, 0, 1, 0, -1, 0, 1, 2, -1, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 2, 0, 2, -1, 1, 1, 0, 0, 1, 1, 0, 0, 2, 0, -1, -2, -1, -1, -1, -1, 1, -1, 0, 1, -1, 1, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, -1, 0, -1, 1, -1, 0, -1, 0, -1, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, -2, 1, -1, 0, 1, 1, -1, 2, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 1, 0, 0, 1, -1, -1, 1, 1, 0, 0, 1, 0, -1, 1, 1, -1, 1, 1, -1, 0, 1, -1, -1, 1, 1, 0, 0, -1, -1, -1, 1, 0, 0, -2, 0, 2, -1, -1, -1, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, -2, -1, 1, 0, 0, -1, -1, -1, 1, -1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 1, 1, 1, 0, -1, -1, 1, 0, 0, 2, -1, 1, -2, -1, 0, 1, 0, -1, 1, -1, 0, 0, -1, -1, 1, -1, 0, -1, 0, 0, 0, 2, -1, 2, 0, 2, 0, 2, 1, 1, 0, -1, 1, 1, 1, 0, 0, 1, -1, 1, 0, 1, 1, -1, 0, 0, 0, 2, 1, -1, 1, 2, -1, -1, -1, 1, -1, 1, 1, 1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, 1, 2, 1, -1, -1, 1, 2, 0, -1, -1, 0, 2, 1, 1, 1, 1, 1, 2, -2, 1, -1, 1, -1, -1, 2, -1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, -1, 0, 1, 2, 2, 0, 0, 0, 1, 2, -1, 2, 0, 0, 1, 0, -2, -1, 0, -1, 0, 0, -1, -1, 0, 0, 1, -1, 0, 0, 2, 1, -1, 0, 1, 0, 1, -1, -1, -1, 0, 0, 1, 2, 0, -1, 0, 0, -1, -1, 0, 2, 0, 0, 2, 0, 0, 0, -1, 0, 2, -1, 1, 0, 0, 2, 0, 2, 1, -1, -1, 1, 0, 0, -2, -1, 0, -2, 1, -1, 1, 0, -1, 1, 2, -1, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 1, -1, 0, 1, 0, 0, -2, 0, 0, -1, 0, 0, 1, -1, 0, -1, -1, 1, 2, 0, -1, -1, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, -1, 1, -1, -1, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, -2, 1, 0, 1, -1, 1, 1, 1, -1, 0, -1, -1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, -2, 1, 0, 1, 0, 0, -1, 0, 1, 2, 0, -1, -1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 0, 2, 2, -1, -1, 0, 0, -2, 1, 1, 1, 1, 0, -1, 1, 1, 0, -1, 2, 1, -1, 0, 0, 2, 0, 1, 1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 1, 2, 0, -1, 0, 0, -1, 0, 0, -1, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, -1, 1, -1, 0, 0, -1, -1, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 1, -1, 0, -1, 1, 1, -1, -1, 0, 2, 0, 0, 1, 0, 0, -1, 0, 1, -1, 0, 1, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 2, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, -1, 1, -1, -1, 2, 0, -1, 0, -1, -1, 0, -1, 0, -1, -1, 1, -1, 0, 0, 0, -1, -1, -1, 1, 1, 0, -1, -1, 0, 1, -1, 0, 1, 1, -1, 0, 1, -1, 1, 1, 0, -1, 1, 0, -1, 0, -1, -1, 0, 0, 1, 0, -1, -2, -2, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, -2, 0, 1, 0, -1, 1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, -2, 0, 0, 0, -1, 1, 0, 0, -2, 0, 0, -1, 0, 1, 0, 1, 0, 1, -1, 2, 1, 0, 0, 1, -1, 2, 0, 0, 1, 1, -2, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, -2, -1, -1, 1, 1, 0, 1, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, -1, -2, 0, 0, 0, -1, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, 0, 0, 1, 0, 2, -1, 1, 0, -1, -2, 0, 0, 0, 1, 2, 2, 0, 0, 1, 1, 1, 2, 0, 0, -1, -1, 0, 1, -1, 0, -2, 0, -1, 0, -2, 0, 0, 1, 0, 0, -1, 0, -1, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, -2, -1, 1, 0, 0, 1, 1, 0, 0, 0, -2, -1, -1, 0, -1, 0, -1, -1, 0, -1, 1, 2, -1, 1, 0, 1, 0, -1, 0, 0, -2, -1, 0, 0, 0, 1, 0, -2, 1, 0, -1, 1, -2, -1, -1, -1, -1, -1, 0, -1, 0, -1, 1, 0, 1, 1, 1, 1, 1, 1, 0, -1, 0, 0, 0, -1, -1, 0, 2, -1, 0, 0, 0, 0, 1, 1, 1, -1, 1, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 2, 1, 0, 0, -1, 0, 0, 0, 0, -1, -2, 1, 1, 2, -1, 2, 1, -1, 2, 1, 0, 0, 0, 1, 2, -1, 0, 0, 1, 0, 1, 0, -1, -1, -1, 1, 0, 0, 0, -1, -1, 0, 1, 1, -1, 0, 0, 1, 1, -1, -1, 1, 2, 1, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, -1, 1, -1, 1, 0, -1, 2, -1, -2, 0, -1, -1, 1, 0, 0, 1, 0, -1, 1, 1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, 1, 0, -1, 0, 0, 0, -1, 1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, -1, 0, 1, 0, -1, 0, 1, 0, 1, 2, -1, 1, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -2, 0, 1, 0, -1, 0, 0, 0, 1, -1, 0, 1, 1, -1, -2, 0, 2, 0, 0, 0, -1, 0, -1, 1, 0, 2, 0, 2, 1, 1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, -2, 1, -2, -1, -1, -2, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, -1, -1, 1, -1, -1, 1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, -1, 0, 1, -1, -2, 1, 0, 1, -1, 2, -2, 0, 0, 0, 1, 1, 0, 0, -1, -1, 1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, -1, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, -1, 1, -1, 1, 0, 0, -1, 1, 1, 1, 0, 1, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 1, -2, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 1, 1, 0, 0, 2, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, -1, 1, -1, 0, 0, 0, 2, 1, 0, 0, 0, 1, -2, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 0, -1, 1, 1, -1, 1, -2, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 1, 0, 1, 1, 2, -1, 0, 1, -1, 0, -1, 0, 1, 1, -1, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 1, -1, 0, -1, 1, 0, 0, -1, 0, 0, 1, 0, 2, -1, 1, 0, 0, 1, 0, 1, 0, 0, 2, -1, 0, 0, 1, 0, -1, -1, 0, -1, -1, 0, 0, -1, 1, 1, 0, 0, -1, 0, 2, 0, 1, -1, 1, 0, 0, 0, 0, 0, -2, 0, -1, -1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, -2, 0, 1, -1, 0, 1, 0, 2, 0, -1, 0, 1, -1, 0, 2, -1, -2, -3, -4, -2, -4, -4, -1, -1, -1, -1, 0, 0, -2, 0, -1, 0, 3, 2, 4, 6, 7, 9, 9, 10, 12, 10, 10, 9, 9, 9, 0, -1, -2, -3, 0, 0, 0, 0, 2, 2, 3, 2, -1, -1, -2, -2, 0, 0, 0, 2, 0, 0, 4, 4, 4, 4, 7, 6, 9, 9, -3, -1, -2, -1, 0, 0, 1, 0, 1, 0, 0, 0, -1, -3, -3, -3, -2, 0, -1, -1, -4, -5, -3, -2, -3, -2, 1, 4, 5, 4, 0, -2, -2, -1, 0, 0, 3, 1, 1, 0, -2, 0, -2, -1, -1, 0, -3, -5, -3, -7, -7, -8, -6, -7, -5, -4, 0, 0, 3, 4, -2, -3, -4, -3, 0, 1, -2, -3, -3, -2, 0, 0, 0, 2, 2, 0, -3, -3, -7, -7, -4, -4, -4, -6, -4, -5, -4, 1, 3, 5, -2, 0, -3, -2, 0, 0, -3, -3, -3, -1, 0, 2, 4, 3, 3, 0, 0, -5, -6, -7, -6, -2, -3, -4, -3, -4, -1, 3, 5, 6, 0, 0, 0, -1, -2, 0, -2, -4, -5, -2, -1, 1, 4, 3, 3, 1, -2, -5, -4, -7, -5, -3, -5, -1, -5, -1, 0, 0, 2, 3, 0, 1, 2, 0, 1, 0, -2, -3, -4, -6, -3, 0, 6, 4, 5, 4, 0, -2, -7, -6, -6, -4, -4, -5, -5, -4, -3, 0, 1, 3, 2, 2, 1, 1, 1, 0, -1, -4, -6, -4, -1, 0, 2, 6, 4, 2, -3, -6, -5, -8, -6, -5, -5, -5, -4, -3, -3, 0, 1, 2, 1, 2, 4, 3, 0, -2, 0, -3, -7, -5, -1, 0, 0, 4, 3, 0, -3, -6, -5, -6, -7, -8, -7, -6, -5, -5, -3, -1, -1, 1, 4, 4, 4, 3, 0, 0, 0, -5, -5, -2, -4, 1, 1, 3, 4, 0, 0, -3, -2, -3, -4, -4, -6, -5, -5, -6, -4, -2, 0, 4, 1, 3, 2, 0, 0, 0, 0, -3, -5, -3, -4, 0, 2, 4, 5, 1, 0, 0, -2, -4, -3, -5, -5, -4, -6, -6, -5, -3, -2, 0, 2, 1, -1, 0, -2, 0, -1, -4, -6, -3, -1, 2, 1, 6, 7, 3, 2, -1, -3, -2, -5, -6, -3, -4, -8, -8, -7, -7, -2, 0, 1, 0, 0, -1, 0, -1, -4, -3, -5, -2, -2, 1, 5, 9, 6, 5, 3, -1, -3, -6, -5, -3, -2, -6, -6, -8, -7, -4, -4, 0, 1, 0, 0, 1, 0, -2, -2, -5, -7, -5, -1, 1, 5, 7, 9, 3, -1, -4, -6, -5, -8, -7, -2, -2, -6, -7, -5, -4, 0, 0, -1, -1, -1, 0, -1, -1, -2, -4, -7, -5, -3, 2, 6, 8, 7, 2, 0, -3, -7, -7, -5, -4, -4, -6, -5, -9, -6, -6, -2, 1, 0, 0, 0, 0, -1, 0, -5, -8, -7, -3, -3, 3, 3, 4, 6, 1, -1, -3, -4, -4, -5, -4, -2, -2, -7, -4, -5, -5, 0, 0, -1, 1, 0, 0, 1, -1, -2, -5, -4, -2, -3, 2, 3, 7, 6, 3, 0, -3, -3, -4, -2, -4, -3, -6, -3, -7, -4, -4, 0, 2, 0, 0, 1, 2, 1, -2, -2, -4, -2, -4, 0, 2, 4, 4, 7, 2, 0, -2, -2, -5, -1, -3, -2, -4, -6, -5, -5, -2, 0, 2, 1, -2, 3, 1, 0, -1, -2, -3, -2, -3, 0, 0, 4, 6, 6, 2, -1, -4, -5, -5, -3, -2, -6, -6, -8, -6, -5, -2, 3, 4, 0, 2, 1, 4, 1, 0, -4, -5, -4, -4, -4, 2, 0, 4, 3, 1, 0, -3, -3, -4, -5, -5, -6, -6, -6, -7, -1, -2, 1, 4, 2, 0, 0, 0, 1, 0, -2, -3, -6, -7, -1, 0, 2, 0, 2, -1, -1, -1, -2, -2, -4, -6, -6, -8, -4, -6, -3, 1, 2, 7, 1, 0, 1, 3, 1, -1, -2, -6, -5, -3, -2, 0, 1, 1, 1, -1, -3, -4, -4, -5, -5, -6, -6, -5, -4, -4, -2, 3, 3, 7, 0, 1, 0, 0, 0, -1, -2, -5, -2, -2, 0, 0, 2, 0, 0, -1, -2, -5, -6, -6, -7, -7, -8, -6, -3, -4, 0, 3, 4, 7, -1, 1, 1, 0, -1, -2, -2, -3, -3, 0, 0, 4, 4, 0, 0, 0, -4, -6, -7, -10, -8, -6, -5, -4, -6, -4, 0, 1, 4, 5, -1, 0, -1, 0, -3, -1, -5, -4, -1, 1, 3, 5, 4, 3, 2, 0, -4, -7, -9, -7, -7, -7, -6, -8, -6, -4, -1, 0, 5, 7, 0, 1, 1, -1, 0, -1, -3, -1, 0, 2, 3, 2, 0, 0, 0, 0, -4, -8, -9, -8, -7, -8, -8, -8, -7, -5, -3, 0, 7, 8, -2, 0, 0, -1, 0, 0, -2, 2, 1, 3, 3, 0, 0, 1, -1, -1, -4, -6, -7, -9, -6, -5, -6, -7, -4, -3, -2, 1, 7, 8, -2, 0, 0, 0, 1, -1, -1, 1, 2, 0, 0, 2, 0, -2, 0, -3, -2, -4, -7, -3, 0, 0, -1, -2, 0, 1, 5, 7, 8, 10, -1, 0, -1, -4, -2, -4, -2, 0, -1, -1, 0, -3, -1, -4, -4, -3, 0, 0, -2, 1, 4, 5, 2, 4, 6, 6, 9, 11, 11, 10, 0, -1, -2, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 1, 3, 1, 1, 3, 3, 0, 2, 3, 4, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 2, 1, -1, -1, 0, 0, 0, 2, 1, 0, 0, 0, 2, 3, 2, 1, 3, 1, 1, 1, -2, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 0, 2, 3, 3, 0, 0, 0, -2, 0, 2, 0, 0, 0, 0, 0, 2, 1, 2, 1, 1, 1, 0, 0, -1, 1, -1, 1, -2, 0, 0, 0, 1, 2, 2, -1, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, 2, 1, 2, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, -2, 0, 0, 2, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 2, 2, 0, 1, 3, 2, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 3, 1, 0, -1, 1, -2, 1, -1, -2, 0, -1, -1, 0, 3, 3, 4, 3, 1, 2, 1, 0, -1, -2, 0, 1, 0, 1, 0, -2, 1, 0, 2, 0, 0, 0, 2, 0, 0, 0, -2, 1, 0, 0, 0, 1, 3, 3, 1, 1, 1, 0, 1, 0, -2, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, 0, -1, 0, 0, 2, 1, 3, 3, 2, 3, 1, 3, -1, 0, 1, -1, 1, -2, -1, 0, 0, -1, 0, 1, 0, 0, 1, 2, 1, -1, 0, 0, 0, -2, 1, 2, 0, 4, 4, 4, 0, 0, 0, 0, 1, 0, 1, 0, -3, -1, 0, 1, -2, 0, 2, 0, 0, 0, -1, 1, -1, 0, 0, -1, 2, 0, 3, 3, 5, 3, 3, 0, 0, 2, 0, 0, 0, 1, -1, -1, -1, -1, 0, 0, 0, -1, 1, 1, 2, 1, 1, 0, 0, 1, -1, 2, 1, 3, 5, 2, 3, 0, 3, 0, 2, 0, -2, -2, 0, 0, 0, 0, -2, 0, 0, 1, 0, 2, 2, -1, 2, 2, 1, 0, 1, 1, 0, 2, 3, 1, 4, 2, 0, 2, 2, 1, 1, -2, -1, -3, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 0, 4, 2, 4, 3, 5, 2, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, -3, -1, 1, 1, 0, 0, 0, -1, 1, 0, 2, 0, 0, 0, 1, 3, 4, 5, 2, 1, 0, 1, 0, -1, 1, -2, -2, 0, -2, -3, 0, -1, 2, -1, 0, 0, 1, 2, 0, 0, 1, 0, 1, 2, 1, 2, 3, 5, 1, 1, 2, 0, 0, -1, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 2, 1, 0, 2, 2, 3, 5, 3, 4, 4, 0, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -1, -1, 2, 2, 1, 1, 0, 2, 1, 0, 3, 1, 4, 1, 1, 0, 0, 2, 1, 0, 1, 0, 0, -2, 0, 0, 0, 2, -1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 3, 3, 4, 4, 4, 3, 2, -1, 1, -1, 0, 2, 0, -1, -1, -2, -1, 0, 2, -1, 0, -1, 1, 2, 1, -1, 0, 1, 1, 2, 1, 1, 3, 1, 3, 1, 1, 0, 0, 1, -1, 0, 0, 0, -2, -1, 0, 2, 0, -2, 0, -1, 0, 1, 1, 1, 1, 1, 1, 2, 1, 3, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -1, -2, 1, 0, 0, 2, -1, 0, 0, 0, 0, 0, -2, 1, -2, 0, 0, 2, 4, 0, 1, 0, 0, 0, 0, 1, 0, -2, 0, -2, -2, -1, 0, 2, 2, 2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, -2, 1, -2, 0, 2, 0, 0, 0, 0, 0, 1, -1, -2, 0, 0, 1, 0, 3, 3, 3, 0, 2, 0, 1, -2, -2, 1, 0, 0, -2, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -2, -1, 0, 0, 0, 3, 1, 1, 3, 2, 0, -1, -2, -2, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, -2, 0, 0, 0, 0, 0, 0, -2, 2, 2, 0, 1, 1, 3, 1, 1, -1, 0, -1, 0, 0, -1, 0, -1, 1, -1, 0, 0, 1, -1, 0, 0, -2, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 0, 2, 1, -1, -2, -3, -1, 0, 0, -2, 0, -1, -1, 0, 2, 2, 1, -2, -1, -1, -2, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, -2, -1, 0, -2, -1, 0, -2, -1, -1, -1, 0, 1, 1, 0, 0, -2, -2, 0, 0, -2, 0, -1, -1, -1, 0, 1, -1, 1, 0, 1, -1, -1, -2, 0, 1, 1, -1, 0, 2, 2, 0, 4, 3, 0, -2, 0, 0, 0, 0, -2, 0, 1, -1, -2, 0, -2, -1, -2, -1, 0, 0, -1, 0, 0, 1, 1, 2, 3, 1, 0, 1, 3, 3, -2, -4, -3, -4, -4, 0, 0, 2, 1, 4, 4, 0, -2, -3, -3, 0, -1, 2, 6, 3, 5, 4, 5, 5, 10, 11, 12, 12, 16, 12, -1, -1, 0, -1, -1, 3, 3, 3, 4, 5, 2, 1, 0, -1, 0, 0, 2, 0, 3, 0, -2, -1, -1, 0, -1, 0, 5, 8, 10, 12, -1, 0, -1, -3, 0, 3, 0, 0, 1, 0, 0, 2, 1, 1, 2, 2, 3, 0, -1, -3, -5, -6, -4, -5, -4, -3, 1, 2, 5, 8, 0, -1, -3, -3, -2, 1, 0, -2, -3, -2, 2, 1, 1, 3, 7, 4, 1, 0, -3, -4, -2, -6, -6, -3, -4, -3, -1, 1, 4, 9, -2, -1, -2, -2, -1, 0, -4, -2, -4, 0, 1, 6, 8, 11, 9, 9, 2, 0, -2, -1, -3, -2, -3, -2, -2, -5, -1, 4, 5, 9, 0, 2, 1, 0, -1, -2, -2, -4, -4, -5, -1, 4, 11, 12, 11, 11, 8, 3, -1, -1, -3, -2, -5, -4, -4, -3, -2, 3, 6, 8, 2, 2, 0, 0, 1, -2, -6, -6, -8, -6, 1, 3, 11, 12, 17, 13, 8, 2, 0, -2, -1, 0, -3, -6, -3, -5, -2, -1, 4, 6, 1, 5, 4, 5, 2, -1, -3, -7, -8, -4, 0, 4, 8, 13, 13, 12, 6, 4, 0, -6, -5, -3, -5, -6, -6, -4, -4, -2, 3, 6, 2, 6, 7, 4, 0, 0, -3, -8, -8, -5, -1, 3, 9, 12, 14, 13, 9, 3, 0, -4, -4, -4, -5, -6, -4, -6, -5, -3, 0, 2, 3, 3, 3, 2, 2, -1, -2, -3, -8, -3, -3, 3, 10, 11, 15, 13, 7, 6, 2, -2, -1, -2, -3, -4, -4, -4, -6, -5, 0, 5, 0, 2, 2, 3, 2, -1, -3, -3, -7, -4, -1, 4, 10, 13, 15, 12, 11, 7, 4, 0, -3, -3, -4, -7, -8, -8, -10, -7, -3, 1, 3, 3, 0, 0, -1, -1, -1, -5, -4, -4, 0, 5, 12, 15, 14, 14, 13, 7, 6, 2, 0, -1, 0, -3, -8, -8, -9, -6, -4, 3, 0, 1, 0, -1, -3, -3, -3, -4, -4, -2, -2, 5, 10, 15, 19, 17, 11, 9, 3, 0, -4, -1, -3, -6, -8, -7, -8, -5, -1, 1, 1, 0, -2, 0, -2, 0, -4, -4, -5, -3, -2, 4, 13, 17, 18, 17, 9, 6, 1, -2, -5, -5, -3, -4, -7, -10, -9, -8, -4, 0, -3, 0, -1, 0, -2, -1, -6, -8, -9, -5, -1, 5, 12, 17, 18, 16, 7, 2, 0, -2, -5, -3, -2, -4, -7, -10, -9, -6, -2, 0, -1, 0, 0, 0, 0, -1, -4, -7, -8, -5, 0, 6, 10, 14, 15, 13, 8, 4, 2, 0, 0, -3, 0, -5, -7, -6, -7, -5, -2, 2, -4, 0, 0, 3, 0, -3, -3, -8, -6, -4, 1, 6, 11, 15, 15, 13, 8, 7, 5, 0, 0, 1, 0, -2, -5, -7, -8, -4, 0, 2, 0, 1, -1, 0, 0, -1, -6, -6, -5, -3, 1, 6, 11, 16, 15, 15, 11, 7, 2, 0, 0, -1, -2, -3, -4, -6, -8, -6, 1, 4, -2, -1, 1, 0, 0, 0, -4, -4, -5, -3, 3, 7, 9, 13, 17, 12, 7, 6, 1, 0, 0, -1, -2, -5, -8, -5, -4, -4, 0, 6, 0, 0, 2, 4, 1, -1, -2, -4, -6, -5, 1, 5, 8, 13, 13, 12, 7, 5, 0, 1, -2, -3, -6, -8, -7, -7, -6, -2, 3, 6, -1, 2, 2, 0, 1, -1, -5, -6, -9, -5, -3, 5, 8, 10, 11, 9, 8, 2, 0, 0, -2, -6, -6, -7, -9, -7, -4, -1, 5, 5, 0, 0, 2, 3, 2, -2, -4, -6, -5, -3, 0, 5, 6, 11, 6, 5, 7, 5, 2, 0, -3, -6, -6, -5, -7, -5, -3, 3, 5, 10, 0, 1, 1, 0, 2, -1, -3, -5, -3, -2, 0, 3, 9, 9, 9, 4, 4, 0, 0, -3, -4, -8, -6, -6, -5, -2, 1, 4, 6, 11, 1, 3, 1, -1, -1, -3, -4, -6, -2, -2, 5, 8, 8, 8, 7, 6, 3, 0, -4, -5, -6, -6, -6, -6, -4, -1, 0, 2, 7, 11, 0, 2, 0, 0, 0, -3, -4, -2, -2, 2, 5, 8, 13, 11, 7, 5, 4, -2, -6, -6, -7, -9, -5, -8, -6, -4, -3, 1, 6, 10, 2, 1, 2, 0, 0, -1, -3, 0, 1, 1, 5, 10, 9, 7, 8, 6, 1, -3, -4, -6, -7, -6, -7, -9, -8, -6, -1, 3, 6, 9, 0, 3, 1, 1, 3, 0, 1, 3, 3, 4, 5, 5, 8, 6, 8, 5, 3, 0, -3, -8, -7, -6, -7, -8, -9, -4, -4, 2, 8, 8, 0, -1, 2, 1, 0, 0, 1, 0, 5, 4, 4, 5, 2, 4, 4, 4, 0, -2, -1, -4, -3, -4, -1, -3, 0, 0, 4, 6, 8, 14, 0, 0, -1, 0, 0, 0, 0, 2, 1, 2, 3, 1, 0, 0, 0, 3, 1, 1, 1, 2, 3, 5, 7, 4, 6, 7, 10, 14, 16, 12, 0, -1, -4, -2, -4, -4, -3, -2, -1, 0, 0, -2, -1, 0, -1, 3, 4, 4, 8, 10, 16, 15, 13, 17, 17, 18, 16, 18, 15, 17, -1, -4, -3, -3, -2, -2, -2, -3, 0, 0, -2, 0, -1, 2, 3, 3, 4, 4, 5, 6, 9, 6, 11, 9, 7, 5, 4, 3, 3, 1, -1, 0, 0, 0, -2, 1, -1, 1, 1, 1, 0, 1, 0, -1, 2, 2, 1, 3, 4, 3, 3, 4, 6, 6, 8, 7, 7, 5, 5, 2, -1, -2, -2, -2, 0, 1, 0, 0, 3, 1, 3, 1, 1, 0, 2, 3, 5, 3, 3, 3, 2, 2, 3, 1, 4, 3, 3, 6, 5, 2, -2, 0, -1, -1, 1, 0, 0, 0, 2, 1, 0, 3, 0, 3, 3, 0, 1, 1, 4, 0, 2, 0, 1, 0, 0, 3, 1, 4, 1, 1, 0, 0, -1, 0, -1, 0, 0, 1, 2, 0, 2, 3, 3, 2, 3, 0, 0, 2, 1, 0, 1, 0, 0, -1, 1, 0, 3, 1, 3, 3, 0, -1, 0, -2, -2, 0, 0, 1, 2, 1, 3, 4, 4, 1, 4, 0, 1, 2, 3, 2, 0, 1, -1, 2, -1, -1, 2, 2, 2, 5, -1, 0, 0, -1, -2, 0, 0, 0, 3, 3, 4, 5, 7, 4, 2, 2, 0, 2, 1, 2, 2, 1, 0, 0, 2, 2, 3, 3, 2, 1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 5, 3, 6, 8, 5, 3, 3, 0, 3, 2, 2, 2, 1, 3, 1, 2, 3, 4, 3, 1, 0, 1, -1, -2, 0, -2, -2, 0, 2, 1, 3, 7, 5, 7, 7, 1, 0, 0, 0, 0, 0, 3, 1, 0, 2, 1, 1, 4, 3, 2, 0, 1, 2, -1, -2, -1, -3, -2, 0, 3, 4, 5, 5, 9, 3, 1, 3, 0, -2, -1, -1, 0, 0, 0, 0, 1, -1, 2, 5, 5, 0, 0, 3, 2, 1, 0, 0, 0, 0, 1, 5, 5, 7, 6, 4, 3, 4, 1, 0, 0, -1, 0, 0, 1, 3, 0, 2, 1, 4, 2, 0, 0, 0, 0, 1, 1, 0, 2, 3, 4, 3, 7, 7, 4, 7, 4, 4, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 3, 5, 0, -2, 0, -2, -1, -1, 1, 0, 1, 4, 3, 3, 7, 6, 6, 5, 5, 3, 0, 0, 2, 1, 0, -1, -1, 0, 0, 2, 1, 4, 1, 0, 1, -1, -1, 0, 1, 0, 1, 6, 7, 7, 9, 8, 6, 3, 2, 3, 2, 2, 2, 1, 2, 0, 1, -1, 0, 3, 3, 2, 0, 1, 0, 0, -1, -1, 0, 0, 1, 5, 8, 7, 9, 9, 5, 2, 3, 3, 2, 0, -1, -1, 1, 0, -1, 0, 1, 0, 0, 4, -1, 0, 0, -2, 1, -1, 0, 0, 4, 6, 5, 8, 8, 9, 7, 3, 3, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 2, 0, 2, 2, -1, -1, 0, 0, 1, 3, 4, 7, 7, 7, 9, 8, 3, 0, 1, 1, 0, -1, 1, 2, -1, 1, -2, 0, 1, 1, 4, 0, 1, 2, 0, 0, -1, 0, 0, 3, 4, 7, 8, 7, 7, 7, 5, 3, 3, 0, 0, 2, 2, 0, 0, -1, 0, -1, 1, 3, 3, -2, 0, 2, 0, -2, -2, -1, 2, 4, 3, 3, 7, 9, 7, 8, 4, 4, 3, 4, 2, 4, 3, 0, -1, 1, 0, 1, 2, 3, 2, 1, 0, 1, 0, 0, 0, 0, -1, 0, 5, 5, 6, 8, 9, 8, 4, 3, 1, 0, 3, 4, 2, 0, 1, 1, -1, 1, 1, 1, 4, 0, -1, 0, -1, 0, 0, 0, 0, 3, 2, 4, 8, 9, 7, 5, 3, 1, 1, 0, 1, 2, 0, 0, 0, -1, 0, 1, 1, 4, 2, 0, -2, 1, 0, -2, 0, -2, 1, 0, 1, 4, 5, 8, 8, 3, 1, 4, 0, -1, 0, 0, 1, 0, 0, -1, -1, 1, 2, 4, 5, 0, 0, 0, 0, -1, 0, 0, -2, 1, 2, 6, 3, 5, 5, 2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 5, 5, -1, 0, 0, 0, -2, -1, 1, 0, 0, 4, 6, 7, 5, 3, 3, 3, 4, 1, 3, 0, 2, -2, 0, -1, 2, -1, 1, 0, 4, 3, -1, 0, 0, 0, -1, 1, -1, 0, 2, 3, 5, 6, 4, 2, 2, 1, 0, 1, 0, 2, 0, 0, -1, 2, 0, 0, 1, 3, 2, 4, 1, 1, -1, -1, 0, -2, -3, 0, 3, 0, 5, 5, 5, 4, 4, 4, 2, 1, -1, 1, 0, 0, 2, -1, 2, 3, 2, 4, 3, 1, 0, 1, 0, -1, 0, -2, -1, -1, 3, 0, 5, 5, 2, 6, 3, 0, -1, -1, 0, 1, 1, -1, -1, 0, 1, 2, 0, 2, 4, 4, 1, 2, 0, 0, -1, -2, -1, 0, 1, 0, 0, 3, 2, 3, 4, 2, 0, -1, 0, -1, -1, 0, -3, 0, 0, -1, 0, 3, 3, 3, 2, 0, 1, 1, 2, 1, 2, 0, 0, 1, 2, 3, 2, 2, 5, 4, 2, 2, -1, 1, -2, 0, -4, -1, -2, 0, 2, 3, 4, 1, 2, 0, -1, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 3, 4, 1, 3, 2, 2, 0, 0, -2, -2, 0, 1, 0, 1, 0, 3, 3, 0, 0, -1, 0, -2, 0, 0, -1, 0, -1, -2, -1, -2, 1, 0, 1, 0, -1, -2, 0, 0, -1, -1, 0, 0, 1, -1, -1, -1, 0, 1, 1, 1, -1, 0, 0, -1, -1, 2, 0, 0, -1, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, 0, 0, -1, 0, 1, 1, 1, -1, 0, 1, 0, -1, 0, 0, -1, 0, 1, 0, 1, 1, 0, 1, -1, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 1, 0, -1, -1, -1, 1, -2, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 2, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, -1, -1, 0, 1, -1, -1, 1, -1, 1, 1, -2, 0, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, 1, -2, 0, 0, 0, -1, 1, -1, -1, 0, 1, -2, -1, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, -2, 2, 0, 1, 0, -1, 1, 1, 0, -2, -2, 1, -1, 0, -2, 1, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 1, 0, 0, -1, 1, 1, 2, 1, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, -1, -1, 1, 0, 0, 1, 0, 0, 1, 2, 0, 2, 1, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, -2, 0, -2, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, -1, -1, -2, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -2, 1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 2, 0, 1, -1, 0, 0, -1, 0, 0, -1, 2, 0, 0, 0, -1, 0, 0, -1, 0, -1, 2, -2, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -2, -2, 0, 0, 1, 1, -1, 0, 0, 0, -1, 2, 2, -1, 1, 0, 1, -1, 1, -1, -1, -1, 0, 1, -1, 1, 0, 1, -1, -1, 1, -1, 0, 2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, -1, 0, 1, -1, 1, -2, 1, 2, 1, 1, 0, -1, 0, -1, -1, 1, 0, 1, 0, 2, -1, 1, 0, 1, -1, -1, 0, -1, 0, 0, 1, -1, 1, -1, -1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, 0, 1, 1, -1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 2, 1, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 2, 2, 1, 1, -1, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, 1, 0, 1, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, -2, 0, -2, 0, 1, -1, -1, -1, 0, 1, 0, 1, 0, 0, -1, -1, -1, -1, -1, 1, -2, 0, 1, 0, 1, 2, 1, -1, -1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, -2, 0, 0, 1, 0, 1, -1, -1, 1, -1, 0, 0, 1, 1, 0, 0, -1, -1, 0, -1, 1, -1, -1, 0, -1, -1, 1, -1, 1, 1, -2, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 1, 0, 1, 0, 0, 1, -1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 1, -1, 2, -1, 0, -1, 2, -1, 1, 0, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 2, -1, -2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 2, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, -1, 1, 0, -2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, -1, -1, 0, 0, 1, 1, 1, 1, -1, 1, 0, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, 0, 0, 0, -1, 0, 0, 1, 0, 0, -2, 1, -1, 1, 0, 2, 0, -1, 2, 0, 1, 1, -1, 0, -1, 2, 2, 0, 2, 1, 1, 1, 2, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, -1, -1, 0, -1, 0, 1, 1, -1, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, -1, -1, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 0,
    -- filter=0 channel=2
    -4, -2, -2, -3, -5, -3, -3, -2, -2, 0, -1, -2, -3, -1, -3, -1, -2, -3, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, 0, 0, -6, -3, -4, -5, -3, -5, -3, -3, -2, -4, -1, -3, -4, -3, -3, -1, -3, -4, 0, -2, -1, 0, -2, -1, -1, -2, -3, 0, -2, 0, -3, -4, -1, -2, -1, -1, -5, -4, -4, -3, -1, -1, -3, -3, -4, -4, -2, -4, -4, 0, -4, -2, -1, 0, -2, 0, -1, -3, -1, 0, -3, -3, -4, -2, -1, -2, -4, -1, -3, -1, -3, -1, -4, -2, -4, -4, -2, -2, -1, -4, 0, -1, -3, -1, 0, -2, -1, -2, 1, 0, -5, -4, -2, -4, -4, -2, -4, -4, -1, -2, -3, -4, -3, -4, -4, -5, -5, -1, -4, -1, -3, -3, -4, 0, -1, 0, -1, -2, 1, 2, -1, -3, -3, -3, 0, -1, 0, 0, -3, -1, -1, -2, -1, -1, -2, -4, -4, -1, -2, -4, -3, -2, -2, -1, 0, 0, 0, 0, -1, 0, -2, -4, -2, -2, 0, 0, -3, -2, -2, -2, -2, -2, 0, -3, -3, -1, -3, 0, -2, -1, -3, -3, -2, 0, -3, 0, -2, -2, 0, 2, -1, -3, -4, -1, -3, -3, -2, -2, 0, -3, -4, -2, -3, -4, -3, -1, -1, 0, -2, -3, -2, -3, 0, -2, 0, -2, -2, -2, 0, 0, -1, -4, -3, -3, -2, -2, -2, 0, -2, -3, -1, 0, -2, 0, -2, -3, -2, -3, -1, 0, -1, 0, 0, -3, 0, -1, 0, 0, 0, 0, -3, -2, -3, -1, -2, -3, -1, 0, 0, 0, -2, -2, -2, -3, -2, 1, 0, 0, -1, -1, 0, 0, -2, -1, -2, -1, 0, -1, -2, 2, -3, -2, -2, -2, -1, -3, -3, 0, -3, -3, 0, -2, 0, 1, 1, 0, 0, 0, -2, -3, -1, 0, -2, -2, -2, -3, -3, 0, 0, 0, -2, -2, -3, -3, -3, -3, -2, 1, -2, -2, 0, 0, 1, 0, -1, 0, 1, -1, -2, -3, 0, 0, -2, -2, -1, 0, -1, 0, 1, 0, -4, -1, -1, -3, -2, -2, 0, -2, 0, 0, 0, 0, 2, 1, 1, 0, -1, 1, 0, 0, -3, 0, 0, 0, 0, -1, -1, 0, 0, 1, -3, -2, -3, -3, -3, -1, 0, -1, -2, 0, -1, -1, 2, -1, 1, -1, 0, 0, -1, -2, -2, -1, -2, 0, -1, 0, -3, -1, 0, 1, -4, -1, -2, -2, -1, -1, 0, 1, -1, -1, -1, 0, 1, 1, 2, -1, -3, -1, 1, 0, 0, -3, 0, -2, -2, 0, -2, 0, 0, 0, -3, -4, 0, 0, 0, -3, -2, -3, 0, -2, 0, 0, -1, 0, -1, 1, -2, -1, 0, 0, -3, -1, 0, -1, -1, 0, -1, -2, -1, 2, -4, -1, -3, -2, -1, -4, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, -1, -1, -3, -2, -3, -3, -1, -2, -1, 2, -1, -5, -3, 0, 0, -2, 0, -1, -2, 0, 0, 1, 0, 0, -2, -1, -1, 0, 0, -2, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, -4, -1, -1, -2, -1, -3, 0, 0, -2, 0, -1, 0, -2, 1, -1, -1, -2, 0, -1, -2, -2, 0, 0, -1, -3, -2, 0, -2, 0, 1, -2, -2, -4, -3, 0, 0, 0, -3, -3, -2, -2, 0, 0, 0, 0, 0, 0, -2, 0, -3, 0, -4, -1, -2, -2, 0, -2, -1, 0, 1, -3, -4, -4, 0, 0, -1, -3, -2, -2, -2, 0, -2, -1, -1, -3, 0, 0, 0, -4, 0, -4, -2, 0, -3, -3, -1, -3, -3, -1, -1, -1, -5, 0, -4, -3, 0, -2, 0, -4, 0, -3, -2, -3, -3, -1, 0, -3, 0, -4, -1, -4, -3, -1, -1, -1, -3, -1, -1, 0, 0, -4, -4, -4, -4, -1, -1, -1, -1, -4, -1, -1, -2, 0, -1, 0, 0, 0, -3, -3, -1, -1, -1, -1, -2, 0, -3, -1, 0, -2, 1, -3, -2, -4, -1, 0, 0, -1, -1, -2, -2, -1, -2, 0, -2, -1, -2, 0, -4, -3, -1, -1, -3, -1, 0, 0, -4, 0, -2, 0, -1, -1, -3, -4, -1, -3, -3, -4, -3, -4, -3, -1, -2, -3, -4, -1, -4, -1, -1, -3, -2, -2, 0, 0, -2, -1, -2, -3, 0, 1, 0, -5, -3, -4, -2, -2, -4, -2, -3, -2, -1, -1, -3, -1, -1, -4, -4, -3, -3, -1, -1, -3, -2, 0, -4, -2, -3, 0, -1, -1, 0, -3, -4, -3, -3, -3, -2, -3, 0, 0, -4, -1, -4, -1, -3, -3, 0, -3, -2, -3, -2, -4, 0, -1, -2, -2, -2, -1, -1, 0, 1, -5, -3, -2, -2, -3, -2, -1, -4, 0, -2, -1, -3, 0, -1, -1, -1, -2, 0, 0, -1, 0, -1, -4, -2, 0, 0, -2, -1, 0, -1, -3, -5, -3, -3, -3, -5, -1, -4, -4, -4, -1, -4, 0, -3, -3, -3, -4, 0, 0, -1, -4, 0, -1, -1, 0, 0, -2, 0, 0, 1, -2, -2, -3, -1, -4, -4, -2, -2, -2, -1, -4, 0, 0, -1, -1, -3, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, -4, -4, 0, -2, 0, 0, -2, 1, 1, -1, 0, 0, -1, -3, -2, -1, -3, 0, 0, 0, -3, -3, -4, -3, -4, -2, -4, -5, -2, -4, -2, 0, 1, 0, -1, 0, -1, 0, 2, 0, -1, 2, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -2, -2, -2, -1, -2, -4, 0, 0, -2, 1, 0, 1, 1, 0, 2, 1, 2, 0, 2, 1, 0, 1, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -3, -3, 0, 0, -1, -1, 1, 1, 2, 1, 0, 1, 0, 0, 1, 1, 1, 2, 3, 3, 2, 3, 0, 2, 0, -1, -2, 1, 0, 0, -1, -3, -2, -2, 0, 0, 1, -1, 0, 2, 4, 3, 1, 2, 2, 0, 2, 4, 2, 4, 4, 0, 2, 2, 2, 0, 1, -1, -2, 0, 0, -2, -2, 0, 0, 2, 1, 0, 2, 2, 1, 4, 1, 1, 4, 3, 4, 4, 4, 5, 4, 5, 3, 4, 0, 1, -1, -1, -1, 0, -1, -4, -2, -1, 0, 0, 1, 2, 4, 3, 3, 3, 4, 2, 5, 6, 6, 3, 3, 1, 5, 3, 2, 1, 3, 2, -1, 0, -1, 1, -2, -4, -3, -1, 0, -1, -2, -1, 3, 3, 4, 4, 5, 6, 5, 6, 3, 6, 5, 4, 3, 2, 5, 3, 3, -1, 0, -1, -2, 0, -1, -3, -2, -1, 0, -2, 0, 3, 3, 2, 6, 5, 5, 3, 4, 7, 4, 5, 6, 3, 2, 3, 4, 2, 3, 0, 0, -1, 0, 0, -1, -2, 0, -1, -2, -1, -1, 0, 3, 3, 4, 3, 3, 5, 3, 4, 7, 4, 2, 2, 2, 3, 3, 1, 3, 2, 0, 0, 0, 0, 0, -3, -2, 1, 0, 0, -1, 0, 0, 3, 1, 3, 5, 5, 6, 5, 5, 5, 0, 0, 0, 2, 3, 3, 1, 1, 1, 0, -1, 0, -3, -2, 0, 0, 0, 0, -1, -1, 1, 2, 0, 0, 2, 2, 1, 3, 4, 2, 1, 1, -1, 0, 1, 1, 0, 0, -2, -1, -1, 0, -2, -3, 0, 0, -1, -1, -1, 0, 2, 0, 0, 0, 0, 1, 4, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, -2, -2, -1, 1, 0, 0, 2, 2, 0, 1, 0, 0, -3, 0, 0, -2, -1, 1, 0, -1, -3, -1, -1, -3, -1, 0, -2, 0, 0, 0, -3, -1, -2, -1, -1, -2, 0, 2, 1, 0, 0, 0, -2, -2, 0, 0, 0, -1, -2, 0, -2, -4, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -3, -1, 1, 1, 0, 0, -1, -1, -5, -3, 0, 0, -2, -2, 0, -3, -2, -2, 0, 0, -2, -1, 0, 0, 1, 0, 0, -1, -3, -2, 0, -2, 1, -2, -1, 0, 1, 0, -3, 0, -2, -1, -1, 0, -1, -2, -1, -3, -3, 0, -3, -3, -1, 0, 1, 1, -1, -1, -1, -2, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, -4, -2, -5, -4, 0, -1, -2, -1, 0, 0, 2, 0, 2, 0, 2, 1, 1, 0, -1, -1, 1, 0, -1, 0, 2, 2, 2, -1, -2, 0, 0, -4, -1, -1, -1, -2, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 1, -1, 2, 1, 0, 2, 1, 2, -1, -2, -1, -3, -4, -1, 0, 0, 0, 0, -2, 2, 0, 3, 1, 3, 3, 3, 1, 1, 0, 0, 0, 0, 1, 2, 3, 1, 0, 1, 1, 1, 1, 0, -1, -2, 1, -2, 0, -1, -2, -1, 0, 0, 1, 5, 2, 4, 5, 3, 0, 1, 0, 2, 1, 2, 2, 2, 1, 0, 2, 0, 0, -2, -1, -2, 0, -1, -3, -3, 0, 1, 2, 4, 3, 2, 2, 6, 5, 3, 1, 2, 0, 1, 1, 2, 3, 1, 0, 1, 1, 0, 0, 0, -1, -2, -2, -1, -1, -2, -2, 0, 0, 0, 3, 2, 2, 3, 4, 3, 4, 3, 1, 4, 3, 3, 4, 0, 1, 0, 1, 0, 1, 0, -3, -3, -1, -2, -2, -1, 0, 0, 1, 2, 0, 3, 5, 2, 5, 3, 2, 0, 3, 3, 4, 3, 4, 0, 1, 0, 0, 1, 0, -2, -4, -3, -3, -2, -1, -1, 0, 0, 1, 0, 1, 2, 0, 3, 2, 2, 4, 3, 2, 4, 5, 5, 1, 0, -1, 0, 0, 2, -1, -1, -3, -3, -1, 0, -2, -1, 0, 0, 1, 0, -1, 2, 1, 1, 2, 3, 3, 3, 2, 1, 2, 3, 2, 0, 1, -1, 1, 0, -1, 0, -2, -1, 0, -2, 0, -1, 0, 0, -1, 0, -1, -1, 2, 0, 1, 2, 0, 1, 0, 3, 1, 3, 0, 2, 0, 0, 0, -1, 0, 0, -1, -2, -2, 0, -3, 0, 0, 0, 0, -1, 0, 2, 0, 1, 0, -1, 0, 0, 2, 1, 0, 2, 1, 0, 3, 2, 0, -2, -3, -3, -3, -4, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -3, 0, -4, -3, -2, -1, -1, -1, -1, -1, 0, -2, 0, -3, -3, -1, -3, -1, -3, -1, 0, -2, -1, -3, 0, -1, -1, -3, -2, -3, -1, -1, -3, -2, 0, -2, -3, 0, -1, -2, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, -3, 0, 0, -2, 0, 0, -1, 0, -2, -3, 0, -1, -3, -3, -2, 0, 0, 0, -1, 0, 0, -2, -1, -1, -1, 0, 0, -1, -2, -1, 0, -3, 1, 0, 0, 0, 0, 0, -2, 0, 0, -1, -3, -4, -3, -1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, 0, -2, -2, 0, 0, 1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -3, 0, -2, 0, 0, -2, -1, 0, 2, 0, 0, -1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, -1, -1, -1, 0, 0, -3, -4, -1, 0, -1, -1, -1, -1, -1, 2, 0, 0, 2, 2, -1, 2, 0, 0, 2, 0, 0, 0, 2, 2, -1, 0, 0, 0, 1, 0, -1, -1, -4, 0, -2, 0, -1, -1, 0, 2, 2, 1, 3, 0, 2, 0, 3, 0, 2, 0, 0, 1, 1, 2, 1, 0, 0, 0, 0, 0, -1, -1, -3, 0, -1, 0, -1, 0, 0, 0, 1, 1, 3, 1, 3, 2, 2, 2, 1, 0, 1, 3, 0, 0, 0, -1, 0, 1, 1, 0, 0, -3, -4, -1, 0, 0, -1, 0, 0, 1, 1, 3, 2, 3, 4, 3, 0, 4, 4, 0, 1, 1, 2, -1, 2, -1, 0, 0, 0, -1, 0, -4, 0, 0, 0, 0, 1, 0, 1, 2, 1, 4, 4, 1, 4, 1, 3, 2, 3, 0, 0, 3, 1, 1, 1, 1, 0, 0, 0, 0, -1, -3, -3, -2, -2, 1, 0, 0, 0, 2, 4, 2, 2, 2, 2, 2, 0, 1, 2, 3, 2, 0, -1, 0, -1, 0, 0, 1, 1, -1, -2, 0, 0, -2, -1, 1, -2, 0, 0, 1, 2, 0, 1, 2, 3, 1, 3, 2, 0, 2, 0, 2, 2, 0, 2, 0, 0, 2, 0, 0, 0, -1, -2, 0, -1, -1, 1, -1, 0, 1, 0, 0, 0, 2, 2, 2, 2, 1, 1, 0, 2, -1, 1, 2, 0, 0, -2, 0, -2, -1, -2, -3, -2, -1, 0, -1, 1, 0, -1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 2, 0, 0, -1, 0, -1, -1, -1, -2, 0, -2, -2, 0, 0, -3, -1, 0, 0, 0, -1, 0, 1, -2, 1, 1, 2, -1, 1, 0, 2, -1, 0, 0, 0, 0, -3, 0, 0, 1, 1, -2, -2, 0, 0, -3, 0, -1, 0, 0, 0, -2, 0, -2, 0, 1, 0, 0, 2, 2, 0, -1, 1, 0, 0, 0, 0, -2, 1, -2, -2, 0, -1, -2, 0, -3, -2, 1, -2, 0, -2, 1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -2, -2, 0, -2, 0, -2, 0, -2, 0, 0, 0, -1, -3, -3, 0, -3, 0, 0, 1, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 0, -1, -2, -1, -4, -2, 0, 0, 0, -2, 0, 0, -1, -1, 1, 0, 1, -1, 0, 1, 0, 1, 0, 0, 1, 0, 1, -1, -1, -1, -2, -2, 0, -1, -3, 0, -2, -2, 0, -1, 0, 1, -1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, -3, -3, 0, 1, 0, 1, 0, 0, 0, 2, 1, 0, 3, 2, 2, 0, -1, -1, -1, 0, 0, 2, 0, 2, 0, 0, -1, -2, -2, 1, -1, -1, 0, -1, -2, -2, 0, 0, 0, -1, 0, 1, 0, 3, 2, 3, 2, 0, 0, 0, -1, -1, 0, 2, 2, 0, 1, 1, -1, -1, -3, 0, 0, -2, -1, 0, 0, -1, -1, 0, 0, 2, 2, 2, 2, 1, 2, 0, 1, 0, 1, -1, 1, 2, 2, -1, -1, 0, 1, 1, -1, -1, 0, -2, -3, 0, -1, 0, 0, -1, 0, 1, 1, 3, 2, 1, 0, 0, 0, 0, 1, 1, 2, 3, 3, 0, 1, -2, 1, 0, -2, -3, -4, -3, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 3, 0, -1, 2, 0, 0, 0, 0, -1, -1, -3, -2, -2, 0, -2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 1, 1, 0, 1, 3, 1, 1, 1, -2, 2, 0, -1, -1, 0, -1, -2, 0, -2, 0, -3, -1, -1, 0, 0, 0, -1, -1, 0, -1, 2, 1, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, -2, -4, -2, -2, -1, -3, -3, 0, 0, -1, 0, 0, 0, -1, 0, -2, 1, 0, 0, -1, 1, 1, 0, 2, 1, 0, 1, 0, 0, 0, -1, -2, -1, -1, -2, 0, -3, -2, 0, -3, -1, -2, -2, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 2, 0, -2, 0, -1, 0, -4, -1, -2, -1, -3, -2, -2, -1, -2, -1, 0, -1, -2, 0, -1, 1, 0, -2, 0, 0, 0, 0, 0, 0, -2, 0, -1, -3, -1, -3, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -2, 1, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, 1, 0, -1, 1, 0, 2, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 1, 1, 0, 0, 0, -1, 1, -2, 1, 1, 0, -1, -1, 0, -1, 0, -1, -2, 1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 1, -1, 0, 0, 0, 0, 1, -1, 0, -2, 0, 0, 0, -2, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 1, 1, 2, 0, 0, 1, -1, -2, -1, 0, 0, -2, 1, -1, -2, 1, -1, 0, -1, 0, -1, 1, 0, -1, 0, 0, 1, -1, 0, 0, 0, -1, -2, 0, -1, 0, -1, -1, -1, -1, -1, 0, -1, 0, -1, -1, -1, 1, 0, -1, 2, -1, 1, 0, 2, 0, -1, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 1, 2, 0, 2, 0, 0, -1, 1, 0, -1, -1, 0, 0, 0, 2, 0, -2, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, -2, 1, -1, 1, -1, 1, -1, 1, 0, 1, -1, 1, 0, 0, 0, 1, 0, -1, 0, 0, -2, 1, -1, 0, 1, 0, -1, -1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, -2, 0, 0, 0, 2, 2, 1, -1, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, -1, -1, 1, 0, -1, 0, 1, 0, -1, 0, 1, -1, 0, 0, 1, 0, 1, 1, -1, 1, 0, 0, -2, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, -2, -1, 1, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, -1, 1, 1, 0, 0, 0, 1, -1, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 1, 2, 1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 1, 1, 1, -1, 0, 0, 0, -1, -1, 1, 0, 2, 0, 0, -1, -2, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 2, 1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, -1, 1, 0, 2, 0, -1, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, 1, 1, 0, -1, -1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, 0, -1, 0, -2, 1, -1, 0, 0, 2, 2, 0, 2, -1, 1, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -1, 2, -1, -1, -1, 0, -1, 0, 0, -1, -1, -1, 0, 2, 0, -1, 2, -1, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, -1, -1, 0, 0, 1, 1, -1, 0, -1, 0, -1, 0, -1, 0, 2, 1, 1, 0, 0, 1, -2, 0, 0, 0, 0, 1, 0, -2, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 1, -1, -1, -1, 1, 0, -1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, -2, -1, 1, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 2, 1, 1, -1, 0, -1, 1, 2, 1, 0, 1, -1, 2, -1, 1, 0, 0, -2, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 0, -2, 0, -2, 0, 0, 0, 0, -1, 0, 1, -2, 1, -2, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 1, 1, -2, 0, -1, 1, 2, 0, 0, -1, 0, -1, 0, -1, 0, 0, -1, 0, 2, 0, -1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, -1, 1, 0, 1, 0, -1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, -1, 1, -1, 1, 0, -1, 1, 1, 1, -1, 2, 1, 3, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 1, 0, 1, 1, 1, 0, 0, -2, -2, 0, -2, 0, 0, 0, -2, 0, 1, 1, 0, 2, 3, 0, 3, 4, 3, 0, 1, 2, 0, 2, 0, 1, 0, 2, -1, -1, -1, 0, -1, 0, -2, 1, 0, 0, -1, -2, 4, 0, 2, 0, 2, 2, 0, 4, 2, 3, 1, 0, 2, 1, 3, 1, 1, 2, 2, 1, 0, 2, 2, -1, 0, 0, 2, 2, 0, -1, 1, 1, 0, 3, 0, 0, 1, 2, 1, 0, 2, 0, 1, 2, 1, 0, 1, 3, 1, 3, 2, 2, 0, 3, 3, 1, 0, 2, 0, -2, 2, 0, 0, 3, 0, 0, 2, 0, 1, 0, 0, 0, -1, 0, 0, 2, 0, 0, 0, 2, 3, 3, 0, 1, 0, 0, 0, 0, 0, 0, -1, 2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 2, 0, 0, 2, 0, 1, 0, 3, 1, 0, 1, 0, 2, 1, -1, 0, -1, 0, 0, 3, 2, 0, 0, 0, -1, 0, 0, 0, -2, -2, -1, 0, -1, 0, 3, 1, 1, 2, 2, 0, 2, 0, 0, 0, -1, 1, 0, -1, 0, 1, 3, -1, 0, -3, -2, 0, 1, 1, 0, -1, 0, -1, -1, 0, 3, 2, 0, 1, 0, 1, 1, 0, 1, 2, 2, -1, 0, -2, 2, 1, 0, 1, -2, -3, 0, -1, 1, 0, -1, 0, -1, 2, 1, -1, 1, 0, 0, -1, -1, 1, 0, 2, 0, 1, -2, 0, 0, -2, 1, 1, -1, -1, 1, 1, -3, 0, 0, 1, 1, 1, 0, 1, 0, 0, -3, 0, -3, 0, 0, -2, 1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, -2, -3, 0, 0, 0, 0, -2, -3, 0, 0, -2, -2, -4, 0, -1, 0, -1, 0, 0, -2, 0, 0, 0, -2, 2, 0, 2, 2, 0, 1, 0, -1, 0, 0, -2, 0, -3, -4, -3, -3, -5, -4, -4, -2, -2, 1, -1, 0, 0, -3, 0, 0, 0, -4, 3, 3, 0, 0, 1, -1, 0, 1, -2, 0, -1, -1, -3, -4, -4, -5, -5, -2, -2, -3, -2, -1, 0, -2, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -2, -1, -1, -1, -1, -2, -2, -4, -3, -5, -4, -2, -3, -5, -3, -5, -1, -1, -2, -2, 1, 0, 0, 0, -3, -4, 0, 1, 2, 1, -2, 0, 0, -2, -2, -3, -3, -3, -7, -5, -3, -5, -5, -4, -4, -6, -2, -3, 0, 0, 0, -1, -3, -1, 0, -3, 2, 1, 1, -1, 0, -1, 0, -1, -4, -2, -4, -3, -3, -3, -6, -5, -3, -3, -4, -4, -4, -2, -1, 0, 1, 0, 0, 0, -2, -1, 1, 1, 1, -1, -3, -1, -2, 0, -1, -2, -3, -5, -5, -3, -7, -3, -5, -2, -5, -2, -2, -2, -1, -2, 1, 1, -2, 0, -1, -1, 0, 0, 0, -2, -2, -1, 0, -2, -1, 0, -1, -4, -6, -5, -5, -2, -3, -5, -1, -2, -1, -1, -2, -2, 1, 0, 0, 0, -3, -3, 1, 1, 0, -1, -1, 1, 0, -2, -2, -4, -4, -2, -6, -3, -5, -4, -1, 0, -4, -3, -1, -2, 1, 0, 0, 0, 0, -2, -2, -3, 1, 2, 1, 1, 1, 0, 0, 0, -1, -1, -2, 0, -2, -5, -4, -5, -2, -1, -2, -2, -1, 0, 0, 0, 3, 1, 1, -1, 1, 0, 0, 2, 0, 2, -1, 0, -2, -2, 0, 0, 1, -1, -1, -3, -1, -1, -3, -6, -3, -2, 1, 1, 0, 1, 1, 2, 0, -1, 0, 0, 0, 0, 2, 0, -2, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, -2, -4, -1, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, -2, -1, 2, 0, 0, 0, -1, 1, -1, 0, 0, 2, 1, 0, 1, 1, 0, 1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, -2, 0, 0, -1, 2, 0, 0, 0, 1, 2, 1, 0, 0, 0, 2, 0, 1, -1, 0, 0, 2, 1, 1, 2, 0, -1, 1, 2, 1, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 3, 0, 2, 2, 0, 1, 1, 2, 2, 4, 2, 1, 0, 0, 0, 2, 1, 0, -1, 0, 0, 0, 2, 2, -1, 0, 0, 1, 2, 3, 1, 2, 1, 0, 2, 3, 2, 1, 3, 3, 3, 0, -2, -1, 1, 0, 2, 1, -1, -1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 1, 1, 1, 0, 2, 0, 2, 2, 1, 2, 1, 2, 0, 1, -2, -1, 0, 0, 1, -1, 0, 1, 0, 2, 0, 0, 2, 3, 2, 0, 1, 0, 0, 0, 2, 2, 3, 1, 2, 0, 0, 1, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 2, 0, 0, 3, 1, 2, 3, 0, 2, 0, 1, -1, 0, 2, 2, 0, 1, 1, 3, 0, 2, 1, 0, 0, -1, 0, -1, -2, 2, 1, 2, 2, 0, 3, 3, 4, 3, 3, 1, 1, 2, 0, 1, 0, 1, 0, 3, 1, 1, 3, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, 0, -2, -2, -1, -1, -1, -2, 0, 0, -1, -2, -1, 0, 0, -1, -2, -2, -2, -2, -1, 0, -2, -1, -2, 0, -2, -1, -2, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -1, -3, -1, -1, 0, -1, 0, -3, 0, 1, 0, 0, 0, -1, 1, -2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, -2, -3, -1, 0, 0, -2, -2, 0, -2, 0, 0, -2, 0, 0, 0, -1, -1, -2, -3, -2, -2, -3, -2, -3, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 1, -2, 0, 2, -1, -2, 0, -2, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, 0, -1, 0, 0, -2, 0, -1, 0, -1, 0, -2, 0, -1, 2, -2, 0, -2, -1, 1, 0, -2, 0, -2, 0, -2, -2, -1, -2, -3, 0, -1, -3, -2, -2, -2, 0, -1, 1, 0, 0, -2, 1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, -3, -1, -1, 0, 0, 0, -1, -1, -2, 0, -1, 1, -1, 1, 0, 0, -1, 1, -2, -1, 1, 0, 0, -2, 0, 0, -1, 0, -2, 0, -3, -1, -1, 0, -3, 0, -1, -1, 0, -1, 0, -1, -1, 0, 1, -2, -1, -1, 1, 0, 1, 0, -2, -1, 0, 0, -3, -2, -1, 0, 0, -1, -3, -2, -1, -2, -1, -1, -1, 1, -1, 0, 0, -2, -1, -1, -1, 0, 0, 0, -1, -1, 0, -2, 1, -1, -2, 1, -1, 0, 0, 0, 0, -2, 0, 0, -2, 0, 0, -1, -1, -1, 0, 0, 1, -1, -1, 1, 1, 1, -1, 0, -1, -1, 0, 0, -1, -2, -2, 0, -1, 0, -2, -1, 0, 0, 0, -1, -1, -1, -2, -2, 0, 0, -2, -2, 0, 1, -2, -1, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, -2, 0, 1, -1, -1, 0, -1, -1, -2, -1, 0, -2, -1, 0, 0, -2, -1, 0, 1, -1, 0, -2, 1, -1, 0, -1, 1, 0, 0, -2, 0, 0, -1, -1, 1, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, -1, 0, -1, -2, -1, -1, 0, 1, -1, -1, -2, 0, 0, -2, -1, -1, -1, -2, -1, 0, 0, -1, -1, -1, 0, 0, -1, 0, 1, 0, -2, -1, 1, 0, 0, 1, -1, -2, 0, 0, 0, 0, -1, 0, -2, 0, -2, -1, 1, 1, 0, 0, 0, -1, -2, 0, -2, 0, -1, 0, 0, 0, 0, 1, -2, -1, 0, -1, -1, -2, 0, -2, 0, -2, 0, 0, 0, -1, -1, 0, 1, -1, -1, 0, -1, 0, 0, 0, -1, 1, 0, -1, -1, 0, -1, -2, -2, -1, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, -1, 1, 1, 0, 0, -2, 0, -2, 0, -1, 0, -2, 1, 0, 0, 0, -1, 0, 1, -1, 1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, -1, -2, 0, -2, -2, 0, 0, -2, 0, 0, 0, -2, 0, -2, -1, -1, -1, 1, 0, -1, 0, 0, -1, 0, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, -2, -2, 0, -1, -3, 0, 0, 0, -2, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 1, -2, 0, -1, 0, 0, -2, -2, 0, -1, -2, -1, 0, -1, -1, -1, 0, -1, 0, -1, 0, 1, -2, 0, -2, 0, 0, 1, -1, -1, 0, 0, -2, 1, 0, 0, -2, -1, 0, -1, 0, -2, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, -2, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 1, 0, -2, 0, -1, 0, -1, -2, 0, -1, -2, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, 0, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -3, 0, -3, -2, 0, -2, -1, -1, -2, 0, 0, -2, 0, -1, 0, -1, -2, -2, 0, 1, 0, 0, -3, -2, 0, 0, 0, -3, 0, -2, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, 0, -3, -1, 0, -1, -1, 0, 0, 0, 0, -3, 0, 0, -1, -2, 0, 0, -2, -2, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -2, -2, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 0, 1, -2, 0, 0, -2, -2, 0, -2, -1, -2, -2, 0, 0, 0, 0, -2, -2, 0, 0, -1, -2, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 1, -1, -2, -2, 0, -2, 0, 0, 0, 0, 1, -2, -1, -1, -2, 0, 0, 0, -2, 0, 0, 0, -2, -1, -1, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 1, 0, 1, -1, 1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, -1, -1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 1, 0, -1, 1, -2, 2, 0, 2, 0, -1, -1, -1, 0, 1, -1, 0, 0, -1, 0, -2, -1, 1, 0, 0, -1, -2, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 2, -1, 0, -2, -1, -2, 0, -1, -1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, -2, 0, 0, -1, -1, 0, 2, 0, 2, 0, 0, 0, 0, -1, -1, 0, -2, -1, 1, -1, 0, 0, 0, 0, -1, 2, -1, -1, 2, 0, 0, 1, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 0, 1, -2, -1, -1, 1, 0, 1, 2, 0, 1, 0, 0, -1, 1, 0, 0, 1, -1, -1, 0, 0, 0, -2, -1, 0, 0, -1, 0, 1, 0, 0, 2, -1, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, -2, 1, 0, 0, -2, 0, 1, 0, -1, 0, 1, 0, 0, 0, 2, 1, -1, 0, 1, 0, -1, -1, 1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -2, -2, -2, 0, -1, -1, -1, 0, 1, 0, 0, 0, -2, -1, 1, -1, 0, 1, 0, 0, -1, -1, 0, 1, -1, -2, 0, 1, 0, -2, -2, 0, 0, 0, -1, -2, 1, 0, 0, 0, 1, 1, -2, 0, -2, -1, -1, 0, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, -2, -2, -2, -2, -1, -2, -1, 0, -1, -1, 0, -1, -1, 0, 0, -2, -1, 0, -1, -2, 0, 0, 1, 0, -1, 0, -1, 0, -1, -2, -1, -1, 1, 0, 0, -1, -1, 1, 0, 1, 0, 1, 1, 2, 0, 0, 0, 0, 1, 0, -2, -1, -2, 0, 0, -1, -1, -2, 0, -1, 1, -1, 0, 0, 1, 0, -1, 0, 1, 1, -1, 0, 0, 1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 1, -1, 0, -2, 1, -1, -1, 0, 1, 1, 0, 0, -2, 1, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, 1, -2, -2, -1, 0, 1, -1, 0, 0, 0, -2, 0, 0, 1, -2, 0, -1, -1, -2, 0, -1, -2, 0, 0, -1, -1, 0, 1, 0, 1, -1, 0, 1, -1, 1, 1, -1, -1, 0, 0, 0, 1, -1, -1, 0, -2, -1, -2, -2, 1, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, -2, 0, 0, -2, -1, 0, 1, -2, 1, -1, 1, -1, 0, 0, 0, -1, -1, 1, -1, -1, -1, 1, 1, 0, -1, 1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, -2, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 1, 0, 0, -1, 1, -1, -2, 0, 0, -2, -2, 0, -1, -1, 0, -3, -2, -2, 0, -2, 0, 1, -1, -1, 0, 1, -1, 0, -1, 0, 1, 0, 0, 0, -2, -2, -1, -1, -1, -1, 0, 1, 0, 0, -2, -2, 0, 1, 0, -2, -1, -2, 0, 0, 1, 2, 0, -1, -1, 0, 0, 2, 2, 0, -1, -1, -2, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, 1, 1, -1, 1, 1, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, 1, 0, 0, -2, 1, -1, 1, 0, -1, -1, 0, 0, 2, 2, 0, 0, 1, 0, 2, 2, -1, 0, 1, 1, 0, 1, -1, -2, 0, 0, -2, 0, -2, -2, -1, 0, 0, 2, -1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 2, 0, -1, -2, -1, 0, 1, 1, 0, 0, 1, -1, 1, 0, -1, 1, 0, 0, 0, -1, -1, 0, -1, 2, 0, 0, 0, 1, 0, 1, 2, 0, 0, 0, 0, 0, 1, -1, 0, -1, 1, 2, 1, 0, 0, -1, 2, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 2, 2, 0, -1, -1, 1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 1, 1, 0, 0, 0, -1, -1, -1, -1, 0, 1, 2, 0, 2, 1, 0, 1, 1, 1, -1, -1, 1, 0, 0, 0, 2, -1, 1, -1, 1, -1, 1, 1, 0, 2, 2, 0, 2, -1, 0, -1, 0, 0, 2, 2, 0, -1, 0, -1, -1, 0, -1, 2, 1, 1, 1, 0, 0, -1, 1, -2, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, 2, 0, 0, 2, 1, 1, -1, 2, 2, 0, -1, 0, 2, 1, 0, 1, 0, -1, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, 2, 1, 2, 0, 0, 1, 2, 2, 0, 0, 4, 1, 3, 3, 2, 2, 3, 2, 2, 4, 2, 2, 0, 2, 2, 2, 1, 0, 3, 3, 3, 1, 1, 1, 0, 0, 2, 0, 1, 0, 4, 3, 3, 1, 3, 2, 0, 3, 2, 2, 2, 0, 1, 1, 4, 0, 4, 2, 4, 3, 3, 3, 3, 3, 1, 0, 2, 0, 1, 0, 4, 2, 4, 1, 4, 4, 2, 1, 3, 3, 3, 2, 3, 2, 2, 4, 3, 4, 4, 4, 2, 3, 1, 1, 0, 1, 2, 0, 0, 1, 0, 2, 3, 1, 0, 0, 5, 4, 5, 5, 1, 5, 3, 3, 3, 1, 2, 3, 5, 4, 3, 1, 0, 2, 3, 0, 2, 2, 0, -2, 4, 3, 0, 1, 3, 3, 2, 1, 3, 0, 2, 2, 3, 4, 2, 4, 4, 1, 3, 1, 3, 2, 1, 3, 2, 0, 0, -1, 0, -1, 1, 4, 0, 3, 0, 4, 1, 3, 2, 2, 3, 2, 1, 3, 3, 4, 3, 4, 2, 3, 2, 2, 3, 0, 1, 0, 0, 0, -1, 0, 2, 4, 2, 2, 1, 4, 2, 3, 4, 3, 5, 1, 5, 1, 5, 4, 1, 4, 4, 2, 4, 0, 3, 2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 4, 2, 3, 4, 3, 4, 3, 5, 2, 2, 0, 3, 3, 3, 1, 0, 4, 2, 3, 2, 0, -1, -1, 0, -1, 2, 3, 3, 1, 0, 0, 1, 3, 3, 3, 2, 1, 2, 2, 1, 0, 0, 4, 0, 2, 1, 1, 3, 0, 2, 0, 0, 0, 0, -3, 3, 3, 1, 2, 1, 2, 2, 3, 3, 4, 3, 2, 3, 0, 2, 1, 3, 2, 0, 3, 3, 0, 2, 0, 0, 2, 0, 0, 0, -4, 4, 3, 1, 2, 0, 3, 1, 1, 0, 0, 0, 2, 2, 3, 3, 2, 0, 2, 2, 3, 3, 2, 0, 1, 1, 1, 1, 0, -2, -4, 3, 3, 0, 0, 3, 3, 1, -1, 0, -1, 0, 0, 2, 0, 3, 2, 1, 3, 2, 0, 1, 2, 0, 1, 0, -1, -1, 0, -3, 0, 2, 3, 1, 2, 2, 0, 0, 1, 2, 0, -1, 0, 1, 1, 1, 0, -1, 1, 0, 0, 0, 2, 2, 0, 1, 1, 0, -2, -2, -2, 2, 3, 1, 2, 2, 0, 0, 1, 1, -1, 0, -2, 1, 0, 0, 2, 2, 1, -1, 0, 1, 2, 0, -1, -1, -2, 0, -2, -2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 1, -1, 0, 2, 0, 0, -1, 0, 0, -1, -1, -1, -2, -4, 1, 2, 1, 0, 2, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, -1, 1, 1, 2, 0, 0, 2, -1, 0, 1, -1, -1, -2, -3, 0, 0, 0, 0, 2, 0, -1, 0, -1, -2, -2, 1, -1, 0, 0, 0, -1, 1, 0, 3, 0, 2, 0, 0, -1, 0, -1, 0, -3, -1, 3, 2, 0, 1, 1, 0, 1, -1, 1, -1, 1, 0, -2, 0, 0, 0, 0, 2, 0, 1, 0, 3, 2, 1, 2, 0, -1, 0, -3, -2, 2, 2, 2, 0, -1, 0, 0, 2, 0, 0, 1, 1, 1, 0, 0, 2, 0, 2, 1, 3, 0, 1, 2, 1, 1, 0, 0, -1, -1, -1, 4, 3, 2, -1, 0, 0, 0, 0, 0, 2, 3, 1, 1, 1, 0, 2, 2, 0, 2, 2, 0, 0, 2, 3, 0, 1, 1, -1, -2, -3, 0, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 1, 3, 3, 4, 0, 0, 4, 3, 4, 1, 3, 2, 0, 3, 0, 0, 1, 0, 0, 0, 3, 1, 2, 1, 0, 1, 3, 1, 0, 3, 1, 2, 0, 3, 1, 1, 0, 2, 3, 1, 3, 0, 1, 0, 3, -1, 0, 1, -1, 3, 3, 1, 0, 0, 0, 4, 2, 2, 4, 4, 0, 3, 4, 2, 0, 2, 4, 1, 2, 2, 3, 0, 1, 2, 1, 0, 0, 0, -2, 4, 2, 2, 2, 0, 3, 1, 0, 4, 4, 2, 4, 2, 2, 5, 4, 2, 2, 0, 3, 0, 2, 3, 3, 0, 0, 1, -1, 1, -3, 2, 3, 2, 3, 3, 2, 1, 1, 4, 3, 4, 2, 1, 5, 1, 4, 5, 2, 2, 4, 1, 2, 0, 1, 2, 0, 0, 2, 0, 1, 1, 4, 1, 1, 3, 2, 1, 3, 4, 4, 4, 3, 4, 3, 5, 5, 3, 1, 3, 3, 4, 1, 3, 2, 3, 0, 0, 0, -1, -1, 2, 4, 0, 0, 2, 4, 3, 4, 3, 2, 4, 4, 4, 4, 3, 1, 1, 4, 2, 4, 2, 1, 2, 3, 2, 2, 1, 0, 0, 0, 3, 3, 2, 1, 2, 4, 1, 4, 5, 3, 1, 2, 0, 4, 4, 5, 2, 1, 0, 3, 4, 4, 2, 1, 0, 1, 1, -1, 1, 0, 2, 1, 1, 4, 3, 4, 4, 2, 1, 1, 4, 1, 2, 2, 1, 2, 4, 0, 4, 2, 1, 2, 2, 1, 1, 1, 0, 1, 1, -1, 4, 3, 0, 0, 3, 4, 1, 2, 1, 0, 1, 3, 2, 0, 2, 3, 1, 1, 2, 1, 1, 0, 2, 0, 0, 2, 1, 0, 0, 2, 10, 10, 7, 8, 5, 7, 6, 8, 6, 6, 5, 3, 3, 4, 3, 2, 5, 2, 4, 3, 0, 0, 1, 0, -1, 0, 0, 1, 1, -2, 9, 9, 10, 8, 8, 5, 7, 8, 6, 5, 6, 4, 4, 4, 5, 5, 6, 4, 3, 3, 2, 2, 3, 0, 3, 3, 0, 3, 0, -1, 7, 8, 8, 8, 7, 5, 7, 8, 6, 5, 4, 3, 5, 3, 3, 7, 4, 4, 4, 5, 5, 4, 2, 3, 3, 1, 2, 1, 3, -2, 8, 9, 8, 6, 7, 3, 7, 5, 7, 4, 3, 1, 2, 4, 2, 6, 3, 5, 5, 4, 6, 4, 6, 3, 3, 3, 2, 1, 3, 0, 9, 5, 7, 6, 4, 6, 4, 4, 4, 3, 3, 3, 3, 1, 2, 2, 4, 3, 6, 7, 4, 7, 6, 5, 3, 2, 4, 3, 0, 0, 8, 8, 6, 4, 3, 3, 3, 3, 4, 2, 2, 3, 0, 3, 3, 1, 4, 4, 5, 6, 5, 4, 5, 3, 1, 3, 1, 2, 1, 0, 9, 6, 6, 5, 1, 1, 2, 0, 0, 2, 1, 2, 2, 0, 3, 2, 1, 0, 3, 4, 4, 5, 5, 4, 3, 4, 3, 1, 2, 0, 6, 8, 3, 3, 3, 0, 0, 0, 1, 0, -1, -1, 0, 1, 3, 2, 1, 0, 1, 2, 4, 4, 5, 1, 1, 2, 2, 1, 0, -3, 7, 5, 3, 2, 3, -1, 1, -2, 0, -1, -2, -2, 0, -2, -1, 1, 1, -2, 1, 0, 0, 1, 0, 2, -1, 0, 1, -1, 0, -2, 6, 3, 1, 1, 1, 0, 1, 0, -1, -2, -2, -2, -1, -3, -3, 0, -3, -3, 0, 1, 0, 2, 1, 1, 2, 2, 0, -2, -1, -6, 8, 4, 1, 1, 0, 0, -2, -1, 0, 0, -1, -1, -2, -1, -5, -3, -7, -5, -1, 0, 0, 2, 0, 1, 0, 1, 0, 0, -4, -6, 7, 6, 1, 1, -1, -2, 0, -1, -1, -4, -4, -2, -4, -6, -6, -8, -8, -8, -4, -2, -1, 2, 0, 2, 0, 0, -1, -2, -5, -7, 6, 2, 1, 2, 1, -1, 0, 0, -1, -4, -4, -4, -6, -7, -8, -10, -7, -8, -4, -2, 1, 1, 0, 1, 0, -2, 0, -1, -4, -4, 4, 3, 0, 0, -1, 0, 0, -2, -2, -6, -5, -5, -8, -9, -10, -9, -6, -6, -3, -2, -1, -1, 0, 2, 0, -1, -1, 0, -5, -7, 4, 5, 2, -1, -2, 0, -1, -3, -4, -6, -4, -6, -10, -7, -8, -9, -7, -5, -4, -3, 0, 0, 1, 1, 0, 0, 0, -2, -5, -7, 3, 6, 3, 1, 0, -3, -4, -4, -2, -5, -7, -7, -10, -10, -8, -9, -8, -4, -4, -3, -2, 0, 1, 2, 2, 0, 1, 0, -1, -7, 4, 3, 1, 0, -1, 0, -1, -1, -3, -5, -8, -9, -11, -7, -11, -7, -7, -6, -6, -3, 0, 0, 0, 2, 0, 0, -1, 0, -2, -4, 7, 4, 1, 0, -1, 0, -2, -2, -5, -3, -6, -9, -9, -7, -9, -8, -6, -4, -3, -3, 0, -1, 0, 2, -1, 1, 1, -1, -3, -4, 5, 5, 2, 0, 1, 1, 1, -1, -5, -3, -6, -8, -9, -6, -8, -5, -6, -6, -3, -4, -1, 0, 2, 2, 1, -1, -2, -2, -1, -5, 4, 3, 4, 4, 0, 0, -1, -2, 0, -1, -4, -5, -6, -7, -5, -5, -3, -3, 0, 0, 0, 2, 1, 0, 3, 2, 0, 0, -2, -6, 8, 3, 2, 5, 2, 0, 0, 0, 1, -2, -1, -2, -4, -6, -5, -7, -3, -3, -3, 0, 1, 2, 2, 1, 3, 1, 1, 0, -3, -5, 8, 4, 4, 1, 1, 3, 1, 2, 3, 0, 1, -2, 0, 0, -4, -3, -6, -2, 0, -1, 0, 1, 2, 1, 4, 4, 3, 0, -1, -4, 8, 4, 4, 2, 1, 3, 2, 1, 1, 1, 1, 2, 2, 1, -2, -2, -1, 0, -1, 0, 2, 5, 3, 2, 4, 5, 2, 2, -1, -1, 7, 7, 5, 5, 4, 5, 6, 3, 2, 1, 3, 4, 4, 1, 0, 3, 2, 3, 2, 3, 3, 3, 2, 2, 2, 5, 2, 0, 1, 0, 6, 7, 5, 4, 5, 5, 6, 6, 5, 7, 4, 5, 2, 5, 4, 2, 1, 5, 2, 3, 2, 3, 1, 0, 2, 1, 1, 3, 0, 0, 5, 7, 4, 5, 6, 8, 6, 6, 4, 5, 7, 6, 3, 7, 7, 6, 6, 4, 4, 3, 4, 3, 1, 2, 3, 2, 0, 2, 0, -2, 8, 6, 5, 5, 6, 8, 5, 5, 6, 6, 3, 5, 3, 3, 6, 7, 4, 6, 5, 6, 1, 4, 1, 2, 3, 2, 1, 1, -1, -2, 9, 10, 4, 4, 6, 8, 8, 5, 6, 8, 5, 4, 6, 4, 4, 5, 6, 5, 3, 6, 4, 2, 5, 5, 4, 3, 2, 1, -1, -1, 9, 9, 6, 4, 7, 8, 6, 6, 7, 6, 8, 5, 3, 5, 4, 5, 7, 4, 6, 3, 4, 4, 5, 2, 1, 0, 0, 1, 0, 0, 10, 10, 10, 7, 9, 7, 11, 9, 9, 6, 7, 4, 6, 5, 5, 4, 3, 6, 2, 3, 3, 1, 2, 2, 0, 0, 1, 0, 1, 1, -1, 0, -2, -1, 0, -1, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 1, -2, 0, -1, 1, -1, 0, -1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, -2, -1, -1, 2, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, -1, -1, 0, -2, 0, -2, -1, 1, -1, -2, -1, 0, 1, 0, 0, 1, 0, 1, 0, -1, 0, 1, -1, 1, -1, 0, -1, 0, 0, -1, 1, -1, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -2, 1, 0, -1, 0, 1, 0, 1, 0, 2, 0, -1, -2, 0, 0, 0, 0, -1, 1, 1, 0, -1, 0, 1, 1, -1, 0, 0, 1, 0, -2, 0, -1, 0, 1, 0, -1, -1, 1, -1, 0, 1, 1, -1, 1, 0, 0, 1, 0, -1, 1, -1, 1, 1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 1, -1, 0, 0, 2, 1, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 1, -2, 0, -1, -2, -1, 1, -1, 0, -1, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 1, -1, -1, -1, -1, -1, 0, -1, -1, -1, 1, 0, -1, -2, 0, 1, 1, 1, 1, 1, 2, -1, 2, 0, 0, 0, 2, -2, 0, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 1, 0, -1, 0, -1, 0, 1, 2, 0, -1, -1, 0, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 1, -1, 0, -1, 0, 0, -2, -1, -1, -2, 0, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, 1, 2, -1, 1, 0, 0, 2, 1, 0, -1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, -1, 1, -1, 0, -1, 0, -1, -1, 0, 0, 1, -1, 0, 0, -1, 1, -1, 0, 1, 1, 0, 0, 1, -2, 2, 0, 0, 1, 1, 0, 2, 2, 0, 2, 0, 0, 1, 0, 1, -1, -1, 2, 0, -1, 0, 1, -1, 0, 1, 0, -1, -2, 0, 0, 0, 2, 2, 1, -1, 1, 0, 1, -1, 0, -1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 1, -1, 0, 0, 0, 1, 1, 0, 1, 2, 0, 1, -1, -1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, -2, -1, -2, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, 1, 1, -1, 2, -1, 0, -1, -1, 0, 1, 0, -1, -1, -1, 0, 1, 1, 0, -1, -2, 1, 1, -1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, -2, 0, 2, 0, 1, 0, 0, 0, 0, 1, 1, -1, 1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, -1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 1, 0, -1, -1, 1, 0, 1, 0, -1, 0, -1, -1, -1, 0, 1, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, -2, 1, 0, -1, -1, 1, -2, 0, 0, -1, -1, 0, 1, -1, 2, 1, 0, 0, 1, 0, -1, 1, 0, 1, 1, -1, 1, 0, 0, 0, 1, 0, 0, -1, -1, 1, -1, 1, -1, -1, 1, 2, 1, 0, 1, 1, 1, -2, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, -1, -1, -1, 1, -1, 0, 0, 1, 0, 0, -2, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, 2, 1, 0, 0, 0, -1, 1, 1, 0, 0, -1, -1, -2, -1, -1, 0, 2, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, 1, 1, 1, -2, 0, 0, -1, -1, 0, 0, 0, 2, -1, -1, 0, -1, 0, -2, 0, 0, 0, 1, -1, 1, 0, -1, -1, 0, 0, -1, 2, 1, -2, -1, 1, -1, -2, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, -1, 0, 2, 1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -2, 0, -1, 0, 0, 0, -2, -1, 1, -1, 0, 0, 1, 1, 0, 0, 0, 1, -1, 0, 0, -1, -1, 2, 0, -1, 2, -1, -1, -1, 1, -1, 0, 1, 0, -1, 1, -1, 0, 1, 0, 1, 0, 1, 1, 0, 1, 1, 1, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, -1, 0, -1, -2, -1, -1, 1, -1, 0, 0, -2, 0, 0, 1, -1, 0, 0, -1, 0, 2, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, 0, -1, -2, -2, 0, 0, -1, 0, 1, 1, 0, -1, 1, 0, -1, 2, -2, -1, 1, 0, 0, -1, 0, -1, 0, 0, -1, -2, 0, 1, 0, 2, -1, 0, -1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, 1, 0, 0, -1, -2, 1, 0, 0, -1, 2, 1, 1, 1, 0, 0, 2, 2, 0, 0, -1, -2, 1, -1, 0, 1, 0, -2, 0, 1, 0, 0, -2, 0, -1, 1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, 1, -1, 0, 1, 0, 2, 1, 0, -2, 1, 0, 1, 0, -1, 1, 2, 0, 0, -1, 1, 0, 0, -1, 0, -1, 1, -1, 2, 0, -1, 0, 1, 1, 1, 0, -1, -1, 1, 0, 0, -1, 1, 0, 1, 0, 0, 2, -1, 0, 0, -1, 1, 1, 0, 0, 0, -1, 1, 2, 0, -1, -1, 1, -1, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 1, -2, 1, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, -1, 0, 2, 1, 0, -1, 0, 0, 0, -1, 2, -1, -1, 1, 0, -1, -1, 0, 0, -1, -1, -1, 1, -1, 1, 0, -1, -1, 1, -1, 0, -1, 1, 0, -1, 0, 1, 0, 0, 0, 0, -2, -1, 1, -1, 1, -1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, -1, 1, 0, -1, 0, -1, 0, -2, -1, -1, 0, 1, 0, 0, 0, 1, -1, -1, 0, 0, 2, 0, 0, 1, 1, 0, 0, -1, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, 2, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 2, 1, -1, 0, 1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 1, -1, 2, 1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 1, 0, -1, 0, 0, 1, -1, 1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, -1, -2, 0, -1, 0, -1, -1, 0, 1, 2, 0, 1, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, -2, 0, 1, 1, 1, -1, 0, 0, 1, -1, -1, 0, 1, -1, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, -1, 1, 1, -1, 0, 1, 0, 0, 0, -1, 0, 1, 0, -1, 1, -1, 1, 0, 2, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, 0, 0, 1, -2, -1, 0, 0, 0, 0, 1, -1, -2, -1, 1, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, 1, 0, 0, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, 1, 1, -1, 0, 1, 0, -1, 0, 0, 1, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, -1, 1, -1, 0, 1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, -1, 1, 1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, -2, -1, 1, 1, 0, 1, 0, 1, 0, 1, 1, -1, 1, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, 1, 2, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 1, 2, -1, 1, -2, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 1, -1, 0, 0, 1, 0, 0, 1, 0, -2, -1, 0, 0, 0, 2, 0, 1, 0, 0, 1, -1, -2, -1, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, 1, 0, 1, -1, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 0, -1, -1, 1, 1, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 1, 0, 0, 0, 1, 1, 1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, -1, 0, 0, 1, 0, 1, -1, 0, 1, 0, 0, 1, 0, -1, 0, -2, 1, 1, 0, 1, 0, 0, 1, -1, -2, 1, 1, 1, 0, 0, 0, -1, 2, -2, 0, 0, 0, 1, 0, -1, 0, 0, 1, -1, -1, 1, 1, 0, 1, 0, -1, 0, 1, 1, 0, 1, 0, -1, -1, -1, 0, 0, 1, -1, 1, 1, 0, 1, 1, 1, 0, -2, -1, -1, 1, 0, 0, 0, -1, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, -1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 1, 1, 0, -1, 0, 0, 1, 0, -1, 2, -1, 1, 0, 1, 0, -1, -1, 0, 0, 1, 3, 5, 1, 5, 5, 2, 3, 3, 0, 1, 0, 0, -1, -1, 1, 0, 1, -1, 0, 0, -3, -1, 0, -1, -1, -2, -2, -3, -5, 2, 4, 2, 2, 2, 4, 2, 3, 4, 3, 1, 4, 0, 1, 0, 1, 0, 0, 2, 3, 2, 0, 2, 2, 0, 0, -1, 0, 0, -5, 2, 2, 1, 1, 3, 2, 3, 1, 5, 2, 1, 2, 3, 2, 1, 5, 3, 2, 4, 5, 3, 4, 1, 2, 0, 0, 0, 0, -1, -1, 0, 1, 4, 3, 2, 0, 3, 2, 3, 3, 2, 4, 3, 3, 3, 6, 7, 4, 7, 7, 5, 7, 6, 2, 3, 2, 1, 1, 0, -2, 0, 1, 4, 4, 5, 1, 4, 3, 6, 2, 1, 4, 3, 4, 5, 4, 5, 5, 7, 6, 5, 7, 5, 4, 1, 1, 1, 2, 0, 0, 0, 4, 4, 4, 1, 0, 0, 3, 4, 3, 4, 4, 5, 4, 5, 7, 7, 4, 5, 7, 8, 5, 7, 1, 1, 4, 2, 0, 0, 0, 1, 3, 0, 2, 0, 0, 2, 4, 2, 3, 3, 2, 6, 6, 6, 7, 7, 7, 7, 6, 5, 6, 4, 3, 2, 4, 4, 3, -1, -3, 1, 2, 1, 0, -2, -1, 2, 2, 2, 3, 5, 5, 5, 7, 6, 10, 6, 4, 3, 6, 3, 3, 5, 3, 1, 3, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 2, 3, 2, 2, 7, 7, 5, 8, 7, 3, 5, 3, 5, 3, 1, 3, 1, 2, 2, 2, 1, 0, 0, -4, 2, 2, 2, 1, 0, -1, 1, 2, 5, 5, 7, 4, 3, 6, 5, 4, 0, 0, 3, 1, 3, 2, 2, 0, 1, 1, 1, 0, 0, -3, 0, 3, 2, 3, 0, 0, 2, 0, 0, 2, 5, 5, 4, 0, 0, -1, 0, -1, 1, 0, 3, 2, 1, 2, 2, -1, -1, 0, -1, -4, 3, 3, 3, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -4, -3, -1, 0, 0, 0, 1, 0, -1, 1, 0, -1, -2, -7, 2, 1, 4, 1, 0, 0, 2, 0, -2, -2, -3, -3, -3, -2, -2, -3, -5, -4, -4, -4, 0, 0, 0, 0, 0, 0, 0, -2, -4, -7, 3, 0, 1, 0, 0, 0, -1, -1, -2, -3, -5, -6, -5, -4, -3, -2, -5, -3, -5, -4, -2, 0, 0, 2, 1, 1, 0, -3, -4, -7, 3, 1, 0, 0, -1, -2, -2, 0, -1, -4, -8, -6, -7, -6, -6, -5, -3, -3, -7, -6, -2, -1, 0, 0, 1, 0, 0, -1, -5, -9, 1, 0, 0, -1, -1, 0, 0, -3, -4, -6, -7, -5, -8, -6, -4, -4, -3, -1, -3, -4, -3, 0, -1, -1, 0, 0, -1, -2, -5, -9, 0, 1, -2, 0, -1, 2, 0, -1, -1, -4, -5, -6, -9, -7, -6, -4, -1, -4, -4, -2, -4, -2, -2, 0, 1, 0, 0, -4, -5, -8, 0, 1, 1, -2, 1, 2, 1, 0, 0, -2, -4, -5, -5, -5, -5, -4, -3, -3, -3, -2, 0, 1, 1, 1, 0, 1, -2, -5, -6, -10, 0, 3, 2, 2, 2, 1, -1, 0, 0, 0, 0, -5, -3, -6, -5, -3, -4, 0, -2, 0, 3, 2, 1, 1, 1, 0, 1, -2, -3, -6, 2, 1, 0, 0, -2, 0, 0, 1, 0, 2, 1, -1, -2, 0, -1, -2, -1, -3, 0, 3, 3, 3, 6, 4, 2, 3, 1, 0, 0, -5, 2, 3, 0, 1, -3, -1, -1, 0, 1, 4, 3, 3, 4, 4, -1, 0, 0, -1, -2, 4, 4, 8, 4, 3, 1, 2, 2, 3, -1, -6, 0, 0, -1, -1, -2, -3, 0, 0, 2, 4, 2, 3, 7, 5, 4, -1, -1, -1, 2, 2, 7, 5, 4, 2, 0, 3, 5, 1, -1, -4, -2, 0, 1, 0, 0, -1, 0, 0, 0, 4, 4, 4, 4, 5, 2, 4, 0, 0, 2, 6, 7, 4, 5, 4, 1, 2, 5, 3, 0, -3, -1, 1, 0, 0, 2, 0, 0, 2, 0, 1, 5, 4, 5, 3, 4, 3, 0, 4, 5, 5, 5, 7, 4, 1, 3, 5, 3, 3, 1, -3, -1, 0, 2, 2, 0, 0, 2, 3, 2, 3, 3, 2, 6, 2, 6, 4, 4, 4, 8, 5, 6, 5, 5, 2, 0, 3, 4, 3, 1, -1, -1, 2, 1, 0, 0, 3, 2, 1, 3, 2, 5, 4, 5, 6, 5, 5, 7, 7, 4, 7, 6, 2, 4, 4, 3, 3, 2, 3, -1, -2, 0, 2, 2, 1, 0, 3, 2, 1, 4, 1, 2, 4, 5, 4, 5, 5, 6, 5, 3, 5, 3, 5, 3, 4, 1, 3, 4, 0, -1, -2, 2, 0, 1, 2, 2, 2, 3, 3, 2, 1, 1, 3, 3, 2, 4, 5, 5, 5, 3, 5, 3, 5, 6, 4, 2, 2, 2, 0, -1, -1, 3, 2, 1, 1, 3, 5, 7, 3, 2, 3, 1, 2, 3, 2, 0, 3, 5, 2, 5, 3, 4, 5, 4, 4, 2, 1, -2, 0, 0, -3, 2, 4, 2, 4, 4, 4, 5, 5, 5, 3, 2, 4, 0, 1, -1, 1, 3, 2, 0, 4, 4, 2, 1, 2, 2, 0, -2, -3, -3, -2, -3, -2, -1, 0, -1, 0, -2, -2, 0, -1, 0, -2, 0, 0, 0, -2, -1, -2, 0, -1, 0, -1, 0, 0, 0, 0, -2, -1, -1, 0, -2, -2, 0, 0, 0, -1, -1, 1, -1, 0, -1, 0, 1, -1, 0, -2, -1, -1, 0, 0, -1, -2, -1, 0, -1, -2, -1, 0, 0, -1, -1, 0, -2, -2, -1, 0, 0, 0, 1, -1, 0, 1, 0, -1, 1, 0, 2, 1, 2, 0, 1, 0, 0, 2, 0, -1, 1, 1, -2, 0, 0, 0, -2, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 0, -1, -1, 0, 0, 0, 0, 0, 2, 0, -1, 1, 1, -2, -1, -1, -2, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 2, 1, 2, 0, 1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -2, -2, -2, 0, -1, 0, 0, 0, 1, 2, 1, 1, 2, 2, 0, 3, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -3, 0, 0, 0, -2, 1, 0, -1, 0, 0, 2, 1, 2, 2, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 2, 2, 0, 2, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, -2, -1, -2, -3, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 2, 2, 0, 0, 0, -1, 1, 0, 1, 1, 1, 0, -1, 1, 1, 1, 0, 0, -1, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 1, 1, -1, 0, -2, 1, 0, -1, 0, 1, -1, -1, 2, 0, 0, 2, 0, 1, 1, -1, 0, -2, -1, -2, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, -2, -2, 0, 0, -2, -1, 0, -1, -1, 0, 1, 1, 0, 1, 1, 0, 0, -2, -2, -2, 0, 1, -1, 1, 0, 2, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 1, -2, -2, 0, -1, 0, -1, -1, -2, 0, -1, 0, -2, -2, -2, 0, 1, 2, 0, -1, 0, 0, 0, 0, -1, 1, -1, 0, -2, 1, 1, -1, 0, -2, 0, -2, 0, -2, 0, -2, 0, -1, 0, -3, -1, 0, -1, 0, -1, 0, -2, 0, -2, 0, 0, -1, -1, 0, 0, 0, 1, 0, -2, 0, -1, -2, -1, 0, -2, -1, 0, -3, -1, -1, -1, 0, -2, 0, -1, -2, 0, -2, -3, 0, 0, 1, -1, 0, 0, 0, 1, -1, -2, -2, 0, 0, -2, -2, 0, -1, 0, 0, -3, -3, 0, -1, 0, 1, 0, 0, -1, 0, -3, -2, -2, -2, 1, 0, -1, 0, 0, 0, 0, 0, -2, 0, -2, -3, 0, -1, -1, -2, 0, -2, 0, 0, 0, 1, -1, 0, -2, -1, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, 0, -3, -2, 0, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, -3, -1, -1, -1, 0, 1, 2, 0, 1, 0, -1, -2, 0, -1, -1, 0, 0, -1, -2, -1, -1, -1, 1, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -2, 0, -2, 0, -1, 0, 0, 1, -2, -2, 0, 0, 0, -1, 0, -2, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, -2, -3, -1, 0, 1, -1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 2, 1, -2, 1, 0, -1, 0, 2, 2, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, -1, -3, -3, -1, 1, 0, 0, 2, 3, 0, 3, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, -2, 0, 2, 0, 1, 3, 0, 0, 2, -1, -2, 0, 0, 0, 0, 2, 0, 0, -1, -1, 1, 0, 1, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, 0, -1, 2, 1, 1, -1, 1, -2, 0, 0, 1, 1, 0, 1, 1, 1, 2, 1, -1, 1, -2, 0, -1, -2, 0, -1, -1, 0, 0, 1, 1, 0, 1, 0, -1, 2, -1, 0, 0, 2, 2, 0, 2, 1, 1, 0, 1, -1, 1, -1, 1, -3, -1, 0, -2, -1, -2, -1, -1, -1, -1, -1, 0, 2, 2, 0, 1, 0, 0, 0, 0, 1, -1, 1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -2, 0, -2, -2, 1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 2, 1, 1, 0, 2, 0, 2, -1, -1, 0, 1, -2, -2, -1, 0, -1, 0, 0, -1, -1, -1, 0, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 1, -1, 0, 0, 1, 0, -1, 0, -1, -1, 1, -1, 2, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 1, -1, 0, 1, -1, 0, -1, 1, -2, 0, -1, -3, -1, 0, 0, 0, 0, -1, 1, -1, 0, 0, 0, 0, -1, -2, -2, 0, -1, 0, 0, 0, 0, 2, -2, 0, -1, 0, 1, -2, -2, 0, 0, -1, -1, 1, 0, 2, 1, 1, -1, -2, -2, 0, -3, 0, -1, 0, 0, 0, -2, -2, -4, 0, -2, -2, -2, 0, -2, -6, -6, -1, -1, 1, 0, 1, 0, 1, 2, 0, 0, 1, -1, 0, -2, -2, 0, 2, 2, 2, 1, 1, 0, 0, 0, 1, 0, 2, 1, 0, -6, -6, -3, -2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, 2, 1, 3, 1, 5, 1, 2, 2, 0, -1, 2, 1, 0, -4, -5, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 0, 0, 1, 2, 3, 5, 4, 3, 2, 3, 3, 1, 1, 1, -1, -1, -4, -4, 0, 0, -3, -1, 0, 1, 0, 1, -1, 0, 0, 2, 2, 2, 3, 3, 5, 5, 4, 5, 4, 3, 1, 2, 0, 0, 0, -2, -5, -2, 0, -2, -3, -5, -4, -1, 0, -1, 0, 0, 2, 2, 4, 3, 3, 2, 3, 2, 4, 3, 3, 1, 1, 3, 0, 0, -1, -4, -2, -2, -3, -2, -7, -5, -3, -2, -1, -1, 0, 1, 2, 3, 3, 4, 5, 1, 2, 2, 3, 1, 4, 1, 0, 2, 0, 3, 1, -1, -7, -5, -2, -6, -3, -5, -3, 0, -1, 2, 2, 4, 4, 2, 5, 4, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 2, 0, -2, -3, -5, -5, -1, -3, -3, -5, -1, 1, 0, 1, 3, 3, 0, 0, 1, 1, -2, -3, -1, 0, -2, 0, 0, -1, 0, 1, 0, -1, 0, -4, -2, -3, 0, -2, -2, -3, -1, -1, -1, 1, 0, 0, 1, -1, 0, -2, -6, -5, -6, -4, 0, -1, 0, -1, -1, 0, -1, 0, -2, -6, -5, 0, 1, -2, -1, -1, -1, -3, -3, -2, -1, -3, -4, -4, -5, -5, -8, -9, -5, -5, -1, 1, 1, 0, 0, -1, 0, -2, -1, -7, 0, 0, -1, -1, -1, 0, -3, -3, -5, -5, -6, -5, -6, -4, -6, -6, -9, -6, -7, -7, -3, -4, 0, -1, 1, 0, 1, -1, -2, -9, -3, -1, -2, -1, -3, -2, -2, -3, -4, -4, -5, -9, -10, -10, -6, -7, -8, -8, -10, -11, -7, -6, -1, 0, 2, 0, -1, -2, -5, -8, -4, -1, -1, -4, -4, -3, -3, -3, -5, -8, -6, -11, -10, -7, -6, -6, -8, -7, -9, -10, -9, -5, -1, -2, -1, 1, 0, 0, -4, -6, -3, -1, 0, -1, -3, -2, -3, -1, -6, -6, -10, -10, -12, -9, -11, -9, -4, -6, -8, -8, -8, -7, -4, 0, 0, 0, 0, 0, -1, -10, -4, -3, -3, -1, -4, 0, 0, -2, -1, -7, -6, -10, -12, -13, -12, -9, -9, -8, -5, -9, -8, -6, -3, -3, 0, -2, -3, -1, -4, -11, -3, -2, 0, -3, 0, 1, 3, 0, -3, -4, -8, -9, -10, -11, -10, -8, -6, -4, -4, -7, -6, -2, -4, -1, -1, -3, 0, -4, -4, -8, -4, -1, -2, 0, -1, 0, 2, 0, -1, -4, -4, -6, -8, -10, -9, -8, -7, -7, -4, -2, -3, 0, 0, 0, 0, 0, -1, -3, -4, -8, -5, -1, 0, 0, 0, -2, -1, -2, -1, -3, -4, -1, -2, -7, -6, -8, -7, -4, -3, -2, 2, 4, 3, 2, 0, 2, 0, 0, -1, -5, -2, -2, 1, -2, -4, -3, -5, 0, 1, 0, 0, 0, 0, 0, -3, -4, -6, -6, -6, -1, 2, 6, 4, 3, 0, 2, 2, 0, 0, -4, -4, -1, -2, -4, -5, -6, -7, 0, -1, 0, 1, 3, 4, 4, 3, 0, -3, -6, -5, -2, 0, 5, 4, 0, 1, 0, 3, 1, 0, -3, -6, -3, -5, -5, -5, -3, -3, -1, 0, 0, 4, 2, 5, 3, 0, 0, -2, -2, -3, 0, 3, 3, 2, 0, 0, 3, 4, 2, 0, -2, -6, -5, -5, 0, -5, -2, -3, -1, 1, 2, 3, 3, 5, 2, 3, 0, -1, 1, 1, 5, 3, 3, 2, 2, 1, 1, 4, 2, 0, -4, -4, -6, -2, 0, 0, -3, -2, -1, -1, 0, 2, 3, 3, 3, 3, 0, 2, 1, 4, 5, 5, 3, 3, 0, 0, 3, 3, 3, 0, -3, -7, -3, -1, 0, -4, -3, -1, -3, -2, -1, 0, 2, 2, 3, 1, 1, 2, 2, 4, 2, 3, 4, 1, 1, 0, 1, 0, 2, -1, -4, -5, -3, -3, -1, -1, -1, -3, -1, -3, 0, 0, -1, -1, 1, 0, 3, 3, 3, 0, 2, 2, 3, 3, 3, 1, 2, 0, -1, -2, -2, -5, -1, -3, -2, -1, -2, 0, 1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 2, 1, 2, 1, 4, 1, 2, -1, 0, -3, -2, -2, 0, 0, 0, 0, 0, 1, 0, 2, 0, -1, 1, 1, -3, -3, -1, 0, 1, 0, 0, 0, 3, 3, 1, 2, 0, -1, -3, -3, -5, -3, -2, -1, 2, 1, 2, 4, 4, 2, -1, -1, 0, -3, -4, -1, -3, -2, 0, 0, -2, -1, 0, 3, 0, 1, -3, -3, -2, -6, -3, -4, -2, 0, -1, 0, 1, 2, 2, 0, -1, -2, -1, -5, -2, -7, -4, -3, -3, -2, -1, -2, 0, -3, -1, -2, -5, -6, -6, -6, -8, -4, -2, -4, -2, -3, -1, -3, -1, -4, -3, -4, -4, -3, -6, -5, -1, -2, -2, -3, -2, -5, -2, -3, 0, 0, -5, -5, -3, -2, -5, -1, -1, -2, -3, -3, -3, -2, -3, -3, -3, -3, 0, -2, -1, -2, -2, -4, -2, -3, -1, -2, -2, -3, 0, -1, -1, 0, -4, -5, -6, -1, -2, -3, -2, -2, -1, -1, 0, -1, -1, -4, -1, -2, -1, 0, -2, -4, -2, -2, -3, -2, -3, -1, -3, -3, -1, -2, -4, -4, -5, -3, -2, -2, -1, -4, -4, -3, 0, 0, 0, -2, 0, 0, 0, -2, 0, 0, 0, -1, 0, 0, 0, 0, -3, -3, 0, -1, -1, -2, -1, -4, -3, -2, -2, -1, 0, 0, 0, -3, -3, -3, -2, -3, -2, -3, -2, 0, -1, -2, 0, 0, -3, -1, -3, -2, 0, -2, 0, -3, -2, -1, -1, -1, -1, 0, -2, -1, 0, -1, -1, -1, -2, 1, 0, -1, -1, -2, 0, 0, 0, -1, -2, -1, -1, -2, -1, -1, -3, -3, -1, -1, 0, -3, -3, -1, -2, 0, -1, -1, -1, 0, -1, 0, 0, 0, -2, 0, 0, 1, 0, 0, -1, -2, -1, -3, -2, 0, -2, -3, -1, -2, -1, -3, -3, -3, -1, 0, -2, -3, -1, 0, -1, 1, 0, 0, -2, -1, 1, -2, 0, -1, 0, -1, 0, -1, 1, -2, 1, 0, 0, 0, -2, -4, -2, -3, -3, 1, -1, -2, 0, 0, 0, 1, -1, 1, -1, 1, 0, 0, 0, 0, -2, 1, -3, -1, -1, 0, 1, -2, -3, -1, -3, -3, -4, -4, -2, 0, 0, 0, 1, 0, 2, 0, 1, 0, -2, -2, 0, 0, 0, -3, -1, -1, 0, 0, -1, -2, -1, 0, 0, -3, -1, -3, -4, -4, -3, 0, 0, 1, 0, 0, 1, -2, 1, 0, 1, 0, 0, -1, -2, -1, -3, -2, 0, -1, 1, 0, 0, 0, 0, 0, -1, -3, -3, -1, 0, 0, -4, 0, 1, 0, -1, -2, 0, -2, 0, 0, -2, 0, 0, -2, 0, -1, 0, 0, -2, 0, -1, -1, -1, -3, -1, 0, -2, -1, -2, -1, -2, 0, 0, 0, 1, 0, 0, 0, -2, -2, 0, -2, -1, -1, -2, 0, -1, -1, 0, -1, 0, -1, -2, -1, 0, -3, -3, 0, -1, -1, -2, 0, -1, -3, 0, 0, -1, -1, -2, 0, -1, -4, -2, -1, -1, -2, 0, -1, -1, 0, 0, -1, -3, -2, -2, -2, -1, -3, 0, -1, -1, -1, 0, -3, -3, -3, 0, -1, -2, -1, -4, -5, -2, -1, 0, -2, 0, 0, 0, -1, -2, -4, -4, 0, -3, -3, -3, 0, 0, -3, -2, -3, -4, -4, -3, -3, -3, -2, 0, -2, 0, -2, -4, -2, -3, 0, 0, -1, 0, -1, 0, -2, -2, -3, -1, -2, -3, 1, -1, -3, -4, -1, 0, -3, -1, -4, -4, -2, -3, 0, -2, -4, -3, -5, -3, -4, 0, -2, -2, 0, -1, 0, -5, 0, 0, -4, 0, -1, 0, 0, -2, 0, 0, 0, -4, -4, -1, 0, 0, -3, -1, -3, -2, -4, -1, -1, -3, -3, -2, 0, -2, -3, -6, -3, 0, -3, -1, -2, 2, 0, -3, -4, -2, -2, -4, -1, -4, 0, -1, -1, -1, -2, -1, -1, -3, -4, -3, -3, 0, 0, -2, -1, -6, -3, 0, 0, -1, 0, 0, 1, -3, -3, 0, -2, -4, -3, -5, -3, -1, -2, -2, 1, -2, 0, -3, 0, -2, 0, 0, -2, -2, -1, -3, -1, 0, -1, -3, -2, 0, 0, 1, 0, -1, 0, -3, -2, -1, -3, -4, -4, -1, -1, 0, 1, 0, -2, 0, 0, 0, 0, -1, -4, -2, 0, -3, -3, -3, -4, -3, 0, -2, 0, 1, -2, -2, 0, -2, -2, -1, -4, -5, -1, -2, -1, -1, -2, -3, 0, 1, -2, -2, -3, -4, -3, 0, -2, -3, -4, -2, -1, -2, 0, -1, -1, 0, 0, -2, -2, -3, -2, -1, -3, 0, 0, 0, -3, -3, -2, 0, 0, -2, -1, -3, 0, 0, -1, -1, -1, -4, -3, -2, -2, -2, 0, -1, -1, -2, 0, -3, -2, -2, -2, 0, 0, 0, -1, -2, -1, 0, 1, -2, -1, 0, 0, -1, 0, -3, -3, -2, 0, -2, -1, -2, -1, -3, 0, -1, -2, -1, -1, -2, 0, 0, 2, -2, -2, -2, -1, 1, 0, -1, 0, -2, -1, -3, -3, -2, -3, -2, -2, -1, -2, -2, 0, 0, -1, -2, -2, -1, -2, 0, -2, 0, 0, -2, -2, 0, -1, 1, 0, -1, -2, -3, -1, -1, -1, -2, -2, 0, -4, -2, -3, -2, -1, -3, -1, -1, -1, -2, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, -1, -1, -4, -2, -1, -2, -2, -3, -4, -2, -1, -1, -1, 0, 0, 0, 0, -1, -3, 0, 0, -1, -1, -1, -2, 0, -2, -2, -1, 0, -3, -3, -2, -3, -2, -2, 0, -1, -4, -3, 0, 0, -1, -1, 0, 0, -2, -1, 0, 0, -1, 0, 0, 0, -1, -3, 0, 0, -2, -3, 0, -1, 0, -3, -1, 0, 0, -1, -1, -1, -2, -3, -4, -3, -1, -3, 0, 0, -3, 0, 1, 1, 1, 0, 0, -2, -3, 0, -3, 0, 1, 0, -1, -1, 1, 2, 1, -1, 0, 0, 2, 0, 0, -1, -1, 0, 1, 1, 0, -1, 0, 1, 0, -1, 0, -1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 1, -1, 0, -1, -1, 1, 0, 0, 1, 0, -1, -1, 0, 1, 0, 1, -1, 1, 0, 1, 2, -1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -2, 0, 0, 2, -1, 0, 0, -1, -1, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, -1, -1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 1, 1, -1, 1, 0, -1, -1, 1, 0, -1, -1, 0, 0, 1, -1, -1, 0, 0, 0, -1, 1, -1, 0, -1, 0, 0, -1, 1, 0, 0, 0, 0, 2, 1, -1, 1, 0, 1, -1, -1, -1, 1, 0, 0, -1, 1, -1, -1, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, -2, 0, 0, 0, -1, -1, 0, 1, 2, 1, 0, 0, 1, 1, -2, 0, 0, 0, -1, 0, -1, 1, -1, 0, -1, -1, -1, 1, 1, 0, -1, 1, -1, -1, -1, 1, 1, 1, 0, 1, 0, -1, 1, 0, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, -1, 0, 0, -2, 2, -1, -1, -1, -1, 0, 1, -1, 0, 0, 1, 1, 0, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 1, -1, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, -1, 1, 1, 0, 0, -1, 1, 0, 1, 0, 0, 0, 1, -1, 0, 2, 0, 0, 0, 0, -1, -2, -1, -2, 1, -1, 0, 1, 1, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 1, -1, 0, -1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, -2, 1, 0, -1, 1, 0, 0, 1, 1, -1, -1, 1, 0, 0, 1, -1, -1, 0, 1, 1, -1, 1, 1, -1, 0, 0, 0, -1, 1, 1, 0, -1, 2, 1, 0, 1, -1, 1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, -1, -1, 1, 1, 1, -1, -1, 0, 0, -1, 2, -1, -1, 1, 1, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, -1, 0, 1, 1, -2, 0, 0, -2, 0, 0, 0, 1, 0, -1, 1, 0, 1, 1, -2, 0, 0, 1, 0, 0, 1, -1, 0, 0, -1, 0, -2, 1, -1, 0, -1, 1, 0, -1, -2, 0, 1, -1, 1, 0, -1, -2, -1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 1, 0, -2, 0, 0, 1, 0, -1, 0, 1, 0, -1, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, -1, 0, 1, 0, 1, 0, -1, -1, 0, 0, -1, 1, 0, 1, 0, 0, 0, 1, 2, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 0, 1, 0, -1, 1, 0, 1, 0, -1, 0, 1, 0, -1, 1, 2, 0, -1, 0, 0, 0, 1, -1, 0, 1, 1, -2, -1, 1, 0, -1, 0, 0, -1, 0, -1, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, -1, 0, -1, 1, 0, 0, 0, 0, -2, -2, 1, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, -1, 1, 0, -1, 0, -1, 1, 1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, -1, 1, 1, -1, 0, 2, 1, 1, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, -1, 1, 1, -1, -1, 2, -1, -2, 0, 1, 1, 1, 1, 1, 0, -1, -1, -1, 0, 1, 0, -1, 1, 0, 2, 0, 0, -1, 0, 1, -1, -1, -2, 0, 1, 0, 1, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, 0, -1, -2, -1, 0, 0, 0, -1, 2, 0, 1, -1, 0, 0, 0, 1, -1, 1, 0, 0, -1, 0, 1, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, -1, 2, -1, 2, -1, -1, 0, -1, 1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 1, 0, 1, -1, 1, 0, 1, -1, 1, 0, 0, 0, 0, 1, 1, -1, 0, 0, -2, 0, 1, 0, 1, -1, -1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 1, -1, 1, 1, -1, 1, -2, 1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 2, 0, -1,
    -- filter=0 channel=3
    1, 1, 3, 2, 0, 2, 3, 3, 0, 0, 1, 3, 0, 2, 3, 1, 4, 2, 3, 2, 3, 3, 3, 1, 1, 1, 4, 4, 4, 1, 1, 3, 2, 3, 0, 0, 2, 0, 0, 2, 1, 3, 0, 0, 4, 0, 3, 3, 3, 0, 0, 2, 4, 3, 0, 3, 3, 4, 4, 1, 0, 1, 1, 2, 1, 2, 0, 2, 0, 2, 3, 0, 3, 0, 0, 2, 2, 0, 2, 2, 3, 1, 2, 1, 2, 2, 2, 1, 1, 0, 1, 2, 1, 1, 0, 2, 1, 0, 1, 0, 3, 2, 4, 2, 1, 1, 2, 3, 2, 2, 3, 1, 0, 2, 2, 1, 0, 2, 2, 1, 1, 3, 1, 2, 0, 1, 3, 0, 3, 0, 0, 0, 2, 2, 0, 3, 2, 0, 2, 3, 0, 1, 4, 1, 1, 0, 0, 0, 4, 2, 1, 0, 2, 2, 1, 0, 1, 0, 2, 2, 4, 2, 0, 1, 1, 2, 3, 3, 2, 0, 2, 3, 2, 3, 1, 1, 0, 3, 3, 3, 2, 1, 0, 3, 0, 2, 0, 0, 0, 1, 0, 2, 3, 1, 3, 3, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 3, 2, 2, 3, 2, 2, 2, 0, 1, 1, 0, -1, 0, 1, 1, 3, 3, 2, 1, 0, 2, 1, 2, 1, 1, 2, 0, 0, 3, 3, 1, 2, 1, 1, 1, 2, 0, 3, 3, 3, 0, 0, 4, 3, 2, 0, 2, 0, 2, 3, 2, 1, 2, 2, 0, 0, 0, 2, 1, 3, 3, 2, 4, 3, 0, 1, 2, 0, 0, 2, 2, 1, 2, 4, 2, 2, 0, 0, 0, 2, 0, 2, 0, 0, 0, 2, 1, 2, 1, 3, 2, 3, 0, 0, 2, 2, 0, 1, 0, 3, 0, 3, 3, 2, 1, 2, 0, 1, 0, 2, 2, 1, 1, 0, 2, 1, 2, 0, 0, 2, 1, 0, 0, 3, 1, 0, 2, 3, 4, 1, 0, 4, 2, 1, 3, 0, 0, 2, 1, -1, 1, 0, 2, 0, 2, 0, 0, 0, 0, 1, 1, 1, 2, 1, 0, 3, 3, 2, 1, 3, 3, 2, 2, 1, 0, 1, -1, 0, 1, 0, 1, 0, 1, 0, 1, 2, 2, 1, 0, 1, 1, 0, 2, 0, 2, 2, 3, 1, 5, 2, 3, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 0, 2, 3, 3, 0, 3, 4, 3, 1, 2, 1, 2, 2, 2, 2, 2, 2, 0, -1, 2, 1, 0, 1, 0, -1, -1, 0, 2, 2, 1, 0, 0, 2, 1, 1, 2, 1, 1, 1, 3, 3, 2, 2, 3, 0, 1, 0, 0, 0, 0, 1, -1, 2, -1, 0, 1, 1, 2, 0, 2, 2, 0, 0, 0, 0, 2, 3, 2, 4, 2, 3, 2, 1, 3, 1, 1, 0, 0, -1, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 2, 1, 2, 0, 2, 0, 1, 3, 1, 3, 4, 0, 3, 2, 3, 1, 3, 1, -1, 2, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 3, 2, 1, 1, 1, 3, 3, 3, 1, 2, 3, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, -1, 0, 1, 2, 0, 0, 3, 0, 1, 3, 0, 3, 3, 3, 2, 1, 0, 1, 3, 2, 0, 1, 3, 0, 0, 0, 2, 1, 0, 1, 1, 2, 0, 2, 0, 1, 2, 0, 3, 2, 2, 1, 0, 0, 3, 0, 0, 2, 0, 1, 2, 2, 2, 1, 0, 0, 0, 0, 3, 1, 1, 3, 1, 3, 3, 1, 0, 2, 1, 0, 0, 1, 2, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 2, 0, 1, 2, 0, 2, 1, 1, 0, 0, 1, 2, 2, 0, 0, 3, 1, 3, 0, 2, 3, 3, 1, 1, 2, 0, 2, 1, 3, 1, 1, 2, 0, 0, 3, 3, 3, 2, 0, 0, 0, 0, 0, 3, 1, 0, 3, 2, 1, 0, 0, 1, 0, 2, 2, 1, 3, 1, 1, 3, 2, 2, 0, 1, 3, 3, 1, 3, 1, 2, 2, 2, 0, 0, 0, 3, 0, 0, 2, 1, 2, 3, 3, 0, 2, 0, 0, 0, 3, 1, 1, 2, 1, 0, 1, 3, 2, 2, 1, 0, 0, 0, 2, 1, 0, 1, 1, 0, 2, 1, 2, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 0, 2, 1, 1, 4, 2, 2, 0, -1, 0, 1, 1, 2, 0, 1, 2, 1, 3, 1, 0, 2, 2, 0, 0, 3, 2, 1, 2, 1, 2, 2, 3, 2, 1, 2, 1, 1, 0, 0, 2, 1, 1, 2, 0, 0, 2, 0, 2, 2, 0, 1, 0, 0, 2, 0, 3, 2, 1, 3, 2, 4, 4, 3, 2, 2, 4, 2, 3, 1, 3, 3, 1, 3, 3, 0, 2, 3, 1, 2, 0, 0, 2, 2, 0, 0, 2, 3, 0, 2, 1, 4, 4, 4, 2, 2, 5, 1, 0, 0, 2, 0, 2, 0, 1, 0, 3, 2, 1, 1, 0, 1, 2, 4, 1, 1, 4, 2, 1, 4, 1, 3, 4, 4, 2, 3, 1, 5, -3, 0, 0, -3, -1, -2, 0, -1, -1, 0, 0, 0, 1, -1, 0, -2, -2, -2, -3, -3, -3, -2, 0, -2, -1, -2, 0, -2, 0, -2, -2, -1, -1, -1, -2, 0, 0, 0, 0, -2, 0, 0, 0, -1, -1, -1, -1, -2, -2, -2, -3, 0, -1, -3, 0, -3, 0, -3, -1, 0, -3, -1, -1, -2, 0, 0, 0, -2, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, -3, 0, 1, -1, 0, -1, 0, 0, 0, 0, -2, -2, -2, -4, -3, -3, -2, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, 1, -1, 0, 0, 0, -2, 0, 0, 0, -1, 0, -1, 0, 0, 1, -4, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, -2, -2, -1, 0, 0, -1, -1, 1, 0, 0, 0, 1, 1, -2, -2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, -3, -1, 1, 0, 1, -1, 0, 2, -1, -1, -2, 0, 0, 1, -1, -2, -2, 0, 0, 0, 0, 0, -1, -1, 1, -1, -2, 0, -2, 0, -2, 0, -2, 0, 1, 0, 0, -2, 0, 1, 0, -1, 0, 1, -1, -4, -1, -2, 1, 0, -2, 0, 0, 0, -2, -2, -1, -2, -1, -2, -3, -2, 0, 0, 0, 1, 1, 1, 0, 0, 2, -1, 1, 2, -2, -4, -3, -2, 0, -1, -2, 0, -1, -2, -2, -2, 0, -2, -2, 0, 0, -1, 1, 0, 2, 2, 0, 0, 0, 0, 2, 0, 3, 0, -2, -2, -1, -3, -1, -1, -2, -1, -1, 0, -1, -1, -1, -2, -1, 1, 0, 1, -1, 2, 2, 2, 1, 0, 1, 2, 0, 1, 3, 1, -2, -3, -2, 0, -3, -2, -2, -3, -1, -2, -1, -3, -2, -1, 0, 2, -1, 1, -1, 1, 0, 1, 0, 0, 0, 0, 2, 3, 1, 3, -3, -2, -2, -1, -3, -1, -4, 0, 0, -2, -3, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 3, 0, 0, 0, 0, 0, 0, 2, 4, -2, -4, -3, -4, -3, -2, -3, 0, -3, -1, -1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 0, 3, 1, 2, 2, 0, 0, 4, 2, 3, -2, -5, -1, -3, -1, -4, -3, -1, -3, -1, 0, -2, 1, 2, 1, 0, 1, 1, 1, 1, 3, 3, 0, 1, 0, 0, 1, 3, 2, 2, -2, -3, -3, -3, -3, -6, -4, -4, -4, -2, -1, -2, 0, 1, 3, 0, 3, 1, 0, 0, 1, 1, 2, 3, 1, 3, 3, 2, 3, 2, -3, -2, -5, -5, -2, -4, -2, -2, -2, -3, -2, -2, 0, 0, 2, 0, 3, 2, 3, 2, 0, 0, 0, 2, 2, 1, 3, 4, 5, 4, -4, -5, -2, -2, -3, -2, -3, -1, -1, -2, -2, 0, -1, 0, 0, 2, 3, 0, 0, 3, 0, 2, 4, 2, 4, 2, 2, 4, 5, 5, -6, -4, -4, -5, -5, -2, -2, -1, -3, -1, -1, -1, 0, 2, 0, 1, 0, 0, 3, 4, 2, 3, 2, 4, 5, 3, 3, 4, 6, 4, -4, -2, -4, -4, -2, -3, -3, -2, -3, -1, -2, 0, -1, 1, 2, 2, 0, 3, 1, 1, 0, 4, 2, 5, 1, 5, 5, 4, 1, 3, -3, -4, -5, -1, -2, -2, -1, -2, -2, -3, 0, -2, -1, 1, 2, 0, 0, 3, 0, 0, 3, 0, 1, 5, 2, 2, 5, 3, 3, 3, -4, -4, -4, -1, -1, -4, -4, -3, -2, 0, -1, 0, 1, 1, 0, 0, 3, 0, 0, 0, 2, 0, 2, 2, 3, 3, 4, 2, 3, 4, -5, -4, -3, -2, -3, -1, 0, -1, -1, -3, 0, -2, 1, 2, -1, 2, 0, -1, 1, 1, 1, 1, 2, 0, 1, 2, 3, 0, 1, 0, -3, -1, -4, -4, -1, -1, 0, -2, 0, -2, -2, 0, 2, 1, 2, 0, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 3, 2, 0, -3, -5, -2, -1, -3, -1, -1, -1, 0, 0, 0, 1, 0, -1, 1, -1, 0, 1, 2, 3, 0, 0, 2, 1, 2, 3, 2, 3, 1, 0, -3, -4, -4, -1, 0, -2, 1, 0, 1, 0, 0, 1, 0, -1, 1, -1, 2, 1, 0, 1, 0, 2, 0, 0, 1, 3, 1, 0, 0, 0, -2, -4, -3, -1, -1, 1, 1, 0, 0, 0, 1, 0, -2, 1, 0, 0, -1, 0, 1, 1, 3, 2, 1, 0, 0, 2, 0, 0, 1, 0, -1, -3, 0, 0, 1, 0, -1, 0, 0, 0, 1, 1, -1, 0, 0, 1, 1, -1, 2, -1, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, -2, -2, -2, -1, 0, -2, 0, -2, -1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, -4, -2, 0, -2, 0, 0, -1, -1, 1, 0, 0, -1, -1, 1, 1, 0, -1, 0, 2, 2, -1, 0, 0, -1, -1, -1, 2, 1, 0, -2, -4, 0, -3, 0, -2, 0, 0, -1, -2, -1, 0, 1, 2, 0, 0, 0, -2, -1, -2, 0, -1, -1, 1, 0, -1, 0, -2, -1, 0, -2, 0, -1, -2, 0, -1, 0, -2, 0, 0, 0, -1, 0, -1, 1, 0, 0, 1, -1, 0, 2, 0, -1, 0, 0, 0, -1, 0, 1, 2, 0, 0, -1, -2, 0, -1, 0, 1, 0, -1, 0, 1, 0, 1, 0, 1, 1, -1, 1, 0, 1, 2, -1, 0, 0, 1, -1, -1, 2, 1, 2, 0, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, -1, 1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 2, 1, 1, -1, 0, -1, -1, 1, 0, 1, -1, 0, 2, 0, 0, 1, 2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 1, 1, -1, 2, 2, 1, -1, 0, 0, -1, -1, -1, -1, 1, 1, 0, 1, 0, -2, 1, 0, 1, 0, 0, 1, 0, -1, -1, 2, 1, 0, 1, 0, 0, 2, 1, -1, 0, -2, -1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, -1, -1, 0, 1, 0, 1, 1, 1, 0, 0, 2, 1, 0, 0, -1, -1, 1, 1, -1, 0, -1, 1, 0, -2, -1, -2, -1, -1, -2, 0, -2, 1, -1, 1, 2, 0, 1, 0, 0, 1, 0, 0, -2, -2, -2, 0, 1, 0, -1, 0, 0, -2, 0, -1, 0, -2, -2, 0, 0, 0, -1, 1, 1, -1, -1, 0, 0, 0, 0, 0, 1, 3, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -3, 0, -2, 0, 1, -1, -1, 0, 0, 0, 2, 1, 0, 0, 1, 1, 2, 0, -2, 0, 0, 1, 1, 0, 0, 1, -1, -2, 0, -1, -2, -1, -2, 1, 0, 1, 1, 0, 0, 0, 1, 1, -1, 0, 0, 1, 0, -2, 0, 0, -2, 0, 0, -2, 0, 0, -1, -2, 0, -3, -2, 0, -1, 0, -2, 0, -1, -2, -1, 1, 0, 1, 0, 0, 1, 2, 2, -2, -1, 0, 0, 1, -2, 0, 0, 0, -1, 0, 0, 0, 0, -2, 1, -1, 0, 0, 1, 1, 1, 0, 0, 2, 0, 0, 1, 0, 1, 0, -3, -1, -1, 0, -2, -1, -1, 0, -2, -1, -3, 0, 0, -1, 0, 0, -1, 1, 1, 1, 1, -1, 0, 1, 1, 1, 0, 2, 0, 0, -1, 0, -2, 0, -2, 0, 0, -1, -2, 0, -1, 0, 1, -2, 0, -1, -1, 0, 2, 0, 0, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 0, -2, -2, -2, -1, -1, 0, 0, -2, 0, 0, 1, 0, 0, 1, 0, -1, 0, 2, 0, 0, 0, -2, 0, -2, -2, -2, -1, -2, -2, -2, 0, -3, -1, -2, 1, 0, 0, 0, 1, 1, 0, -1, 2, 0, 1, 1, 3, 0, 2, 0, 1, -1, -3, -3, 0, -1, -1, -3, -1, -2, 0, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 2, 2, -1, 2, 0, 0, 3, 2, 0, 0, -2, -2, -1, -1, 0, -1, 0, 0, -3, 0, 0, 0, 1, 0, 1, -1, 2, 0, 0, 2, 0, 0, 1, 0, 2, 0, 1, 3, 0, -3, 0, -3, 0, 0, -1, -2, -2, 0, -2, -1, 0, -1, -1, -2, -1, 0, 1, 0, -1, 1, 2, 0, 2, 2, 0, 1, 1, 3, 2, 0, -1, -2, 0, -1, 0, 0, -1, 0, 0, 0, 0, -2, -1, 0, 0, -1, 1, 0, 2, 1, 1, 0, 0, 2, 3, 0, 1, 3, 1, 0, -1, 0, 0, -3, -2, -2, -3, -3, 0, 0, 0, 0, -2, 1, 1, 2, 0, -1, 1, 0, -1, 0, 2, 0, 1, 0, 0, 3, 1, 0, -3, -2, -1, -1, 0, -2, -3, 0, 0, 0, 0, -2, 1, 1, 0, -1, 1, 0, 0, -1, 0, 1, 0, 2, 2, 1, 2, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, 0, -1, -2, 0, -1, 1, -1, 0, -1, -1, 0, -1, 0, 2, 2, 0, 0, 0, 2, 0, 0, 1, 0, -3, -1, 0, -1, 0, 0, -1, 0, 0, 0, -2, 0, 1, -1, 0, 0, 1, -1, 0, 2, 2, 1, 0, 2, 0, 2, 2, 0, 0, 0, -3, 0, -2, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 2, 2, 0, 0, 0, 3, 0, 2, 0, 0, 1, -2, -1, -1, 0, 1, 1, 0, 1, 0, 0, 1, 1, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 2, 0, 1, 0, 0, 1, 1, -1, -1, 0, -1, 1, -2, 0, 0, 2, -2, 0, 0, -1, 0, 0, -1, -2, -1, 0, 1, 2, 1, 0, 0, 2, 0, 0, 2, 0, 2, -2, -2, 0, 0, -1, -1, -1, 0, 1, 0, -1, 0, 1, 0, -1, -1, -1, 1, 2, 0, 1, 0, 2, 0, 1, 0, 1, 2, 0, 0, -2, -2, 0, -1, -1, 0, 1, 1, 1, 0, -1, 0, 0, 2, -1, 0, 1, 0, 2, 0, 0, -1, 0, 1, -1, 0, 0, 1, 0, 1, 0, -2, 0, -1, 0, -1, 0, 0, 0, 2, 0, 1, 0, 1, 1, 0, 0, 0, 2, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -2, 2, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 1, 0, 0, 0, -1, -2, 0, 1, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 1, 1, 1, -1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, -2, -1, 2, -1, -1, -1, -1, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 1, 1, -1, 0, 1, -1, 1, 1, 1, 0, -1, 0, -1, 1, -1, 1, 1, -1, 0, 1, 0, 1, 0, 1, -1, -1, 0, 0, -1, 0, 1, 1, 1, 1, 0, 1, 0, -1, 1, 2, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, -1, 1, -1, 0, 1, 0, 1, -1, -1, 1, -1, 0, 1, 1, -1, -2, 1, 1, -1, -1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 0, 0, -1, -1, 0, 2, 0, -2, -1, -2, -1, 1, 1, 1, 1, 0, -1, -2, 1, 0, 0, -2, 0, 1, 0, 1, 1, 2, 0, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, -1, 0, -1, 0, -1, 0, -1, -1, 0, -1, 1, 0, 1, 1, -1, -1, 2, 2, 1, 1, 1, 1, 1, -1, -1, 1, -1, 1, 1, 0, -1, 0, 0, 0, 1, 0, 1, 1, -1, -1, 0, 0, 0, 1, 0, 1, -2, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -2, -2, 0, -1, 0, 1, -1, 0, -2, -1, 0, -1, 1, 0, 2, 0, -1, 1, 1, 0, 0, 1, -2, 1, 0, 0, -1, -1, 0, 1, 0, -1, 0, 0, 1, -1, -1, 0, 1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, 1, 1, 1, 0, 1, 0, 1, -1, 0, -1, 1, 0, -1, 0, 2, 0, 1, 0, -1, -1, 1, -1, 0, 0, -2, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 1, -1, -1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 1, 0, 1, -1, 0, 2, 0, 0, 0, -1, 2, -1, 1, -1, 0, 0, -1, -1, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, -1, 2, 0, 0, 0, 1, -2, 0, 2, 2, -2, -1, 0, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 2, 2, 1, 0, 0, 1, 2, 0, 0, 0, 1, 0, 1, 1, -1, 0, 0, -1, 0, -1, 1, 2, 0, -1, 0, -1, -1, 0, -1, 1, 0, 0, -1, 0, -2, 1, -1, -1, 0, -1, -1, 2, 0, 1, 0, 0, 0, 0, -2, -1, -1, -1, 1, -1, 1, 0, 0, 1, -1, -1, 1, -1, 0, -1, 0, -1, 1, 1, -1, 1, -2, 0, -1, 1, 0, -2, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, -1, 2, 1, 1, 0, -1, 0, 2, 0, 0, 1, 0, -1, -1, 1, 1, 1, 0, 1, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, -1, 0, -1, 1, -1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, -1, 0, 1, -1, 0, -1, 2, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -2, -2, 1, -2, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 1, 0, -1, -1, 0, 1, 0, 2, 2, -1, 1, 0, 1, 1, 1, -1, -1, 0, 0, -1, 0, -1, 1, 0, -1, 1, 0, 0, 1, -1, 0, -2, 0, -1, 0, 0, -1, 1, 0, 2, 1, 1, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 1, 0, -1, 1, -1, -1, -1, 0, 1, 0, 0, 0, -2, 1, -1, 1, 0, -1, 0, -2, -1, -1, 1, 0, 2, 0, 1, 0, -1, 0, 1, 1, 0, -1, 1, -1, 0, -1, -1, 0, 0, 1, -1, 0, 1, 0, 0, 0, -1, 2, 1, 0, 1, -1, 1, 0, 2, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, -1, 0, 0, 2, 1, 1, 1, 0, -1, 0, 1, 1, 1, 0, 0, 1, -1, 0, 0, -1, -1, -1, 0, 1, 2, -1, 0, -1, 0, -2, 1, -1, 0, -2, 1, 1, 0, -1, 0, 1, 1, -1, 0, 1, 1, 0, 2, 0, 0, 2, 1, 1, 0, 1, -1, 2, 0, 0, 1, 0, 0, 0, 1, -1, 0, -2, 0, -2, -3, -1, -3, 0, -2, -1, 0, 0, 1, 0, 2, 0, 0, 2, 1, 0, 0, 2, 0, 0, 0, -1, 1, 1, 0, -2, -2, 1, 0, -2, -1, -3, -2, 0, 0, -1, 0, 0, 2, 3, 3, 2, 1, 0, 0, 1, 0, 3, 1, -1, 2, 1, -1, 1, -1, 0, -1, 1, -3, 0, -1, 0, 0, 0, -3, -1, -2, 2, 1, 3, 0, 3, 1, 1, 1, 2, 0, 2, 0, 3, 0, 1, 1, 0, -2, 1, 1, 0, 1, 1, -2, -2, -2, 0, 0, 0, 0, 0, 2, 1, 0, 2, 0, 0, 1, 0, 2, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, -2, -1, 0, -2, 0, 0, 0, -2, -1, 1, -1, 0, 3, 1, 0, 0, 2, 0, 2, 0, 0, 1, 0, 0, 0, 0, -2, -1, 1, 0, 0, -1, 0, -1, -1, 0, 1, 0, 1, -2, 2, 1, 2, 2, 0, 0, 2, 3, 2, 1, 3, 0, 1, 0, -1, -2, 0, -2, 0, 0, -1, -1, 2, 1, 0, 0, 0, -2, 0, 0, 1, 2, 2, 0, 0, 1, 0, 1, 3, 2, 0, 0, 0, 1, 0, -2, 0, -1, -1, 0, -1, -1, 0, 0, 2, -1, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 3, 1, 0, 0, -1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 2, 2, -1, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 1, 0, 1, 1, 0, -1, 0, -1, 2, 1, 1, 1, 1, -1, 1, 0, 1, 0, 1, -1, 0, 1, -1, 1, -1, 0, 0, 0, -1, 0, 1, 1, 0, 2, 0, 0, 1, 0, 0, 2, 1, 2, 0, -1, 2, 0, 1, -1, 1, 1, 0, 0, 0, 0, 0, 2, 0, -1, 0, 2, 0, 2, 0, 0, 1, 0, 0, 3, -1, 0, -1, 2, 1, -1, 2, -1, -2, 1, 1, -1, 1, 0, 2, -1, 0, 0, 0, 0, 0, 1, 2, 2, 1, 1, 0, 2, 0, -1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 0, 2, 1, 1, 0, 2, 1, 0, 3, 1, 2, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, 1, -1, -1, 0, 0, -2, -1, -1, 2, 2, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 1, 2, 3, 1, 3, 0, 0, -1, 0, 0, -1, -2, 0, 0, 1, 0, 0, -2, 0, 2, 0, 0, 0, 1, 0, -1, 0, 3, 0, 3, 0, 0, 3, 2, 2, 2, 2, 2, -1, 1, 0, -1, -1, 0, -1, -1, -1, 0, -1, 1, 0, 1, 0, -1, 2, -1, 0, 3, 3, 3, 3, 1, 2, 3, 0, 0, 1, 0, 0, 0, -1, 1, -2, -2, -2, 0, 0, 1, 0, 0, 1, 1, -1, 1, 2, 1, 1, 0, 3, 2, 1, 4, 2, 2, 0, 1, 0, 1, 2, 1, 1, 0, 0, -2, -1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 3, 2, 4, 4, 0, 4, 2, 0, 1, 0, 1, 0, 0, 0, 1, -1, -2, -1, 0, -2, -1, -1, 0, 0, 0, 1, 0, -1, 1, 2, 0, 0, 2, 3, 1, 0, 3, 2, 1, 1, 0, 0, 1, 2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 2, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 2, 2, 0, 1, 2, 1, 0, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, -1, 1, 2, 2, 2, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 0, 0, -1, 1, 0, 1, -1, 1, 0, 0, 0, 0, -1, 0, 2, 0, 1, -1, 1, 2, 0, 2, 2, 0, 2, 0, 0, 0, 1, 1, 0, 0, 0, -1, 2, 0, 0, 1, 2, 1, 0, -1, 0, 3, 0, 0, -1, -1, 1, 2, 1, 0, 3, 3, 2, 3, 2, 2, 2, 1, 0, 0, -1, 0, -1, 0, 2, 1, 0, -2, 1, 0, 2, 0, 0, 0, 0, 1, 1, 3, 1, 3, 3, 1, 1, 1, 0, 0, 0, 0, 2, 0, 2, 0, 0, -1, 1, 0, 0, 0, -2, 0, 0, 0, 2, 0, 0, 0, 3, 4, 1, 0, 0, 2, 0, 2, 1, 2, 0, 0, 1, 0, -1, 2, 0, 2, 0, 1, 0, 1, 0, 0, 0, -1, -1, 2, 0, -1, 3, 1, 3, 3, 0, 1, 3, 2, 1, 1, 1, 0, 1, 0, 0, 2, 1, 1, -1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 2, 0, 1, 0, 1, 1, 3, 2, 2, 1, 3, 2, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 2, 3, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 2, 1, 0, 1, 0, 2, 0, 0, -1, 1, 0, -2, -1, 0, -1, 0, 0, 0, -1, 0, 1, -1, -1, 1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 2, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, -1, -1, 2, 1, 2, -1, 0, 1, 0, 1, 0, -1, 1, 1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, -1, 1, 1, 1, 0, 1, -1, 0, 0, 1, -1, 0, 0, -1, 0, 1, 1, 0, 2, 1, 0, 1, 0, -1, 1, -1, 0, 0, -1, -1, -1, 2, 1, 0, 0, 0, 0, -1, -1, 2, 0, 0, 0, 1, -1, 0, 1, 0, 1, -1, 1, 1, 1, 0, -1, 1, 1, 1, 0, 1, 0, 1, 0, 0, -1, -1, 1, 1, -2, 1, 1, 0, 0, -2, -1, -1, 0, 1, 0, -1, -1, -1, 0, 1, -1, 1, 0, 2, 1, 1, 0, 2, 0, 0, 2, 0, 0, 0, 1, -2, 0, 0, 2, -1, 2, 0, 0, -2, 1, 0, 0, -1, 1, 0, 1, 1, 0, 0, 1, 2, 2, 1, 0, 0, 2, 0, -2, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, 1, -1, 2, 0, -1, 0, 0, -2, -1, 1, -2, -1, 0, 1, -1, 0, -1, 0, 1, 0, 0, -1, 0, 1, 0, -1, 0, 1, 2, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 1, 2, 1, 0, 1, 1, 0, 0, 2, 0, 1, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, -1, 0, -2, -1, 1, 0, -1, -2, 1, 0, 1, 1, 0, -1, 0, 2, 0, 0, 0, 1, 1, -1, 1, 0, 1, 2, -1, 0, 0, -1, 0, 0, -1, -2, 0, 0, -1, -2, 0, 1, -2, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 1, -2, 0, 0, -2, 0, 0, 0, -2, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 1, 1, 1, -2, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, -1, 1, 0, 1, 1, -1, -1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 1, -1, -1, 0, 1, 0, 2, 2, 0, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, -1, 1, 1, 0, -2, 0, 0, 0, 1, -2, -2, -1, 0, 0, 1, 1, 0, 1, 2, 2, 1, 0, -1, 0, 0, 0, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, -2, 0, 0, 0, 1, 1, 0, -1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, -1, 0, 1, 1, 0, 1, 0, 1, -1, -1, -1, -2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 2, 0, 1, -2, 1, 1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, -1, -1, 1, 0, -1, 1, 0, 0, 1, 2, 2, 0, 0, -2, 0, 0, -1, -1, -2, -2, 1, -1, 0, -1, 0, 1, 1, 1, 1, 0, 0, 2, 0, -1, 0, 0, 0, -1, 2, 0, 0, 0, -2, 1, 1, 0, 0, 1, 1, 0, -2, -2, 0, -2, 0, -1, -1, 0, 0, -1, -1, -1, 2, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 2, -1, 0, 0, 0, 0, -2, -1, 1, 0, -2, 0, 1, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 0, -1, 1, 0, -1, -1, 1, 0, 1, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, -1, 0, 1, 1, 0, 1, 0, 1, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, -1, 0, -1, -1, 0, -1, 0, 1, 0, 1, 1, 1, -1, -1, 0, 1, 0, -1, 0, 0, -1, 0, 1, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 1, 2, 1, 0, -1, 1, 1, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 1, -1, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, -1, 1, -1, 1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, -1, -1, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, -1, -1, 1, 0, 1, 0, -1, -1, 0, 2, 1, 2, 1, 0, 2, 0, 2, 1, 1, 2, 0, 0, 1, 1, 0, 0, 2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, -1, 2, -1, 0, 2, 0, 1, -1, 0, 0, 1, 1, 0, 2, -1, 2, 1, 2, -1, 1, 0, 1, 1, 0, 1, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, -1, 1, 0, 0, 2, 1, 0, -1, 0, 1, -1, 2, 1, 0, 2, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 2, 1, 2, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, 2, 0, 1, -1, -1, 2, 0, 0, -1, 1, 1, 0, 2, 1, -1, 0, 1, 0, 1, 0, 1, -1, 0, 0, 1, 1, -1, 2, 0, 1, 2, 1, 1, 1, 1, -1, 2, 1, 0, 2, -1, -1, 0, 2, 1, -1, 2, 1, 0, 0, 0, 2, 2, -1, 2, 0, 0, 1, 1, -1, 1, 1, 2, 0, 1, 1, -1, 1, -1, 0, 0, 2, 1, 2, 0, 0, 2, 0, 0, 0, 1, 0, 2, 2, 0, 1, 2, 1, 0, 0, 1, 0, 1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 2, 2, 0, 2, -1, -1, 1, 0, 0, 1, 2, 0, 1, 2, 1, 2, 0, 2, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, -1, -1, 1, 0, 2, 1, -1, 1, 0, 2, 1, 0, 2, 2, 1, -1, 0, 0, -1, 0, 2, -1, 0, 0, 0, 0, 1, 2, 1, -1, 0, 1, 1, 0, 1, 2, 0, 1, 2, 1, 1, 0, 1, 2, 0, 0, 0, 1, 1, 1, 0, 0, -1, 2, 0, 2, -1, 1, 1, 0, 0, 2, -1, 1, 0, 1, 1, 2, 2, 2, 0, 0, 2, 2, -1, 0, 0, 0, -1, 0, 1, 2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 2, 0, 0, -1, 0, 1, 1, 0, -1, 1, -1, 1, 0, 0, 1, 1, 1, 1, -1, -1, 0, -1, 1, 0, 0, 2, 0, 1, 2, 0, 0, 0, 1, 2, 0, 1, -1, -1, 0, 2, 1, 2, 0, 1, -1, 0, 1, 0, -1, -1, 0, -1, 1, 0, 1, 2, 0, 1, 0, 0, 1, 2, 2, 2, 1, 1, 0, 2, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 1, 2, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 0, 2, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 1, 0, 1, 0, 1, 2, 0, 0, 0, -1, -1, 2, 0, 2, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 2, 1, 0, 2, 1, 0, 0, 0, 0, -1, 1, 2, 0, -1, -1, 0, 0, 0, -1, 0, 1, -1, 0, 2, 0, 0, 1, 1, -1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, 0, 2, 0, 0, 2, 1, 0, 2, 0, 0, 0, 1, 0, 1, 0, -1, 1, 1, 0, 0, 2, 0, 1, 0, 0, 0, 2, 0, 1, 1, 0, 2, 1, 0, -1, 1, -1, 0, 0, 0, -1, 1, 0, 1, 2, 2, 0, 1, -1, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 2, 0, 1, 1, 1, 0, 2, 0, 1, 1, 1, 0, 1, 0, 0, 0, -1, 2, 1, 0, 0, 1, 0, 0, -1, -1, 0, -1, 2, 2, 1, 1, 1, 2, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, -1, 0, 0, 1, 2, -1, -1, 2, 1, 0, 0, 1, 1, 0, 2, 1, -1, 0, 0, -1, 2, 0, -1, 2, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 1, 0, 0, 2, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 2, 0, 2, 1, -1, -1, 0, 0, 0, 1, 0, 1, -1, 0, 1, 0, 0, 0, -1, -1, 0, 2, 1, 2, 0, 0, -1, 0, 1, 0, -1, 2, 0, 1, 1, 0, 1, 1, 1, 2, 2, -1, 0, 0, 0, 2, 2, -1, 2, 0, -1, 0, 2, 0, 1, 0, 0, 1, -1, 2, 0, 0, -1, 0, 2, 1, 0, 0, 1, 2, 0, 1, 2, 0, -1, 1, 0, 1, 0, 2, 1, 0, 0, 1, 2, 0, 1, 1, 0, 2, -1, 0, 0, 0, 0, 0, 0, 2, -1, 0, 2, -1, 0, -1, -1, 1, 1, 2, 0, 2, 0, 2, 0, 0, 1, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 2, 0, 2, 0, 1, 1, 2, 2, 2, 1, 0, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 2, 2, 2, 0, 0, 1, 1, 0, 2, 0, 1, 0, 1, 2, 0, 1, 2, 1, 0, 1, 1, 0, 1, 1, 0, 1, 2, 2, 1, 0, 2, -2, -1, 0, -1, 0, 1, 0, -2, 0, 1, 0, -2, -2, 0, -1, 0, -3, 0, -1, -3, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, -1, 0, -1, -2, 0, 1, 0, 0, 1, 0, 0, -2, 0, 0, 0, -3, -2, -1, -2, 0, -1, 0, 0, 0, 0, -1, 0, -3, 0, -1, 1, 0, -1, 0, -1, -1, -1, 1, 0, 0, 0, 0, -2, -1, -3, -2, -2, 1, -2, 0, -2, 0, 0, -1, 0, -2, -3, 0, -2, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 1, -2, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, -2, 0, 0, -1, 0, 1, 0, 0, 1, -1, -2, -2, 0, -2, 0, -1, 0, -1, -1, -1, 0, 1, 1, -1, -2, -1, -1, 0, 1, -2, -2, -2, 1, 0, 0, -1, 1, -2, 0, 1, -2, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, 0, 0, -2, 1, -1, 1, -2, 0, 0, -2, 0, -2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, -2, 0, -1, -1, 1, 1, -1, 1, -2, 0, -1, 0, 0, 0, -1, 1, 0, 0, -2, -1, 0, 0, -2, -2, 1, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, 1, 0, -1, 1, 0, -2, -1, 0, 0, 1, -2, -1, 0, 0, -1, 0, -2, 0, 0, 1, -1, 0, -1, -1, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 1, -1, -1, 1, -1, 0, 0, 2, 1, 1, 0, 0, 2, 0, 0, 1, 0, 1, 1, -1, 0, -2, -1, -2, 0, -3, -1, -2, 0, 0, -1, 0, 2, 0, -1, 1, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 1, -2, 0, -1, 1, 1, -3, 0, -2, -2, -2, 0, -3, 0, 1, -2, 1, 2, 1, 2, -1, 0, 0, 2, 0, 1, 1, 1, 0, -1, -1, 0, 1, 1, 0, 0, -1, -2, -2, -1, -2, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 2, 2, 0, 1, 0, -1, 0, 0, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, -1, -2, -1, -2, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, -1, 1, 0, 0, 1, -3, -3, 0, -1, -2, -3, 0, 0, 1, 0, 0, 2, 2, 2, 1, 0, 2, -1, 1, 0, 0, 0, 0, 0, 0, -1, 1, -1, -1, 0, -3, 0, 0, -1, -2, 0, 0, -1, -2, -1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 1, 1, 2, -1, 0, -1, 0, -1, -2, -2, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, 0, 1, 0, 1, 1, 2, 2, 2, 0, 2, 0, 2, 0, 2, 0, -1, 0, 1, -2, 0, -1, -2, -3, -1, -1, 0, 0, 1, 1, 2, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 2, 0, 0, 0, 1, 0, 0, -1, 1, 1, 1, 2, 1, 0, -1, -1, 0, -1, 0, -2, 0, -2, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 2, 0, -1, -1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -2, 0, -1, 1, 0, -2, -1, 1, 0, 1, 0, -1, 2, 0, 0, -1, 1, -1, 0, -1, 1, 1, -1, -1, 0, 0, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, 2, -1, 0, 0, 0, -1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, 1, -1, 1, -1, -1, 0, -1, 0, 0, -2, 0, 0, -2, 1, 0, 1, 2, 1, -1, 0, 2, 0, 1, -1, 1, -1, -2, -1, -1, -1, -2, -1, -1, -2, 0, -1, -1, 0, -1, -1, -2, 1, -1, -2, 0, -1, 0, -1, 0, -1, 0, 0, 1, 1, -1, -2, 0, 0, -1, 0, 0, -1, 0, 0, -1, -1, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, -2, 0, 0, -2, -3, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, -1, 0, 1, -1, -1, -2, 1, 0, 0, 0, -1, 0, -2, -2, -1, -2, -1, -1, -1, -2, -1, 0, -1, 1, -1, 0, 0, 0, -1, 0, 0, -1, -2, 1, -2, -1, -1, 0, 1, -1, -2, -2, -2, -1, -2, 0, -2, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -3, 0, 0, 0, -2, 0, -1, -2, -2, 0, -3, 0, 0, 0, -2, 0, -2, -2, -2, -2, -2, 0, -1, 0, -2, -2, -1, -1, -3, 0, -1, -1, -2, -1, -2, 0, -2, -2, -2, 0, 0, 0, 0, -2, 0, -2, -1, -2, -1, -2, -1, -3, -1, -2, -3, 0, -3, -3, -3, 0, -3, -1, 0, -1, -1, 3, 1, 1, 1, 1, 2, 4, 2, 1, 2, 3, 0, 0, 2, 1, -1, 0, -1, 0, -1, -1, 0, 0, -3, -4, 0, -2, -2, -1, -4, 2, 2, 3, 2, 2, 2, 2, 3, 2, 2, 3, 2, 1, 1, 0, 0, -1, -1, 0, -1, -1, -1, 0, -3, -1, -3, -3, -4, -3, -3, 1, 3, 2, 4, 5, 1, 1, 1, 3, 3, 4, 0, 0, 0, 0, 1, -2, -2, 0, 0, -2, -1, 0, -3, -3, -1, -3, 0, -4, -4, 3, 2, 4, 4, 3, 5, 4, 3, 3, 1, 3, 0, 0, 2, 0, -1, -1, -2, 1, -2, -1, -2, -1, 0, -1, -2, -2, -1, -2, -1, 3, 4, 5, 4, 4, 4, 4, 3, 4, 2, 0, 1, 2, 0, 1, 0, 0, -1, 0, 1, -2, 0, -2, -1, -3, 0, -3, -2, -3, -1, 5, 4, 1, 3, 4, 3, 3, 4, 2, 3, 2, 0, 1, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 5, 2, 5, 2, 2, 1, 5, 5, 4, 3, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, -2, 0, -2, 0, -3, -1, 2, 2, 2, 5, 2, 1, 4, 2, 4, 4, 1, 3, 1, 2, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, -1, -1, 1, -2, 0, -2, 3, 3, 2, 2, 2, 2, 2, 5, 2, 1, 0, 2, 3, 2, 1, 0, 1, 1, 2, 1, 1, 1, -1, 0, 0, 1, 1, -1, 0, -1, 5, 1, 2, 3, 4, 4, 3, 2, 0, 3, 3, 1, 0, 1, 0, 0, 0, 1, 2, 2, -1, 1, 2, 0, 2, 0, 0, 0, 0, 0, 3, 1, 4, 3, 2, 3, 3, 0, 3, 3, 3, 2, 0, 2, 0, -1, 0, -1, -1, 0, -1, 0, 1, 0, 2, 2, 2, 0, 0, 0, 2, 2, 3, 0, 3, 3, 0, 0, 2, 1, 0, 1, 2, -1, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, 3, 1, 2, 0, -1, -2, 2, 2, 4, 1, 3, 2, 3, 0, 0, 0, 0, 1, 1, -1, -1, 0, -1, 1, 0, -1, -1, 1, 0, 2, 2, 1, 1, 1, 0, -2, 1, 3, 3, 1, 3, 0, 0, 3, 0, 3, 2, 2, 0, 0, 1, -1, 2, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, -1, -2, 1, 1, 2, 3, 2, 0, 0, -1, 0, 0, 1, 2, 1, 2, 0, 0, 0, 1, 0, 0, 2, 2, 0, 2, 2, 0, 0, 1, -2, 0, 4, 1, 1, 1, 2, 1, 0, 2, -1, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 2, -1, 0, 0, 2, 3, 2, 0, -2, -2, -1, 2, 2, 2, 4, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 2, 0, 2, 2, 1, 0, -1, 0, -1, 0, -1, 1, 2, 4, 2, 0, -1, 1, 2, 0, -1, 0, 2, 2, 1, 0, 2, 2, 0, -1, -1, 1, 2, 3, 3, 3, 0, -1, 2, 0, 0, 2, 2, 1, 3, 2, 0, 0, -1, 0, 0, 1, -1, 1, 0, 0, 1, -2, -1, 0, 0, 0, 2, 3, 2, 0, 1, 0, 0, -1, 1, 3, 4, 2, 3, 1, 0, 0, 1, 1, 0, 0, 1, 1, -1, 0, -1, -1, 0, 0, 1, -1, 1, 0, 2, 0, 1, 0, 0, 0, 0, 5, 3, 1, 4, 3, 2, 0, 0, 2, 2, 1, 0, 0, 1, 0, -2, 1, -2, 0, 0, 1, 0, 2, 0, 1, 0, -1, -1, 0, 1, 6, 2, 3, 3, 2, 2, 3, 2, 1, 2, 2, 0, 1, 0, 0, -1, 0, -3, -2, -1, -1, 0, -2, 1, 1, 0, 1, -2, -1, -2, 4, 3, 6, 2, 5, 4, 3, 1, 1, 0, 3, 3, 1, 2, 0, 0, -2, 0, 0, -2, 0, 0, -2, 0, 0, 1, 1, -1, 1, 0, 7, 4, 4, 3, 6, 4, 2, 3, 1, 2, 4, 2, 1, 1, 0, 0, -1, -3, -1, -2, 0, 0, 1, -2, 0, 0, 0, 0, 0, -2, 7, 4, 3, 3, 4, 1, 4, 2, 2, 3, 3, 3, 0, 2, 2, -1, 0, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, 5, 3, 6, 3, 3, 3, 2, 3, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, 0, 0, -1, -2, 0, -2, 3, 6, 3, 5, 2, 4, 2, 2, 3, 4, 3, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -1, -3, 0, -3, 0, 0, 5, 4, 3, 4, 5, 4, 4, 3, 3, 1, 0, 3, 1, 0, 2, 2, 0, -1, 1, 1, 1, -1, 0, -1, -3, -2, 0, 0, -2, 0, 5, 6, 5, 4, 2, 1, 4, 1, 4, 3, 1, 0, 2, 1, -1, -1, 1, 0, 2, 0, 0, -2, -1, 0, -2, 0, -1, 0, 0, -1, 2, 4, 2, 4, 4, 3, 1, 3, 1, 2, 0, 0, 2, 0, 0, 0, 2, 0, 1, 0, 0, -2, -2, -2, -3, -1, -3, 0, -3, -3, 1, 1, 2, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, -1, 2, 1, -1, 1, 0, 0, 1, 1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 0, 0, -1, 0, 0, 0, -2, 2, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 2, 1, -2, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 2, -1, 1, 1, -1, 1, 1, 0, 1, 2, 0, -1, 1, 0, 1, 0, 0, -1, -1, 0, 0, 1, 0, -1, -1, 0, 1, 0, -1, 0, -1, 1, 0, 2, 1, 0, 0, 1, 1, 0, -1, 0, 2, 0, -2, 0, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, -1, 1, 2, 0, -1, 2, 0, 0, 0, -1, 0, -1, 1, 1, 0, 1, 0, -1, 1, -1, -2, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, -1, 0, -1, -1, 1, 0, 0, 0, -1, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 2, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, 1, -2, 1, -1, 0, -1, -1, -1, -1, 1, 0, 0, 1, 1, 0, -1, 1, 1, 1, 1, 1, 0, 0, 0, 1, -1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, -1, 0, -1, 1, -1, 0, 0, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, -2, 0, 2, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, 1, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -2, 1, 0, 0, -2, 1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, -1, 1, 0, 1, -2, -1, -1, -1, 1, 0, 1, 0, 1, 0, -2, 0, 0, -1, 2, -2, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, -1, -1, 0, -1, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 1, -1, 0, -1, -2, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 2, -1, 1, 0, -1, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, -1, -1, 0, -1, -2, 1, -1, -2, -1, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, 1, 2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 0, -1, -2, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -2, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 1, 1, -1, 1, 1, 2, -1, 0, 1, 0, -1, 1, -1, 1, -1, 1, 0, -1, -1, -1, -1, 0, -1, -1, -2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 1, 1, 0, 1, 1, 0, 0, -2, 0, -2, -2, 0, 2, 0, 0, 0, -1, 0, 0, 0, -2, 0, -2, 0, 0, 0, -1, -1, 0, -1, 2, -1, 1, 1, -1, -1, 1, 0, 1, 0, -1, 1, 0, -1, 1, 2, 1, 0, 1, 0, 0, 1, 0, -2, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, -2, 1, 1, -1, 0, 1, -1, 1, 1, -1, 2, 0, 0, 1, -1, -1, 0, -1, 0, 0, -1, -2, 0, 1, 1, 1, -1, 0, -1, -1, 1, 1, 0, 1, 1, 0, 1, 0, -1, 2, -1, 0, 1, 1, 0, 2, -1, -1, -1, -1, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 1, -1, 0, -1, -1, 0, 1, -2, 1, 1, -1, -1, 0, -1, 1, 1, 0, 1, -1, -1, -1, 1, 2, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, -1, -1, 0, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -1, 1, -1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 0, 1, 0, -1, 1, 0, 0, 0, -2, 1, 1, 1, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 1, 0, 1, 0, 0, 1, -2, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, -1, 1, 0, 0, 2, 0, 1, -1, 0, -1, 1, -1, 0, -1, 1, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 1, -1, 0, -1, 0, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 1, -1, 0, 1, 0, 1, 0, 1, -1, 1, -1, -1, 1, 1, -1, 1, 0, 0, 0, -1, 1, 1, 0, 0, -1, 1, 0, 0, 1, -1, 0, 1, 0, -1, -1, 0, 1, 0, -1, 0, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, 2, 0, 0, 1, -1, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, -1, -2, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, -1, -1, -1, -1, 0, -1, -1, 0, 0, -1, 1, 1, 1, 0, -1, 0, 0, 1, 0, -1, 1, -2, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, -1, -1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, -2, 0, -1, 0, 0, 0, 1, 1, 2, 0, 0, -1, 0, -1, 1, 0, 0, 1, 0, 1, -1, 2, 1, -1, 1, 1, 1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, -1, 2, 0, 0, 1, -1, 0, -2, 1, -2, 0, -1, -1, -1, 1, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 1, -1, 1, 0, -2, 1, 0, -1, -1, -1, 2, 0, 1, 0, 0, -1, 2, -2, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, -1, 1, -1, 2, 0, -1, 1, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, 1, 1, -1, 0, 0, 0, 1, -1, 0, 1, -1, 0, 1, 0, -1, 1, 1, 1, 0, 0, 0, -1, -2, 0, -1, -1, 0, 1, -1, -1, -1, 0, 0, 0, -1, 2, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, -1, 1, 0, 0, -1, 0, 1, 1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 1, -1, 0, 0, 1, -1, 0, 0, 0, 0, -2, 0, 0, 1, 0, 0, 1, 1, 1, -1, 1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, 1, 1, 0, 0, 1, -1, -1, 0, -1, 0, -2, 0, 0, 0, -1, 1, 0, -1, 1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, -1, 1, -1, 0, -1, 1, -1, 0, 1, 0, 1, -1, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, -1, 1, -1, 1, 2, 0, 1, 0, 0, -2, 0, 0, 1, 2, 1, 1, 0, 0, -1, -1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, -2, -1, 1, -1, 1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, -2, 1, 2, 2, 1, 1, -2, 0, 1, 1, 0, 0, 1, 2, -1, -1, -2, 0, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, 1, -1, 0, 0, 0, -1, 1, 0, 0, 1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 1, 0, 0, -1, 1, 1, -1, 1, 1, -1, 0, 0, 1, 0, 0, 1, -1, 1, 1, -2, 0, 1, 0, -1, 0, 0, -1, 0, 1, 0, -1, 0, 0, 1, -1, -1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, -1, -1, 1, 0, 0, 0, -2, -1, 0, -1, 1, 0, -1, 0, 0, 0, 0, -1, -1, -2, 1, 1, 1, 0, 0, 2, 0, 1, 2, 0, 0, -1, 1, -1, 1, 2, -2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 0, -1, 0, 1, 1, 1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 0, -1, 1, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 1, -1, -1, 1, -1, -1, 1, 0, -1, -1, -1, 1, 0, 0, 0, -1, 2, 2, 1, -1, 0, 0, -1, 0, 2, -1, 0, 0, -1, 1, -1, 0, -1, -1, 0, -1, 2, 1, 0, 0, -1, -1, 0, -1, -1, 0, 1, -1, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 0, -2, 1, 0, 1, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, -1, 1, -1, 1, 0, 0, 1, 1, -1, 1, 1, 1, 1, -1, 1, -1, 0, 0, -2, 1, 0, -1, 1, 0, 1, 0, 1, 0, 0, 1, -3, -1, 0, 0, -1, -1, 0, 1, -1, 0, 0, 0, 0, -1, -2, 0, -1, -3, -3, -2, -4, -5, -6, -6, -4, -3, -5, -6, -6, -2, -3, 1, 0, 0, 1, 1, 2, 2, 0, 3, -1, -1, 1, -2, 0, 0, -3, -5, -3, -4, -2, -6, -6, -4, -3, -4, -6, -5, -6, -4, 0, 0, 1, 1, 2, 2, 3, 2, 0, 1, 2, 0, 0, -2, -2, -3, -3, -4, -5, -1, -2, -5, -1, -5, -5, -4, -5, -3, -3, -2, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 1, 0, 1, 0, -1, -2, -4, -1, -2, -4, -3, -2, -2, -3, -5, -3, -5, -5, -3, -3, 0, 0, -2, 2, 0, 1, 1, 1, 3, 2, 0, -1, 0, 0, -1, -3, -5, -2, -2, -2, -3, -2, 0, -3, -2, -4, -4, -1, -2, -4, -2, 0, 1, 0, 3, 1, 2, 1, 2, -1, -2, -1, -2, -2, -2, -1, -1, -3, -1, -1, -1, 0, -2, -2, -1, -3, -1, -2, -1, -2, -3, 1, -1, 0, 0, 2, 0, 3, 1, -1, 0, -1, -3, -4, -4, -2, -4, -1, -3, 0, 0, -1, 0, -1, 0, 0, 0, -2, 0, -2, -1, 0, 0, 0, 1, 1, 1, 0, 0, -1, -3, -2, -2, -1, -4, 0, 0, 0, -1, 1, -2, 1, 0, 0, 1, -1, -2, -1, -2, 1, -1, 0, -1, -1, -1, -2, 0, 2, 1, 0, -1, -1, -2, -1, 0, -3, -2, -2, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 2, -1, -2, -4, -3, -2, 0, 0, -3, -2, -1, 0, -3, -2, -4, 0, 0, 0, 0, 0, 0, 0, -1, 2, 0, 1, 0, 0, 0, 0, 0, 1, -5, -5, -1, -4, -1, -3, -3, -1, -4, -2, -3, -3, 0, -1, 0, -2, -1, -1, -1, -1, 2, 1, 0, 1, 2, 0, 1, 2, 2, 3, -3, -5, -2, -4, -5, -5, -5, -2, -4, -2, -2, -3, -1, 0, 0, -1, -1, 0, 0, 0, 3, 2, 1, 1, 2, 2, 2, 1, 2, 3, -2, -4, -4, -3, -5, -3, -6, -4, -5, -2, -4, 1, 0, 0, 1, 0, 1, 1, 0, 1, 3, 1, 2, 2, 2, 1, 2, 2, 1, 0, -3, -5, -4, -4, -5, -6, -4, -6, -4, -4, -1, 0, 0, 1, 1, 3, 1, 1, 1, 1, 3, 0, 0, 2, 1, 4, 3, 2, 4, 2, -3, -3, -4, -2, -3, -7, -3, -3, -4, -2, -2, 1, 3, 3, 1, 3, 2, -1, 2, 3, 3, 3, 4, 2, 5, 3, 2, 4, 3, 2, -3, -5, -6, -6, -6, -7, -5, -3, -3, -4, -2, 0, 1, 2, 1, 2, 0, 3, 0, 2, 1, 2, 4, 4, 5, 4, 3, 4, 7, 2, -2, -4, -3, -7, -4, -4, -7, -6, -5, -1, 0, -2, 2, 0, 1, 1, 3, 2, 3, 1, 1, 4, 3, 4, 6, 7, 5, 8, 4, 5, -4, -2, -4, -5, -4, -5, -6, -7, -3, -1, 0, -1, 0, 3, 2, 2, 1, 0, 4, 2, 3, 5, 6, 4, 6, 4, 4, 6, 5, 1, -2, -3, -3, -4, -2, -4, -6, -3, -2, -2, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 1, 3, 3, 4, 6, 6, 5, 5, 1, 1, -4, -1, -2, -4, -4, -5, -5, -2, -4, -2, 0, 0, 1, 0, 3, 2, 0, 1, 0, 2, 2, 4, 3, 2, 2, 4, 2, 2, 3, 2, -1, -2, -3, -2, -2, -2, -1, -5, -4, -1, -3, 1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 2, 0, 3, 0, 1, 2, 0, 0, 0, -2, -2, 0, -2, 1, -1, -2, 0, -2, -2, 0, 1, -1, -1, 0, 0, 1, -1, 0, 0, -1, 1, 1, 1, 2, 1, 0, 0, -1, 0, -3, -3, 0, -1, 0, 1, 1, -1, 0, 0, 0, 2, 1, 1, -1, -2, 1, 0, 0, 2, -1, -2, -2, 0, 2, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 2, -1, 0, 1, 2, -1, 0, -1, 0, 1, 1, 2, 2, 1, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 1, 2, 2, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -2, 0, 0, 0, -1, 0, 2, 3, 0, 4, 2, 2, 0, 2, 2, 1, 0, 0, -1, 0, 1, 1, 0, 0, -2, -1, -2, 0, -2, 1, 0, 0, -2, -1, 0, 0, 2, 3, 3, 0, 3, 3, 3, 3, 0, 0, -1, 0, -1, 0, 0, 1, -1, 0, -2, 0, 0, 0, -3, -1, 0, 0, 0, -2, 1, 1, 0, 1, 3, 0, 0, 3, 0, 1, 1, 2, 0, 0, 1, 0, -1, -1, 0, 0, -2, -2, -1, -3, 0, 0, 0, -1, -4, -1, 0, 1, 0, 0, 0, 2, 2, 2, 0, 0, 2, 1, 1, -1, 0, -1, 1, 1, 0, -3, -2, -1, 0, 0, -1, -4, -4, -4, -5, -2, 0, -2, 0, 0, -1, 1, 1, 2, 2, 0, -1, -1, 1, 0, 0, -1, -1, -1, -1, -2, -2, -1, -3, -4, -2, -5, -3, -3, -3, -3, -2, 0, 0, 0, 2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, 0, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -2, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 1, -1, -1, 0, 0, -1, -1, -1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, -1, 2, 1, 1, 0, -2, -1, 0, 2, 0, 0, 0, 1, 0, 0, -2, 0, -2, 0, 1, 1, 2, -1, 0, 0, 0, 0, 2, -1, 1, 0, 0, -2, 0, -2, 0, 0, 1, 0, 0, -1, 0, -1, -2, -1, 2, -1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -2, 0, 0, -1, 0, -1, 0, 0, -1, -1, 1, -1, 0, 0, 1, 0, -1, -1, 1, 0, 1, 1, 0, 0, 2, 0, -1, 0, 0, -2, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, -1, 1, -1, 0, -2, 2, 1, 0, 2, -1, 0, 0, 0, 2, 2, 1, 0, -1, 1, -1, 0, 0, 1, 0, 0, 0, -2, -1, 1, 0, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 2, 0, 0, 1, 2, 0, -2, -2, 0, 1, -1, 0, -2, 1, -2, -2, 0, 0, -1, -2, -1, 1, 0, 1, 0, 0, 2, -1, 0, 1, 1, 0, 2, 0, 2, 0, 0, 0, 0, -1, -1, 0, -2, -1, 0, 0, 0, -2, -2, 0, -1, -1, -1, 0, 1, 0, 0, -1, 0, -1, 1, 0, 0, 0, 2, 2, 0, -2, 0, 0, -3, 0, 1, 0, -1, 0, -1, 1, 0, -1, 1, -1, -1, 0, 0, 0, 2, 1, 0, 0, 2, 0, 0, 3, 1, 0, -2, -1, 0, -1, 1, -3, 0, 0, 0, 0, -1, -2, -2, -1, 1, -1, -1, -2, 0, -1, 1, -1, -1, 0, 0, 2, 0, 0, 1, 3, 0, -2, -1, -2, -3, -1, 0, -2, 0, 0, -2, 1, 1, 0, 1, 0, 2, 0, 1, -1, 0, -1, 0, 1, 0, 0, 2, 2, 2, 3, -1, -2, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 1, 3, 2, -2, 0, 0, 0, -2, -1, -2, -2, -3, 0, 1, -1, 2, 1, -1, 1, 0, 0, 0, 0, -1, 0, 3, 0, 1, 0, 0, 0, 1, 1, 0, -1, -2, -2, 0, -1, -2, 0, 1, -2, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 0, 3, 2, 2, 1, 2, 2, 1, -2, 0, -3, -1, -1, 0, -1, 0, -1, 0, 0, 0, 1, -1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 2, 0, 1, 1, 3, 3, 1, 0, -2, 1, -1, 0, -1, -1, 0, 0, -2, -2, -1, 1, 0, 2, 1, -1, 0, 0, -1, 2, 0, 0, 0, 0, 0, 3, 0, 2, 0, 0, -2, -1, 0, 1, -2, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 2, 0, -2, 0, -1, 0, -1, -2, 0, -2, 0, 1, 0, 0, 1, 0, 1, -1, -1, -1, 1, 0, 0, 0, 2, 2, 1, 1, 0, 1, 1, -1, 0, -2, -1, 0, 1, 0, 0, -1, 1, 1, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 2, 2, 0, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, 1, 0, -1, -2, 0, 0, -1, -1, -1, -1, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, 1, 1, 2, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 1, -1, 0, 1, 0, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 1, -1, 0, -1, 1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, -1, 1, 0, 0, 1, 2, 0, -1, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 2, 0, 1, 2, -1, -1, -1, 2, 2, 1, 1, 0, 2, 0, 0, 0, -1, -1, 0, 0, 2, 0, -1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 2, 0, 0, -1, 0, 0, 1, 2, 0, 0, 1, 0, 1, 1, 1, 0, 0, 2, 0, 0, -1, -1, -1, 2, 2, 0, 2, 0, 0, 1, 0, -1, 2, 2, 0, 0, 0, 0, 0, 1, 0, -1, 2, -1, 0, -1, 1, 1, 0, -1, 0, 0, 0, -1, 2, -1, -1, 0, 0, 2, 0, 2, 0, 1, 0, 0, 2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 2, 0, 0, 0, 0, 1, 0, 3, 0, 1, 2, 1, 3, 3, 2, 0, 1, 2, -1, -2, 0, 0, -2, -2, -5, -2, -5, -5, -1, -3, -1, -3, 1, 0, 0, 1, 4, 3, 4, 3, 4, 3, 2, 5, 1, 1, -1, 1, -1, -2, -3, -3, -4, -4, -4, -1, -4, -5, -4, -2, 0, -4, -1, -1, 0, 2, 4, 4, 5, 2, 2, 1, 3, 1, 0, 2, 0, -3, -3, -2, -3, -3, -1, 0, -3, 0, -2, -1, -1, -1, -1, 0, 1, -1, 1, 0, 4, 2, 2, 3, 4, 2, 3, 1, -2, -1, 0, -1, -3, -1, -1, 0, -1, -1, 0, 0, 0, -2, -1, 0, 0, -2, 0, 1, 0, 1, 3, 5, 4, 3, 5, 3, 0, 0, 0, 0, -2, -3, -4, -1, -2, 0, -1, 0, 1, 0, 1, -2, 0, -1, 0, 0, 0, 0, 1, 3, 1, 4, 3, 5, 3, 1, 0, 0, -1, -4, -3, -4, -1, 0, 0, -1, 0, 0, -1, 1, 2, 2, 0, 0, -1, 0, 0, 1, 0, 2, 3, 4, 1, 2, 1, 0, 1, -1, -3, -1, -3, -2, -3, -2, -2, -1, 2, 1, 0, 1, 0, 1, 0, 3, 0, 0, -2, -2, 0, 2, 2, 2, 0, 3, 2, 0, -1, -4, 0, -1, -3, -2, -1, -2, 0, 1, 0, 3, 1, 1, 0, 0, 1, 1, 0, 3, -4, 0, -2, -3, 0, -2, 1, 0, 1, -2, -4, -1, 0, -3, -1, -3, -1, 0, 0, 1, 0, 0, 2, 4, 0, 2, 0, 1, 3, 1, -5, -4, -4, 0, -1, -1, -2, -3, -1, -1, -2, -3, -1, -3, -2, -2, -3, 0, -2, -2, 0, 2, 4, 3, 1, 3, 4, 5, 4, 2, -3, -3, -2, -4, -2, -2, -1, -2, -5, -5, -3, -1, -3, -3, -3, 0, 0, -2, 0, 0, 0, 2, 1, 4, 1, 1, 4, 5, 5, 4, -4, -4, -1, -2, -5, -5, -3, -6, -3, -5, -3, 0, 0, -1, 0, 1, 1, 0, 3, 2, 2, 4, 2, 5, 5, 5, 5, 5, 5, 2, -4, -1, -4, -2, -6, -5, -4, -6, -6, -5, -4, 0, 0, 2, 0, 0, 0, 0, 0, 0, 4, 5, 3, 5, 5, 4, 6, 6, 7, 5, -5, -4, -1, -3, -6, -7, -7, -5, -3, -2, -2, -1, 0, 2, 2, 0, 0, 1, 3, 0, 3, 3, 2, 4, 5, 5, 7, 7, 7, 5, -3, -3, -2, -3, -4, -8, -7, -6, -3, -4, -1, -2, 0, 3, 0, 1, 0, 0, 1, 1, 5, 3, 6, 8, 8, 9, 9, 10, 6, 7, -5, -2, -4, -4, -7, -8, -5, -7, -4, -4, -2, 0, -1, 1, 3, 0, 0, 4, 5, 4, 5, 3, 7, 6, 8, 10, 10, 9, 8, 8, -2, -3, -3, -2, -3, -6, -6, -5, -3, -4, -2, -3, -2, 1, 0, 2, 0, 3, 2, 2, 3, 8, 7, 6, 9, 7, 9, 10, 8, 6, -3, -2, -3, -5, -2, -3, -6, -6, -3, -1, -1, 0, -1, 0, 1, 1, 0, 2, 1, 1, 5, 8, 6, 10, 9, 6, 8, 8, 5, 7, -4, -2, -1, -4, -3, -4, -4, -4, -2, -3, -2, 0, 0, 2, 0, 3, -1, 0, -1, 0, 3, 4, 7, 7, 7, 4, 6, 6, 5, 4, -2, -1, -1, -3, 0, -1, -3, -2, -5, -2, -2, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 1, 3, 1, 4, 5, 4, 2, 3, 2, -3, 0, -1, 0, 0, -2, -3, -3, -2, -1, 0, 0, 1, 0, 0, -1, -3, 0, 1, 0, 0, 0, 0, 3, 2, 2, 4, 4, 0, 1, -2, 0, 0, 0, 2, 1, 2, 2, -1, -1, 0, -1, 0, -1, 0, 0, -1, -2, 0, 0, 2, 0, 0, 1, 3, 0, 1, 3, 3, 1, 0, 0, 2, 2, 1, 2, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, 0, 1, 0, 2, 1, 2, 4, 2, 2, 1, 2, 0, 0, 1, 5, 4, 4, 5, 1, 4, 2, 1, 0, 2, 0, 0, -1, 0, 2, 2, 3, 0, 1, 0, 0, 2, 2, 0, 2, 2, -1, 1, 3, 2, 2, 5, 5, 6, 2, 5, 5, 1, 1, 2, 0, 2, 2, 0, 0, 2, 3, 2, 0, 0, 0, -1, 0, 2, 0, 1, 1, 0, 3, 2, 5, 3, 3, 6, 4, 3, 1, 4, 4, 3, 1, 2, 2, 3, 3, 3, 0, 2, 1, -1, -1, 1, -1, 0, 2, 2, 1, 0, 4, 1, 5, 2, 4, 2, 3, 4, 2, 2, 1, 2, 1, 2, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, -1, 0, 2, 2, 1, 2, 4, 3, 5, 5, 5, 5, 2, 4, 2, 1, 0, 2, 2, 2, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 1, 2, 1, 1, 4, 3, 2, 1, 4, 2, 3, 1, 1, 1, 3, 0, 0, 0, 0, -2, 0, -3, -1, -1, -3, -4, 0, -2, -4, 0, 1, 1, 2, 0, 2, 1, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, -3, -4, -3, -4, -3, -2, -2, -4, -2, -3, -1, 0, 0, -1, 0, 2, -1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 2, 0, 0, 2, 0, 0, 1, 0, 0, -1, 0, 0, 2, 2, 0, 0, 1, 0, -1, 2, -1, 1, 1, -1, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, 2, 2, 0, 1, 1, 2, 0, 0, 0, 0, -1, 0, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, -2, 1, -1, -1, 0, 2, 1, 2, 2, 0, 0, 0, 2, 2, 0, 0, 2, 0, -1, 1, 0, 1, 0, -1, -1, 1, -1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 3, 0, 2, 2, 0, 0, 2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 2, 0, 1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, -1, -2, -1, -1, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 0, 2, 2, 1, 0, 2, 0, 0, 2, 0, 0, 1, 2, 2, -1, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, -1, 2, 2, 0, 0, 1, 0, 1, 1, 2, 1, 0, 0, 2, 0, 1, 1, 0, 1, -1, 1, -2, -2, 0, 1, -1, 0, 2, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, 2, 0, 2, 0, 0, 1, 0, 1, -1, -2, 0, -1, 1, 0, 0, -1, 1, 0, 0, 2, 2, 0, 0, 1, 0, 0, 2, 0, 1, 0, 0, 2, 2, -1, -1, 2, 1, -1, -2, 0, 0, 1, 1, -1, 0, 0, 0, 0, -1, 2, 0, 1, -1, 2, 0, 0, 0, 2, 0, -1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -2, -1, -1, -1, 0, 0, 1, -1, 0, 0, 1, 0, 3, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, -1, 1, 1, 0, 1, 0, 0, -1, -1, 2, 2, -1, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, 2, 0, 0, -1, -1, 0, -2, 0, 1, 0, -1, -1, -2, -1, 1, -1, 0, 1, 0, -1, 0, 2, 2, 2, 0, 0, 0, 1, 0, 0, 0, -2, -1, -2, 1, -1, 0, -1, 0, 0, 0, 2, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 3, 0, 1, -1, -1, 1, 0, 0, -2, -1, 1, 2, 0, 0, 1, 0, 0, 1, 1, 0, 2, 1, 0, 1, 3, 1, 2, 1, 0, 3, 2, 0, -2, 0, 0, -2, 1, 0, -1, 0, -1, 0, 0, 0, 2, 1, 0, -1, -1, 0, -1, 3, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, 1, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 3, 2, 1, 3, 2, 3, 0, -3, 0, -1, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 3, 0, 0, 1, 0, 2, 1, 0, 2, 2, 4, 0, 3, 1, 0, 1, -2, 0, 0, -1, -1, 0, 0, -1, -1, 1, 2, 2, 0, 1, 1, 3, 3, 0, 3, 3, 0, 1, 3, 2, 1, 3, 1, 0, 0, 0, -2, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 2, 3, 3, 0, 2, 2, 1, 1, 0, 0, 3, 3, 3, 0, 1, -1, -2, 0, -2, -1, 0, -1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 2, 3, 0, 0, 0, 0, 3, 0, 1, 0, 1, 1, -1, -1, -1, 0, -2, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 1, 2, 3, 2, 2, 1, 1, 1, -1, 1, 0, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, 2, 2, 2, 0, 3, 1, 0, 1, 3, 3, 0, 1, 1, 1, 0, 2, 0, 0, 1, 0, 1, -1, -1, -2, 0, 1, 0, 1, -1, 0, -1, -1, 0, 0, 3, 2, 3, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 1, 1, -1, 0, 1, 1, 0, 0, -1, -1, -1, 1, -1, -1, 1, 1, 2, 0, 2, 1, 0, 2, 2, 0, 0, 2, 0, 2, 0, 1, 2, 0, 1, 0, 1, 0, 2, 1, 1, 0, 0, 0, -1, 0, 1, 0, 2, 0, 1, 3, 0, 1, 0, 2, 0, 0, 2, 2, 0, 0, 0, 2, 1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 0, 2, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 0, 0, 0, 0, 1, -1, 2, 0, 0, 1, -1, 1, 0, 1, 0, 0, 3, 0, 2, 1, 0, 0, 2, 0, 0, 0, 0, 1, 0, 1, 2, 3, 0, 3, 1, 0, -1, 0, 0, 0, 1, 2, 2, 2, 2, 0, 0, 2, 1, 0, 0, 0, 0, 1, 1, 1, 0, 2, 2, 1, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 3, 1, 0, 2, 3, 0, 0, 2, 0, 1, 1, 0, 0, 0, 1, 0, 0, -1, 1, 0, 1, 0, 0, -1, 0, 0, 1, -1, 0, 2, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 2, 1, 1, 0, 0, 1, -1, 0, 0, -2, 0, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 2, -1, 0, 1, 0, 2, 1, -2, 1, -1, 0, 0, 0, 0, 0, -1, 1, 0, 0, -2, -1, 0, 0, 0, 1, 0, 1, 0, 1, 1, -1, 0, 1, 0, -1, 1, 1, 0, 1, 0, -1, 0, 2, -1, -1, -1, -1, 0, 0, 1, 2, 2, -1, 1, 2, -1, -1, 0, 0, -1, -2, -1, 1, 0, 0, 0, 0, -1, -1, 1, -1, 0, 1, 1, -1, -1, 0, -1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, -1, -1, -1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, -1, 0, -2, 0, 0, 1, -1, 1, -1, 0, -1, 0, 1, 2, 2, -1, 0, 0, 1, 0, 1, 0, 1, -1, 0, -1, 0, 2, 0, 0, 0, 0, 2, 0, 0, -1, -1, -1, -1, -1, 1, -1, -1, 1, 2, 1, 2, -2, 0, 0, -1, 0, -1, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 1, 0, 0, -1, 1, 0, 0, -1, -2, -1, 0, -1, 0, 0, -1, 1, 1, -1, -1, 0, 0, 1, 0, 1, 1, -1, 0, 1, 1, 1, -1, 0, -1, 0, -1, 0, 1, -1, -2, 0, 1, 0, 0, 0, 0, 0, -1, -1, 2, -2, -1, 1, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 1, 1, 0, 0, 1, 0, 2, -1, 0, -1, -1, 1, 0, 0, -1, 0, -1, 1, 1, 0, -1, 0, 0, 1, 0, 0, 2, 0, 0, -1, 1, 0, 1, -1, 1, 0, 0, 0, -1, -1, 1, 1, -1, 1, 0, 0, 1, 0, -1, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, -2, 0, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, -1, -1, 1, -1, 0, 0, -1, 1, 0, -1, 1, -1, 0, 1, -1, -1, 1, 0, -2, 1, 1, 0, 0, 1, 0, 1, 0, 0, -2, 0, -1, 0, 0, 0, -1, 1, 1, -1, -1, 1, -1, 1, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -2, -1, 0, -1, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, -2, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, 1, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, -2, 0, 0, 0, -1, -1, -1, 0, -1, 0, -1, 0, 1, 0, 1, 0, -2, 1, 1, 0, -1, -1, 1, 0, -1, 0, 1, -1, 1, 1, 0, 0, -1, -1, 1, 1, 1, 1, 1, -1, 1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 1, 1, 0, 0, 1, 0, 0, 1, -1, 2, 0, 1, 0, 0, 0, -2, 1, 1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, -2, 0, 0, 0, -1, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, -1, 0, 2, -1, -1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, 1, 0, 1, 0, 2, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -1, 2, 0, -1, 1, -1, -1, -1, 1, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 1, -1, -1, 0, 0, 0, 0, 1, 2, -1, 0, 0, 0, -1, 1, 0, -1, 2, -1, -1, 0, 0, -1, 1, 0, -1, 1, -1, -1, -1, 1, 1, -1, -1, 2, 1, -2, 0, 1, 1, 1, -1, 0, 0, 1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, -1, 1, 0, 1, 0, 0, -1, 2, -1, 0, 0, -1, -1, 0, 1, -1, -1, -1, 0, 1, 0, 1, 0, 0, 2, 0, 0, 1, -2, 0, -1, 0, -1, -1, 0, 1, 0, 0, 1, 1, -1, -1, 1, 1, -1, 0, 0, 1, 1, 0, 1, -2, 1, 0, 0, -1, 1, 0, 1, 0, 0, -2, 0, 1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, -1, -1, -1, 1, 0, -1, 0, 1, 0, -1, -1, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, -1, 1, 1, 0, -1, 0, -1, 0, 1, -1, 0, 0, -1, 0, 0,
    -- filter=0 channel=4
    1, 0, 0, 0, -1, 0, 0, 0, -2, -2, -2, -1, -2, -1, -2, 0, 0, -3, -1, 0, -2, -1, 0, -1, -3, -1, -3, -2, -4, -1, 1, 1, -2, -1, 1, -2, -1, -2, -2, -2, 0, 0, -2, -1, 0, -3, -2, 0, -1, -1, -2, -2, 0, -2, -3, 0, -2, -2, -2, -1, 0, 0, 0, 0, 0, -2, -2, 1, -1, 0, 0, -1, 0, 0, -3, 0, -3, 0, -4, -2, -4, -4, 0, -1, -4, -1, -1, -2, -3, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -2, -3, 0, -3, 0, -4, -3, -2, -2, -4, -5, -1, -4, -1, -3, -3, -3, 1, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, -2, -2, -1, -1, -3, -2, -2, 0, -4, -3, -4, -1, -1, -4, -3, -4, -1, -4, 0, 0, 0, -2, -2, -1, -1, 0, -1, -2, -1, -2, -1, -1, -2, -2, 0, -2, -2, -1, 0, 0, -3, -2, -1, -4, 0, -4, -4, -3, -1, 0, -3, -3, -1, -3, -2, 0, -1, -1, -2, -2, -1, 0, 0, 0, 0, -1, -1, -3, -2, 0, -2, -4, -2, -1, -2, 0, -2, -2, -1, -1, -1, -2, 0, -2, 0, -3, -2, -3, -3, 0, -2, -2, 0, -1, -1, 0, -3, -3, -3, -2, -2, 0, 0, 0, -2, -3, -3, -5, -5, -3, -2, -2, -2, -1, -2, -1, -3, -3, -3, -3, -2, -2, 0, 0, -1, 0, -1, -3, -2, -4, -1, -1, -2, -3, -1, -3, -3, -5, -5, -2, -1, -1, -1, -3, -4, -3, -3, -3, -2, 0, 0, 0, -2, 0, -3, -1, 0, 0, -4, -4, 0, -1, -2, -1, -3, -4, -3, -5, -1, -3, -1, -2, 0, -1, 0, -4, 0, -1, 0, 0, 0, -2, -1, -1, -1, -3, 0, -3, 0, -3, -1, 0, -1, -1, -2, -4, -4, -4, -5, -2, -3, -1, -3, -1, 0, -2, 0, 0, -4, -1, 0, -2, 0, -1, 0, -1, 0, 0, -2, -3, 0, -3, -1, -4, -5, -4, -3, -2, -4, -2, -1, -2, -1, 0, 0, -1, -1, 0, -2, -1, -3, -3, 0, -3, 0, -1, 0, 0, 0, -2, 0, -1, 0, -1, -2, -5, -3, -5, -2, 0, -1, -2, -3, -2, 0, -2, -2, -1, 0, -2, -3, 0, 0, -1, -2, -1, 0, -2, 1, 0, 0, -3, 0, 0, -4, -5, -2, -4, -5, -1, 0, 0, 0, 0, -1, -1, 0, -2, 0, -1, -2, 0, 0, 0, -3, -1, 0, 0, -1, -2, -2, 0, 0, 0, -2, -5, -2, -4, -1, 0, 0, 0, -1, -2, -1, -2, 0, -3, -2, -1, 0, 0, -1, -2, -3, -1, 0, -2, 1, 0, -1, -3, -3, -2, -4, -3, -5, -2, -5, 0, -1, -1, 0, -3, 0, 0, 0, 0, -3, 0, -1, 0, -1, -3, -3, -2, 1, -1, -2, -2, -2, -3, -1, -3, -4, -4, -4, -3, -4, -1, 0, 0, -2, -3, 0, -2, 0, 0, -1, 0, 0, -2, 0, -3, -3, 0, -1, 1, 0, 0, 0, 0, -1, -1, -2, -3, -2, -4, -4, 0, -2, 0, 0, 0, -1, 0, -1, -3, -1, -3, -1, 0, -2, -1, -4, -2, -1, 0, -1, -1, 0, -2, -1, -3, -4, -3, -4, -1, -2, 1, -1, 0, 0, -3, -1, 0, 1, 0, 0, -1, -3, -1, -3, 0, -1, 0, -3, 0, -1, -3, -1, -2, -4, -4, 0, -2, -2, -4, -4, 0, -2, 0, -2, 0, -2, -2, -1, -1, -3, 0, -2, 0, -3, -1, -4, 0, 0, 0, 0, 0, -1, -3, -2, -2, -2, -2, -3, -3, -2, 0, 0, -4, -1, 0, -2, -1, 0, -2, -1, 0, 0, 0, -2, 0, -2, 0, 0, 0, -1, -3, 0, -4, -2, -2, -3, -2, -5, -4, 0, -3, -1, -1, -2, 0, -1, -1, 0, -1, 0, 0, -3, 0, -2, 0, -4, -3, 0, -2, -3, -2, -1, -2, -3, -3, -2, -5, -2, -1, -3, 0, 0, -2, -3, -1, -3, 0, 0, 2, -1, -2, -1, 0, -1, -2, -1, -3, -3, 0, -3, 0, -2, -2, -3, 0, -2, -4, -3, -1, -2, -3, 0, 0, 0, -1, -2, 1, 0, 0, 0, 0, -2, 0, -3, 0, -3, -1, -3, 0, 0, 0, -1, -3, -3, -2, -3, -4, -4, -3, -3, 0, -2, 0, 0, -1, 0, -1, -1, -2, -1, 0, -1, -1, 0, 0, -1, -4, -1, -1, -4, -4, -4, -2, 0, -2, -3, 0, -3, -1, -3, -2, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -2, 0, -2, -2, 0, -3, -4, -3, -1, -2, -3, -3, 0, -1, -2, -4, -1, 0, 1, -1, -1, -2, 0, -1, 0, -2, 0, 0, 0, -2, -1, -1, -1, -1, -1, 0, -1, -1, -1, -2, -2, 0, 0, -3, -3, -4, -2, 0, 0, -1, -2, -2, 1, 0, -1, 0, 0, 0, 0, -2, 0, -1, -2, -2, -1, -1, 0, 0, -1, -3, 1, -2, -1, -2, -1, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, 0, -1, -1, 0, -1, -2, 1, 0, 0, -2, 0, -1, 1, 0, 0, 0, -1, -2, -1, -1, -1, -1, -5, -4, -4, 0, -2, -2, 0, 3, 3, 2, 3, 3, 3, 4, 1, 4, 1, 4, 2, 0, 1, 2, 0, 0, 1, 0, 1, -1, 2, 1, -2, -1, -4, -2, -1, 0, 0, 1, 2, 1, 2, 5, 2, 3, 2, 2, 5, 4, 2, 3, 1, 3, 3, 2, 0, 2, 0, 0, -1, 0, -2, -2, 0, 0, 0, 0, 1, 2, 2, 3, 5, 3, 4, 4, 4, 4, 2, 4, 5, 4, 3, 3, 2, 3, 1, 1, 0, 0, 2, 0, -2, -2, -1, 1, 2, 3, 1, 3, 1, 3, 3, 5, 1, 5, 2, 3, 5, 2, 4, 6, 5, 6, 2, 4, 3, 0, 0, 0, 0, 3, -2, 0, 1, 0, 3, 4, 4, 2, 3, 1, 0, 1, 1, 3, 3, 5, 4, 4, 3, 2, 3, 5, 1, 4, 3, 2, 3, 1, 0, 5, -1, 0, 1, 3, 2, 4, 1, 1, 3, 0, 2, 1, 2, 1, 2, 2, 4, 3, 2, 5, 5, 1, 3, 4, 2, 1, -1, 0, 3, 2, 0, 1, 0, 0, 4, 3, 1, 2, 3, 4, 4, 0, 0, 0, 0, 0, 2, 3, 3, 3, 3, 3, 1, 3, 2, 1, 2, 1, 2, 1, 0, 0, 0, 3, 4, 4, 5, 2, 5, 2, 4, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 3, 2, 1, 3, 1, 1, 0, 0, 1, 1, 1, 2, 2, 1, 2, 2, 3, 3, 3, 1, 0, 0, -1, 0, -2, -2, 0, 0, 0, 3, 1, 1, 3, 1, 0, 2, 3, 4, 0, 1, 2, 3, 3, 3, 1, 2, 3, 2, 3, 1, 1, 0, 0, -2, -2, -2, 1, 0, 0, 1, 0, 2, 0, 0, 0, 1, 2, 4, 1, 1, 2, 1, 3, 1, 5, 3, 4, 5, 2, 3, 2, 0, -3, -2, -2, 0, 0, -2, 1, 0, 4, 2, 1, 0, 3, 0, 3, 3, 1, 1, 0, 1, 5, 5, 4, 3, 3, 3, 0, 1, -2, -1, -3, -3, -3, -3, -1, 1, -1, 1, 1, 1, 0, 4, 1, 1, 2, 0, 1, 2, 4, 2, 4, 2, 3, 1, 4, 3, 0, -2, -1, -3, -3, -6, -3, -3, -1, -1, -2, -2, 0, 1, 0, 3, 0, 3, 0, 0, 0, 0, 2, 2, 5, 3, 0, 2, 0, 1, 2, 0, -1, -2, -3, -4, -4, -5, -2, -6, -5, -2, -2, 0, -1, 2, 2, 1, 2, 0, -1, 0, 1, 2, 4, 1, 3, 2, 0, 3, -1, 1, -3, -1, -6, -7, -6, -6, -5, -3, -5, -4, -1, -1, 0, 1, 1, 0, 2, 2, 0, 0, 4, 4, 1, 2, 1, 1, 1, 0, -1, 0, -2, -4, -7, -7, -7, -7, -8, -6, -8, -4, -4, -2, -1, 2, 0, 2, 1, 3, 1, 3, 2, 0, 5, 2, 0, 2, 2, 2, 0, 0, -2, -4, -6, -5, -5, -5, -4, -8, -9, -7, -3, -2, -1, -1, 0, 2, 0, 2, 0, 2, 2, 3, 5, 4, 2, 2, 2, 0, -1, -2, -1, -5, -6, -3, -3, -5, -4, -7, -4, -5, -4, 0, 0, 0, 1, 1, 1, 1, 0, 1, 0, 2, 5, 3, 5, 4, 1, 1, 2, 0, -2, -4, -5, -3, -3, -5, -6, -4, -5, -1, 0, 0, 3, 1, 0, 2, 4, 3, 1, 0, 0, 4, 3, 4, 4, 4, 3, 3, 1, 0, 0, -2, -3, -4, -2, -2, -4, -1, 0, 1, 0, 0, 4, 2, 3, 3, 1, 0, -1, 0, 1, 2, 2, 5, 1, 3, 1, 0, 1, 0, 0, 0, -2, -1, 0, -2, -2, 0, -2, 0, 0, 0, 1, 3, 2, 0, 1, 3, 0, 2, 4, 3, 2, 5, 5, 3, 5, 1, 3, 1, 3, 0, 0, 0, -1, 0, 1, 0, 0, 0, 2, 0, 2, 3, 1, 1, 0, 2, 0, 1, 0, 3, 6, 5, 3, 5, 3, 2, 1, 1, 0, 0, 0, -2, 0, 0, 0, -2, -1, 0, 0, 3, 4, 4, 0, -1, 1, 0, 0, 0, 4, 2, 2, 4, 4, 4, 4, 5, 1, 3, 1, 0, 0, 1, -1, 0, 2, 0, 0, 0, 0, 3, 1, 0, -1, -1, 2, 3, 0, 0, 4, 4, 2, 4, 5, 2, 3, 4, 2, 0, 2, 3, 4, 1, 1, 2, 0, 1, 2, 0, 1, 3, 0, 0, 1, 0, 0, 2, -1, 2, 2, 5, 2, 3, 3, 4, 1, 4, 1, 3, 3, 3, 3, 4, 4, 1, 1, 4, 4, 2, 0, 2, 2, 2, 0, 2, 0, 0, -1, -1, 2, 1, 1, 2, 3, 3, 2, 2, 3, 1, 1, 0, 4, 0, 4, 2, 2, 4, 3, 4, 4, 5, 4, 3, 3, 1, 0, 0, 0, 0, 2, 3, 2, 3, 2, 3, 3, 2, 1, 4, 4, 4, 1, 3, 3, 6, 6, 3, 3, 2, 2, 2, 1, 0, 3, 1, 0, 0, -3, 0, 1, 3, 1, 4, 4, 2, 3, 5, 3, 0, 1, 3, 3, 2, 5, 4, 6, 6, 4, 5, 3, 2, 2, 0, 2, 1, 0, 1, -3, -3, 0, 0, 0, 0, 0, 1, 0, 4, 2, 5, 0, 5, 3, 3, 5, 5, 5, 6, 6, 4, 2, 0, 0, 0, 0, 2, 2, 1, -1, 0, 0, 0, 0, -2, 0, 0, 0, -1, 1, 2, 0, 1, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, -2, -1, 0, 2, -2, 0, -2, -3, 0, 0, 0, -1, -1, 1, 0, 2, 0, 2, 0, 0, 2, 3, 3, 0, 2, 3, 0, 2, 1, 0, -1, 1, 1, 1, 1, 0, -2, 0, -2, 0, 0, 0, 2, 0, 0, 3, 0, 0, 0, 2, 1, 2, 2, 2, 1, 2, 1, 0, 2, 1, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, 1, 0, 1, -1, 1, 0, 2, 3, -1, 0, 3, 0, 0, 0, 1, 2, 0, 2, 3, 0, 1, 1, 2, 1, 2, 0, -2, -2, 0, 0, 1, 0, 2, 0, 0, 0, 1, -1, 0, 1, 2, 3, 0, 0, 1, 0, 0, 0, 0, 1, 2, -1, 0, -1, -1, 1, 1, -2, 1, 1, 1, 0, 0, 2, 1, 0, 1, -1, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 2, 1, 1, 2, 1, 2, 0, 2, -1, 0, 0, 2, 0, 0, -1, 1, 0, 0, 0, 0, 1, -2, 0, 0, -1, -1, 2, 0, 0, 0, 2, -1, 1, 0, 0, 0, 1, 1, 0, 1, 1, 1, 0, -1, 2, -1, 0, 1, 1, 0, 1, -2, 1, 1, 0, -2, 1, 1, 1, 0, 1, 0, -1, 1, -1, -2, 1, 1, 0, 2, 0, 2, 0, 0, 2, 1, 1, 2, 0, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, 1, 2, -1, 0, 0, 0, 0, 0, 2, 1, 1, 3, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 1, 0, 0, 0, 2, 1, 1, 2, 0, -1, 0, 0, 0, 3, 0, 3, 1, 0, 0, 0, -1, -2, 0, -2, -2, -3, -2, 0, -1, 1, 0, 1, 0, 0, 0, -2, 0, 2, 0, 2, 0, 2, 2, 0, 2, 0, 0, 0, -1, -1, 1, 0, 0, -3, 0, -4, -2, 0, 0, -2, 1, 1, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -4, -3, -4, -3, -2, -2, -1, -2, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, -2, -3, -4, -4, -4, -2, -5, -2, -2, 0, -2, -2, 0, -2, -1, 1, -2, -1, -1, 0, 1, 2, 0, 2, 0, 1, 1, -1, 0, -1, -1, -2, -1, -4, -2, -5, -5, -1, -1, -2, 0, -2, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, -3, -2, -1, -4, -4, -6, -4, -4, -2, -4, -4, -1, -2, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 1, 0, 1, -1, -3, -5, -5, -4, -2, -5, -1, -3, -3, -3, -2, -1, 0, -1, 0, -1, -1, 1, -1, 0, 1, 2, 0, 3, 1, 1, 2, -1, -1, 0, 0, -2, -3, -3, -1, -1, -3, -4, -4, -4, -1, -1, -1, 0, -2, 1, 0, -1, 1, 1, 2, 1, 2, 1, 1, 2, 1, 0, 1, 0, -3, -1, -2, -1, -2, -1, -4, -2, -1, -1, 0, -2, 2, 1, -1, -1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -3, -1, -2, -1, -2, -2, -4, -2, -3, -1, 1, 2, -1, 0, 0, -1, 1, 1, 0, 0, 1, 0, 2, 1, 1, 1, 0, 0, 0, 0, -2, -2, 0, -1, -2, -3, 0, -2, -2, 1, 0, 0, -1, 0, -1, -2, 1, -1, -1, 0, 0, 1, 1, 2, 0, 0, 1, 2, 1, 0, 1, 0, 0, -1, -1, -2, -1, -2, -1, -1, -1, 0, -1, 2, -2, -1, 1, 2, 0, 0, 1, 1, 0, 3, 2, 3, 1, 0, 0, 3, 0, -2, -2, 0, 0, 1, -2, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, -1, 3, 0, 0, 0, 0, 4, 3, 2, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 1, -2, -1, 0, 0, 0, 0, 1, 1, 0, 2, 3, 0, 0, 0, 0, 1, 1, 1, 1, -1, 1, 1, -1, -1, -1, 0, -1, -1, 1, 1, -1, 0, -1, 0, 0, 0, 1, 2, 2, 2, 0, 1, 1, 2, 1, 0, 1, 0, 0, 2, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 1, 0, 2, 0, 3, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 3, 0, 2, 1, 1, 2, 1, 0, 0, -1, -1, -1, 0, 0, -2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 1, 1, 3, 3, 0, 2, 2, 2, -1, 0, -1, 0, 0, 0, 0, 2, 2, 1, 0, 0, 1, 0, 1, 0, 2, 1, 1, 0, 3, 1, 1, 2, 3, 1, 0, 3, 1, 0, 1, 1, 1, -1, 0, 0, -2, -1, 1, -1, 0, 0, 2, 0, 3, 3, 2, 1, 1, 1, 3, 3, 0, 3, 3, 1, 0, 2, 1, 0, -2, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 1, 1, 1, -1, 1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, -1, 1, 1, -2, 0, -1, 0, -1, -1, 1, 0, 0, -1, -1, 1, 0, -1, -1, 0, 2, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, -1, -1, 1, 1, -1, 0, 0, 0, 0, 0, -1, 1, 0, 1, -1, 0, 0, -1, 0, 1, -1, -1, -1, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 2, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 2, -1, 0, 0, -2, -1, 0, 0, 1, -1, 1, 1, -1, 0, 0, 0, 0, -1, -1, 1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 2, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, -1, -1, -1, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 1, 0, 1, -1, 0, 0, 1, 0, 1, 0, 0, 1, 2, 0, 0, 0, 1, 0, -2, 0, 1, 0, 0, 1, -1, 1, -2, -1, 0, 1, 1, 1, 1, 0, 1, -1, -2, 0, -1, 1, 0, 2, 1, 0, 0, 0, -2, 0, 1, -2, 0, 0, 0, 1, 0, -1, 0, -1, 1, -1, -1, -1, -1, 0, 0, -1, -1, 1, -1, 0, 0, -1, 0, 1, -1, 0, 1, -1, -1, 0, 0, 1, 2, 0, 0, 0, 0, 1, -1, -1, 1, 0, -1, 0, 0, 1, 0, -1, 0, 0, -2, 1, -1, 1, 1, 1, 0, -1, 1, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, -1, 1, 0, 0, -1, 1, 1, 0, 1, 1, 0, 0, -1, 0, 1, 0, 1, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -1, 1, -1, -1, -1, 0, -1, -2, -1, 1, 0, 1, 0, 1, 1, -1, 1, 1, 0, -1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, -1, 1, -1, 2, -1, -1, 0, 0, -2, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, -1, 1, -1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, 1, -1, -1, -1, 0, 1, 0, 0, 0, 1, -1, -1, 0, -1, -1, 1, -1, 0, 0, -1, 1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, -1, 0, -1, 1, 0, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, -1, 2, 1, -1, 1, -1, 0, 1, 0, 0, 0, -1, 0, -2, 0, 1, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, -2, 0, 0, -1, -1, 1, 0, -2, 1, 1, -1, 1, 1, 1, 0, 1, 1, 0, 0, 1, -1, 0, 1, 1, 1, 0, -1, 0, 1, 0, -1, -2, -1, 0, -1, 0, 0, -1, 1, -1, 1, -1, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 1, -2, 1, 1, -1, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, 1, 1, -1, -1, -2, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, 0, 1, -2, -1, -1, -1, -1, 1, 1, -1, -2, -1, 0, -1, -1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 1, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, -2, 0, -1, -1, -2, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 1, -1, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 1, 1, 0, 1, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 0, 1, 1, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, -1, 0, 2, 0, -1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 2, -2, 1, -1, 1, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, 1, -1, 0, -2, -1, 0, -1, 1, -1, -1, -2, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 2, -1, 1, 2, -1, 0, 0, 0, 1, 0, -1, 0, 1, -1, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, -2, 0, 0, -2, 0, 0, 0, 1, -1, 0, 1, 2, 0, 1, -1, 1, -2, 1, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -6, -2, -4, -4, -3, -1, -2, -2, -1, -3, -1, 0, 0, -2, -1, -1, -3, -2, 0, -1, 0, 0, 0, 0, 1, 2, -1, -1, -1, 1, -2, -3, -4, -3, -2, -2, -4, -2, 0, -1, 0, -1, 0, -1, -2, 0, 0, 0, 1, -1, 0, 0, 1, 2, 2, 2, 0, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, 2, 1, 0, 3, 0, 1, -1, 1, 1, 2, 3, -1, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, -1, -1, -1, 2, 0, 0, -1, 1, 2, 0, 3, 3, 0, 3, 2, 3, 1, 2, 4, 0, -3, -1, 0, -2, -1, 0, -2, 0, -2, -1, 0, 1, 0, -1, 0, -1, 1, 2, 0, 1, 3, 2, 3, 1, 0, 0, 2, 1, 4, -2, -2, -1, -1, 0, 1, 0, -1, -1, -2, -2, -1, 0, -1, 0, -2, -1, 1, 0, 1, 2, 0, 4, 1, 1, 3, 0, 1, 0, 4, 0, 0, -2, 1, -1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 0, 0, 2, 2, 0, 0, 2, 1, 2, 1, 0, 3, 5, 0, -1, -1, 0, 0, 0, 0, 2, 1, 1, -1, 1, 0, 2, 2, 1, 0, 1, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, 3, 3, -2, -1, 0, 1, 1, 2, 0, 0, -1, 0, 0, 1, 0, 1, -3, 0, -2, 1, 0, 1, 1, 3, 2, 1, 0, 0, 1, 0, 3, 2, -3, 0, 0, 0, 0, 0, 1, 0, 1, 0, 3, 2, 2, 0, 0, 1, 2, 0, 1, 2, 3, 0, 0, 0, 1, 3, 1, 0, 5, 5, -1, -2, -1, -1, 1, 0, -1, 2, 2, 1, -1, 0, 0, 0, 0, 1, 0, 2, 2, 1, 0, 1, 3, 1, 0, 3, 0, 4, 5, 2, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, -1, -2, -2, 1, 1, -1, 2, 3, 3, 2, 1, 3, 0, 2, 1, 3, 4, 5, 3, 3, -2, 0, 0, 1, -1, -3, -1, -2, -2, 1, 2, 1, 0, -1, 0, 0, 0, 2, 0, -1, 2, -1, 0, 0, 0, 3, 4, 6, 2, 4, -2, 0, -1, 0, 1, 0, 0, -1, -2, -1, 0, 0, 1, 0, 0, 0, 0, -2, -2, 0, -2, 0, -1, 1, 0, 2, 2, 1, 2, 3, -3, -1, 0, 0, -1, 0, 0, -1, 1, -1, -1, 0, -1, 0, 0, 0, 1, 0, -1, -3, -2, -3, -3, 1, 2, 2, 3, 1, 5, 2, 0, 0, 0, 1, -2, -3, 0, -1, 0, -2, 1, -2, -1, 0, 1, 0, 0, -1, 0, -1, -5, -3, -3, -2, -1, 3, 1, 1, 4, 2, -2, 0, 0, -1, 1, -2, 0, -1, -1, -2, 0, 0, 0, 1, 2, 1, 2, 1, 0, -1, -2, -4, -1, -3, -2, 0, 2, 4, 2, 4, -2, 0, -1, 1, 1, -2, -2, 0, -2, 1, 0, 1, 1, 1, 0, 2, 2, 1, 0, -4, -3, -1, -2, -1, 0, 0, 0, 1, 4, 2, -1, -1, 0, -1, 0, 0, -2, -3, -1, -2, 0, 0, -1, 0, 1, 2, 1, 1, -1, -3, -1, -1, 0, 1, 1, 1, 4, 1, 3, 2, -2, 0, 0, -2, 0, 0, -1, -1, -3, -1, 0, 0, 0, -1, 2, 3, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 3, 3, 1, 4, -4, 0, 1, 1, 1, -1, 0, -2, 0, -2, -1, 0, 2, 0, 0, 2, 1, 3, 0, 1, 0, 1, 0, 0, 2, 0, 1, 2, 1, 4, -2, -1, 0, 0, 1, 2, 0, 0, -2, -4, -2, 0, 1, 1, 0, 3, 3, 3, 1, 1, 1, -1, 0, 3, 4, 0, 0, 2, 3, 3, 0, -3, 0, 0, 0, 0, 1, 0, -2, -3, -1, -1, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 2, 2, 1, 0, 4, 3, 4, -1, 0, 2, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 2, 4, 0, 0, -1, 0, 2, 0, 2, 0, 1, 1, 2, 2, 0, 0, 0, 0, 2, 1, -1, -1, -3, 0, -2, 0, -1, 1, 0, 0, 0, 4, 1, 1, 3, 0, 2, 1, 0, 3, 2, 2, 1, 2, 0, 0, 1, 0, 1, 0, 0, -1, -2, -2, 0, -3, -2, 0, 0, -1, 0, 2, 1, 0, 2, 0, 2, 1, 4, 2, 1, 3, 1, 4, -1, -2, -1, 0, 0, 2, -1, 1, 0, 0, 0, 0, -3, -2, 0, -2, 0, 1, 3, 1, 4, 2, 0, 1, 4, 0, 0, 2, 2, 3, -1, 0, -1, 2, -2, 0, -1, -1, 1, 0, -3, -3, -1, -1, -1, -1, -1, 3, 3, 3, 2, 3, 0, 2, 0, 1, 1, 1, 0, 1, -4, 0, -1, 0, 1, -1, -1, -2, -2, -1, -1, -3, -3, -1, -1, 0, -1, 0, 2, 2, 0, 1, 2, -1, 1, -1, 0, 1, 2, 2, -3, -1, 0, -2, -2, -1, -1, -1, 0, -1, 0, 1, 1, 0, 1, -2, 0, 0, 0, 3, 1, 1, 1, 0, 0, 0, 0, 0, -1, 0, -1, -2, 1, 0, 0, 0, 0, 0, -1, -2, -1, -1, 0, -2, -1, 0, -2, 0, -2, -2, -2, 0, -1, 1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 1, 0, -2, 0, 0, 0, 0, -2, -2, -2, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, -2, 1, 0, -1, 0, 1, -1, 0, 1, -2, 0, 0, -2, -1, 0, -1, -1, 0, -2, -2, -2, 0, -2, -1, -1, 0, 0, 0, -2, -2, 1, 0, 0, 0, 0, -2, -1, -1, 0, -1, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, -2, 1, 1, -2, 0, -1, -1, 0, -1, 1, 0, 0, -2, -1, -3, 0, -2, -1, -1, 0, 0, -1, -3, -1, -2, 0, -1, -1, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, -3, -2, 0, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 1, -1, 0, 0, 0, -1, -3, -2, -3, 0, 0, 0, -3, 0, -3, 0, 0, -1, -3, 0, 0, -1, 0, -1, -2, 1, 0, 1, 0, 0, -1, -1, 0, 0, -2, 0, -2, 0, 0, -1, -2, -3, 0, 0, 0, -1, 0, -2, -3, -2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, -2, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, 0, 0, 0, -2, 0, -1, 0, -2, -2, 0, -2, 1, -1, 1, -1, 0, -1, -2, 0, 0, -1, -1, -2, 0, 0, 1, -2, -1, -1, -2, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, -2, -1, -2, 0, 0, -2, -2, 0, 0, -2, 1, 0, -3, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, -3, 0, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, -2, 1, 0, 0, 0, 1, -1, -3, -1, 0, 0, 0, 1, -2, 0, 0, -1, 0, 0, 0, 1, -2, 1, -2, -1, 0, 0, 0, -1, 0, -2, 0, 0, -2, -1, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, -2, 0, 0, 0, 0, -2, 0, 0, 0, -2, 0, 1, -2, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, -1, -1, 1, -1, -2, -1, -1, 0, -2, 1, -2, 0, -1, -1, 0, 0, -2, 0, -2, -2, -2, 0, 0, -1, 0, 1, 0, -2, 0, -2, 0, 0, -3, 0, -2, -2, 0, 0, -2, 1, -2, -1, -1, 0, 0, -2, 0, -3, -2, -1, -1, -2, 0, 0, 0, -2, -2, 0, 0, 0, -1, 0, -2, -3, -2, -2, 0, -1, 0, -1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, -2, 0, -1, -1, -2, 0, -1, -2, 0, -2, -2, -1, 0, 0, -1, -2, -1, 1, -1, 0, 0, 0, 1, -2, -2, -1, -3, 0, 0, 0, -1, -2, 0, 0, -1, -1, -2, -2, -1, 0, 0, 0, -1, 0, 0, 1, -2, 0, 0, 0, -1, 0, 1, -1, -2, 0, 0, 0, -1, 0, -2, -2, -2, 0, -2, -3, -2, -2, -2, 0, -1, 0, -1, 0, 0, 0, 0, 1, 0, -2, -1, -2, 0, 0, 0, -2, 0, 0, 0, -1, 0, -2, -1, 0, 0, -2, -2, 0, 0, 0, -3, -3, -1, -2, 0, 0, 0, 0, 0, 1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, -1, -3, -2, -1, -1, -1, -2, -3, -2, -3, 1, -1, -2, 0, 0, -1, -1, 1, -2, 0, 0, -3, 0, 0, 0, 0, -2, 0, 0, -2, -2, 0, 0, -2, -1, -1, -1, 0, 0, 0, -2, 1, -2, -1, -1, -1, 0, -1, -2, 0, 1, -2, 0, 0, 0, 0, -2, -2, 0, -2, 0, 0, 0, -2, -1, -2, 0, -1, 0, -2, 0, -2, 0, 0, -1, 1, -1, 1, 0, -3, -2, -1, -2, 0, -2, -1, -3, -1, 0, 0, -3, 0, 0, -2, -2, -1, -2, -2, -2, 0, 0, 1, -2, -1, -1, 1, 0, -1, -1, 0, 0, -3, 0, -1, 0, -1, -2, 0, -1, 0, 0, -1, -2, -3, 0, -1, -2, -2, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, 0, -2, -3, 0, -3, 0, -3, 0, -2, -2, 0, 0, -2, 0, -1, 1, -1, 0, 0, -1, 0, 0, -2, 0, 0, -1, 1, -1, -3, -2, -1, -1, 0, -1, -2, 0, -3, 0, -3, -2, -1, 1, 0, -2, -2, 1, -1, 0, -2, 0, -1, 1, 0, -2, -1, -2, 0, 0, -2, 0, 0, 0, 0, -2, -1, 0, -2, -1, 0, 0, 1, 0, -1, 0, -1, 1, 1, 0, -1, 0, -2, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, -1, 0, -2, -2, -2, 0, 0, 0, -2, 0, -2, -3, -2, -2, -2, -3, -3, -2, -2, -1, 0, -2, -3, 0, 0, 0, 0, -2, -1, 0, -3, -2, -2, 1, 0, 0, -2, 0, -3, 0, 0, 0, 0, -3, 0, 0, 0, 0, -3, 0, 0, -3, 0, -1, -3, 0, -2, -2, -2, -2, -1, 0, -2, 1, 0, -1, 0, 0, -1, -1, -2, 0, 0, -2, -2, -1, -1, 0, -1, -1, 0, -3, -2, -2, -1, -1, 0, 0, 0, -2, -2, 0, -1, 0, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, -1, 0, -2, -2, -3, 0, 0, 0, 0, -2, 0, -1, -3, 0, -2, 1, -1, -2, 1, -1, 0, 0, -1, -1, -1, 0, -2, -2, 0, -1, 0, -3, -1, -2, 0, -2, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -3, -3, -1, 0, -2, -3, -1, -2, -1, -2, 0, 0, -3, -1, 0, -1, 1, 0, 1, 0, -1, -1, 0, 0, -1, 1, 0, -1, 0, -1, -2, -3, -2, -2, 0, 0, -2, 0, -1, -2, -1, -2, -1, 0, 0, -1, -1, -1, -2, 0, -2, 0, 0, -1, 1, 0, 1, 0, -1, -1, -3, 0, 0, -3, -3, 0, -1, -2, -2, -2, -2, -2, -2, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, -3, -1, -2, -3, -2, -3, -1, 0, 0, 0, -1, -2, -2, 0, -2, 0, 0, 0, 0, 0, -1, -2, -2, -1, -2, 0, 1, -1, -2, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, -1, -1, -1, -1, 0, -2, 0, -3, -1, -1, 0, 0, -2, -2, 0, -1, -1, 0, -1, -2, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, -2, -3, -2, 0, -1, -2, 0, 1, 1, -1, 1, 1, -3, 0, 0, -2, 0, -3, 0, 0, -2, 1, 0, 0, -2, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, -1, 0, 0, -1, -2, -1, -2, 0, -1, -1, -2, -3, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 0, 1, 0, 1, -1, 0, 1, 1, 0, -2, -3, -3, -2, -1, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, -2, -2, 0, -2, 0, 0, 0, -1, 1, 0, 1, 1, 1, -1, 1, 0, 0, -2, 0, -3, -1, -2, 0, 0, 1, -2, 0, -2, -2, -2, 0, -2, 0, 1, -2, 0, 1, -1, 0, -2, 0, 0, 0, -1, 0, 0, -2, -1, -3, -2, -3, -1, 0, 0, -1, -2, -1, 0, -1, 0, -2, 0, -2, 0, 0, 1, 0, -2, 0, 1, 0, 0, 0, 1, -1, -2, 0, -3, 0, -3, 0, -1, -1, -1, -1, -2, 0, -1, 0, -1, 0, -1, 0, -1, -2, -1, -1, 0, 0, -2, 1, -1, -1, 0, -1, -3, 0, -3, 0, 0, -3, -1, 0, -1, 0, 0, -2, 0, 0, 0, -2, 0, -2, 0, -1, 0, -1, 0, 0, -1, 0, -1, 0, 1, 1, -1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, -1, -2, -1, -3, -1, 0, -2, 0, -1, -3, 0, 0, 0, 0, 1, 0, -1, -2, -3, -1, 0, 0, -1, 0, -3, 0, 0, -1, -3, -1, -1, -3, -3, 0, 0, 0, -2, 0, 0, -1, 0, -2, 0, 0, 1, -3, 0, 0, -2, 0, -1, -2, -1, 0, -3, -2, -2, 0, -3, -2, -3, -2, -3, -2, -1, -3, -2, -3, 0, -1, -1, -2, 1, 0, 0, -2, -1, -1, -1, 0, 0, -3, -1, -2, -3, -1, 0, 0, 0, 0, -2, -1, 0, -2, -1, -2, -1, -2, -2, -1, -1, 0, 1, -1, -2, 0, -1, 0, -3, 0, -2, 0, 0, -1, -3, -2, -2, 0, -3, -2, -1, -3, -2, -2, 0, -1, -1, -1, 0, 0, -2, -1, 0, 0, 0, 0, -2, -3, -2, -1, 0, 0, 0, -2, -3, -1, 0, 0, -1, -1, 0, -2, -2, 0, 0, -2, -1, -2, -1, 0, -1, 0, -1, 0, -1, 0, -2, -2, -1, -1, 0, -2, -1, 0, 0, -1, -2, 1, 0, -2, 0, -1, -3, -3, 0, -2, 0, -2, -3, -1, -1, 0, 0, 0, 1, -2, -1, -1, 0, -3, -3, -2, 0, -2, -3, 0, -1, -2, 0, -2, 0, -2, -3, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -2, -2, 0, -1, -1, -1, -1, -3, 0, 0, -2, 0, -2, -1, 0, 0, -3, -2, -2, -1, 0, -1, 0, 0, -2, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -2, -2, 0, -2, -2, -1, 1, 1, 0, 0, -2, 0, 0, -1, -2, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 0, -3, -2, 0, -3, 0, -3, -1, -1, -1, 1, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, -2, -1, 0, -2, -1, -1, -1, 0, -1, 0, -3, 0, -3, -2, 0, 0, -2, -1, -1, 0, -1, 0, 1, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, 3, 1, 2, 4, 3, 1, 4, 1, 1, 1, 3, 2, 3, 2, 1, 3, 4, 5, -1, 0, 0, 0, 0, 1, 2, 3, 0, 2, 1, 0, 4, 3, 2, 2, 4, 2, 1, 2, 4, 4, 1, 4, 4, 4, 3, 5, 2, 5, 2, 1, 2, 2, 2, 0, 3, 0, 2, 1, 0, 4, 2, 2, 3, 3, 3, 2, 3, 1, 4, 2, 1, 2, 4, 3, 1, 4, 5, 2, 1, -1, 0, 0, 0, 2, 3, 1, 0, 3, 3, 3, 3, 3, 1, 4, 3, 4, 2, 2, 1, 1, 2, 3, 2, 2, 3, 4, 1, 4, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, 1, 4, 0, 0, 3, 4, 2, 4, 4, 2, 3, 3, 2, 2, 3, 1, 1, 5, 2, 3, 0, 3, 0, 2, 0, 1, 1, 2, 0, 1, 0, 3, 4, 0, 3, 3, 0, 3, 3, 3, 0, 4, 1, 1, 1, 4, 1, 5, 2, 3, 0, 0, 1, 0, 3, 2, 3, 0, 1, 0, 3, 2, 0, 1, 0, 2, 0, 1, 2, 0, 4, 2, 1, 0, 0, 5, 2, 4, 5, 2, 0, 4, 2, 0, 3, 1, 3, 2, 1, 0, 0, 3, 3, 1, 2, 0, 0, 0, 0, 2, 2, 0, 2, 1, 3, 2, 3, 3, 3, 6, 2, 3, 0, 2, 3, 0, 2, 2, 3, 1, 0, 1, 2, 2, 0, 1, 1, 1, 0, 1, 0, 1, 0, 3, 1, 5, 2, 5, 6, 6, 0, 0, 3, 0, 0, 2, 0, 1, 1, 1, 3, 1, 0, 0, 0, 2, 0, 1, -1, -1, 0, 1, 2, 3, 3, 3, 5, 2, 6, 6, 3, 2, 2, 3, 1, 3, 1, 3, 2, 2, 0, 1, 0, 1, 1, 1, 0, 1, -1, -1, 0, 0, 1, 3, 1, 5, 3, 2, 3, 5, 0, 2, 1, 0, 2, 1, 3, 2, 2, 3, 0, 2, 2, -1, 0, 0, -1, -1, 0, -2, -2, -1, 1, 2, 2, 3, 5, 3, 3, 4, 1, 2, 1, 1, 1, 1, 1, 0, 2, 4, 2, 0, 0, 2, 0, 0, -1, -4, 0, -1, -3, -3, -1, 0, 1, 0, 1, 2, 5, 4, 0, 2, 1, 0, 0, 1, 1, 2, 1, 3, 0, 0, 0, 0, -2, -2, -4, -2, -1, -4, -2, -3, 0, -1, 0, 1, 3, 5, 4, 5, 2, 1, 0, 0, 0, 2, 3, 0, 1, 2, 2, 0, 1, -1, -1, 0, 0, -4, -1, -2, -3, 0, -2, 0, 0, 0, 3, 3, 2, 5, 0, 2, 0, 2, 1, 1, 2, 1, 2, 4, 3, 2, 1, 0, -1, -2, -1, -2, -5, -2, -2, -3, 0, 0, -1, 2, 1, 5, 6, 2, 2, 0, 3, 2, 1, 2, 0, 3, 2, 4, 4, 3, 0, 0, 0, -1, -3, -1, -4, -1, 0, 1, -1, 1, 0, 1, 5, 3, 5, 4, 1, 2, 2, 1, 3, 3, 3, 3, 2, 2, 0, 0, 0, 0, -3, -2, -3, -1, -2, 0, -1, -1, 0, 2, 0, 3, 1, 1, 2, 5, 0, 2, 0, 2, 2, 0, 2, 2, 2, 3, 2, 3, 3, -1, 0, -2, 0, -3, -3, -3, 0, -1, 2, 1, 2, 1, 2, 3, 6, 2, 1, 2, 1, 2, 1, 1, 4, 3, 2, 4, 1, 1, 0, 0, -1, 0, 0, -2, -1, 0, 1, 0, 1, 0, 0, 2, 3, 2, 4, 3, 2, 0, 3, 1, 0, 4, 2, 3, 0, 2, 1, 2, 2, 2, 1, 1, 0, 0, -2, 0, 0, 0, 1, -1, -1, 4, 2, 2, 4, 3, 2, 0, 1, 2, 0, 0, 2, 2, 3, 4, 0, 3, 3, 1, 0, 0, 1, -1, 0, 0, 0, 1, 1, 0, -1, 1, 4, 2, 4, 1, 2, 1, 0, 1, 3, 4, 2, 0, 0, 4, 2, 1, 3, 0, 1, 0, 1, 1, 0, -1, 3, 2, 0, 0, 1, 3, 5, 4, 5, 2, 1, 3, 2, 2, 4, 2, 2, 2, 3, 0, 1, 4, 2, 1, 0, 3, 0, 0, 1, 0, 0, 0, 2, 2, 1, 3, 5, 5, 2, 4, 3, 1, 0, 0, 0, 2, 3, 3, 2, 2, 3, 0, 2, 2, 3, 2, 3, 3, 3, 1, 1, 2, 0, 1, 1, 1, 2, 4, 2, 4, 1, 2, 0, 0, 1, 1, 3, 2, 0, 2, 0, 0, 3, 0, 2, 3, 4, 1, 2, 2, 2, 2, 1, 3, 0, 0, 4, 5, 4, 2, 2, 2, 3, 1, 0, 0, 1, 3, 1, 1, 2, 0, 3, 4, 0, 4, 4, 2, 2, 4, 0, 3, 0, 0, 4, 0, 3, 2, 3, 4, 1, 0, 0, 2, 1, 0, 2, 1, 3, 0, 0, 3, 3, 3, 3, 3, 3, 4, 2, 3, 1, 2, 3, 1, 1, 1, 3, 3, 5, 1, 1, 0, 0, 2, 1, 1, 1, 2, 4, 2, 3, 2, 3, 3, 2, 0, 3, 1, 3, 0, 2, 2, 1, 0, 2, 3, 1, 4, 3, 3, -1, 2, 2, 2, 0, 0, 1, 2, 1, 0, 2, 0, 0, 3, 0, 1, 1, 2, 0, 0, 1, 3, 1, 0, 2, 2, 2, 3, 2, 0, -4, -3, -4, -4, -3, -5, -7, -7, -4, -2, 0, -1, -4, -5, -3, -2, -1, -3, -3, 0, 0, 0, 2, 3, 3, 2, 2, 5, 7, 6, -5, -3, -1, -3, -2, -5, -5, -3, -4, -4, 0, 0, -2, -3, 0, 0, -2, -2, 0, 1, 2, 2, 4, 3, 3, 4, 6, 4, 7, 5, -5, -3, -4, -4, -3, -2, -3, -2, -3, -2, -1, -3, -2, 0, 0, 0, 0, -1, 0, 0, 1, 4, 3, 4, 3, 5, 5, 5, 5, 5, -3, -5, -2, -2, -2, -2, -4, -4, -2, -1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 1, 5, 3, 6, 7, 4, 7, 6, 6, 7, 7, -5, -4, -2, -2, -4, -1, -4, -2, -4, -4, -1, 0, 0, 2, 1, 0, 1, 0, 2, 4, 1, 6, 3, 7, 8, 4, 7, 7, 8, 7, -2, -2, -4, -1, -3, -2, -2, 0, 0, -4, -2, 0, 1, 2, 0, -1, 2, 0, 1, 2, 5, 5, 7, 6, 8, 5, 7, 9, 8, 6, -4, -2, -2, -1, 0, -2, -1, 0, -2, 0, 0, 1, 2, 0, -2, 0, 2, 0, 0, 1, 1, 3, 2, 4, 6, 6, 6, 6, 8, 11, -4, 0, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, 2, 0, 0, -1, 2, 0, 1, 0, 0, 2, 5, 3, 6, 4, 7, 7, 10, 8, -3, -2, 0, -1, 0, 0, 1, 2, 0, 0, 0, 2, -1, 1, 1, 0, 1, 2, 0, 3, 0, 3, 2, 3, 2, 5, 8, 11, 9, 10, -2, 1, -1, 0, 0, 1, 1, 2, 2, 2, 2, 2, -1, -1, 0, 0, 2, 0, 1, 0, 1, 2, 0, 1, 4, 5, 7, 8, 10, 11, -4, -2, -1, 0, -1, 0, 0, 3, 0, 2, 0, 1, 0, 0, 0, 1, 1, 2, 0, 1, 0, 1, 0, 1, 6, 6, 6, 10, 11, 11, -2, 0, 0, -1, -2, 0, 1, 1, 1, 0, 0, 0, 0, 0, 3, 2, 4, 3, 2, 0, 0, -1, 0, 2, 4, 5, 8, 12, 12, 13, -3, -2, -1, -1, -2, -2, 0, 2, 2, 1, 0, 0, 0, 1, 1, 3, 0, 3, -1, 1, -2, 0, 0, 1, 5, 6, 11, 10, 14, 14, -3, -1, 0, 0, 0, -3, -1, 0, 0, 1, 3, 3, 2, 0, 3, 0, 1, 0, 0, -1, -2, -3, 0, 3, 6, 7, 10, 12, 14, 14, -3, 0, -1, -2, 0, 0, 1, 0, 1, 1, 2, 0, 4, 4, 2, 2, 4, 1, -1, -1, -4, -2, -1, 2, 2, 5, 7, 12, 13, 12, -2, -2, -2, -1, -3, 0, 1, -1, 0, 3, 3, 4, 2, 3, 5, 2, 1, 0, -2, -4, -5, -2, -2, -1, 3, 5, 8, 12, 13, 11, -1, -3, -3, 0, -2, 0, -3, -2, 1, 2, 3, 1, 3, 6, 5, 4, 3, 3, -1, 0, -1, -2, -2, -2, 2, 4, 8, 12, 10, 10, -3, -1, 0, 0, -2, -1, 0, 0, -1, -1, 1, 3, 4, 3, 5, 4, 2, 2, 0, -1, -3, -2, -3, -2, 2, 2, 9, 8, 11, 12, -4, 0, -3, -1, 0, 1, -1, 0, -1, 0, 0, 1, 3, 2, 4, 2, 2, 4, 2, 1, 0, -2, -1, 0, 2, 3, 6, 11, 12, 8, -2, 0, -4, -3, -1, -2, 0, -3, 0, 0, 0, 1, 3, 2, 1, 5, 5, 5, 1, 2, -2, 0, 0, -1, 2, 4, 7, 9, 11, 12, -2, -3, -3, -1, -1, 0, 0, 0, 0, 0, 0, 1, 3, 3, 2, 5, 3, 6, 1, 0, -1, 0, 0, 1, 1, 6, 7, 11, 10, 11, 0, 0, 0, 1, 0, -1, -2, -3, -5, -1, 0, 2, 0, 1, 2, 3, 5, 3, 2, 2, 0, 1, 0, 2, 5, 3, 5, 11, 11, 8, -2, 0, -1, 1, 1, 1, 0, -1, -3, -3, -1, 2, 0, 0, 0, 4, 4, 6, 1, 2, 1, -1, 4, 4, 6, 5, 8, 11, 9, 8, -2, -3, 0, 1, 0, 1, -2, -2, -2, -1, 0, -1, 0, 0, 0, 1, 6, 3, 2, 3, 3, 1, 3, 4, 3, 4, 6, 8, 9, 8, -1, -2, 1, 0, -1, 0, -3, -1, 0, -1, 0, -2, 0, 0, 0, 0, 3, 6, 3, 4, 5, 2, 2, 2, 4, 5, 7, 9, 8, 10, -1, -3, 0, -2, -2, -3, -3, -3, 0, -1, -1, -3, 1, 0, 0, 3, 3, 2, 6, 4, 2, 6, 4, 6, 6, 6, 6, 6, 10, 8, -4, -3, -2, -1, -1, -1, 0, -3, -2, -3, 0, -1, -1, 0, 1, 2, 4, 2, 6, 4, 3, 2, 6, 4, 2, 4, 5, 6, 7, 10, -5, -3, 0, -1, -3, 0, -2, -2, -1, -2, -3, 0, 0, 0, 0, 0, 3, 2, 3, 3, 4, 3, 3, 3, 5, 5, 7, 5, 5, 6, -5, 0, -3, 0, -2, -2, -2, -3, -2, -1, 0, -1, -2, -1, -1, 0, -2, 0, 1, 2, 1, 1, -1, -1, 2, 1, 2, 3, 4, 6, -6, -2, -3, -4, -4, -5, -3, -6, -2, -4, -2, -2, -3, 0, -3, -2, -2, -3, 0, 0, 0, 0, 0, -2, 0, 0, 2, 3, 5, 6, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 1, -2, 1, 1, -2, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, 1, -2, 0, 0, -2, 0, 1, -1, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, -1, 1, -1, -1, -1, 0, -1, -1, 1, 0, 1, -1, 0, -1, -2, 0, 0, -2, -2, 0, -1, -1, 0, 0, -2, -1, 0, 1, 0, -1, 0, 0, -1, -1, -1, 0, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 2, 0, -2, 1, 0, 0, 0, -1, -1, 1, -2, 0, 0, -2, -1, 1, 0, 0, -1, 0, 0, -1, 1, 0, -2, 0, -1, 0, 0, -2, -2, 0, 0, -1, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 1, 1, -1, -1, 1, 1, -2, -1, 0, 1, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -2, 0, 0, -1, -1, 0, -1, 0, -1, 1, 1, 0, 1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -2, -2, 1, 1, -2, 0, 0, 0, 0, -1, 0, 1, -2, 0, -1, 1, 1, -2, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -2, -1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, -1, 0, 1, -2, 1, 0, -1, -1, 0, 0, -1, 1, -1, 0, 1, 0, 0, -1, 0, -1, 0, -2, -1, 0, 0, 0, 0, 1, 1, -1, 1, -1, -1, 1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, -2, 1, 0, 0, 0, 0, -2, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 1, 1, -1, 0, 0, 0, -2, 1, 0, 0, 1, 0, 0, -1, -1, -1, -1, 1, -2, 0, 0, 1, 0, -1, 1, -2, -1, 1, 1, 1, -1, -2, -1, -1, -1, -1, 1, 0, 1, -1, -2, -1, -1, 1, -1, 0, 1, -1, 0, 0, 1, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 1, -2, 0, 0, -1, -1, -1, 1, 1, -1, 0, -1, 0, -1, 0, 1, -1, 0, -1, 1, 1, -1, 0, 0, 0, -1, 0, -1, -2, -1, -1, 0, -1, 1, 0, 0, 0, -1, 0, 0, 1, 1, -2, 1, 0, 1, 0, -1, 0, 0, -2, 0, -1, 0, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, 1, -2, -1, -1, 0, 0, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, -1, -1, 1, 0, 1, 0, -2, 1, -1, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, -1, -2, 0, 0, 0, 1, -1, 0, 0, 0, -2, 1, 0, 0, 1, 1, -1, 0, -1, -1, 1, 0, 0, 1, 1, 0, -1, -1, -2, 0, 0, -1, 0, 0, 0, 0, -1, 1, -1, 0, -1, -1, 2, 0, -1, 0, 1, 0, 1, 0, -1, 0, 1, 0, 0, 1, -1, 1, 1, 1, 0, -1, 0, -1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, -1, 1, -1, 0, -1, 0, -2, 0, -1, 0, 1, -1, 0, -1, 0, 1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 1, -1, 0, -1, 1, 1, 0, 0, -1, 0, 0, -1, 0, 1, -2, 0, -2, 0, 1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -2, -1, 1, -1, -2, -1, -2, -1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 1, 0, -2, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, 1, 0, 0, 0, 1, -2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, -1, -1, 1, 1, -2, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 1, 0, 1, -2, 0, 1, 0, -2, -2, 1, -2, 0, 0, -1, -2, -1, 1, 0, 0, 1, 0, -1, 0, -1, 1, -1, 0, 1, -1, -2, 0, 1, 1, -1, -1, 1, -1, 0, 1, 1, 1, -1, -1, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -2, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, 0, -2, 0, -1, 0, -1, -2, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, -2, -1, 1, 1, -1, 1, -2, 1, 1, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 1, 0, -2, -1, 1, -1, 0, 1, 0, 0, 1, -1, 0, 1, 1, -1, 1, 0, -1, 0, -1, 1, -1, -1, 0, 1, -1, -1, 1, 1, -1, 1, -1, -1, 0, 0, -1, 1, 0, 1, -2, 0, -1, 0, 0, 1, 0, 1, 0, -1, 1, 1, -1, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, -1, 0, 1, 0, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, 1, 0, -1, 1, -2, -1, 1, -1, -1, 0, 0, 1, -1, -1, 1, 0, 1, -1, -1, 1, 0, -1, 0, 1, 1, 1, 0, 1, -1, 1, 0, 1, 1, -1, 1, 1, 1, -2, 0, -1, 0, 0, 0, 2, -1, -1, 0, -1, 1, -1, 0, -1, -1, 0, 1, 1, -2, 1, 0, 0, -1, 0, 1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, 1, -1, 0, 2, 0, 1, 1, -2, 0, 0, 0, 0, -2, 0, -1, -1, 0, 1, 1, 0, 0, 0, 1, 0, -1, -1, 0, 1, 1, 0, 0, -1, 0, -1, 1, -1, -2, 0, 0, -1, -1, 0, 1, 1, 1, 0, 1, 1, -1, -1, -1, -1, 0, 2, -2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -1, 1, 0, 0, -1, 0, 0, 0, -1, 1, 0, -1, 0, 2, 0, -1, 0, 0, 0, 1, -1, 1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, 1, 1, 0, -1, 0, 0, -2, 0, 0, -1, 1, 0, 1, 0, 0, 2, 0, 1, 2, -1, 0, 0, 0, 1, 0, 0, -1, 0, -1, -1, -1, 0, 2, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, -1, 1, -1, 1, 0, 0, -1, -2, 0, 0, 0, 1, -1, -1, 0, -2, -1, 1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, 0, 1, 2, 0, 0, -1, 0, 0, -1, -1, 0, -2, 0, -1, 0, 0, -2, 0, 0, 1, 0, 0, 0, 1, -1, 1, 1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 1, -2, 0, 1, -1, 0, 0, 0, 0, -1, 0, 1, 1, 2, 0, -2, -1, -1, 1, 0, 0, -1, 0, 0, 0, 2, 0, -1, -1, 1, 0, 0, -1, 1, 0, 0, -1, 0, 1, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 1, 1, -1, -1, 0, 0, -1, -1, 1, 0, -1, 1, 0, 0, 1, 0, 1, 0, 0, 1, -1, -2, -1, -1, 1, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 1, 0, -1, 0, 0, 0, 0, 1, -1, -2, 0, 1, -1, 1, 0, 0, -1, 0, 0, -2, -1, 1, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, -2, -1, -1, 0, -1, -1, -2, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 0, 1, 0, 1, -2, 0, 1, -1, 0, 0, 0, 0, 1, -1, 0, -1, 1, -1, 1, 1, -1, 0, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, -2, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, 1, -2, 1, 1, 1, 0, 2, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 1, 2, -1, -2, 0, -2, 0, -1, -1, 0, 0, 1, -1, -1, 1, 1, -1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, -1, 1, 0, 0, 1, 2, 1, 0, 1, -1, -1, 0, 0, -1, 1, 0, -1, 0, 0, 1, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 0, 1, 2, 1, 1, -1, -1, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, -1, 1, 0, 1, 1, 0, 0, 0, 0, -2, 0, 0, 0, -1, 1, 0, 0, 1, -1, -1, 2, 0, 0, 1, -1, 1, 1, 0, 1, 0, 0, 1, 1, 1, -1, -2, 0, 0, 0, 0, -1, 1, 1, -1, 1, 0, -1, 0, -2, 0, -2, 1, 0, -2, -1, 1, 0, 1, 0, -1, 0, -1, 1, 0, 1, -1, 0, -1, 2, -1, -1, 1, 2, 0, 0, 0, -1, 0, 0, -2, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 2, 1, 1, 0, 1, -1, 0, 1, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, -1, -1, -2, 1, 0, -1, -1, 0, 0, 0, 0, -1, -2, 1, 0, 0, -1, 1, -1, 1, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, -2, 0, 1, -1, -1, 0, -1, -2, 0, 1, -2, -1, 1, 1, 1, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, -2, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, -1, 0, 1, 0, -1, 1, 1, 0, -1, 0, -9, -8, -6, -5, -8, -7, -6, -3, 0, 1, -1, 1, -2, 0, -1, 0, -2, 0, 0, 0, 0, 2, 0, 0, 2, 0, -2, 0, 1, 2, -10, -7, -5, -3, -3, -4, -4, -1, 1, 2, 2, 1, 0, 0, 0, 0, 0, 1, 2, 5, 5, 3, 2, 2, 0, 0, 1, 0, 2, 2, -4, -3, -3, 0, -1, -3, -3, 0, 2, 1, -1, 0, 0, 0, 3, 1, 2, 1, 3, 3, 4, 6, 2, 1, 1, 2, -1, 1, 2, 5, -5, -3, -3, -1, 0, 0, 0, 0, -1, 1, 0, 2, 0, 0, 4, 2, 4, 3, 6, 6, 6, 7, 6, 3, 2, 0, 1, 4, 4, 2, -4, -5, -1, -1, 1, 0, 0, -1, 0, -2, 1, 0, 2, 1, 2, 0, 1, 5, 3, 4, 7, 5, 7, 3, 1, 2, 1, 0, 2, 4, -5, -2, 1, 0, 0, 2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 2, 5, 3, 6, 2, 2, 4, 3, 4, 0, 2, 2, 4, 4, -1, -1, 0, 2, 0, 3, 0, 4, 0, 3, 2, 1, 1, 0, 1, 0, 2, 1, 3, 1, 5, 3, 3, 3, 0, 1, 0, 2, 4, 3, 0, 0, 0, 4, 3, 1, 1, 1, 3, 1, 3, 3, 1, -1, 0, 0, -1, 0, 0, 2, 0, 5, 2, 2, 1, 1, -1, 1, 3, 3, -1, 0, 4, 3, 1, 1, 3, 3, 2, 4, 3, 0, -1, 0, -2, 1, 0, 0, 0, 2, 2, 4, 5, 0, 0, 0, 1, 3, 4, 5, -1, 2, 1, 1, 1, 0, 3, 0, 2, 3, 0, -1, 0, -3, -3, 0, 3, 0, 1, 2, 4, 4, 0, 3, 2, 0, 2, 4, 4, 7, -2, 2, 2, 0, 2, 2, 1, 1, 3, 4, 0, 2, -3, -3, -1, 0, -1, 1, 1, 1, 2, 3, 4, 2, 2, 3, 4, 4, 5, 6, -2, 0, 2, 0, 0, 0, 2, 0, 0, 0, 2, -2, -2, -2, -2, 0, -1, 0, 0, 0, 2, 0, 4, 1, 5, 6, 4, 3, 4, 7, -3, -1, 1, 1, -1, -2, 0, -1, 1, 1, 0, -2, -4, -1, -3, -3, 0, 0, -2, -2, -3, 0, 1, 0, 3, 5, 3, 5, 8, 4, -1, 0, 1, 0, 0, -3, -3, -1, 1, 0, -2, -2, -2, -4, -5, -2, -4, -4, -3, -8, -7, -4, -3, -1, 4, 2, 4, 3, 4, 7, -1, 0, 3, 2, 1, -1, -2, 0, -2, -2, -1, 0, -3, -4, -2, -4, -5, -3, -8, -8, -6, -8, -4, -1, 0, 0, 4, 3, 5, 6, 0, -1, 0, 2, -1, -2, 0, 0, 0, -1, -3, -3, -3, -4, -2, -4, -4, -6, -11, -11, -11, -7, -5, -2, -1, 0, 1, 3, 5, 5, 0, -1, 0, 1, 2, 1, -2, -1, 0, -2, -2, 0, -2, -1, -2, 0, -3, -5, -9, -10, -10, -6, -2, -3, -1, -1, 2, 2, 6, 2, -3, 0, 0, 3, 0, 2, 0, -1, -3, -1, -1, -4, 0, -2, -2, -2, -3, -4, -8, -7, -6, -3, 0, -2, 1, 0, 3, 3, 4, 5, -1, -1, 2, 0, 0, 0, -1, 0, -3, -1, -3, -3, -2, 0, -4, -4, -3, -1, -2, -5, -5, -3, 2, 2, 2, 1, 4, 5, 4, 4, -1, 0, 0, 2, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, -3, 0, 0, 0, 1, 3, 2, 5, 5, 4, 6, 0, 0, 0, 1, 0, 1, 3, 0, 0, -1, -1, 1, 0, 0, -1, 2, 1, 1, -1, -1, 0, -2, 0, 3, 3, 3, 2, 3, 7, 6, -1, 0, 4, 2, 3, 3, 0, 1, -2, -1, 2, 0, 1, 1, -1, 0, 3, 2, 0, 1, 0, 0, 4, 4, 3, 2, 3, 6, 6, 3, -4, 1, 3, 1, 2, 3, 0, 2, -1, 1, 0, 2, 3, 0, 1, 1, 3, 1, 0, -1, 0, -1, 3, 1, 3, 0, 3, 3, 2, 4, -1, 1, 3, 3, 2, 1, 2, 2, -1, 0, -2, 0, 0, 0, 0, 2, 4, 2, 3, 0, 2, 1, 3, 2, 2, 3, 2, 5, 3, 3, -2, 0, 1, 3, 4, 3, 2, 0, 0, 1, -3, 0, 0, 0, 2, 1, 1, 2, 4, 4, 0, 4, 5, 5, 4, 2, 1, 3, 2, 1, -2, -2, -1, 1, 3, 2, 2, 2, 1, -1, 0, -1, -1, 2, 0, 0, 1, 5, 5, 4, 6, 4, 5, 6, 4, 1, 4, 0, 0, 0, -6, -2, -1, 1, 1, 2, 2, 2, 0, 0, -1, -1, 0, 1, 0, 3, 3, 4, 5, 4, 5, 6, 6, 5, 3, 3, 3, 1, 1, 0, -7, -2, 1, 0, 1, -1, 0, 0, -1, 0, 1, -2, 1, 2, 0, 2, 3, 3, 5, 7, 6, 3, 4, 1, 0, 2, 3, 2, 2, -1, -5, -3, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 1, 2, 0, 1, 2, 5, 5, 6, 3, 2, 0, 1, -2, 1, 0, 0, 0, -1, -9, -7, -5, -1, -3, -4, -1, -3, 0, 2, 0, 2, 0, 2, 1, 0, 2, 1, 2, 0, 0, 0, -2, -4, -3, -3, -1, 0, 0, 0, -2, -3, 0, -1, -1, -1, 0, -2, -3, -1, -2, -1, -2, -3, 0, -2, 0, 0, -2, -1, -3, -2, 0, -1, 0, -1, 0, -3, -2, -1, -1, -1, -4, -1, -3, -1, 0, 0, 0, 0, -1, 0, -1, -2, 0, -1, -2, 1, -1, -1, 0, -1, 0, -1, -2, 0, 0, -2, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -2, -1, -1, 0, 0, -2, 0, 1, 0, 0, -1, 0, -2, -1, 0, 0, -3, 0, -1, -1, 0, 0, -2, -1, -1, 0, -3, -2, -2, 0, -1, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, -2, -1, -2, 0, 0, -3, -1, -3, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, -2, -1, -1, -1, 0, -2, 0, -2, -3, -4, -1, 0, 0, -3, 0, 0, 0, -1, -2, 0, -1, -2, 0, 0, -1, -2, -1, -2, 1, 2, -1, -1, -1, -3, 0, -1, -2, 0, -3, 0, -2, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, -3, 0, -3, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, -2, -1, 0, 0, -2, -2, -2, 0, 0, -2, 0, -1, 0, -3, 0, 1, -2, -2, -2, -1, 0, 0, -2, 0, 0, 0, 0, -2, 0, -2, 0, -1, -1, -2, 1, 0, 0, -2, 0, -2, -2, -1, 0, -1, 0, -2, -1, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, -2, 0, 0, -3, -1, 1, 0, -2, 0, -2, -2, -1, 0, 0, 0, 0, 2, 0, -2, 0, 0, 0, 0, -1, -2, 0, 0, -1, 0, -3, -2, -2, -2, -1, -1, 0, 0, -1, -2, -3, -2, -3, -2, 0, 0, 0, 0, -1, -1, -2, -1, 0, 0, 0, -2, 0, 0, 0, -2, -1, -1, 0, -1, 0, 0, 0, 0, 0, -3, -1, -1, 0, -2, 0, 0, -1, 0, 1, -1, -2, 1, -2, 0, -1, -2, 0, -1, 0, 0, 0, -2, -2, 0, -2, 0, -1, -3, -1, -1, 0, -2, -2, -3, -2, -1, -2, 1, 0, -1, 0, -1, -1, 0, -1, -1, 0, 0, 0, -3, -2, 0, 0, -3, 0, 0, -1, -2, -3, -3, -1, -4, -2, -3, 0, 0, 0, 0, -1, -1, -1, -1, -1, 0, 1, -2, 0, 0, 0, -1, -1, 0, -2, -2, -2, -3, -1, -4, -3, -2, -2, 0, -2, 0, 0, 0, -1, 0, -4, -2, 0, -1, 0, -3, -2, 0, 0, -3, -1, -1, -1, -1, -3, 0, -3, -2, -2, -2, -2, -4, -2, -4, -2, 0, 0, -1, -3, -3, -3, -3, -3, -1, 0, 0, 0, -2, -2, -3, -3, -2, -3, -3, -2, -2, -2, -2, -1, -1, -1, -1, -1, -2, -3, 0, -3, -3, 0, -1, -1, -1, -3, 1, 0, -2, -1, -1, -1, -3, -2, 0, 0, -1, -1, 0, -3, 0, -2, -2, -3, -2, -2, -1, -1, -3, -1, 0, -2, 0, 0, 0, -2, -2, 0, -1, -1, 0, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, -3, -1, -2, 0, 0, -2, 0, 0, -1, 0, -3, -3, -2, -2, -1, -2, 0, -2, 0, 0, -2, -2, -3, -1, -1, 0, 0, 0, -2, -1, -2, -1, -3, 0, -3, -1, -1, -3, -2, -2, -2, -3, 0, -2, 0, 2, 1, 1, -2, -1, 0, -1, -1, -1, 0, -1, -2, -2, -3, 0, -2, -2, -1, 0, 0, -2, -2, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, -3, -2, -2, 0, -4, -2, 0, -1, 0, 1, -1, -1, 0, -3, 0, -2, -2, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -3, -3, -3, 0, 0, 0, -2, -1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 0, 0, 0, 1, 0, -2, 0, 0, -2, -3, 0, 0, 0, -1, -1, -2, -1, -1, -1, -1, -1, 1, -1, -1, 0, -1, -1, -2, 0, -1, -2, -2, 0, -1, 0, 0, 1, 0, 0, -3, 0, -2, -1, 0, 0, -1, -2, -2, 0, 0, -1, -2, 0, -1, -1, 0, 0, 0, -1, -1, 0, -2, 1, 1, -1, 0, 0, -2, -2, 0, -2, -2, -3, -2, -2, 0, 0, 0, -1, 1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, -2, 1, -1, 0, -2, -1, -1, -2, -1, -2, -1, -2, -1, -2, 0, 0, -2, 0, -2, 0, 0, -2, 0, -2, 0, -1, 0, -2, 1, -2, -1, 0, -1, 0, -1, 0, -1, 0, -1, -2, -3, 0, -2, -1, -2, 0, -2, 0, 0, -1, 0, -2, 0, 0, 0, 1, 0, 2, 1, 1, 0, 1, 0, -1, -2, 0, -3, -1, -1, -5, -1, -3, -1, -2, -1, 0, -2, -3, 0, 0, 0, -2, 0, 0, -2, 0, 0, 1, 0, 0, 0, 0, -3, 0, -2, -1, 0, -1, -1, -3, -4, -3, 0, -1, -3, 0, -3, -3, -2, -1, 0, -2, 0, 1, 0, 1, 0, 0, 0, 1, -3, 0, -3, 0, -1, -3, -3, -2, -2, -13, -13, -9, -8, -8, -9, -8, -6, -5, -3, -1, -3, -2, -3, -6, -6, -5, -4, -4, -1, 0, 0, -2, -3, -6, -7, -5, -8, -6, -5, -12, -9, -5, -6, -5, -5, -6, -5, -4, 0, -1, -2, -4, -3, -3, -5, -2, -3, 0, 0, 1, 0, 1, -1, -3, -3, -7, -5, -3, 0, -10, -9, -4, -5, -5, -3, -2, -3, -6, -3, -4, -2, -2, -2, -2, -3, -2, 0, 1, 2, 3, 3, 2, 0, -3, -4, -4, -4, -3, 1, -9, -6, -3, -4, -3, -2, -4, -3, -2, -5, -5, -3, -4, -2, -3, -1, 0, 0, 3, 1, 3, 0, 0, 2, -1, -2, -4, -1, -3, -3, -10, -8, -5, -4, 0, -3, -2, 0, -1, -4, -4, -3, -5, -5, -3, -4, 0, -1, 0, 4, 2, 1, 0, -1, -2, -2, -7, -4, -4, -2, -8, -4, -5, -3, 0, -2, 0, -1, 0, -3, -2, -2, -4, -3, -2, -3, -5, -4, -3, 0, 0, 0, 0, 0, -5, -4, -3, -2, -3, 0, -8, -4, -1, 0, -1, -1, -1, 1, 0, 0, -1, 0, -4, -5, -3, -6, -4, -1, -1, -1, -2, -1, -1, 0, -5, -7, -7, -5, -1, -2, -4, -1, 0, 1, 0, -3, 0, -3, -1, 1, 1, 0, -4, -6, -5, -3, -2, -3, -2, -1, 2, 0, -1, 0, -3, -6, -3, -5, -3, 0, -4, -3, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -2, -2, -5, -4, 0, 1, 3, 0, 1, 4, 0, 0, -1, -3, -3, -1, 0, 0, -4, -2, 0, 1, 0, -3, -1, 0, 0, -1, -1, 0, -3, -4, -4, 0, 1, 3, 3, 3, 2, 3, 2, 2, -3, -3, -1, -3, -1, -1, -7, -4, 0, 0, -4, -5, -4, -1, -1, 0, -3, -6, -3, -6, -3, -1, -1, 2, 2, 0, 3, 3, 1, 1, 0, 0, -1, 0, -3, 0, -6, -3, -1, 0, -2, -6, -9, -4, -4, -1, -3, -6, -7, -6, -6, -4, -2, 0, 1, 0, 0, -1, 0, -1, 2, 0, 0, 2, -1, 0, -7, -5, -3, -3, -3, -7, -8, -7, -6, -6, -2, -5, -3, -6, -4, -4, -3, -3, -3, -1, -2, -2, -2, -2, 2, -1, 1, -2, -1, -2, -4, -5, -2, -1, -4, -7, -5, -4, -4, -8, -4, -3, -4, -3, -2, -1, -1, -4, -6, -8, -7, -8, -6, -1, 0, 0, -2, 0, 0, -1, -4, -3, -4, -4, -5, -5, -9, -8, -7, -5, -4, -5, -3, -2, -1, -1, -1, -3, -7, -10, -14, -10, -7, -3, -4, -1, -3, 0, 0, -3, -7, -6, -4, -1, -3, -3, -7, -6, -8, -7, -7, -5, -4, -2, 0, 0, -2, -1, -9, -13, -15, -9, -5, -5, -3, -4, -1, -1, 0, 0, -7, -3, -2, -4, -3, -5, -6, -8, -9, -7, -7, -5, -5, -3, 0, 0, -2, -3, -7, -8, -10, -7, -4, -1, -1, -3, -1, -2, 0, -2, -6, -4, -5, -4, -2, -4, -3, -6, -9, -9, -6, -5, -6, -3, -3, -1, -4, -1, -2, -4, -4, -3, 1, 1, -1, 0, -2, 0, 0, -1, -5, -7, -4, -2, -2, -5, -5, -6, -8, -7, -4, -4, -5, -2, -4, 0, 0, 1, 1, -3, -1, -1, 0, 0, 0, -2, 0, 0, -3, -3, -8, -3, -1, 0, -2, -1, -5, -6, -8, -8, -4, -1, 0, -2, -1, 1, 2, 4, 2, -1, -3, -2, 1, 1, 2, 0, -3, 0, 0, 0, -8, -5, 0, 1, 0, -3, -1, -3, -7, -4, -4, -2, 1, 0, 0, -1, 2, 3, 1, 0, 0, -3, 2, 3, 0, -1, -4, -3, -1, -1, -8, -6, -2, 1, 0, 0, -2, -4, -3, -4, -6, 0, -2, 1, 0, -1, 0, 2, 0, -1, -4, -4, 0, 2, 0, -1, -4, -4, -3, -5, -6, -6, -2, 1, 0, 1, 0, -1, -3, -2, -6, -2, 0, -2, -1, 1, 2, 0, 0, 1, -2, 0, -1, 0, 0, 0, -4, -2, -2, -2, -9, -4, -3, 1, -1, -1, -2, -3, -6, -4, -7, -4, -5, -1, 0, -2, 0, 1, 1, 1, 0, 0, 2, 1, 2, -1, -2, -1, -5, -5, -11, -6, -5, -1, -2, 0, 0, -2, -3, -6, -6, -4, -7, -4, -3, 0, 1, 1, 3, 0, 1, 4, 3, 4, 2, 0, -3, -1, -5, -4, -10, -5, -3, -1, 0, 0, -1, 0, -2, -6, -4, -6, -7, -2, -1, 0, 0, 1, 4, 4, 1, 5, 1, 2, 2, 0, -1, -5, -6, -4, -11, -9, -2, -3, -4, -3, -2, -3, -1, -5, -4, -5, -3, -6, -4, -1, -1, 0, 3, 3, 2, 2, 0, 0, -1, -4, -4, -5, -5, -5, -11, -8, -3, -4, -3, -5, -5, -2, -2, -5, -3, -6, -6, -5, -4, 0, -3, -2, 0, 2, 2, 2, 0, -4, -5, -4, -3, -2, -7, -8, -15, -10, -7, -4, -4, -7, -5, -8, -4, -4, -2, -1, -3, -3, -5, -2, -2, -4, 0, 0, 0, -1, -2, -7, -7, -6, -4, -3, -5, -4, -18, -12, -8, -5, -7, -9, -7, -7, -9, -4, -5, -2, -2, -3, -7, -4, -6, -6, -5, -4, -4, -7, -9, -11, -8, -10, -8, -4, -4, -7, -3, -3, -2, -3, -3, -2, -1, 0, 0, -1, 0, 0, -2, -4, -4, -1, -2, 0, -3, -1, -4, -2, -2, -4, -3, -1, -4, 0, -1, 0, -2, -2, -2, -3, -3, -2, 0, -1, 0, -1, -2, -1, -2, -2, -4, -2, 0, 0, 0, -1, -3, -3, -1, 0, -5, -3, -2, 0, 0, 0, -2, -2, -2, -2, -4, -1, -1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, -1, -2, 0, 0, 0, -2, -1, -1, -2, -2, -2, -1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, -2, -2, -3, 0, 0, -2, -2, 0, -1, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, -3, -4, -2, -2, -2, -1, 0, -1, 0, 0, -1, -1, 0, -1, 0, 0, -4, -3, -3, -2, 0, 0, -3, 1, -1, 0, 1, 0, 0, -2, -1, -2, -3, -1, -2, -3, -2, 1, 0, -1, -1, 0, 0, 0, 0, 0, -4, -1, -4, -3, -3, -1, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, -1, 0, -1, 1, 0, 1, -1, 0, -1, -4, -4, -4, -1, 0, 0, -1, -2, 1, -2, -1, -1, 0, -1, 0, -2, -1, -1, -1, -3, -1, -3, -3, -3, -2, 0, 0, -2, -2, 0, -3, -4, -3, -2, 0, -3, 0, 0, 1, -1, 0, -1, -3, 0, 0, -1, 0, 0, -2, 0, 0, -2, 0, -1, -3, -2, 1, -2, -3, -1, -3, -5, -4, 0, -1, -1, -2, -2, 0, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, 0, -3, 0, -1, -1, 0, 0, 0, 1, 0, -3, -4, -1, -1, -4, -1, -2, 0, 0, -1, -2, -2, -2, -1, 0, 0, 0, -2, -1, -2, 0, -2, 0, 1, 1, 0, -1, -1, 0, 1, 0, 0, -1, -2, -2, -4, -4, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, -2, -1, 0, -1, 1, 1, 2, 0, 2, 2, 2, 0, 0, -2, -3, -1, -1, -2, -2, -3, 1, -1, -1, -3, -1, -1, -1, -2, 0, -1, -1, -5, -3, -1, -3, 0, -1, -1, 0, 1, 2, 0, -1, -2, 0, -1, -2, -1, -4, -1, -1, -2, 0, -3, -4, -4, -2, -1, -3, 0, 0, -1, -3, -3, -2, -2, 0, -2, 0, 1, 2, 0, -1, 0, -1, -2, -2, -1, -3, -3, 0, -1, -2, -2, -3, -4, 0, 0, -3, -2, -2, -1, 0, -1, 0, -2, 0, -3, -1, -1, 1, 1, 2, 2, -1, -1, -1, 0, -3, -2, -1, 0, 0, 0, -4, -1, -1, -2, -1, 0, -2, -1, -3, -2, -3, -3, -1, -5, -4, -1, -1, 0, -1, 1, 0, -3, -2, -2, -3, -2, -1, 0, -2, 0, -1, -5, -2, -3, -1, -1, 0, 0, 0, 1, 0, -1, 0, -2, -3, -3, -1, 0, -3, -2, -2, -3, -2, 0, -3, -4, -1, 0, 1, 1, -2, -1, -4, -3, -1, -3, -3, 0, 1, 1, 0, 0, -1, -2, -5, -2, -3, -1, 0, -3, -3, -3, -3, 0, -1, -1, -1, -1, -2, 0, -2, -1, -1, -2, 0, -2, -1, -2, -2, 0, -2, 0, -2, -4, -3, -2, -3, 0, -1, -2, -2, -2, -1, 0, -4, -5, 0, 1, -3, -1, -3, -1, -4, -2, -2, -2, -2, -2, -2, 0, -3, 0, -2, -3, -3, -4, -1, 0, 0, -2, 0, -2, 0, -4, 0, -4, 0, 0, -2, -1, 0, 0, -4, -4, -1, -1, 0, -2, -2, -3, -3, -1, -1, 0, -2, -1, 0, -1, 2, -2, -4, -1, 0, 0, -2, -1, 0, 1, -1, -3, 0, -3, -3, -2, -3, -3, 0, 0, 0, 0, -1, 1, 1, 1, 0, -2, -3, 0, 1, 2, 0, -1, -3, -2, -2, -2, 0, 1, 1, -2, -1, -2, -1, -1, -3, -1, 0, -1, 0, -2, -3, 0, 0, -2, -1, -2, 0, 0, 0, 1, -3, -1, -2, 0, -3, -5, 1, -1, 0, 0, -2, -3, 0, -1, -1, -3, -1, -1, 1, 0, -1, 0, -1, -1, -3, -5, -3, 0, 0, 0, -2, -3, -3, -1, -4, -2, 0, 0, 0, 0, 0, -2, -2, -3, -5, -3, -4, -2, 0, -1, 0, 0, 0, -2, 0, -1, 0, 0, -2, 0, -3, -4, -2, -4, -2, -3, -1, 2, -1, 0, 1, 0, -3, -4, -1, -4, -1, -3, -3, 0, -3, -2, -2, -2, 0, -2, -3, 0, 0, -1, -3, -4, -4, -1, -4, -3, 1, 0, 0, 1, -1, 0, -1, -3, -3, -4, -2, -1, -1, -3, -2, -1, 0, 0, -2, -2, -3, 1, -2, 0, 0, -3, -3, -2, -4, -1, 1, 2, 0, 0, -2, 0, 0, 0, -3, -3, -2, -4, -1, -1, -3, 0, 0, -1, -1, -1, 1, 0, -2, -3, 0, -3, -4, -2, -2, -1, 0, 1, 2, 0, 0, 1, 0, 0, 1, -3, -3, -3, -3, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, -2, -1, -2, -1, 0, 0, -1, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, -3, -1, 0, 1, 1, 0, 0, 1, -2, 0, -3, 0, -1, -4, -4, -3, 0, 1, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, -1, -1, -1, 0, 0, 0, 1, 1, -2, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 1, -1, -2, 0, -1, -1, -1, -1, -1, -1, 0, 1, 0, 0, 0, -1, 0, 1, -1, 1, 1, -1, -1, 0, -1, 1, -1, -1, 0, 1, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 1, 1, 1, 0, -1, -1, -1, 0, 0, 1, -2, -1, -2, -1, 0, 0, 0, 0, 1, 1, 1, -1, -2, -1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, -1, 1, 0, -1, 0, 0, -1, 1, 0, -1, 0, 1, 0, 1, 2, 1, -1, 0, 1, 0, 1, -1, 1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -2, 1, 0, 0, -1, 1, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, -1, 1, 1, 0, 2, 0, 0, -1, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, 1, -1, -1, 0, 1, 1, 1, -1, 2, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, 2, 0, -1, 1, 1, 0, -1, 0, 1, 0, 0, -1, 0, -1, -1, 0, 1, -1, 1, -1, 0, -1, 0, 0, -1, 1, -1, 2, 0, 0, 0, 0, -1, -1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, -2, 0, 0, -1, 1, 0, 1, 0, 0, 0, -1, 1, -1, -1, 0, 1, -1, 0, 1, 1, 0, 1, 1, 1, 0, -2, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 1, 1, -1, 1, -1, 0, -1, 0, 1, 2, 0, 0, 0, 0, 1, 1, -1, 1, 1, 0, 2, 0, 1, 0, 0, 1, -1, 0, 0, 0, -1, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -1, 1, 1, 1, 0, -1, 0, 0, 0, -1, 1, 1, 1, -1, 0, -1, 1, -1, 1, 1, -1, -1, 1, -1, 0, 0, -2, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, -1, -2, 0, 1, 1, 0, -1, 0, -1, 0, 0, -1, -2, -1, 0, -1, -1, 2, 0, -1, 0, -1, -1, 0, 1, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 2, -1, -1, 0, 0, 0, 1, 0, -1, -2, 1, 1, -1, 1, 0, 0, 0, 1, -1, 0, -1, 0, 0, 1, -1, 0, 0, -1, 0, 0, 1, 1, -1, 0, 1, 1, -1, 0, 0, 2, 1, -1, 1, -1, 1, 1, 0, -1, -1, 0, -1, 1, 0, 1, 2, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 1, 2, 0, 0, 0, -1, -1, 1, -2, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 2, 1, 0, 0, 1, -2, 0, 0, 2, -1, 0, 0, 1, 1, 0, -1, -1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, -2, 0, 0, 1, 0, 1, -2, 1, 2, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, -1, 1, -1, 0, -1, 1, 1, -1, 1, 1, 0, 0, 1, 1, 0, 1, 0, -1, -1, 0, 0, 0, 2, 1, 0, -1, 1, 1, 0, -1, 1, -1, 0, -1, 0, 0, 1, 0, -1, 0, 1, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, -1, -1, -2, 0, 0, 0, 1, 0, 1, 0, -1, 1, -1, 1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 1, 1, 1, 0, 1, -1, -1, 0, -1, -1, 0, 1, 1, 0, 0, 0, 0, -1, 1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 1, -1, -1, 0, 1, 0, 0, 1, -1, 1, 1, 0, 0, -1, 0, -1, 1, 0, -1, -1, 0, 1, 1, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, 2, -1, 0, 1, 1, 0, 0, 1, 1, -1, -1, -1, -1, 0, -1, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 0, 1, 1, -1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, -1, 1, 0, 0, 0, 1, 0, 1, 0, -1, -1, 0, 0, -1, 0, 2, 0, -1, 1, -1, 0, -1, -1, 0, 1, -1, 0, -1, -1, 1, -1, 1, 0, 1, -2, -1, -1, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 2, -1, -1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, -1, 1, -1, 0, 0, 0, 2, 1, 1, -1, 0, -1, 0, 0, 1, 1, 0, 0,
    -- filter=0 channel=5
    0, 0, 0, 1, -1, 0, 0, 1, -2, 0, -2, 0, 0, -1, 0, -1, -2, -2, 1, 0, 0, 2, 0, -2, -1, -1, 1, -1, 1, 0, 0, 1, -1, 0, 0, -1, -1, 0, 1, 0, -2, 0, -1, 1, -2, 0, 0, -1, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, -1, 0, 1, -1, -1, 1, 0, 0, -2, -2, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, 0, -2, 0, -2, 0, -2, 1, 0, -1, -2, 0, 0, 0, -2, -2, 1, 0, -2, -2, -1, 0, 0, -2, -1, -2, -1, -2, -1, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, 1, 0, 0, 0, 0, -2, -2, 0, -1, 0, -2, 0, 0, -2, -3, -2, -1, 1, 0, -1, -1, -2, 1, 0, 0, 0, -2, 1, -2, 1, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, 0, -1, 0, 0, 0, 0, 0, 0, -2, -2, -2, 1, 0, 0, -1, -1, 0, 1, -1, 2, 1, 2, 0, 1, -2, -1, 0, -2, -2, 0, 0, -2, -3, -3, -3, -1, 0, 0, -2, 0, -1, -2, 0, 0, 0, 0, 2, 2, 0, 0, 2, 2, 0, 0, -1, -2, 0, -2, 0, 0, 1, 0, -1, -2, -3, -1, 0, -1, -3, 0, -2, 0, -2, 0, 2, 2, 0, 2, 2, 1, 2, 1, 0, 1, -1, -3, -3, 0, -2, 0, 0, 0, -1, 0, -2, -2, 0, -1, -1, -3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, -2, -3, -1, -3, 0, -2, -2, -2, 0, -2, -2, -3, -1, -1, 0, 0, 1, 1, -1, 1, 0, 1, 1, 2, 0, 0, -1, 1, 0, 0, 0, 0, -3, 0, -2, -3, -3, -3, 0, 0, -3, -3, -1, 0, 1, 1, -2, 1, 0, 0, 1, 2, 0, 0, 0, 0, 2, -2, -2, -2, -1, -2, -1, 0, -2, -1, 0, 0, -1, -1, 0, -1, -2, -1, 1, 0, 1, 1, -1, -1, 0, 0, 0, 0, 2, 0, 0, 1, -2, -2, 0, -1, -2, 0, -2, -1, 0, -1, 0, -2, -2, -1, 1, 0, -2, 0, 1, -1, -1, 1, 2, 0, 0, 2, 2, 1, 0, -1, 1, 1, -1, -1, -1, 0, -1, 0, -2, 0, -2, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, 2, 2, 0, -1, 0, 0, 1, -1, 0, 2, -1, 0, -2, -2, 0, -2, 0, -2, 0, 0, -1, 0, -1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 1, 1, 1, 0, -1, 1, -1, -1, -2, 0, 0, 0, -3, 0, 0, 0, -2, 0, -3, -2, 1, -1, 0, 0, 0, 1, 0, 0, 1, 2, 2, 0, 0, -2, 0, -2, 1, -2, 0, -1, -2, -3, -2, 0, -2, -2, -2, -2, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 1, 2, 2, 2, -1, 0, 1, 0, -2, -1, 1, 0, 0, 0, -2, -3, 0, 0, -2, -1, -1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, -1, -1, 0, -2, -2, -1, -3, -2, -1, -2, 0, -1, 0, -1, -1, 1, -1, 0, -1, -1, 1, 1, 1, 0, 0, -1, 2, 1, 1, 1, -2, 0, -1, -2, 0, 0, 0, 1, -1, -3, 0, -1, -1, -1, 0, 0, 2, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -2, -1, -1, -1, -2, -1, 0, -1, -1, 0, -1, -1, -1, -1, 1, 1, -1, 1, 2, 1, -1, 0, 1, 1, -1, -1, 0, 0, 0, -3, -1, 0, -3, -2, 0, -3, -1, -3, -1, 0, -2, -1, -2, -1, 1, 0, 1, -1, 0, -1, 0, 0, 1, 0, -2, -1, 0, -1, -2, -3, -2, -2, 0, 0, -1, -1, -3, 0, 0, 1, -2, -2, -2, -2, -1, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -2, -3, 0, -2, -2, -1, -1, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, 2, 0, -1, 0, 0, 0, 0, 0, -2, -1, -1, -2, -2, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, -1, 0, 0, 1, -1, -1, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 1, -2, -1, -3, 0, 0, 0, 1, 0, 1, 0, 0, -1, -1, -1, 1, 0, 0, 1, -1, -1, 0, 1, -1, 0, -2, 0, 0, -1, 0, 0, -1, -2, -3, -1, 0, 1, 2, -1, -1, 2, 0, -1, 0, 0, -2, -2, 1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, 0, 2, 0, 1, 0, 1, 0, -1, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, -9, -5, -6, -5, -3, -6, -5, -6, -3, -4, -6, -6, -3, -4, -5, -2, -5, -2, -6, -5, -3, -7, -6, -6, -5, -4, -4, -7, -4, -5, -9, -8, -7, -6, -5, -4, -6, -5, -7, -6, -3, -2, -4, -3, -2, -2, -4, -3, -4, -6, -5, -6, -5, -7, -5, -4, -5, -4, -4, -5, -7, -8, -4, -5, -7, -7, -5, -3, -4, -4, -3, -3, -4, -4, -5, -4, -5, -4, -3, -5, -4, -3, -4, -2, -2, -1, -3, -1, -2, -4, -7, -5, -5, -4, -6, -6, -7, -5, -2, -5, -4, -2, -2, -5, -4, -4, -4, -3, -4, -2, -3, -2, -2, -4, -2, -3, -1, 0, 0, -4, -9, -7, -6, -5, -7, -5, -4, -4, -4, -4, -5, -3, -2, -3, -6, -4, -4, -3, -3, -1, -2, -4, -2, 0, 0, -2, -1, 0, -3, -2, -8, -7, -6, -5, -4, -6, -5, -5, -3, -5, -3, -3, -5, -4, -2, -3, -5, -4, -1, 0, -1, -1, -1, 0, -3, 0, 0, 0, -1, 0, -9, -9, -5, -6, -3, -3, -4, -6, -5, -3, -4, -2, -4, -2, -1, -3, -1, -1, 0, -1, 0, -3, -2, 0, 0, 0, -1, -3, 0, 1, -8, -8, -7, -3, -2, -3, -6, -6, -5, -5, -4, -2, -2, -5, -3, -2, 0, -1, 0, 0, 0, 0, -3, -2, -2, -1, -1, 0, -2, -2, -7, -6, -4, -5, -4, -6, -4, -2, -6, -2, -2, -5, -5, -2, -3, -2, -1, -2, 0, 0, 0, -1, 0, -3, -1, -2, 0, 0, 0, 0, -10, -7, -3, -3, -1, -1, -1, -6, -3, -5, -2, -5, -5, -3, -2, -3, -2, 1, 1, 0, -1, 1, -2, -2, -3, 0, 1, 0, 2, 1, -8, -4, -5, -3, -1, -3, -4, -3, -3, -5, -2, -3, -6, -5, -3, 0, 0, 0, 1, 2, 0, 0, -1, 1, -1, 0, 0, 1, 1, -1, -7, -7, -4, -2, 0, 0, 0, -3, -1, -2, -4, -3, -2, -3, -1, 0, 1, 0, 1, 3, 1, 0, 1, 0, 0, -2, 1, -1, 0, 0, -7, -3, -3, -2, 0, 1, -1, -1, -2, -4, -4, -1, 0, -4, -2, -1, 0, 2, 2, 2, 2, 3, 0, 0, -1, 0, 0, 0, 2, 2, -5, -3, -3, -2, 0, 0, 0, -1, 0, -1, -1, -2, -3, -2, -2, 0, 2, 0, 1, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, -7, -3, 0, 0, 0, 1, 1, 1, 0, -1, 0, 0, -3, -1, 0, 1, 2, 3, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -5, -2, -3, 0, 2, 2, -1, 0, 0, 0, -1, -1, 0, -2, -1, 2, 2, 0, 0, 0, 2, 0, -1, 0, -2, -2, 0, 0, 0, 0, -7, -3, 0, 0, 2, 0, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 1, 0, -2, -2, 0, -3, -4, -3, -1, -1, 0, 0, 0, 1, -1, 0, -3, -4, -1, -3, 0, 0, -1, -1, 1, 0, 0, -1, 0, 1, 1, 0, 1, 0, -2, 0, -5, -2, 0, 0, 0, 2, 1, 1, 0, 1, -1, -2, -1, -5, -3, -2, -1, 1, -1, -1, 0, -1, 1, 0, 1, 1, 0, 0, 0, -1, -6, -3, 0, 1, 1, 0, 1, -1, -2, 0, 0, -3, -4, -2, -5, -1, -2, 0, 0, 0, 0, -2, 2, 1, 1, -1, 0, -1, 0, 0, -7, -5, -3, 0, -2, 1, -1, -1, -2, -1, -1, 0, -1, -3, -6, -6, -4, 0, -2, -1, -2, 0, -1, 1, 1, -1, 0, -1, 1, -1, -8, -3, -2, -3, -2, -2, -1, 1, 0, -2, -2, -2, -4, -2, -5, -2, -3, -2, 1, 0, 0, -1, -2, 1, 0, 0, 1, 0, 1, 0, -7, -7, -4, -4, -1, -1, -1, -1, -1, -1, -2, -1, -3, -1, -1, -4, -1, -2, 0, 0, 0, -2, -1, -2, -2, 0, 1, 0, 1, 0, -8, -5, -3, -5, -1, -4, -1, -2, -4, -3, -5, -4, -1, -3, -2, -2, 0, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 1, 1, -6, -6, -6, -5, -5, -2, -5, -2, -1, -3, -3, -5, -3, -2, -1, 0, 0, -2, 0, -2, -1, -1, 1, 2, 2, 2, 0, 1, 1, 0, -10, -7, -8, -6, -5, -4, -4, -4, -2, -5, -5, -4, -4, -2, -3, 0, -2, 0, 0, 0, 0, -2, -1, 1, 2, 0, -1, -2, 0, 0, -8, -10, -6, -6, -6, -4, -3, -2, -1, -3, -2, -4, -4, -3, -1, -3, 0, -1, 0, -2, -1, -2, -2, 0, -1, 0, 0, 0, 0, -2, -10, -8, -6, -8, -5, -4, -1, -3, -3, -3, -3, -4, -3, -3, -2, -3, -2, -3, -2, -1, 0, -3, -1, 0, -2, 0, 0, -1, 0, -2, -8, -8, -8, -7, -3, -2, -4, -4, -6, -2, -4, -5, -2, -5, -1, -4, -2, -4, -1, -3, -3, -5, -2, -2, -1, -3, -1, -2, -3, -3, -7, -5, -7, -5, -6, -3, -4, -4, -1, -3, -5, -2, -4, -4, -2, -2, -4, -3, -3, -4, -2, -4, -5, -3, -4, -4, -2, -2, -4, -3, -1, -1, -1, -2, -1, -3, -1, 0, -1, -2, -3, -1, 0, 0, 0, 1, -1, 0, 0, -2, 0, -2, -1, -2, -1, -2, 0, 0, 0, 0, -1, -3, -2, -1, -1, -2, 0, -3, 0, -3, -1, -1, -2, 0, -2, 0, 0, -1, -1, 0, -1, -2, 0, 0, -2, -2, -2, -2, 0, 1, -5, -1, -1, -1, 0, -2, -3, -3, 0, 0, -2, 0, 0, 0, -3, -2, 0, 0, -1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 2, 1, -5, -3, -3, 0, 0, 0, 0, -3, -1, -3, 0, -1, 0, 0, -3, 0, -1, 0, 0, -1, -1, 0, -1, -1, 1, -1, 1, -1, 0, 0, -1, -2, -3, -1, 0, -3, -3, -2, -1, 0, 0, -2, 0, 0, 0, 0, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -4, -1, -3, -3, -3, -2, -3, 0, -1, -2, 0, 0, -2, 0, -2, -1, -2, -2, 0, -2, 0, 1, -2, -1, 1, 0, 0, 1, 1, 2, -4, -2, -2, -1, -1, 0, 0, -2, -1, -2, -2, -3, -3, 0, -2, 0, 1, -1, -1, 0, 0, 0, 1, 0, -2, 0, 0, -1, 1, -1, -3, -3, -1, -2, 0, 0, -2, 0, -2, 0, -1, 0, -2, 0, -2, -1, 0, 1, 0, 0, -2, -1, 0, -2, 0, -2, 0, 0, 1, -1, -4, -4, 0, -3, -2, 0, 0, -3, -1, 0, 0, 0, 0, -2, -1, 0, -1, -2, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -2, -3, -4, -3, -3, -1, 0, 0, -2, -1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, -2, 0, 1, 1, 0, 0, -1, 2, -1, -3, -3, -1, -1, -1, -3, 0, -2, 0, -2, 0, -2, -2, -2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, -3, -1, -4, -1, -3, -2, -2, 0, -3, -1, -1, -2, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -1, -3, -2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 2, -1, -1, 0, 1, 1, 0, 0, -1, 1, 0, -2, 0, -1, 0, -1, 0, -2, -1, -1, 0, -3, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, -4, -3, -2, 0, 0, 0, -1, 0, 0, -2, -1, 0, -1, 0, 0, 2, -1, -1, 2, 2, 0, 0, 0, 1, 0, 1, -2, 0, 0, 0, -3, 0, -1, 0, 0, 1, -1, -2, 0, 0, -2, 0, -1, -1, 2, 0, 2, 1, 0, 2, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, -2, 0, 0, -2, 0, -2, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -2, 0, -1, 0, 1, 0, 0, 0, 0, 1, -2, -1, 0, -2, 0, 2, 1, -1, -1, 0, -1, 0, -2, 0, 0, -2, -2, 0, 1, -1, -2, -1, -1, -1, 1, 0, 0, 1, 1, -1, -2, -1, -1, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, -1, -2, -1, 1, 1, 1, 0, -1, 0, 0, 1, 0, -1, -1, -1, 1, 0, 0, 1, 1, -2, 0, 0, 0, -2, -1, 1, 0, -1, -1, -1, 0, 1, 0, -1, 0, 1, 0, -3, -2, 0, 0, -1, 0, 1, 1, -1, 0, -2, -1, -2, -1, 0, 0, 0, 0, -2, -2, -1, -1, -2, 1, 1, -1, -1, -1, 0, 0, -3, -2, -2, 0, 1, 2, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, -1, -2, 0, -2, 0, 0, 0, 1, -1, 2, -1, 0, 0, -1, -3, -1, -1, -1, -2, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, -1, 1, -2, 0, -1, -2, 1, 0, -1, 1, -1, -3, 0, 0, -2, 0, -2, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, -3, -1, 0, 0, 0, -2, 0, -2, -1, -2, -1, 0, -2, -2, 0, -1, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4, -3, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -2, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 1, 1, -5, 0, -4, 0, 0, 1, 1, 0, -2, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 1, 1, 1, 0, 2, 0, 0, -2, 0, -1, -2, 0, 0, 1, 0, 1, -2, -2, 1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 1, -1, -1, 0, 0, -1, 0, 1, 0, 0, -3, -1, 0, -2, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, -2, -1, 0, 1, 1, 0, 0, -2, 0, -1, -1, 0, 1, 1, 0, 0, -3, -1, 0, 0, 1, -2, 0, 1, -1, 0, 0, -2, -2, 0, -1, 0, 0, -2, -2, -1, 0, -1, 1, 0, -1, 0, 1, -1, 0, 0, 0, 0, -2, 1, 1, 1, -1, 1, 0, 1, 0, -1, -2, 0, 0, 1, -1, -2, 1, 0, 1, 0, -2, -1, -2, 1, 0, 0, 0, 1, -1, 1, -1, 0, 0, 0, -1, -1, 1, -1, 0, -1, -1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, 0, 0, 1, 1, 0, 1, -1, 1, -1, 0, 0, 1, -1, 1, 1, -1, -1, 0, -1, -1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, -1, 1, -1, 0, 1, -1, 0, -1, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 0, -2, -2, -2, -1, -1, 1, 0, 0, 1, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, -1, -1, 0, 0, 0, 1, -1, 0, 1, 0, -1, 0, 0, 1, -1, 0, 1, 0, 1, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, -1, -2, 0, 0, -1, 0, -2, -1, 0, 0, 0, 1, -1, -1, 0, -1, 1, 0, 0, 0, 1, -1, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 1, -1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 2, 1, -1, -1, -1, 1, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, -1, -1, -2, 1, 1, -1, -2, -1, -1, 0, -1, -1, -1, -1, -1, 0, -1, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 0, 2, 1, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, -1, 1, 1, 0, 0, 1, 0, -1, 1, -1, 0, 0, -1, 0, -1, 1, 1, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, 2, -1, 1, -1, 0, -1, 1, 0, -1, -2, 0, 1, 0, 0, -1, -2, -1, -1, 1, 0, 1, -2, -1, 1, 0, 1, 1, -1, 0, 0, 0, 1, 2, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, 0, -2, 1, 0, 1, 1, 1, 1, -1, -2, -1, 0, 1, -1, -1, 0, -1, 0, 1, 0, 2, -1, -1, 0, -1, 0, 1, 1, -1, 0, -1, 0, -1, -1, 0, -1, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, 0, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -2, 1, -1, 1, 0, 1, -1, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 2, 0, 1, 0, 0, -1, 1, -1, -1, -1, 0, 1, 1, -1, 1, -1, 1, -1, 0, 1, -1, 1, 0, 0, 0, -1, 1, -1, 1, 0, -1, 0, 2, 0, -1, -1, 0, 1, 1, 0, 0, 1, 0, -1, 0, -1, 0, 1, 1, 1, 1, -1, 1, -2, 0, 1, 0, 1, -1, 0, 0, 0, -1, 0, 1, 1, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, -1, 2, 1, 1, -1, 1, 0, -1, -1, 1, -2, -1, 0, -1, 0, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, -2, -1, 0, 0, -1, 1, -1, -1, -1, -1, 0, -1, 0, 0, 1, -1, -1, 1, 0, -1, 0, -1, 0, -1, 1, -1, 0, 1, 0, -1, 0, 0, 0, -1, -2, -1, -2, 2, 0, 0, -1, -2, 0, 0, -1, 0, -2, 1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, 0, 1, 0, 0, -1, 1, 1, 1, -2, 0, -2, 0, 1, 0, 1, 0, -1, 0, 2, 0, 0, 0, 2, 0, -1, 1, 0, 1, 1, -1, -1, 0, 1, 1, 0, 2, 0, 0, 1, -1, 1, -1, -2, 1, 0, 0, -1, 0, 1, -2, 0, 1, -1, -1, -1, 0, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, -1, 1, -1, 0, 0, -2, -1, 0, 0, 1, -1, 0, 0, 0, 1, 0, 0, 1, 1, -1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 1, 2, 1, -1, 0, 0, 0, 1, 0, 1, -1, 1, -2, 1, 0, -1, -1, 1, 1, 0, 0, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, -1, 1, 0, -1, -1, 0, -1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, -1, 0, 0, 1, 0, 0, 0, -2, 1, -2, -1, -1, 0, 0, 1, 1, 0, 1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 1, 1, -1, 0, 1, 0, 0, 0, 2, -1, 0, 0, -1, 1, -1, 1, -2, -3, 0, -4, -1, -3, -1, -4, -3, -1, -3, -1, -1, 0, -1, -2, -2, -4, -3, -2, -2, -6, -3, -4, -6, -8, -3, -4, -5, -4, -6, -4, -1, -2, -2, -2, -3, -3, 0, -2, 0, -3, -2, -1, 0, -1, -2, -4, -2, -3, -3, -3, -2, -5, -2, -2, -5, -6, -5, -4, -3, -3, -4, -2, -2, -2, -1, -2, -1, -1, -1, 0, -3, 0, -2, -2, -1, -1, 0, -2, -2, -3, -5, -4, -2, -4, -1, -3, -5, -3, -2, -2, -2, -3, -3, -1, -1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -2, -3, 0, -2, -3, -2, -2, -3, -4, -1, -2, -3, -3, -2, -2, -3, 0, -2, 0, -1, 0, -1, 0, 1, 1, -1, 0, 0, -1, -2, -2, -4, -3, -1, -2, -2, 0, -3, -1, -3, 0, -2, 0, -2, 0, -3, 0, -1, -2, 2, 1, 1, 1, 0, -2, 1, 0, 0, -2, 0, 0, -2, -2, -2, 0, -2, 1, -2, 0, 0, -2, -1, -2, -2, -2, 0, 1, -1, 0, -2, 1, -1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 2, 0, 2, 0, 2, 1, -2, 0, 0, 0, 0, -2, -1, 2, 0, 0, 1, 0, 0, 1, 0, 2, -1, -2, -2, 0, 2, 0, 0, 0, 2, 1, 0, -1, 0, 0, 1, 0, 0, 2, -2, 0, 1, 0, 2, 1, 0, 2, 0, 1, 0, 1, 0, -3, -2, -1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 3, 1, 2, 2, -1, -1, -2, 0, 2, 2, 2, 2, 1, 0, 1, -1, 0, -1, -2, 0, -2, 0, 0, 2, 3, 0, 0, 2, 2, 0, 1, 1, 1, 1, 0, -1, 0, 0, 2, 0, 1, 0, 0, 1, 0, 1, -2, -2, 0, -3, 1, 1, 0, 1, 2, 1, 1, 0, 0, 2, 0, 0, 0, 0, 2, -1, 0, 2, 1, 1, 1, 2, 2, 0, 1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 4, 4, 1, 2, 0, 1, 2, 1, 0, 2, 1, 2, 1, 1, 5, 2, 4, 1, 0, 0, 0, -2, -3, 0, 0, 0, 1, 1, 1, 0, 2, 4, 2, 3, 2, 2, 5, 4, 2, 3, 1, 1, 1, 2, 4, 3, 4, 3, 4, 1, -1, -1, -1, 1, 0, 0, 1, 2, 2, 2, 1, 2, 3, 1, 1, 2, 4, 1, 3, 1, -1, 1, 1, 3, 5, 4, 2, 4, 4, 2, 2, 0, -1, 0, 0, -1, -1, 0, 0, 2, 2, 1, 0, 0, 3, 0, 1, 2, 2, 0, -1, 2, 2, 5, 4, 4, 3, 2, 2, 1, 0, 2, 0, -1, -1, -1, 0, -1, 0, 0, -1, 0, 2, 2, 2, 1, 2, 0, 3, 1, -1, 0, 1, 2, 4, 4, 5, 3, 4, 1, -1, 0, 1, 1, -1, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 2, 0, 0, 2, 0, 0, 0, 2, 5, 3, 2, 4, 5, 5, 2, 0, 0, 0, -1, 0, -1, 1, 2, 1, 1, -1, 0, 1, 2, 3, 3, 3, 0, 2, 0, -2, 0, 4, 4, 2, 5, 1, 4, 3, 2, 0, 2, 0, -1, -3, 0, 0, 0, 1, 2, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 3, 2, 2, 4, 0, 4, 2, 0, 3, 2, -1, -3, -3, -2, 0, -1, 1, 0, 1, 1, 3, 0, 0, 2, 4, 2, 1, 2, -2, 1, 3, 1, 2, 1, 3, 3, 3, 1, 0, 1, 0, -2, -1, -3, -1, 0, 3, 1, 0, -1, 2, 0, 0, 3, 1, 0, 1, 0, -4, 0, 1, 0, 0, 3, 3, 1, 4, 2, -1, 2, 0, -1, 0, -1, 0, 0, 3, 2, 3, 1, 0, 2, 1, 0, 1, 0, 1, 2, -1, 0, -1, 1, 1, 1, 2, 3, 0, 0, 0, -1, 1, -2, -3, 0, -1, 0, 0, 0, 2, 2, 1, 0, 2, -1, 1, 0, 0, 0, -4, -3, -2, -2, -1, 1, 2, 0, 0, 1, 0, -1, 0, -1, 1, 0, 2, 2, -1, 1, 1, 0, 2, 0, 3, 0, -1, 0, 0, -2, -1, -4, -3, -1, 1, 0, 0, 0, 1, 1, -3, 0, -1, -2, 0, 1, 0, 1, 3, 2, 3, 0, 2, 0, 0, -1, 1, 0, 0, 0, -4, -1, -3, -3, -1, 0, 0, 1, 1, -3, 0, 1, 0, -1, 0, -1, 1, 0, 0, 0, 1, 1, 2, 0, 0, 0, 1, -3, 0, 0, -6, -1, -4, -3, -4, 0, -1, 0, 0, 0, -3, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, -1, 1, 0, 2, -1, -1, 0, 0, -5, -3, -4, -2, -2, -2, 0, -3, 0, -2, -1, -1, 0, -2, 0, -3, -1, -3, 0, -1, -2, 0, 0, 0, 0, 1, -2, -2, -2, -2, -4, -5, -1, -4, -2, -4, -1, 0, -2, -4, -3, -2, -1, -4, -2, -2, -3, -3, 0, 0, -2, -2, -2, -3, -1, 0, -3, -3, -3, 0, -4, -3, -1, -1, -1, -3, -4, -3, -2, -1, -2, -2, -2, 0, -1, -4, -1, -2, 0, -4, -2, -1, 0, 0, -1, -3, -2, -3, -1, -1, 0, 1, 0, -1, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, -1, 0, 1, 0, -1, 0, -1, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 1, -2, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, -2, 0, 1, 0, -1, -1, 1, 1, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, 0, 0, 1, -1, 1, -1, 0, 0, 0, -1, 1, 0, -1, 0, 0, -2, -1, -1, 0, 1, -1, 0, 0, 0, -1, 0, -1, -1, -1, -2, 1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 1, 0, 1, 0, 0, -2, 0, -1, -1, -2, 0, -2, -2, 0, -2, 1, 1, 0, -1, 1, 1, 0, 0, -1, -1, 1, -1, 2, 0, 0, 1, -2, -1, -1, 0, 0, 0, -2, 0, -2, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -1, 1, 2, 0, 0, 1, -2, 0, -1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, 0, -1, 2, -2, -1, 0, 0, 0, 2, 0, -1, 0, -1, 0, 1, 0, -2, 0, 1, 2, 0, 1, -1, -2, 0, 0, 0, -1, 1, 0, 0, -1, 0, -2, 0, 0, -1, 2, 2, 0, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 1, 2, 2, 2, 2, 0, 0, -1, 1, 0, 0, -2, 0, 0, -2, -1, 0, 0, 1, 0, -1, 0, 0, 1, -2, 0, 0, 1, 0, 0, 0, 1, 2, 0, -1, 0, 0, -1, 0, 0, 0, -2, 0, 0, 0, -1, -1, -2, 0, 1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 1, -1, 0, 1, 1, 1, 0, 2, 0, 0, 0, 0, 1, 0, -2, 0, -2, -2, 0, 0, -2, -1, 0, -1, 0, -1, 0, 1, -1, 1, 2, 0, 1, 0, 0, 1, 0, 1, 0, 1, -1, 0, 0, 1, -1, 0, 0, 0, 0, -2, -2, 0, -1, 0, -1, 0, 1, -1, 0, 0, 0, 1, 3, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0, -1, -2, 0, -1, 1, -1, 0, 0, 1, 2, 0, 0, -1, 0, 0, 0, 1, 2, 0, -1, 1, 2, 1, 1, 1, 1, 0, -1, 0, 0, 0, -1, 0, 0, 1, -1, 1, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, -1, 0, 1, 1, -1, 1, 0, 1, 0, 0, 0, 1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 1, 0, 0, -2, 1, 1, -2, 0, -1, 0, 1, 0, 1, -1, 0, -1, 1, 1, 1, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, -2, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, -2, 1, 0, 1, 1, -2, 0, 0, 0, 1, 0, 0, 0, 1, 0, -1, -1, 0, 1, 0, 0, -1, 2, 0, 0, 1, 2, 1, 1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, -2, 0, 0, 1, -1, -1, 2, 2, 0, 0, 1, 1, 0, -1, -2, 0, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 2, 0, -1, 0, 0, 2, 0, 0, 0, 0, -1, -2, -2, -1, -1, -1, -2, 0, 0, 0, -1, -1, 0, -2, 1, -1, 1, 1, -1, 0, 1, 2, 0, 0, -1, -1, -1, 1, -1, 0, 0, 1, 0, 1, 0, 0, 1, -1, -2, -1, -2, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, -1, 0, 0, -2, 0, 0, 1, 0, -1, -2, 0, -1, -1, 0, 0, 0, 0, -1, -1, -2, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, -2, 0, 0, 1, 1, 0, 1, -1, 0, 0, -1, -1, -1, -1, -1, 1, 2, 0, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 0, -1, 1, -1, 0, -1, -1, 0, 1, 0, 0, -2, 0, 1, 1, 0, 1, -1, -1, 1, 0, 1, 0, 0, -1, 1, 0, 0, 0, -2, -1, -1, -1, -1, 0, -1, 2, 0, -1, 0, 0, 0, 0, 1, -1, -1, 0, 1, 0, -1, 0, 1, 0, -2, 0, 1, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 1, -1, 0, -1, 0, 1, 1, 1, -1, 0, -1, -1, 0, -2, -1, 0, -1, 1, 0, 0, -2, -1, 0, -1, 0, 0, -1, -1, 0, -1, 1, 0, 0, -1, 1, 0, 1, 1, 0, 2, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, -1, 0, 2, 0, 2, 0, 0, -1, 0, 1, 1, 2, -1, 0, -1, 0, 0, 0, 2, 2, 2, 0, 1, -1, -1, 0, 0, -1, 2, 0, -1, 0, -1, 0, 1, -1, 0, 2, 0, 1, 1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 2, 0, 0, 0, 0, 2, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 2, 0, 1, 0, 1, 0, -1, 1, 0, 0, 0, -1, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 2, 1, 1, 1, 0, 1, 0, 2, 0, 2, 0, 1, 1, 0, -1, -1, 0, 1, 2, 1, 1, 1, 0, 1, 1, 0, 2, 2, 0, 0, 0, 1, 0, 0, 0, 3, 1, 0, 0, 2, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 2, 0, -1, -1, 1, 0, 2, 0, 0, 0, 0, 0, 0, 1, 3, 0, 1, 3, 3, 1, 2, 0, 0, 1, 0, 0, 1, 0, -1, 0, 1, 0, -1, 1, 0, 0, 2, 1, 0, 0, 1, 0, 1, 3, 2, 1, 0, 0, 3, 0, 0, 2, 0, 0, 0, -1, 0, 0, 0, 2, 1, 0, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 3, 1, 2, 0, 0, 1, 2, 0, 1, 1, 2, -1, 0, -1, 0, 1, 1, 1, -1, 0, 1, 1, -1, 0, 1, -1, -1, 1, 2, 0, 0, 0, 1, 1, 0, 0, 1, 2, 0, 0, 0, 1, -1, 1, 1, 0, -1, 0, 1, -1, 0, 0, -1, 2, 1, 0, -1, 0, 0, 2, -1, 2, 1, 1, 1, 0, -1, 1, 0, 0, 0, 0, 1, -1, 0, -1, 0, -1, 0, 1, 0, -1, 1, -1, 0, 0, -2, 1, 0, 0, 0, 2, 0, -1, -1, 2, 2, 0, 2, -1, 1, 0, 0, -1, -1, -2, 1, 0, 1, 1, 0, 0, 1, -1, 0, -1, -2, -1, -2, -1, 1, 0, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, -1, 1, 0, 1, 0, 0, 1, -1, 0, 0, -2, -1, 0, 0, -1, 1, -1, 0, 0, -1, 2, 2, 0, 0, 2, -1, 0, -1, 1, 0, -2, 1, 0, 0, 0, 0, -1, -1, 2, -1, 0, 2, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 2, 2, 0, 0, -1, 2, 1, 0, 0, -1, 0, 1, 0, -1, -1, 0, -1, 0, 1, -2, -1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 0, -1, -1, 0, 0, 1, 0, -1, 1, 0, -1, 0, -1, -2, 2, 0, 1, -1, 0, 0, 0, 0, 1, 1, -1, -1, 0, 0, 3, 1, 1, 0, -1, 1, 0, 0, -2, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, 1, -1, 1, 0, 0, -1, 2, 2, 2, 2, 3, 0, 1, 0, 0, -1, 0, 1, -1, 1, 1, -2, 0, 0, -2, 1, 0, 1, -1, 1, 0, 0, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, -1, 0, 0, -1, -1, 0, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, -1, 1, 1, 0, 1, 1, 2, 0, 0, 0, 1, 0, -2, 0, 1, 1, 0, 0, 1, 1, 0, 1, 0, -1, -1, -1, 1, 0, 0, 0, 0, 2, 0, 2, 0, 1, 0, 0, 1, 1, -1, 0, 2, -1, 1, 1, 0, 0, 0, 1, 1, 1, 0, -1, 1, 0, 1, 2, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, -1, 0, 0, 2, 2, -1, 0, 1, 2, 0, 2, 2, 2, 2, 2, 1, 0, 1, 0, -1, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 2, 2, 0, 0, 0, 0, 2, 0, 1, 2, 0, 2, 1, -1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 2, 0, -1, 1, 2, 1, 1, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 2, 0, 2, 2, 0, 0, 0, 0, -1, -1, 0, -1, 2, 2, 0, 2, 0, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, 0, 0, 2, -1, 1, -1, -1, 1, 1, -1, 1, 0, 1, 0, 2, -1, 0, 0, -1, 0, -1, 1, 0, 0, 2, 0, 2, 1, 1, -1, 1, 1, 0, 1, 2, 0, 1, 2, -1, 0, 0, 0, 0, 2, 0, 2, -1, 0, 0, 1, 1, -1, 0, 0, 1, -1, 0, -1, 1, 0, 2, 0, 1, -1, 0, -1, 0, 2, 2, 0, 0, 1, 2, 0, 2, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, -1, 0, -1, 0, 0, -1, 1, 1, 1, 0, 2, 0, 2, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, -1, -1, 2, 0, 1, -1, 1, -1, 2, 0, 0, 0, -1, 2, 1, 0, 0, 1, 2, 2, -1, 0, -1, -1, 0, 1, -1, 0, 1, 0, 0, 1, 1, -2, -2, 0, -3, 0, -2, -2, 0, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, -1, 1, -1, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, -2, -2, 1, 0, -1, -2, 0, -3, 0, -1, 1, -1, -1, 0, -1, 0, 0, -2, -2, -1, -1, 1, -3, -2, 0, -2, -2, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, -3, 0, 0, 0, 0, 0, 1, 1, 1, 0, -3, -2, -1, 0, -2, -1, 0, -1, 0, -2, 0, -1, 0, -2, 0, 0, -2, 0, -3, 0, -2, 1, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1, -2, 0, 0, -2, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, 0, -1, -2, -1, -2, -2, 1, -1, 1, -1, -1, 0, 0, 0, 0, -1, -2, -1, -2, -1, 0, -2, 0, -2, -1, -2, -1, -2, -3, 0, 0, 0, -1, 0, 0, -1, -1, -2, -1, 0, -1, 0, 0, 0, -3, -3, -2, -1, 0, -1, -2, -2, 1, 0, -1, -2, 0, -1, 0, -1, -2, 0, -1, -1, 0, 0, -1, 0, 1, 1, 0, 0, -2, -1, -3, -1, -1, 0, -1, -2, 0, -1, 1, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -2, -1, -3, -1, -1, 0, 0, 0, 0, 0, -1, -2, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, -2, -2, -1, -3, -1, -2, 0, 0, -2, -2, -1, 1, -1, 1, 0, 1, -1, -3, 0, 0, -3, -3, -2, 0, 0, -1, -1, 0, 0, -1, 0, -3, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, -3, -2, 0, 0, -1, 0, -3, -3, -2, 0, -3, -2, 0, -1, -1, -3, -1, -1, 0, 0, 0, -1, -1, 0, 1, -1, 1, 0, -1, -3, -2, 0, -1, -1, 0, -3, -3, -3, 0, 0, 0, 0, -1, -2, -1, -3, -2, -1, 0, 0, 0, -2, -3, -2, 1, -1, 0, -1, -1, 0, -3, -2, -3, -2, -2, -1, 0, -1, 0, -1, 0, 0, 0, -2, -2, 0, -3, -3, -1, -3, 0, 0, -3, -3, -1, -2, -1, 0, 0, 0, 0, 0, 0, -3, -2, -2, -1, 0, -1, -3, -2, -3, -2, -1, 0, -2, -1, 0, 0, 0, -1, 0, -3, -1, -2, -1, 1, -2, -2, -2, 0, -1, -2, -2, -1, -1, 0, 0, -2, -2, 0, -2, -1, -2, -1, -1, -1, -1, -1, -3, 0, -3, -2, -3, 1, 0, 0, 0, 0, 0, -2, -2, -4, 0, -2, -1, -3, 0, -2, -3, -3, -3, 0, -2, -2, -2, -1, 0, 0, -3, 0, 0, -1, -2, -1, 1, 0, 0, -1, -2, -2, -3, -2, -3, -2, -4, -1, -2, -3, -2, -2, -1, -2, 0, -3, -3, 0, 0, -2, 0, -1, 0, -1, -1, 0, 0, -2, -2, -2, -1, -2, -2, 0, -1, -4, 0, -1, -1, 0, 0, 0, -2, -3, -2, -2, 0, -2, -2, -2, -1, -4, 0, 0, -3, -2, 0, -1, 0, 0, -3, -2, 0, 0, -3, -1, 0, -3, -1, 0, -2, 0, -1, 0, -3, -2, -1, 0, -3, 0, 0, -1, -1, 0, -2, 0, -2, -1, -2, -2, 0, 0, -2, -1, -4, 0, -4, -3, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, 0, 0, 0, -2, -1, 0, -2, -1, -1, -2, -2, -2, -2, -3, -1, 0, 0, 0, -3, -2, -1, 0, -2, -2, 0, 0, -2, -2, -3, 0, 0, 0, -2, -2, 0, 0, -1, 0, 0, -2, 0, -3, -1, -3, -3, -4, 0, 0, -2, -2, -1, 0, 0, 0, -1, 0, -3, -2, -3, -2, -1, 0, 0, 0, -3, -3, 0, -3, -1, 0, -2, 0, 0, -2, 0, -2, -2, -3, -1, -1, -2, -1, 0, 0, -2, 0, 0, 0, 0, -2, -1, 0, 0, -2, 0, 0, -2, -2, -1, 0, 0, -2, -1, -3, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 0, -2, -2, 0, -1, 0, -3, 0, 0, -1, -3, 0, -2, -3, 0, 0, -1, -1, -3, -2, 0, -1, 0, -2, 0, -1, -1, 0, 0, 0, -2, -3, -3, -1, 0, 0, -2, 0, -2, -1, -1, -4, -3, -1, 0, 0, -2, 0, 0, -1, -2, 0, 0, 0, -3, -1, 0, 0, 0, -1, -2, -1, -2, -3, -2, -3, -3, -1, 0, -1, -2, 0, -2, 0, -2, 0, 0, 0, -3, 0, -1, -1, -2, -2, -3, -2, 0, 0, -2, -2, -1, -3, -3, -1, -2, -2, -2, -2, 0, -1, -2, -1, 0, -1, 0, -2, -1, -2, 0, -1, 0, 0, -3, -3, -3, 0, -2, -1, 0, -3, -2, 0, -3, -2, -3, 0, -2, -3, -2, -2, 0, -1, -1, 0, -1, -1, 0, -2, -1, 0, -1, 0, -2, -1, -1, 0, -1, 0, -2, -1, -4, 0, -2, -4, -2, -1, -3, 0, -2, -1, -3, 0, 0, 3, 1, 0, 2, 2, -1, 0, 2, 2, 0, 2, 1, -1, 1, -2, -2, -1, -1, -1, 0, -4, -3, -6, -6, -4, -4, -4, -6, -4, 1, 0, 3, 0, 1, 2, 0, 1, 0, 0, 3, 1, 3, 1, 0, 0, 0, -2, 0, -2, 0, -1, -3, -1, -5, -5, -5, -3, -5, -6, 3, 2, 0, 1, 0, 2, 0, 0, 1, 3, 3, 0, 2, 0, -1, -2, 0, -1, -1, -3, -1, -2, -2, -1, -3, -3, -1, -3, -4, -3, 0, 1, 2, 0, 0, 1, 3, 0, 2, 2, 1, 2, 0, -1, 0, 0, -3, 0, 0, -1, -2, 0, 0, -3, -3, -1, -2, -2, -4, -1, 1, 4, 2, 2, 4, 3, 3, 3, 2, 1, 1, 3, 0, 0, -2, 0, -1, -1, 0, 0, 0, -1, -1, -2, 0, -3, 0, -1, -4, -2, 3, 2, 3, 4, 4, 6, 4, 2, 3, 3, 4, 2, 0, -1, 0, -2, 0, -1, -2, -1, -1, 0, 0, 1, 0, -1, 0, -2, -3, -2, 3, 2, 2, 6, 5, 5, 4, 5, 3, 4, 1, 4, 0, 0, -1, 0, -2, 0, 1, 0, -2, -2, 2, 2, 1, 1, 0, 0, 0, 1, 2, 5, 2, 6, 4, 4, 3, 2, 6, 5, 4, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, 3, 0, 0, 2, 3, 4, 5, 6, 5, 5, 5, 6, 2, 3, 5, 3, 2, 1, 1, -1, -2, 0, 1, -1, 0, 1, 0, 1, 2, 2, 1, 0, 0, 1, 1, 3, 3, 6, 5, 7, 7, 6, 3, 4, 3, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, -1, 1, 1, 2, 3, 3, 3, 3, 1, 2, 3, 3, 6, 5, 7, 3, 4, 4, 4, 2, 0, 0, -3, -2, -1, -1, -2, -1, 0, 2, 2, 1, 1, 0, 2, 1, 4, 3, 1, 2, 4, 3, 7, 6, 7, 5, 6, 5, 4, 0, -1, 0, 0, -2, -2, -3, -1, -2, 0, 1, 1, 2, 2, 0, 1, 3, 1, 2, 3, 0, 5, 3, 5, 6, 8, 4, 4, 4, 2, 0, 0, 0, 0, -3, 0, 0, -1, 0, 0, 0, 1, 3, 1, 3, 4, 2, 5, 2, 3, 0, 5, 3, 4, 8, 8, 4, 3, 4, 1, 0, -1, 0, -1, -3, -3, -4, -2, -1, -4, -3, -1, 1, 1, 1, 2, 3, 3, 1, 1, 1, 2, 4, 6, 6, 4, 4, 4, 4, 3, 1, 0, -2, -3, -1, -4, -2, -1, -3, -3, -3, 0, 0, 1, 0, 0, 2, 3, 5, 3, -1, 3, 4, 4, 5, 4, 7, 4, 4, 2, 0, 2, -1, 0, -2, -1, -3, -2, -3, -3, -2, 0, -2, -2, 0, 0, 0, 0, 2, 2, 1, 5, 6, 3, 5, 5, 6, 4, 2, 3, 1, 1, -2, -2, -1, -1, -3, -2, -2, -2, 0, -2, 1, -1, 0, 3, 2, 3, 0, 1, 2, 3, 6, 5, 3, 5, 6, 6, 6, 0, 2, 0, 0, 0, 0, -5, -5, -3, -4, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 2, 0, 3, 4, 5, 3, 3, 7, 6, 6, 1, 1, -1, -1, 0, -3, -2, 0, -3, -2, -1, -1, -1, 0, 0, 0, 2, 4, 1, 3, 2, 1, 4, 3, 4, 5, 6, 2, 3, 3, 3, 4, 3, 0, -3, -4, -5, -2, -2, 0, 0, 0, 0, 0, 0, 2, 1, 3, 0, 0, 0, 2, 5, 5, 5, 5, 5, 2, 2, 3, 3, 1, 1, 0, -3, -2, -1, -1, -1, 0, -1, 2, 2, 0, 3, 0, 1, 2, 2, 3, 1, 0, 3, 3, 3, 5, 2, 5, 5, 4, 3, 2, 0, 0, 0, -2, 0, 0, 0, 3, 1, 2, 3, 0, 0, 2, 0, 1, 0, 2, 1, 0, 1, 0, 2, 4, 3, 2, 5, 2, 2, 2, 1, 1, 1, 0, -1, 1, 0, 2, 3, 3, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 4, 1, 3, 3, 5, 4, 3, 4, 2, 2, 0, 0, 0, -1, -1, 2, 2, 0, 0, 1, 0, 1, 1, 0, 0, -2, 0, 0, -1, 0, 2, 3, 4, 1, 1, 2, 1, 0, 3, 0, 0, 0, 0, 0, 1, 0, 1, 1, 2, 0, 2, 1, 1, -2, 0, -1, 0, -2, -2, 1, 0, 1, 2, 3, 3, 3, 0, 3, 2, 3, 2, 1, -1, -1, 0, 0, 0, 2, 1, 1, 0, 1, 0, 0, -1, 0, 0, -3, 0, 0, 2, 2, 2, 4, 2, 1, 0, -1, 1, 0, 0, 0, 0, 0, 1, -1, 0, 2, 1, 0, 0, 2, -1, 1, -1, -2, 0, -1, -1, 0, 0, -1, 1, 0, 2, 2, 2, 1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 2, 0, -1, -2, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, -1, -1, 0, 0, -2, 0, 0, -2, 0, -2, -1, 0, -1, -1, 0, -2, -2, -3, -3, 1, 1, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, -3, 0, -3, -1, -3, -2, -2, -3, -2, -2, -3, -1, 0, -3, -2, -1, -3, 0, -1, 0, -1, -1, 0, 0, 0, 1, 0, 0, 1, -1, 2, 1, 0, 1, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, 1, -1, 2, 0, 0, -1, 1, 0, -1, 2, 0, 1, 1, 0, 1, -1, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 0, 1, 2, -1, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 1, -1, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, 1, -1, 0, 2, -1, -1, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, -1, 0, 1, 0, 1, 1, 2, -1, 0, 0, 0, 0, 0, -1, 1, -1, -1, 0, 1, 1, -2, 0, 0, 2, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 1, 1, -1, 1, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, -1, 1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 2, -1, 0, 0, 0, -1, 0, 1, 1, -1, -1, 0, 1, 0, 1, -2, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, 2, -1, 2, -2, -1, -2, 1, -1, -1, 0, -1, -1, 1, 1, 1, 0, 2, 1, 2, -1, -2, 0, -1, 0, -1, -1, 1, -1, 0, 2, 0, 1, -1, -1, -1, 0, -1, 0, -1, -1, 2, 1, -1, 0, -1, -1, -1, 1, 1, 0, 1, 1, 0, 0, 1, 0, -1, -1, 1, 1, -1, 0, -1, 1, -1, 1, 0, 0, -1, 1, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 1, 0, -1, 1, 0, -1, 0, 1, 2, 0, 0, -1, -1, -1, 0, 1, 0, 1, 0, -1, -1, -2, 0, 1, -1, 0, -2, 0, 0, 1, -2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, -1, 1, 0, 1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, -1, -1, 0, 1, -1, 2, 1, -1, -1, 1, -1, -1, 2, 0, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 2, -1, 0, 0, 0, 1, 1, 0, -2, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 2, 0, 0, -1, 0, 1, -1, -2, 0, 1, -1, -1, 0, 0, -1, 1, -2, 0, -1, -1, 1, -1, 0, 2, 0, 0, -1, 1, 2, -1, 0, 0, 2, 1, 0, -1, 1, 1, 0, 0, 1, 0, -1, 0, 1, 0, 0, -1, 0, -1, -1, 1, -1, 1, 1, 0, -1, 1, 2, 0, 0, 0, -1, 1, 1, 1, -1, -1, -1, -1, -1, 1, 0, -1, -1, 0, 1, 1, -1, 0, 0, 1, 2, 1, 0, 2, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -1, -1, 0, -2, -2, -1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, -1, 2, -1, 1, 0, 0, -1, 0, 0, -1, 0, 2, 0, -1, -1, 0, 0, 0, 1, 1, 1, 0, -2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 2, 2, 1, 0, 1, 0, -1, 1, 0, -1, 0, 1, 0, 0, -1, 2, -1, 0, 1, -1, 1, 0, 0, 0, -1, 2, 1, 0, 1, 0, 0, 0, 1, 1, 1, 1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 1, -1, -1, 0, 0, -1, 0, 0, -1, 0, 2, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 1, 1, -1, 1, 1, 1, 2, 1, 0, -2, -1, 1, 0, -1, -1, -1, 0, 0, -1, 1, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 1, -1, 1, -1, 1, -1, -1, 1, 2, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, -1, 1, 0, 0, 0, 0, -1, 1, -1, 1, -1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 2, 1, 1, 0, -2, 1, 0, 0, -2, -1, 0, 1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, -2, -1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, -1, 1, 2, -1, 0, 1, 0, -1, 0, 1, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 0, -1, -1, 1, 0, 1, -1, 0, 0, 0, -1, -1, 1, -1, 0, 0, 0, 0, -1, 0, 1, -1, 1, -1, -1, -1, -1, 0, 0, -1, -1, 0, 0, -2, 1, 1, 1, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, -1, 0, 1, 0, 0, 1, 0, -1, 1, 1, 1, 0, -1, 0, 0, 0, 1, 1, 0, 0, -1, 0, -1, 1, 0, -1, 0, 1, 0, 1, 0, -1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 1, 1, 0, 0, 0, 1, 0, -1, -1, -1, 0, -1, -2, 0, 0, -1, 1, 0, 1, 0, 1, -1, 1, 1, -1, 0, 0, 1, -2, -1, 0, 0, -1, 1, -1, 1, 0, 0, 1, -1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, -1, 0, -1, -1, 1, -2, 0, -1, 0, 0, 1, -1, 0, 0, -2, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 1, 1, 0, -1, 1, 0, 0, -1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 1, 0, 1, -1, -2, 1, -1, -1, 0, 1, 1, 1, 1, -2, 0, -1, -1, -1, 0, 0, 0, -1, 1, 0, 0, -1, -1, -1, 1, -1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, -2, -1, 0, 0, 0, -1, 0, 1, -1, -2, 0, 1, 1, -1, -1, 1, -2, 0, 0, 0, 1, -1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, -1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 0, 1, -1, 2, 1, 0, -1, -1, 0, 0, 0, 0, 0, 1, -2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, -1, -1, 0, -1, -2, 1, -1, -1, 0, 0, -1, 0, -1, 0, 0, 2, -1, -1, 2, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, 1, -2, 1, 1, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 0, 1, -1, -1, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, -1, 1, 0, 0, -1, -1, 1, -1, 0, 0, 0, 2, -1, 1, 1, -1, 0, 0, 1, 0, -1, 1, 0, 1, 1, 1, 0, -1, -2, 1, -1, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 1, 0, 1, -1, 1, 0, 0, 0, -1, 0, 0, 1, -1, 2, 1, 0, -1, 1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 0, 2, -1, 0, 1, 1, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, -1, 2, 0, 1, 0, 0, 0, -1, -1, -1, 2, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, -1, 1, -1, 0, 0, -1, 1, 1, 0, 1, 0, -1, -1, 1, 0, 0, 1, -1, -1, 2, 0, -1, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, 1, 2, 0, 0, 0, 1, 0, 0, 1, -2, 2, -1, 0, -1, -2, 1, 1, 0, 0, 0, 1, 0, -1, 0, -2, 0, -1, 1, 0, 0, 0, 0, -1, 0, 1, 0, -1, 1, 0, 0, 2, 0, 0, 0, 1, -1, 1, -1, 2, 1, 0, 2, 1, -1, 0, 1, -2, 0, 0, 1, 0, -1, 0, -1, 0, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 2, -1, 1, 1, -1, 2, -1, 1, 1, -1, 0, 0, -1, -2, -1, 0, 0, -1, -1, 0, 0, 1, -1, 0, 1, 2, 0, -1, 0, 0, 1, -1, 0, -1, 0, 1, -1, 0, -1, 0, 1, 0, 1, 0, 0, 1, 1, 0, -1, -1, 0, -1, 1, 0, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -2, 0, 2, 0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, -1, -1, 0, -1, 0, -1, 0, 1, 0, -1, 1, 0, -2, 0, 1, 0, 1, 1, -1, 0, 0, -1, -1, 1, 0, -1, 0, 1, -1, 1, 1, 0, -1, -1, 0, 1, -1, 0, -2, 0, 1, -2, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, -1, -1, 2, 2, -1, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, 1, -1, 1, -1, -1, -1, 1, 0, 1, 1, 2, -2, 0, 1, -1, -1, 0, 1, 1, -1, 0, 0, 1, 0, 0, 1, -2, 1, 0, 0, -1, 0, 1, -1, 0, 1, 0, -2, 0, -1, 0, -2, 2, 0, -2, -1, 0, 0, 0, -6, -6, -2, -2, -6, -4, -4, -2, -5, -2, -1, -3, -2, 0, -2, -2, -3, -5, -4, -6, -6, -10, -10, -11, -9, -10, -7, -10, -8, -8, -9, -3, -2, -5, -6, -4, -3, -2, -2, -3, -3, -1, -3, -2, -3, -2, -4, -4, -5, -2, -5, -6, -8, -5, -6, -5, -5, -5, -8, -6, -8, -5, -6, -6, -6, -5, -3, -2, -1, -2, -4, -3, -3, -4, -4, -4, -2, -5, -3, -4, -4, -5, -3, -4, -5, -5, -3, -4, -5, -7, -8, -4, -5, -3, -6, -1, -2, -3, -1, -1, -3, 0, -3, -3, -2, -4, -5, -4, -3, -4, -4, -4, -1, -3, -4, -2, -2, -3, -3, -3, -6, -2, -1, -2, 0, 0, 0, -2, -3, 0, -2, 0, -2, -4, -3, -2, -1, -1, -3, -3, -2, 0, -3, -1, -1, 1, 0, 0, -2, -5, -5, -5, -4, 0, 0, 0, -1, -1, -2, -1, -2, -1, -1, -2, 0, 0, -1, -1, 1, -1, -1, 0, 0, 0, 1, -1, 0, 0, 0, -3, -6, -2, 0, -2, -1, 0, 0, 0, 0, 0, 1, -2, -1, -1, -1, 1, 1, 2, 1, 1, 3, 0, -1, 0, 0, 2, 0, 1, 0, 0, -4, -1, -1, 0, 0, 0, 1, 1, 0, 2, 0, -2, -3, 0, 0, 0, 0, 2, 3, 2, 1, 0, 0, 2, 0, 4, 1, 3, 0, 0, -7, -3, 1, 1, 0, 3, 1, -1, -1, 0, 1, -1, -3, 0, 0, 0, 3, 3, 3, 1, 3, 0, 0, 0, 1, 4, 5, 1, 2, 0, -4, 0, 2, 4, 2, 3, 3, -1, -1, -1, -1, 0, 0, -1, 2, 1, 4, 4, 3, 5, 5, 1, 2, 1, 3, 4, 5, 3, 5, 3, -4, 1, 3, 4, 3, 3, 1, 1, 0, 0, -2, -1, -2, -2, 3, 3, 3, 6, 7, 7, 2, 2, 1, 1, 5, 4, 5, 4, 3, 2, -1, 2, 3, 7, 7, 7, 5, 1, 0, -1, 0, 0, 1, 0, 0, 1, 4, 3, 4, 4, 7, 4, 1, 4, 4, 4, 4, 5, 5, 3, -1, 2, 5, 6, 8, 8, 7, 1, 1, 0, 0, 1, 0, 3, 2, 3, 2, 4, 4, 3, 3, 5, 6, 4, 5, 7, 5, 2, 1, 0, 0, 4, 8, 8, 10, 8, 8, 4, 4, 2, 0, 1, 0, 0, 2, 2, 1, 3, 4, 2, 4, 3, 4, 4, 2, 3, 4, 4, 3, 2, 1, 4, 8, 9, 8, 8, 6, 6, 4, 2, 4, 1, 0, 0, 1, 1, 4, 2, 3, 3, 4, 5, 5, 1, 1, 4, 3, 0, 3, 0, -2, 3, 9, 8, 8, 7, 7, 4, 6, 4, 3, 0, 1, 0, 2, 1, 3, 4, 3, 2, 2, 2, 1, 0, 1, 0, 1, 3, -1, -1, 0, 7, 9, 10, 8, 7, 9, 6, 3, 4, 0, -1, 0, -1, 3, 1, 1, 1, 1, 2, 4, 2, 1, 3, 3, 3, 0, 0, -1, 0, 1, 5, 8, 6, 9, 8, 7, 7, 3, 4, 0, -1, -1, 0, -1, 1, 3, 2, 1, 2, 2, 2, 3, 3, 2, 1, 1, 2, 0, 0, 1, 4, 4, 7, 7, 9, 7, 4, 4, 3, 2, 0, 0, -4, 0, 0, 3, 0, 3, 3, 3, 0, 2, 2, 3, 4, 2, 1, 1, 1, -2, 2, 2, 6, 5, 6, 4, 3, 4, 5, 0, -2, -1, -3, -2, -3, -1, 2, 0, 3, 1, 3, 2, 1, 5, 5, 3, 0, 1, 2, -4, 0, 4, 6, 5, 7, 5, 5, 3, 1, 1, -1, -2, -3, -5, -1, -1, 1, 3, 2, 2, 2, 3, 0, 4, 2, 0, 2, 2, 1, -3, -3, 2, 0, 3, 5, 3, 5, 1, 0, 0, 0, -3, -1, 0, -1, 2, 2, 4, 0, 3, 3, 1, 3, 1, 3, 0, 0, 1, 0, -6, -2, 0, 0, 3, 1, 3, 2, 0, -2, 0, -2, -1, -2, 0, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 2, 0, -1, -2, -6, -4, -3, -1, 0, 1, 3, 1, 0, 0, -2, 0, -1, -2, -1, 1, 0, 0, 1, 3, 4, 5, 4, 6, 1, 2, 1, 1, -1, 0, -7, -7, -3, -3, -2, 1, 0, 1, 0, -2, 0, -2, -1, 0, 1, 1, 2, 0, 1, 3, 2, 3, 4, 4, 2, 0, 0, 0, 1, -3, -10, -8, -3, -4, -2, -1, 0, -1, -2, -3, -1, -1, -1, 0, -2, 0, 2, 1, 1, 2, 4, 0, 1, 4, 0, 0, 0, 0, -1, -3, -8, -8, -6, -5, 0, -2, -1, -2, -2, -4, 0, -2, -3, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, 2, 0, -1, -1, -3, -2, -4, -9, -5, -5, -4, -3, -2, -4, -5, -4, -2, -3, -4, -4, -4, -4, -1, -1, -3, -2, 0, 0, -1, -1, 1, 0, -3, -1, -4, 0, -4, -7, -8, -6, -5, -4, -2, -3, -5, -5, -2, -4, -3, -3, -4, -1, -4, -4, 0, -3, -3, -5, -5, -3, -1, -1, -4, -4, -2, -3, -6, -7, -5, -5, -3, -3, -5, -6, -4, -3, -5, -5, -2, -5, -3, -3, -2, -3, -6, -3, -3, -5, -6, -6, -4, -5, -5, -8, -6, -6, -7, -4, 0, 0, 0, 0, -2, -1, 0, -2, 0, 0, -1, 1, 0, 1, 0, -1, 0, -1, 0, -1, 0, -3, -3, 0, 0, -1, 0, 0, -3, 0, -1, -2, -1, -1, 0, 0, 0, 0, 0, 1, -1, 1, 0, -1, 1, -1, -2, -2, 0, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -1, 0, 0, -1, 0, 0, -1, 0, 1, 0, 0, 1, 0, -1, -1, 1, -1, 0, 0, -2, 0, -1, -1, 0, 0, -1, -2, -2, -3, -2, -1, -2, -1, 0, 0, 0, 1, 1, 1, -1, -2, 0, -1, -1, -2, 0, 0, 1, 0, -2, -1, 0, 1, 0, 0, 0, -1, 0, -2, -1, 0, -1, -1, 0, 0, 1, 1, -1, 1, 1, 1, 0, -1, 1, 0, -1, 0, -1, 0, 0, -1, 0, 1, -1, -1, 1, -1, -1, -4, 0, -1, -1, 0, 1, -1, -1, 0, 1, 1, 0, 0, 1, 2, 0, 1, 1, -1, 0, 0, 2, -1, 0, 2, 0, 1, 0, 0, 1, -3, -1, 0, -1, 1, 1, 1, 1, -1, 0, 0, -1, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 2, 0, 2, 1, 0, 0, 1, 1, -1, -1, -1, 1, 1, 0, 1, 0, 0, 2, 1, 1, 0, 0, 2, 2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 3, 1, 0, 2, 0, -2, -1, 0, -1, -1, 1, 0, 0, 0, 1, 1, 0, 2, 1, 2, 0, 0, 1, 1, 1, 0, 0, 1, 0, 1, 2, 3, 0, 3, 0, 0, 0, -1, 2, 1, 1, 0, 0, 2, 0, -1, 0, -1, 1, 0, 1, 3, 2, 0, 1, 0, 1, 1, 2, 0, 0, 3, 1, 2, 0, 0, 1, 1, 0, 0, 2, 0, 1, 1, 0, 0, -1, 2, 0, 3, 1, 1, 0, 0, 0, 3, 2, 2, 0, 0, 3, 2, 0, 0, 2, -1, -1, 0, 2, 0, 0, 2, 0, 3, 0, 2, 0, 3, 2, 0, 0, 2, 1, 3, 1, 2, 1, 1, 3, 1, 0, 0, 1, 2, 1, -2, 1, 0, 1, 0, 0, 2, 0, 0, 2, 0, 0, 1, 0, 3, 2, 1, 0, 1, 2, 2, 2, 0, 2, 0, 0, 1, 3, 3, 0, 0, 1, 2, 4, 2, 1, 1, 1, 1, 1, 0, 3, 0, 2, 1, 2, 2, 1, 3, 2, 2, 1, 1, 3, 3, 1, 1, 0, 2, 2, 0, -1, 0, 3, 2, 0, 3, 2, 3, 1, 0, 2, 0, 3, 0, 1, 3, 1, 2, 0, 3, 3, 0, 0, 3, 0, 0, 0, 0, 2, -2, 1, 3, 4, 4, 3, 3, 4, 1, 0, 1, 0, 2, 1, 1, 4, 3, 0, 3, 2, 0, 1, 2, 0, 0, 1, 2, 1, 0, 0, -1, 1, 2, 1, 3, 2, 3, 0, 1, 0, 3, 1, 0, 2, 1, 2, 1, 2, 0, 0, 3, 3, 1, 3, 2, 1, 2, 0, 1, 0, -1, 0, 0, 1, 4, 2, 4, 4, 2, 0, 1, 1, 3, 2, 0, 1, 0, 1, 0, 0, 2, 1, 0, 2, 0, 0, 1, 2, 0, 2, -2, -1, 1, 0, 0, 2, 3, 3, 1, 0, 0, 0, 1, 0, 1, 0, 2, 1, 0, 1, 1, 1, 3, 1, 1, 2, 2, 0, 0, 0, 0, 0, 2, 3, 2, 3, 1, 1, 2, 2, 0, 2, 1, 0, 2, 0, 0, 0, 2, 2, 0, 0, 1, 2, 1, 2, 2, -1, 2, 2, -1, 1, 0, 1, 0, 3, 3, 2, 1, 2, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, -2, -2, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 2, 2, 1, 0, 1, 2, 0, 1, 2, 0, 2, 0, 0, -3, 0, -2, 2, 1, 1, 0, 0, 2, 0, 1, 2, 1, 2, -1, 1, -1, 2, 1, 0, 1, 0, 2, 0, 2, 3, 1, 2, 1, 1, -4, -3, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 2, 0, 0, 0, 0, 1, 2, 0, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 1, 1, 1, 2, 0, 0, 2, 1, 0, 2, 2, 0, 1, 2, 0, 0, 1, 1, 0, 1, -4, -4, 0, -1, 0, -1, 0, 1, 0, 0, 1, 2, 0, 2, 1, 1, 0, 1, 2, 2, 2, 2, 0, 2, 2, 2, 1, 1, 2, 0, -1, -4, -1, 0, -1, 0, 1, 0, 1, -1, 0, -2, -1, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, -1, 0, 1, 2, -3, -2, -3, -1, -1, -1, -1, 0, -2, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, -1, 0, -1, 1, 0, 0, -1, 0, -1, -1, 0, 0, -2, -2, 0, 0, -2, -1, 0, 0, -1, -1, -1, 0, 0, -1, -2, 0, -2, 0, -1, 0, 1, -1, 0, 0, -2, -1, -1, -1, -2, -2, -3, -3, -2, 0, -3, 0, 0, -1, 0, 1, 0, -2, 0, 0, 0, -1, 0, 0, -2, -3, -2, -1, -3, 0, -2, 0, 0, -2, -12, -9, -6, -6, -4, -7, -4, -4, -5, -3, -2, -1, -4, -2, -1, -4, -7, -6, -5, -7, -8, -8, -11, -11, -11, -8, -8, -9, -11, -8, -10, -10, -7, -9, -6, -7, -6, -2, -4, -2, 0, -3, -2, -4, -4, -2, -7, -6, -4, -5, -4, -6, -9, -7, -6, -3, -5, -7, -7, -7, -12, -9, -4, -6, -4, -6, -1, 0, 0, -2, 0, 0, -2, -3, -6, -3, -5, -3, -2, -5, -4, -5, -2, -2, -2, 0, 0, -4, -5, -8, -11, -7, -4, -2, -3, -2, 0, 0, 0, -2, -2, -3, -3, -2, -2, -4, -2, -2, -2, -1, -1, -2, -2, 0, 0, 0, 0, 0, -2, -3, -9, -4, -5, 0, 0, -2, 1, 0, -1, 0, 0, 0, -2, 0, 1, 0, 0, 2, 3, 0, -1, 2, 0, 2, 1, 3, 1, 1, -1, 0, -9, -4, -3, -2, -1, -2, 1, -1, 2, 1, 3, 1, 0, 2, 1, 1, 4, 4, 2, 3, 6, 1, 2, 2, 5, 3, 4, 1, 1, 0, -8, -2, -1, 0, 0, 1, 0, 0, 1, 3, 4, 1, 0, 2, 0, 3, 2, 3, 3, 5, 5, 4, 4, 3, 6, 6, 5, 7, 5, 1, -9, -6, 0, 3, 2, 2, 2, 0, 2, 2, 2, 1, 0, 0, 0, 3, 4, 7, 6, 5, 6, 3, 3, 5, 5, 8, 8, 9, 6, 4, -8, -3, 0, 6, 5, 3, 6, 4, 4, 1, 3, 1, 1, 0, 1, 4, 6, 8, 9, 7, 5, 8, 6, 7, 6, 11, 8, 10, 7, 5, -6, -1, 3, 7, 6, 9, 7, 5, 5, 3, 0, 0, 0, 2, 4, 4, 8, 11, 11, 11, 10, 9, 7, 7, 5, 7, 8, 9, 8, 2, -2, 0, 3, 9, 11, 11, 10, 5, 3, 0, 1, 0, 4, 4, 4, 7, 10, 9, 8, 10, 13, 11, 7, 7, 6, 9, 7, 7, 9, 5, 0, 5, 10, 10, 12, 14, 12, 7, 6, 2, 2, 0, 2, 4, 4, 7, 8, 8, 7, 10, 10, 9, 10, 10, 7, 10, 9, 10, 9, 5, 0, 5, 8, 12, 13, 15, 11, 10, 9, 7, 5, 4, 1, 2, 3, 5, 8, 6, 5, 9, 7, 9, 9, 10, 10, 9, 10, 7, 8, 5, -2, 4, 11, 14, 15, 15, 12, 12, 9, 7, 9, 7, 2, 5, 3, 4, 8, 9, 5, 7, 9, 9, 6, 6, 7, 5, 7, 5, 6, 1, 0, 4, 10, 12, 14, 15, 14, 11, 10, 7, 6, 4, 1, 4, 6, 5, 7, 6, 4, 7, 7, 6, 7, 8, 5, 6, 5, 5, 2, 2, -1, 5, 11, 13, 16, 15, 17, 12, 11, 6, 3, 5, 2, 1, 2, 7, 7, 6, 3, 5, 5, 7, 6, 5, 7, 8, 3, 6, 2, 2, -2, 8, 13, 13, 16, 17, 15, 14, 13, 8, 5, 4, 3, 0, 2, 6, 5, 6, 4, 6, 8, 7, 7, 7, 7, 7, 7, 5, 1, 0, -3, 6, 9, 13, 13, 15, 15, 13, 8, 8, 5, 6, 1, -2, -1, 3, 4, 3, 4, 6, 7, 7, 9, 8, 5, 6, 8, 6, 4, 2, -3, 4, 7, 11, 10, 9, 10, 9, 9, 8, 7, 6, 0, -4, -4, -2, 3, 6, 6, 4, 6, 5, 9, 9, 6, 7, 5, 5, 1, 0, -5, 1, 6, 9, 8, 10, 10, 10, 7, 6, 5, 1, -1, -2, -2, 0, 2, 6, 5, 4, 3, 6, 7, 6, 6, 5, 8, 5, 3, 1, -7, -2, 3, 5, 6, 9, 10, 8, 7, 6, 2, 3, 3, 1, 1, 0, 4, 6, 7, 6, 6, 3, 6, 4, 5, 5, 6, 5, 3, 3, -9, -2, 0, 3, 7, 5, 8, 7, 3, 1, 0, 2, 1, 0, 0, 4, 4, 3, 4, 4, 4, 5, 4, 3, 4, 4, 2, 4, 2, 2, -11, -7, -1, 0, 0, 5, 2, 3, 1, 1, -1, 0, 1, 1, 4, 5, 3, 4, 2, 2, 6, 7, 7, 7, 6, 4, 3, 4, 2, 0, -12, -7, -3, -2, 1, 3, 2, 2, 1, -1, -3, 0, 0, -1, 1, 5, 3, 5, 5, 8, 5, 5, 6, 9, 9, 7, 3, 3, 0, 1, -14, -11, -9, -5, 0, 0, 0, 0, -2, -3, -2, 0, 0, 0, 1, 1, 2, 5, 7, 6, 4, 4, 5, 6, 5, 6, 3, 1, 3, 0, -13, -11, -11, -7, -5, 0, 0, 0, -3, 0, -2, -2, -1, 0, 0, -2, 1, 0, 2, 2, 5, 4, 3, 6, 3, 1, 0, 2, 0, 0, -10, -9, -8, -7, -7, -4, -2, -4, -4, -4, -1, -2, -3, -2, -1, -4, -3, -1, -1, 0, 0, -1, 1, 1, 3, 0, 1, -2, -2, -3, -11, -8, -8, -6, -5, -6, -3, -5, -4, -3, -3, -3, -2, -3, -4, -5, -3, -2, 0, -1, -2, -2, -3, -2, -1, 0, -4, -4, -3, -2, -9, -9, -11, -8, -6, -9, -7, -4, -6, -3, -3, -5, -6, -2, -5, -4, -4, -4, -5, -7, -6, -6, -7, -7, -8, -8, -5, -8, -5, -8, -9, -9, -8, -10, -6, -6, -6, -7, -5, -5, -6, -4, -6, -2, -5, -5, -6, -8, -7, -11, -9, -11, -10, -10, -12, -12, -12, -11, -12, -9, -2, -1, -1, -3, -1, -1, -1, -1, -1, -2, 0, -2, -2, -1, 0, -3, -4, -4, -1, -3, -4, -6, -6, -4, -3, -2, -4, -3, -2, 0, -4, 0, -2, -2, -2, -1, -4, -3, -1, -4, -3, 0, 0, 0, 0, 0, -3, -4, -3, -3, -5, -3, -3, -4, -3, -3, -3, -5, 0, -2, -2, -3, -4, -1, -3, 0, -2, -3, -4, -1, -4, 0, -2, -3, -2, -2, -4, -2, -3, -2, -3, -2, -4, -2, -3, -4, -4, -3, -4, 0, -2, -2, -2, -3, -3, -1, -3, 0, -2, -3, 0, -1, -2, 0, 0, -1, -2, -2, 0, -1, -1, -2, -1, 0, -1, 0, 0, -3, -2, -2, -2, -1, 0, -4, -1, -1, -2, -1, -2, 0, -2, -4, -1, -1, -4, -2, -3, -3, -4, 0, -3, -2, 0, 0, -2, -1, 0, -3, -3, -2, -3, -2, -1, 0, -2, 0, -2, 0, -1, -1, 0, -3, -1, -2, 0, -3, -1, 0, -3, -3, -2, -1, -2, -2, -2, 0, -2, -2, -1, 0, -2, 0, -3, 0, 0, 0, -1, -3, -2, 0, -3, -1, -2, -2, -2, 0, -1, 0, 1, -2, -1, 0, 0, 2, -1, 0, 0, -2, -1, -1, 1, -2, 0, -1, -4, -2, 0, 1, -2, 1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, -2, -1, -1, -1, 1, 0, -2, 1, 2, 1, -1, -1, 0, 0, 0, 0, 1, -1, 2, 2, 0, 0, -2, 0, 0, -1, 0, 0, 0, -2, 0, -1, 1, 0, 0, 0, 0, -1, 0, 2, 0, -2, 0, 0, 0, 1, 0, 1, 3, 0, 1, -2, 0, 0, 1, 0, 1, 0, 0, -1, -2, 1, -1, 0, 0, 0, -1, 0, 1, 0, 2, 1, 1, 0, 1, -2, 0, 2, 0, 2, 0, -1, 0, 1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 3, 0, 0, 1, 3, 2, 1, 1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 0, 3, 0, 3, 1, 0, -1, -2, -1, 0, -1, 2, 3, 3, 4, 3, 0, 2, 0, 2, 0, 0, 0, 3, 2, 0, -1, 0, -1, 1, 3, 1, 2, 1, 0, 3, 1, 1, 2, 0, -1, 0, 2, 0, 3, 0, 1, 0, 2, 3, 0, 0, 0, 2, 3, 1, 1, 0, -2, 1, 1, 2, 2, 3, 1, 2, 1, 3, 1, 3, 2, 0, 0, 1, 2, 2, 2, 0, 0, 0, 0, 1, 2, 2, 0, 2, 2, 1, 0, 0, 2, 3, 1, 1, 0, -1, -1, 3, 2, 1, 0, 0, 2, 1, 2, 0, 1, 0, 0, 3, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 3, 0, 0, 1, -1, 2, 0, -1, 0, 2, 1, 1, 2, 0, 0, 1, 1, 0, 0, 1, 0, 1, -1, 0, -2, 0, 3, 3, 1, 1, 4, 5, 1, 1, -1, 2, 0, 0, 0, 2, 4, 3, 2, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 1, 5, 3, 1, 1, 2, 4, 3, 3, 1, 3, 0, 0, 0, 3, 2, 1, 1, 0, 1, 2, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 3, 4, 2, 3, 3, 3, 0, 0, 3, 1, -1, 0, 0, 0, 2, 1, 0, 0, 0, -1, 0, 1, 0, 2, 1, 0, 0, 0, 1, 0, 2, 2, 2, 2, 3, 0, 2, 2, 0, 0, -1, -2, -3, 0, 1, 2, 2, 0, 0, 0, 2, 0, 2, 2, 3, 1, 2, 1, 0, 1, 3, 3, 2, 1, 3, 4, 0, 0, 1, 2, 1, 0, 0, 1, 0, 0, 0, 3, 1, -1, 0, 0, -1, 0, 1, 2, 0, 2, -1, -1, 1, 1, 1, 1, 2, 2, 3, 0, 0, 0, 0, -1, 0, 1, 1, 2, 0, 2, 1, 0, 0, 0, 1, -1, 0, 1, 2, 0, 0, -2, 1, 0, 1, 2, 0, 3, 2, 0, -2, 1, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, -2, -1, 1, -1, 1, 1, 1, 0, 0, -1, -1, 0, 0, -2, 2, -1, 2, 1, 0, 2, 2, 0, 1, 0, 1, 0, 1, 0, 0, 2, -2, 0, -2, -1, 0, 0, 0, 0, -1, 0, -2, 0, 2, 0, -1, -1, 2, 1, 0, 1, 2, 1, 2, 3, 0, 1, 0, 0, 0, 2, -2, -1, -3, -2, -1, 0, -1, -1, 0, -1, 0, -1, 1, 1, 0, 2, 0, 2, 3, 0, 0, 1, 1, 1, 3, 0, 1, 0, -1, 0, -2, -5, -4, -3, -2, 0, 0, 1, 0, 1, -1, 0, -1, 1, 0, 0, -1, 0, 0, 1, 0, 1, 1, 2, 1, 2, 0, 1, 0, 0, -2, -2, 0, -1, 0, 0, 0, -3, -2, 0, -1, 0, -2, 0, 0, -1, -1, -2, -2, 0, 0, 1, -1, 0, -1, -1, -1, -1, 0, 1, -2, -5, -2, -1, 0, 0, 0, -1, -1, 0, -2, 0, -3, 0, 0, -1, 0, -2, 0, -1, -1, -1, 1, -2, -1, 0, 0, 2, 1, -1, 0, -2, 1, 1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, 1, 1, -1, 1, -1, 0, -1, 0, 0, 0, 1, 0, 1, 0, 1, -2, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 1, 1, 0, -1, 0, 2, -1, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, 0, -1, 1, -1, 0, -1, 1, 1, 2, 0, 1, 0, 2, 0, 1, 1, 1, 0, -1, 0, -2, 1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, -1, 0, 1, 0, 1, -1, -1, 0, -1, 0, 1, 2, 0, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, -1, 0, 0, 1, -1, -1, -2, -2, -1, 0, 2, 0, 1, 0, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, 0, 0, 1, 1, 0, -1, 0, 0, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -1, 1, 1, 2, 1, 0, 1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 0, -2, -1, -1, -1, 1, 0, -1, 0, 0, 1, 0, 0, -1, 1, -1, 1, 0, 0, -1, 0, 0, -1, 0, -1, 2, 1, 0, -2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 1, -1, 0, -1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 1, -1, 0, -1, -1, -1, 1, 0, -1, -1, -1, 2, -1, 0, 1, 0, 0, 1, -1, 1, 0, -1, 1, 1, 1, 0, 0, 1, 0, -1, 1, 0, 0, -1, 0, -1, -1, 0, 1, -1, -1, 0, 1, 1, 0, 0, 1, -1, 1, 0, 0, -1, 0, 1, -1, 0, 1, 0, -1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, 2, -1, 0, 1, 0, -1, -2, 0, 0, 0, -1, 1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -1, 1, 0, 2, 0, 0, 0, 1, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 0, 0, -1, -1, 1, 0, 0, 1, 0, -1, 1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 1, 0, 1, -1, 0, -1, -1, 0, -1, -2, -2, 1, 0, 0, 0, 0, 1, -2, -1, 1, 0, -1, -2, 0, 1, -1, 1, -1, -1, 0, 1, 0, -1, -2, 1, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, -1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 1, -1, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, 0, -2, 0, 1, 0, 1, -1, -1, -1, 1, -1, 2, 1, -1, -1, 1, 1, -1, 0, 1, 0, 0, 1, 0, -1, -1, 0, -1, -1, -1, 0, 1, 0, -1, 1, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 1, -1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 0, 1, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 1, -1, 0, 1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, -2, 0, 0, 0, -1, 1, 0, 0, 0, 1, -1, 0, 1, -1, 0, 1, -1, 1, -1, 0, -1, -1, 1, -1, -1, 1, 1, 0, -1, 1, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, -1, -2, 2, 1, 0, 0, 1, 1, 0, 0, 0, 0, -2, 0, 1, 0, 0, -1, 0, 0, 0, 0, 2, -1, 0, -1, 1, 1, 1, 1, -1, 0, -1, -1, 1, -1, 0, 1, 1, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 1, 1, -1, 0, -2, 1, -1, 0, 1, 0, -1, 0, 0, -1, 0, -1, 1, -1, -1, 1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, -1, 0, 0, 0, -1, 0, 1, 1, -1, -1, 0, -1, -1, -1, -1, -1, 0, 1, 0, 1, 1, 0, -1, 0, 0, -1, 1, 0, -1, -1, 1, 0, -1, -1, 0, -1, -1, 1, 0, 0, 0, 1, 0, -1, -1, 0, 1, -1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 2, 0, 0, 1, 0, 1, 0, 0, -1, 0, -1, -1, 0, 0, 1, -1, 1, -1, 0, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, 1, -2, 0, 1, 0, -1, -1, 0, 1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0,
    -- filter=0 channel=6
    -2, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 1, 0, 2, 0, 1, 3, 3, 1, 1, 0, 0, 0, 0, 0, 3, 0, 0, 1, 2, 0, 0, 2, 1, 1, 0, 1, 1, 2, 0, 2, 1, 3, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, 0, -1, 2, 0, 0, 0, 2, 0, 2, 1, 2, 1, 0, 2, 2, 2, 0, 1, -1, -1, 0, 0, 0, 1, 2, 2, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, 2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 1, 0, 0, -1, -2, 1, -1, -1, 2, 0, 0, 0, -1, 2, 0, -1, 0, 0, -2, 0, -2, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, 1, 2, 0, -2, 0, 0, 1, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 1, -1, 1, 0, 0, 0, 0, 0, -1, 0, 1, -1, -1, 0, 1, 0, 2, 0, 0, 2, 0, 0, 1, -2, -2, 0, 0, -2, 0, 0, 0, 0, -1, -1, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 2, 0, 1, 1, -1, 0, -2, 0, 1, 0, 0, -3, -1, 0, -2, -2, -1, -1, -1, 1, 1, 0, 0, 0, 1, -2, -2, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -4, -2, -1, -1, -3, 0, -2, 0, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 1, -1, 0, 2, 1, 0, -2, -2, -2, -2, -1, -4, -1, -4, -3, -4, -2, -2, -2, -1, 1, 0, 0, 1, 0, -1, -1, 0, 1, 2, 0, 2, 1, 1, 0, -1, -1, -3, -3, -3, -1, -2, -5, -3, -4, -5, -3, -3, -2, 0, 1, 0, -1, 0, 0, 0, 0, 0, -1, 3, 0, 0, 2, 0, -1, -1, -2, -2, -3, -4, -3, -2, -2, -5, -5, -6, -3, -1, -4, -1, 0, -1, 2, 0, 1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, -2, -1, -4, -2, -3, -3, -3, -5, -4, -2, -4, -4, -1, 0, 0, -1, 1, 0, 0, -1, -1, 0, 0, 1, 2, 0, -1, 0, 0, -3, -2, -2, -2, -3, -5, -4, -2, -4, -3, -5, -3, -2, 0, -3, -1, 0, 1, 1, 0, -2, 0, 1, 1, 3, -1, 2, -1, 0, 0, -3, -2, -3, -4, -3, -2, -5, -5, -3, -3, -3, -3, -3, -1, 0, 1, 0, 1, 0, -1, -1, 0, 2, 2, 0, 0, 1, -1, -1, 0, -1, -2, -2, -2, -4, -3, -3, -4, -2, -4, -2, -4, -3, -1, 0, 1, 0, 1, 1, 0, 1, -1, 0, 0, 2, 0, 0, 1, -2, 0, 0, -2, -3, -2, -1, -1, -2, -2, -3, -4, -2, -2, -1, -2, 0, 2, 1, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, -3, 0, 0, -2, -1, -2, -2, -5, -2, -3, -3, -4, 0, 1, 0, 0, 1, 0, -1, -2, 0, -1, 1, 0, 2, 3, 0, 2, 1, -2, -1, 0, 0, -4, -2, -2, 0, -1, -3, 0, -1, -3, 1, -1, 0, 1, 0, 2, -1, 0, -1, 0, 0, 1, 2, 1, 0, 0, 0, 0, 0, -1, 0, -3, 0, -3, -1, -3, -2, -3, 0, -1, 0, 0, 1, 0, 2, 2, 1, 0, -1, -1, 0, 0, 0, 0, -1, 2, 0, -1, -2, -2, 0, -1, -3, 0, -2, -2, -3, -2, 0, 2, 2, 0, 1, 1, 0, 2, 1, 0, 0, 2, 1, 0, 1, 3, 0, 2, 0, 0, 0, 0, 0, -1, -2, -2, -2, 0, 1, 0, -1, 0, 3, 2, 1, 0, 0, 0, 1, -1, 0, 0, 2, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, -1, 0, -1, 1, 2, 3, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, 0, 1, 1, -1, 1, -1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, -1, -1, -2, -2, 1, 1, 0, -1, 0, -1, 2, 1, 1, 2, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 3, 1, 0, 2, 0, -1, 1, 1, 1, 1, 0, 1, -1, -1, 0, 1, 1, 2, 1, 0, -1, 2, 1, 2, 1, 0, 1, 0, 0, 2, 0, 0, 2, -1, 1, -1, -1, 0, 0, 0, 1, 1, 1, 1, -1, 1, 1, 1, 1, 2, 2, 0, 0, 0, 0, -1, 0, 1, 0, 1, 3, 0, 2, 0, 0, 2, 2, 2, 2, 1, 2, 1, 1, 0, 1, 2, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, -1, 1, 3, 0, 1, 3, 2, 0, 2, 1, 1, 0, 2, 2, 0, 2, -1, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, -1, 0, 0, 0, 1, 0, 1, 2, 2, 2, -1, 0, 0, 0, 0, 2, 1, 2, 1, 1, 0, -1, -1, 1, -2, -3, -1, -1, 1, 1, 1, 0, 0, 0, 4, 6, 2, 5, 4, 7, 5, 4, 5, 4, 1, 0, 1, 0, 3, 3, 1, 3, 0, 2, -1, -3, -1, -2, -1, -1, 0, 1, -1, 1, 2, 1, 0, 3, 1, 4, 2, 2, 2, 1, 0, 0, 0, 2, 0, 1, 0, 1, 0, 0, -2, -1, -1, -2, 0, 1, -1, 0, -1, -2, 0, 1, 0, 0, 1, 0, 2, 0, 0, 1, 0, 1, 2, 2, 1, 1, 2, 2, 1, 2, -4, -2, 0, -1, 1, 1, -1, 1, 0, 1, -1, 0, -1, -1, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, -2, -1, 1, 0, 1, 0, -7, -4, 0, 0, -1, 0, 0, 0, 2, 1, 0, 0, 0, -2, 1, 0, -1, -2, -1, 0, 0, 1, -1, -3, 0, -1, -1, 0, 1, -1, -4, -2, -1, 0, -1, 0, 0, -1, 0, 0, 2, 0, -2, -1, -1, 0, 1, -2, -1, -1, -1, 1, -1, -1, -1, 0, -1, 0, 0, 0, -4, -4, 0, 0, -1, -1, 0, 1, 0, 2, 1, 1, 0, -2, 0, -1, 1, 1, 0, 0, 0, 1, 1, 0, -1, -2, 0, -1, 0, -2, -4, -1, -3, 0, -3, 0, 1, 0, 0, -1, -1, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, -2, 0, -2, -2, 0, -1, 0, -3, -5, -3, -1, -2, 0, 0, 0, 0, 0, 1, 0, -1, 0, 2, 2, 2, 1, 0, 0, 0, -2, 0, 1, 0, -1, -1, -2, -3, -3, -2, -4, -1, -1, -2, -3, 0, 0, 1, 0, -1, 0, 1, 2, 3, 2, 3, 2, 1, 0, 0, 0, -2, 0, 0, -1, -2, -1, -1, -2, 0, -2, 0, -1, 0, -1, -1, -2, -3, -1, -3, -3, -1, 3, 5, 4, 4, 2, 4, 1, -1, 0, -3, -4, -1, -1, 0, -1, -1, 0, -3, -1, 0, 0, -2, -4, -2, 0, -4, -1, -2, 0, -1, 2, 5, 5, 4, 6, 3, 1, 1, -1, -1, -2, -4, 0, -3, -1, -1, -3, -3, -3, -1, 0, -1, -4, -4, 0, 0, -2, -1, -2, 0, 1, 3, 5, 7, 6, 4, 4, 2, -1, -4, -4, -3, -2, -2, -4, -1, -1, -2, -2, -1, -2, 0, -4, -1, -5, -2, -3, -2, -1, 1, 3, 3, 8, 6, 6, 7, 2, 1, 2, -1, -2, -4, -4, -5, -3, -1, -1, -2, -2, 0, 0, -3, -1, -5, -4, -5, -5, -2, -2, 1, 0, 5, 5, 7, 6, 5, 5, 2, 0, -3, -3, -3, -3, -2, -2, -3, -5, -2, -5, 0, -1, -2, -1, -3, -2, -6, -5, -2, -3, 0, 3, 3, 4, 8, 6, 3, 2, 5, 1, 0, -1, -4, -4, -3, -5, -1, -4, -3, -5, -1, 0, 1, -3, -1, -2, -7, -3, -1, -2, -1, 3, 3, 4, 5, 7, 5, 2, 4, 2, 0, -2, -3, -3, -6, -4, -1, -3, -3, -3, -1, -2, -2, -4, -4, -5, -6, -3, -2, -2, -1, 0, 2, 2, 6, 6, 8, 4, 4, 1, -1, -5, -3, -6, -3, -3, -1, -3, -2, 0, 0, -3, 0, -2, -5, -4, -6, -3, -3, 0, -2, 1, 4, 3, 7, 6, 8, 5, 2, 0, -2, -3, -4, -6, -5, -6, -3, -3, 0, 0, -3, -2, -3, -1, -3, -5, -1, -4, 0, -1, 0, 2, 5, 5, 4, 5, 6, 3, 0, 1, -5, -5, -5, -6, -4, -3, 0, -2, -1, -3, 0, -2, -3, -3, -1, -1, -3, -1, -1, -1, 0, 2, 2, 4, 3, 3, 5, 3, 0, 0, -3, -4, -3, -2, -1, -3, -3, 0, 0, -5, -3, -2, -3, 0, -1, -1, -1, -2, 1, -1, 1, 0, 2, 4, 4, 1, 2, 0, 1, -1, 0, -1, -4, -3, -2, -2, -3, -3, -3, -5, -1, -1, -2, 0, -1, 0, -2, -1, -1, -1, -1, 1, 1, 3, 0, 2, 0, -3, 0, -3, -3, -1, -1, -2, -4, -2, -2, -1, 0, -6, -4, 0, -2, -1, 0, 0, 0, 0, -2, 0, 2, 1, 0, 2, 3, 2, 1, -1, 0, 1, 0, -3, 0, 0, -3, -2, -1, 0, -1, -2, -1, -3, 0, -2, 1, 2, 0, 2, -1, 0, 1, 1, 0, -1, -2, 0, -2, 0, -2, 0, 0, 0, -1, 0, -1, -1, 0, 2, 0, -5, -3, 1, 0, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, 1, 0, 0, -1, 1, 2, 1, 0, -5, -3, 0, -1, 0, -1, 0, 0, 0, 0, 0, 1, 2, 0, -2, 0, -2, 0, -1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 0, -5, -2, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, 0, 2, 0, 0, -2, 0, 0, 0, -1, 1, -2, 0, -1, 0, 0, 2, 1, 3, -2, -2, -2, -1, 0, 0, 1, 0, 0, 0, 3, 2, 3, 0, 2, -3, -1, 0, -2, 0, 0, 0, -1, 2, 0, 1, 2, 1, 2, 1, -3, -2, -3, 0, 0, 0, 1, 2, 0, 2, 3, 3, 2, 3, 1, 1, 1, 0, 1, -1, -1, 0, 1, 2, 1, 1, 0, 0, 1, 1, -5, -3, -2, 0, 0, 0, 1, 0, -1, 1, 0, 3, 2, 4, 1, 2, 2, 4, 0, 3, 2, 3, 1, -1, 2, 0, 1, 0, 0, 1, -5, -4, 0, -2, 0, -1, 1, 1, -1, 0, 0, 2, 2, 1, 3, 0, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, -5, -2, -2, 0, -1, 0, 0, -2, -1, -1, 0, -1, 0, 1, 1, 1, 2, -1, -1, -1, -2, -2, 0, 1, 0, -1, -1, 0, 0, 0, -3, -3, -3, 0, -1, -1, 0, 1, -3, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, -1, 0, -1, 1, 1, 1, 0, -1, -1, -2, -1, 0, -1, 0, -2, -1, 0, -1, -1, -2, -2, -1, -2, -2, -1, -1, 0, -2, -2, -2, -1, -2, -1, 0, 0, -2, -2, 0, 0, -3, -3, 0, -1, 0, -3, 0, -2, 0, 0, 0, 0, 0, -2, -2, -1, -2, -3, -1, 0, -2, 0, -1, 0, 0, 0, 0, -1, 1, 0, -5, -1, -2, -1, 0, 0, -2, -2, -3, -3, -1, -3, -3, 0, -4, -4, -3, -1, 0, -2, -2, -1, -2, -2, 0, 0, 0, 0, 0, -2, -2, -3, -1, -2, -1, -2, -1, 0, -4, -3, -1, -3, 0, -1, -4, -1, -1, 0, -3, -3, -2, -1, -2, -2, -2, -1, 0, -1, 0, -2, -5, -2, -3, -4, -1, -3, 0, -2, -2, -4, -4, -4, -3, -3, -3, -4, -3, 0, -2, 0, -3, -2, -1, -2, -1, -2, 0, 0, -1, 0, -1, -1, -2, -2, -2, 0, 0, -4, -4, -2, -4, -4, -4, -4, -2, -2, -2, 0, -4, -1, -1, -1, -1, -3, -3, 0, -2, -4, 0, 0, -3, -1, -2, -3, -3, -4, -2, -2, -4, -3, -5, -2, -1, -1, -2, 0, -2, -1, -3, -2, -1, -3, -2, 0, -3, -2, 0, 0, 0, -2, -1, -3, 0, -2, -3, 0, -3, -3, -4, -5, -3, -6, -5, -4, -2, -1, -2, -3, -4, 0, -3, -2, 0, -3, 0, -2, 0, -3, 0, 1, -3, -1, 0, -3, -1, -4, -3, -1, -2, -5, -5, -3, -1, -4, -2, -2, 0, -3, 0, -2, -1, -2, -2, -1, 0, -2, -1, 0, 0, -1, -2, -2, -1, -2, 0, -1, -4, -4, -2, -5, -4, -3, -3, -1, -3, 0, 0, -2, -3, -2, 0, -2, -3, 0, 0, -3, -2, -1, -1, -2, -2, -2, 0, 0, 0, -3, -3, -4, -6, -3, -4, -5, -5, -2, -2, 0, -1, 0, -3, -1, -3, -2, -4, -1, 0, -1, -3, 0, 0, -2, -1, -2, -1, 0, -2, -2, -2, -6, -6, -4, -5, -2, -2, -1, -1, -3, 0, -3, 0, 0, -2, -1, -3, -4, -4, -4, -1, -3, 0, 1, -1, 0, 0, 0, -1, -3, -4, -6, -6, -3, -3, -5, -3, -3, 0, -2, -2, -2, -1, -3, -2, -1, -3, -3, -4, -3, -2, -3, -2, -2, -1, 0, -2, 0, 0, -2, -2, -3, -2, -3, -2, -1, -3, -4, -2, 0, -3, 0, 0, 0, -2, -2, -3, -2, -3, -2, -2, -2, -2, 0, -2, 0, -2, -2, -3, -4, -4, -3, -5, -3, -3, -2, -5, -5, -2, -2, -3, -2, 0, 0, 0, -3, -2, -4, -4, -1, -4, -1, 0, 0, -2, 0, -2, 0, -4, -3, -4, -2, -5, -4, -5, -5, -1, -4, -3, -1, -2, 0, 0, -3, -2, -1, -1, -2, -3, -4, -3, -1, -1, 0, -2, -2, -1, 0, -2, -3, -2, -5, -5, -3, -2, -4, -2, -2, -1, -2, -2, 1, 0, -3, -4, -2, 0, -4, -3, -2, 0, -2, -1, -1, -4, -1, 0, 0, -1, -2, -2, -4, -4, -3, -3, -4, -1, -4, -2, 0, 0, -2, 0, -3, -3, 0, 0, -2, 0, 0, -2, 0, -1, -2, -1, -3, 0, 0, -2, 0, -3, -1, -5, -2, -1, -2, -1, -3, -2, -2, -1, -1, -1, -3, -1, 0, -1, -4, -1, -1, -2, -2, -2, -2, -1, -3, 0, 0, -2, -1, 0, -1, -3, -2, -2, -3, -1, -2, -1, 0, -1, -3, -2, -1, 0, 0, -1, 0, -2, -3, 0, 0, 0, 1, 0, -1, -1, 0, -2, -1, -2, -2, 0, -2, -2, 0, 0, 0, -2, -2, 0, -2, -2, 0, -2, -3, 0, 0, 0, 0, -1, -1, 0, 1, -1, -3, -2, 0, -1, -1, -2, 1, -2, -1, 0, 0, -2, -3, -3, -3, 0, 0, -2, 0, -1, 0, -1, -2, 0, 0, 0, -1, 0, 2, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, 0, -2, 0, -2, 0, -2, -1, -3, -2, -2, 0, 0, -1, 0, -1, 0, 1, -1, 2, 2, -1, -3, -1, 0, -1, 0, -2, 0, 0, 1, -2, 0, 0, -1, -1, -2, -3, -2, -1, -2, 0, -1, -1, 0, 0, -2, 2, 1, 1, 0, -1, -1, 0, 0, -2, 1, 0, 0, -1, 1, 0, 2, 0, 0, 0, 0, -2, 0, 1, -1, 0, 1, 1, 0, 0, -1, -1, 0, 0, 2, -2, -2, -2, -2, 0, -1, 0, 0, 1, -1, 1, 1, 0, 0, 2, 1, 0, -2, -2, 1, -1, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 1, -1, 1, 0, -1, 1, 0, 2, 0, 0, -1, 1, 0, -1, 0, -1, 0, 0, 1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 1, -1, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 1, 0, -1, 2, 1, 1, -1, 0, 1, 0, -1, -1, -1, 1, 0, 1, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, -1, 0, -2, 1, 0, 1, 0, -1, -2, 2, -1, 0, 0, 0, 1, 1, 0, -1, 1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 1, -1, -1, 1, -1, 0, 1, 0, -1, 0, -1, 0, 0, 2, 1, 0, 1, 1, 0, 0, 0, 0, -2, -1, -1, 0, 0, -1, -2, -1, 1, -1, 0, 2, 1, 1, 0, 0, 0, 0, 1, -2, 0, -1, 0, 0, 0, 1, -1, 0, 1, 1, -1, 0, 1, 0, 2, 0, 1, 0, -1, 1, 1, 0, -1, -1, -1, 0, 0, 0, 1, -2, 2, 0, 0, 0, -1, -1, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, 1, -1, 1, 0, 0, 0, -1, -1, 0, -1, 1, 0, 0, -2, 0, -1, 0, 1, 1, 0, 0, -1, 0, 2, 1, 0, 0, -1, -1, 0, 0, 0, 1, -1, 2, 0, 1, 0, 0, 0, 1, 0, 1, -2, 1, 0, -1, 1, -1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 0, 1, 0, 1, 1, -1, 1, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, 0, 1, 0, 1, -1, 1, 0, 1, 0, 0, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, -1, 1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, -1, 0, 0, -1, 0, 1, 0, -1, 0, 0, -2, 0, 1, 1, -1, 0, 0, 0, 0, -1, -2, 1, 0, -1, -1, 0, 0, -1, -1, 0, 1, 1, 0, -1, -2, 1, 0, -1, 0, -1, -1, 0, -1, -2, 1, 1, 0, 0, 0, 0, 1, -2, 1, 0, -1, 1, 0, 0, -1, -1, 1, 1, 0, -1, 0, -1, 0, 2, 0, -1, -1, 1, 0, 0, -1, 1, -2, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 0, 1, 1, 1, -1, 1, 1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, 0, 1, 0, 2, 1, 1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, -2, -1, -1, 0, 1, 0, 2, -1, -1, -1, -1, -2, -1, 0, 0, 0, 1, -1, 0, 0, 1, 0, -1, -2, 1, 1, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, -1, 1, 1, 1, 0, 1, 1, 0, 1, -1, 2, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 1, -1, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 1, 0, 1, 0, -1, -1, 0, -1, 1, 0, -1, 0, 1, 1, 2, 0, -1, 1, 1, 0, 2, 0, 1, -1, 1, -1, 1, 0, -2, 0, 1, 1, 1, -2, 0, 0, 0, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 2, -1, 0, 0, -1, 0, -1, 2, -1, 0, 1, 0, 0, 0, -1, 0, 1, -1, 0, 1, -1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 1, 1, -1, 1, 1, -2, 0, 0, 0, 2, 1, -1, 0, 0, 0, 0, 0, 1, -2, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, 1, -1, -1, 1, -1, 0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 2, 0, 1, -2, 0, 1, 0, -1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, 2, 0, 1, 1, 0, 0, 0, 1, -1, -1, 1, 0, 0, 0, 1, -1, 0, 1, 2, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 0, 2, 0, -2, 1, 1, -1, 0, 0, -1, -1, 1, 0, 1, 0, 0, -2, -1, 2, 1, 0, 2, 2, 1, 1, 2, 0, 1, -1, 0, 0, 1, 1, 0, 0, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, 0, 0, -1, 1, 0, 0, 1, 1, 3, 5, 1, 3, 1, 1, 3, 4, 3, 0, 2, 3, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 0, -1, 2, 2, 2, 0, 0, 0, 3, 1, 3, 1, 1, 3, 0, 0, 0, 0, 0, 1, -2, 0, 1, 0, 1, -1, 0, -2, 0, 0, 0, 1, 2, 0, 0, 2, 2, 0, 3, 1, 2, 2, 3, 0, 0, -1, 1, 0, -2, 0, 0, 0, -3, -2, -1, -3, -1, -2, -2, 1, 2, -1, 1, 2, 4, 0, 0, 3, 1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, -1, -1, -3, 0, -3, -3, -3, 0, -1, 0, 0, 0, -1, -1, 2, 0, 3, 0, 3, 3, 0, 1, 1, 2, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, -1, 0, 1, 1, -1, 1, 0, 2, 2, 0, 3, 3, 1, 1, 0, 2, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -2, -1, 0, -2, -1, -2, 0, -1, 1, 2, 3, 1, 2, 1, 2, 3, 2, 0, 0, 1, 0, 0, 0, 2, 0, -1, -2, 0, -1, -1, -2, -2, -3, -2, 0, 0, 0, -1, 2, 0, -1, 1, 2, 1, 3, 3, 1, -1, 2, 0, 1, 0, 1, 3, 1, 0, 1, 0, -1, -1, 0, 0, 0, -2, -1, -3, -2, 0, 0, 0, 1, 2, 0, 0, 0, 0, 1, 0, 2, -1, 0, -2, -1, 0, 1, 0, 2, 0, 0, 0, 1, 1, 0, -1, 0, -4, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 1, 1, 2, 0, -2, -1, 0, 0, 2, 1, 0, 0, 2, 0, 2, 1, 0, 1, 0, 0, -3, 0, 0, -2, 2, 3, 1, 2, 0, 0, 1, 1, 0, 1, 0, 0, 2, 0, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, -1, -2, 0, 2, 3, 1, 2, 2, 2, -1, 1, 2, 0, 0, -1, 1, 0, 0, 3, 3, 1, 4, 4, 3, 1, 1, 0, 0, 0, 0, -2, 0, 1, 0, 3, 2, -1, 2, 2, -1, 0, 1, 0, 0, -1, 0, 0, 3, 3, 4, 2, 2, 4, 2, 4, 5, 5, 2, 2, 3, 0, -3, 0, -1, 0, 0, -1, 1, 1, 0, 2, 0, 0, -2, 0, -3, 1, 1, 3, 0, 3, 3, 5, 1, 3, 5, 5, 2, 6, 4, 2, 0, -1, 0, -1, 0, 3, 0, -1, 0, 1, -1, 0, -2, -1, 1, 2, 0, 0, 1, 3, 2, 1, 4, 5, 4, 5, 3, 2, 3, 0, 0, 1, 1, 1, -1, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 2, 3, 4, 5, 5, 3, 2, 4, 5, 2, 1, 4, 3, 0, 0, 2, 0, 0, 1, 2, 2, 0, 0, -2, 0, 0, -1, 0, 0, 1, 0, 2, 3, 5, 5, 5, 4, 2, 3, 3, 1, 3, 2, 3, 0, 0, 0, 0, 0, 1, 2, 1, 0, -1, -3, 0, 0, 0, -2, -1, 2, 2, 4, 1, 5, 5, 2, 4, 3, 6, 4, 5, 3, 2, 1, -1, -1, 0, 3, 0, 0, 2, 0, 2, -1, -3, -1, 1, -1, 1, 3, 1, 1, 1, 3, 2, 3, 2, 1, 3, 5, 2, 4, 2, -2, -1, 0, 0, 0, -1, 3, 3, 0, 1, -1, -3, -1, 0, 1, 1, 2, 1, 1, 3, 0, 5, 6, 4, 3, 3, 5, 3, 0, -1, -1, 0, 0, 0, -1, 1, 1, 2, 0, 0, 0, 0, -1, 0, 1, 0, 0, 2, 4, 0, 0, 0, 4, 2, 3, 2, 0, -1, -2, 0, -3, -1, 2, 0, 3, 0, 2, 1, 0, 0, 1, 0, 0, 0, 2, 1, 1, 3, 3, 1, 1, 1, 0, 0, 2, -2, -4, -3, -2, -3, 0, -1, 0, 1, 2, 0, 3, -1, 1, -1, -1, 0, -2, -1, 0, 0, 0, 1, 2, 0, 0, 1, 2, 0, 0, -1, -4, -2, -2, -1, 1, 0, 0, 0, 3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, -2, -2, -3, -2, -5, -2, 1, 1, -2, -1, 0, 2, 0, 2, 1, 2, 2, 2, 0, 1, -2, 0, 0, 0, -1, 2, 2, 0, -2, -1, -3, -5, -5, -5, -4, 0, -1, -1, 0, 0, 1, 0, 3, 3, 0, 0, 3, 0, 1, 2, 1, 0, 0, 2, 1, 0, -1, 0, -1, -2, -2, -3, -4, -5, -2, -2, 0, 2, 2, 3, 0, 1, 0, 1, 4, 4, 2, 3, 1, 1, 0, 0, 1, 0, 1, -1, 0, 0, 0, -2, -3, -2, -5, -1, -3, 0, 2, 3, 2, 2, 1, 0, 2, 5, 5, 2, 2, 0, 0, 3, 0, 1, -1, -1, 0, 1, 0, 0, -1, 0, -1, -4, -4, -2, 0, 0, -1, 1, 2, 3, 3, 0, 1, 1, 5, 1, 4, 3, 3, 3, 0, 0, -1, 1, 0, 0, 0, 0, 1, -1, -1, -3, -3, -3, 0, -2, -1, 0, -1, 2, 2, 3, 3, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 1, -2, -1, -2, -1, -3, -2, 0, -2, -1, -2, 0, 0, -1, 2, 1, 1, 1, 0, 3, 1, 2, -1, 0, 0, 0, 1, 1, 0, 0, 0, 2, 0, 1, 1, 0, 0, 1, 0, 3, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 0, -1, 0, 2, -1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 0, 1, -1, 2, 1, 0, 2, 2, 1, 2, 0, 3, 0, 2, -1, 0, 0, -1, 0, 1, 2, 0, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 2, -1, 2, 2, 0, 1, 1, 0, 2, 0, 1, -1, 1, 0, 2, 1, -1, 0, 0, 2, 0, 1, 0, 3, 0, 0, 0, 0, 1, -1, -1, 1, 1, 0, 0, -1, 1, 3, 2, 2, -1, 0, 0, 1, 0, 0, 1, 1, 0, 2, 2, 0, 0, 1, 1, 1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, 2, 0, 0, 1, 0, 1, -1, 1, 0, 2, 3, 2, 1, 0, 0, 2, 2, 2, 0, 1, 0, -1, 1, 1, 0, 0, 0, 0, 1, 1, 0, -1, 0, 2, 0, 2, 2, 2, 1, 2, 1, 2, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 2, -1, -1, 0, 1, -1, -1, 0, 0, 0, -1, 0, -1, 2, -1, -1, 0, 0, 1, 0, 2, 0, 2, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 1, 1, 1, 2, 1, 2, 1, 1, 0, -1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 0, 3, 2, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 1, 0, 2, 2, 0, 0, 1, 0, 2, 0, 0, 1, 2, 1, -1, 0, 2, 0, -1, 0, 0, 0, 1, 0, -1, -1, 1, 2, 2, 1, 1, 0, 1, 0, 0, 2, -1, -1, -1, -1, -1, 0, 1, -1, 2, 0, -1, 1, 1, -2, 1, -2, 1, 0, -1, 0, 2, 0, 1, 0, 1, 3, 2, 2, 0, 1, 0, -1, 1, -1, -1, 0, 1, 1, 0, 0, -2, -2, 0, 1, 0, -2, -2, 0, -1, -1, 0, 0, 0, 1, 2, 1, 0, -1, 3, -1, 2, -1, 1, 2, 0, -2, 0, 1, 0, 1, 1, -2, -2, 0, 0, -1, -1, 0, 0, -2, 2, 0, 1, 0, 0, 3, 1, 2, 1, 2, -2, 2, 0, 1, 1, -2, 0, 1, -2, -1, 0, 0, -2, -3, 0, 1, 1, -2, 2, -1, 0, 0, 0, 0, 1, 2, 1, 2, 1, 0, 1, 1, 1, 2, 0, 0, 0, 0, 0, -2, 0, -1, -2, 0, -1, 0, 0, -1, -1, -1, 2, 2, 3, 1, 1, 0, 1, 0, 0, 1, 0, -2, 2, -1, 2, 2, 1, -1, 0, 0, 0, -2, 0, 0, 0, 0, -2, 1, 0, 2, -1, 0, 1, 0, 1, 3, 3, 0, 3, 2, 0, 1, 0, 2, -1, 0, 1, 0, -2, 1, -1, 0, -1, 1, -2, 0, 0, 0, 2, 2, 0, 0, 0, 0, 2, 1, 0, 2, 1, 2, 0, 0, 1, 0, -1, 1, -2, 0, -1, -2, 0, -1, 0, 0, -1, -1, 0, 0, 2, 0, 2, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 3, 0, 1, 1, 1, 0, 0, 0, 3, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, -1, 0, 0, 0, 2, 0, 0, 0, 0, 2, 0, 0, 2, 3, 0, 2, 0, -1, -1, 0, 1, 2, 1, 0, 0, 1, 0, 0, 1, 1, 2, 2, 1, 0, 0, 2, 2, 0, 0, 1, 2, 0, 2, 0, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 1, 2, 1, 0, 0, 2, 0, 1, 2, 1, 0, 1, 2, 0, 0, 0, 3, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 2, 2, 0, 0, 1, 1, 0, 0, 0, 0, 1, 1, 0, 1, 3, 2, 2, 0, 0, 1, 1, -1, 0, -1, 0, 0, 0, -1, 1, 0, 0, 3, 0, 1, 0, 2, 0, 0, 2, 0, 0, 2, 0, 3, 0, 0, 0, 3, 1, 1, -1, 0, 0, 0, -1, 1, 1, 2, 0, 3, 1, 1, 0, 0, 1, 2, 2, 2, -1, 0, 2, 0, 1, 1, 0, 1, 0, 1, 3, 1, 0, 2, 2, -1, 1, 0, 0, 1, 0, 1, 2, 0, 1, 1, 2, 0, 0, 2, 0, 0, 0, 2, 2, 0, 3, 2, 0, 0, 3, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 2, 2, 0, 2, 2, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 2, 3, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 2, 1, 0, 0, 0, 1, 2, 0, 0, 2, 0, 0, 2, 1, 2, 0, 0, 0, -1, 1, 1, 2, 0, -1, 0, 1, 0, 1, 0, 1, 1, 2, 2, -1, 0, -1, 0, 1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 2, 1, 0, 0, -1, 2, 1, 0, -1, 0, 0, -1, 1, 1, 1, 0, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, -2, 1, -1, -2, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 2, -1, -1, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, -2, 0, 0, 0, 0, 0, 1, 1, 1, -1, 2, -1, 0, 2, -1, 2, 0, -1, 0, 0, -1, -1, 0, 1, -2, 0, -1, 0, -2, -2, 0, 0, -1, 0, -1, 1, 1, -1, 1, 0, 1, -1, 1, -1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 1, -1, 0, 1, 1, 2, -1, 0, 0, 0, -1, 1, 1, 0, 0, 1, 1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, -1, 1, 0, 0, 0, -1, 0, 0, -1, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 1, -2, 0, 0, 0, -2, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 2, 0, -1, 0, 1, 0, 0, -1, 0, 0, 0, -2, -1, 0, 0, -1, 1, -3, 0, 0, 1, -1, 0, -1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 0, 1, 1, -2, -1, 2, 0, 1, -1, 0, 1, 0, -1, 0, 0, -2, 0, -1, 1, 0, -1, 0, 2, -1, 2, 0, -1, 0, 0, 1, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -3, -2, -3, -1, 0, 1, 0, 1, 1, -1, -1, -1, 0, 0, 2, 0, 1, 2, 2, 1, -2, 0, -2, 1, 0, 0, 0, -2, -1, 0, -2, -2, -3, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 0, -1, -2, -1, 0, 0, 0, -1, 0, 1, 1, 0, 2, -1, 0, 0, 0, 0, 0, 1, 2, 1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, 0, 0, -1, 1, 0, 1, 0, -1, 0, 0, 2, 0, 0, -1, 1, 1, 2, 0, 0, 0, -1, -1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 2, 0, 0, 2, -1, 0, -1, 1, 0, 0, 0, -1, -1, 0, 1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 2, 0, -1, 2, -1, 0, 1, 2, 2, 2, -1, 0, -1, 2, -1, -1, -1, 1, 0, -2, -1, 0, -2, -1, 1, -1, 2, 2, 2, 2, 1, 0, 0, 1, 2, 2, 0, -1, 0, 0, 2, 2, 2, 0, -1, 0, 1, 0, 0, -1, -2, 0, -1, 0, 1, 2, 1, 1, 1, 1, 2, 0, 2, -1, 1, -1, -1, 0, 2, -1, -1, 0, -1, 0, 0, 0, 1, -1, 0, 0, -1, 0, 1, -1, 0, 2, 0, 1, 1, 2, 2, 0, 1, -1, 0, 0, 1, 1, 1, 1, 1, 0, 0, 0, 1, 1, -1, 0, 0, -1, 0, 1, -1, 0, 1, 0, 2, 0, 2, -1, 1, -1, 1, 2, 1, 0, -1, 0, 0, -1, 0, -1, 1, 2, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, 0, 2, 0, -1, 0, 0, -1, 0, 2, 1, 2, 1, 1, 1, 1, -1, -1, 0, 0, -1, -1, 0, 2, 0, 0, 2, 1, 0, -1, 0, 2, 1, -1, -1, 0, 2, -2, -1, 0, -1, 1, 1, 1, 1, 2, 0, 0, 1, 1, 1, 0, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, 2, -1, 0, -1, -1, 1, 1, 0, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, 1, 0, 0, -1, -1, 0, 0, 2, 1, 1, -1, 0, 0, -1, -1, 0, 2, 1, 0, 2, 0, -2, 0, 1, 1, 2, 1, 2, -1, 0, 2, 1, 1, 2, 1, 0, 0, 0, 1, 0, -1, 0, -1, -1, 1, 1, -1, -1, 1, -1, -2, 0, 0, 0, 1, -1, 2, 1, 0, -1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, -1, 1, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, 2, -1, 1, 2, -1, 1, -1, 2, 0, 0, 1, 0, 2, 0, 1, 0, 0, -2, 0, -1, 0, 1, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 2, -1, -1, 0, 0, 1, 0, -1, -1, 1, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 1, 0, 1, 0, 0, 2, 1, 1, 0, 0, 2, 2, 0, 1, 1, -1, 2, 0, -1, -1, -1, 1, -1, -1, -2, 0, 0, -1, 0, 0, 1, 0, 0, 0, 2, 1, 2, -1, 1, 2, -1, 0, 1, -1, 0, -1, 0, 0, -2, 0, -2, 1, 0, 0, 0, -1, -3, 0, -1, -1, 0, -2, -2, 0, -1, -1, 1, 0, 1, -1, 2, 0, -1, 0, 1, 2, 0, 0, -1, -2, 0, -3, -1, 0, -4, 0, -1, -2, -3, -1, -1, -2, -1, -3, -2, -1, -1, -3, 0, -2, -1, -1, -2, 0, 0, 2, 0, 0, -1, -1, -2, -3, -3, -2, -1, -4, -1, -3, -3, -2, 0, 0, -3, 0, -3, 0, -2, -2, 0, 0, -1, -2, 0, 1, 2, 0, 1, 0, 0, 0, -1, 0, -2, -1, -1, -1, 0, -3, -2, 0, -1, -3, 1, 0, -1, -1, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, 0, -1, 0, -1, -1, -2, -2, -1, -1, 0, 0, -1, 0, -1, 1, 1, 1, 0, 0, 0, -1, 1, -2, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -2, 0, 0, -1, -2, -1, 0, 1, 0, 0, 0, 0, -1, -1, 1, 2, 0, 0, 1, 2, -1, 1, 0, 2, 2, -1, -2, -2, -2, -1, 0, 0, 0, 0, -1, -3, 1, -1, -1, 0, 2, 2, 0, 0, 0, 0, 0, 2, 0, 3, 1, 0, 1, 1, 0, 1, 1, 1, 0, -2, -2, -1, -3, 0, -1, -1, 0, 0, 0, 2, 2, 0, 2, 0, 2, 0, 0, 2, 1, 2, 3, 4, 2, 3, 0, 0, 0, 0, 1, 0, -2, 0, -1, -2, -3, -2, 2, 0, 0, 2, 0, 0, 1, 0, 0, 2, 1, 3, 5, 3, 4, 6, 3, 2, 3, 1, 0, 0, 0, -1, -2, -2, 0, -3, -2, -2, 1, -1, 0, 0, 0, 0, 1, 1, 4, 4, 3, 4, 5, 5, 6, 5, 6, 4, 3, 2, 2, 3, 0, 2, -3, 0, 0, -2, -4, 0, 0, 1, 1, 0, 0, 0, 1, 2, 3, 4, 3, 7, 7, 5, 8, 6, 6, 4, 6, 1, 3, 0, 1, 0, -2, -1, 0, -1, -3, -1, 0, -2, 1, -1, 0, 0, 2, 2, 3, 2, 4, 6, 4, 5, 6, 9, 8, 5, 4, 1, 4, 1, -1, 0, 0, 0, 0, -1, -2, 0, -2, 1, -1, 1, 2, 0, 0, 1, 1, 2, 3, 5, 8, 8, 7, 7, 8, 5, 4, 5, 0, 0, 0, 0, 0, -2, -1, -1, -2, 0, 1, 1, 1, 2, 2, 2, 2, 3, 2, 4, 4, 8, 7, 9, 10, 6, 7, 5, 3, 3, 1, 3, 0, 0, 1, -1, -3, 0, -1, 0, 0, 0, 1, 2, 2, 2, 1, 5, 4, 3, 6, 8, 8, 7, 10, 7, 6, 9, 5, 6, 2, 3, 1, 0, 0, 0, 0, 0, -2, 0, 2, 0, 0, 1, 2, 0, 1, 5, 6, 5, 5, 9, 8, 6, 10, 9, 7, 8, 8, 3, 4, 1, 2, 0, 2, 0, -1, -1, -2, -2, 1, 0, -1, 1, 0, 3, 2, 5, 2, 5, 5, 9, 6, 8, 11, 10, 8, 6, 7, 4, 3, 3, 0, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 5, 1, 4, 7, 8, 7, 5, 9, 7, 7, 7, 3, 4, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, -1, -2, 1, 0, 0, 1, 1, 3, 4, 5, 4, 4, 9, 7, 6, 9, 5, 3, 6, 3, 2, 3, 1, 0, 1, 0, -1, 0, 0, -3, -1, 0, 1, 0, 2, 2, 3, 4, 3, 3, 5, 5, 5, 6, 5, 7, 3, 2, 2, 4, 2, 3, 3, 1, -1, 0, -1, 0, -1, -2, 0, 0, -1, 0, -1, 0, 1, 3, 4, 4, 3, 4, 3, 5, 7, 4, 5, 5, 5, 2, 2, 0, 2, 1, -1, 1, 0, -1, -2, -1, 0, -1, 0, 1, -1, 0, 2, 3, 4, 4, 2, 5, 5, 5, 5, 5, 4, 4, 4, 2, 2, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 3, 3, 1, 2, 4, 1, 1, 1, 0, 1, 4, 2, 1, 2, 1, 1, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, 2, 4, 2, 1, 2, 2, 1, 4, 0, 2, 0, 1, 0, 0, -1, 1, -1, -1, -1, -2, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 3, 0, 0, 3, 0, 0, 0, 0, 2, 0, 1, 1, 0, -1, 0, 1, 0, 1, -2, -3, 0, -1, -2, 0, -1, 0, 2, 0, 0, -1, 0, 3, 0, 2, 0, 0, 1, 0, 2, 1, 2, 2, 1, -1, 0, 0, 0, -2, -1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 2, -1, 1, 1, -1, 1, 0, -1, 1, -1, 0, 1, 1, 2, 1, 1, 1, -1, 0, 0, 0, -1, 0, -2, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, -2, -1, 0, 1, 1, -1, 0, -1, -2, -2, -2, -2, 1, 0, 0, -1, 1, 1, -1, 1, 0, 1, -1, 0, 0, 0, -1, -2, 0, 0, -1, 1, 0, -1, 0, -1, 1, 0, -2, -1, 0, 0, -1, 1, 1, 0, 1, 0, 0, 0, 1, 0, -1, 1, -1, -2, 0, -1, 0, 0, 2, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 10, 6, 8, 3, 2, 2, 4, 1, 2, 1, -1, -2, -3, -2, -2, -3, -5, -5, -4, -4, -6, -2, -4, -3, -3, 0, -3, -1, -2, -1, 9, 7, 5, 1, 1, 0, 0, 3, 1, -1, -1, -5, -6, -7, -5, -7, -8, -5, -6, -6, -3, -3, 0, -2, -1, 0, 1, 1, 1, -2, 9, 5, 3, 4, 1, 1, 0, 0, 0, -3, -2, -5, -3, -4, -8, -5, -8, -3, -4, -3, -3, -1, -2, -2, 0, 2, 0, 2, 0, 0, 5, 7, 2, 0, 0, 0, 0, 1, -1, 0, -4, -4, -5, -5, -6, -9, -4, -3, -1, 0, -2, 0, -1, 0, -1, 0, 3, 1, 0, -1, 7, 6, 2, 1, 0, 0, 2, 2, 0, 0, 0, 0, -1, -5, -5, -5, -4, -3, -2, 0, 1, 0, -1, 1, 2, 1, 3, 3, 1, 0, 7, 6, 3, 4, 1, 3, 0, -1, 0, 2, 2, 0, -2, -1, -3, -2, -6, -5, -3, 0, 3, 2, 0, 0, 0, 2, 1, 4, 0, 1, 6, 5, 2, 4, 4, 1, 0, -1, -1, -1, 1, 0, 1, 0, -3, -2, -2, -3, -3, -1, 1, -1, 2, 0, 2, 1, 1, 0, 2, -1, 5, 4, 4, 2, 2, 1, 1, 1, 1, 2, 1, 0, 2, 2, 0, -4, -2, -5, 0, 0, 1, -1, 1, 2, 0, 0, 3, 0, 0, 1, 6, 3, 0, 1, 2, 2, 3, 2, 3, 4, 2, 4, 5, 2, 2, -1, -2, 0, -3, 0, 0, 0, 0, 3, 3, 0, 0, 0, -1, -2, 4, 3, 0, 2, 0, 2, 5, 7, 6, 5, 8, 7, 7, 5, 5, 2, -1, 0, -1, -1, -1, 1, 1, 4, 3, 1, 4, 2, 1, -1, 4, 5, 4, 1, 2, 6, 3, 9, 10, 9, 9, 7, 8, 8, 5, 3, 2, 1, 3, 0, 0, -1, 0, 2, 2, 4, 4, 2, 1, 0, 3, 4, 2, 2, 2, 4, 7, 7, 9, 13, 11, 11, 11, 9, 6, 8, 6, 2, 3, 2, -1, 0, 4, 3, 3, 1, 4, 4, 1, -2, 4, 2, 0, 2, 3, 6, 6, 11, 11, 12, 14, 13, 14, 10, 11, 9, 6, 5, 5, 5, 1, 2, 3, 2, 3, 2, 2, 0, 0, -3, 4, 3, 1, 1, 2, 6, 5, 11, 12, 14, 14, 16, 14, 12, 10, 12, 8, 10, 7, 4, 5, 4, 4, 3, 5, 4, 2, 0, 0, -1, 2, 1, -1, 1, 1, 6, 7, 12, 13, 15, 14, 14, 15, 14, 12, 9, 8, 7, 8, 5, 3, 2, 3, 5, 3, 4, 1, 2, 2, 0, 3, 0, 2, 0, 2, 5, 7, 12, 14, 15, 17, 14, 13, 12, 9, 7, 7, 8, 9, 7, 5, 2, 4, 6, 7, 4, 4, 2, 0, -1, 1, 0, 0, 1, 5, 9, 11, 11, 14, 16, 17, 16, 16, 10, 10, 7, 6, 6, 5, 8, 6, 3, 4, 3, 4, 5, 5, 2, 1, 0, 0, 0, 0, 2, 5, 7, 8, 13, 16, 16, 16, 14, 14, 11, 11, 9, 10, 6, 5, 6, 3, 2, 6, 8, 4, 4, 6, 5, 1, 0, 2, -3, 0, 3, 2, 6, 7, 13, 14, 11, 13, 15, 14, 11, 9, 7, 7, 4, 7, 6, 5, 3, 2, 6, 3, 6, 4, 3, 2, 2, 1, 0, -1, 0, 2, 4, 7, 10, 13, 13, 13, 11, 12, 10, 8, 6, 7, 2, 2, 3, 1, 1, 4, 3, 5, 5, 3, 3, 0, -2, 1, 0, 1, 0, 2, 2, 7, 10, 12, 12, 10, 9, 9, 9, 5, 2, 4, -1, -1, 0, 2, 0, 0, 3, 5, 4, 4, 0, 2, 1, 4, 0, 0, 3, 0, 1, 6, 5, 8, 7, 7, 5, 8, 5, 1, 1, -2, -1, -2, 0, 1, 1, 0, 3, 5, 5, 4, 3, 0, 0, 2, 1, 2, 0, 0, 0, 0, 3, 2, 5, 5, 3, 4, 3, 0, -2, -6, -5, -4, -3, 0, 0, 1, 3, 1, 4, 1, 0, 2, 0, 2, 4, 0, 1, 1, -1, 0, 0, 3, 1, 0, 0, -1, 0, -3, -6, -5, -6, -5, -2, -1, 0, 2, 1, 1, 4, 2, 3, 3, 0, 6, 2, 0, 0, 1, 1, -1, 0, 0, 2, 0, -2, -2, -4, -7, -7, -7, -5, -2, -2, 0, 0, 0, 3, 3, 4, 3, 4, 2, 0, 6, 3, 2, 2, 0, 0, 0, -1, 0, -1, -3, -4, -2, -6, -8, -8, -7, -3, -3, -1, 0, 3, 4, 3, 2, 2, 4, 2, 1, 0, 5, 3, 1, 0, 0, -1, 0, 0, -2, -3, -1, -5, -3, -7, -6, -6, -7, -4, -2, 0, 0, 2, 1, 0, 2, 2, 4, 5, 3, 2, 6, 3, 3, 3, 0, 2, -1, 0, -2, -1, -3, -3, -7, -9, -6, -5, -3, -1, -2, 0, 1, 2, 2, 1, 1, 2, 4, 4, 3, 0, 5, 5, 0, 1, 0, 1, 0, 0, -2, -2, -1, -5, -7, -7, -6, -6, -2, -4, -1, 0, 1, 0, 3, 2, 2, 3, 0, 3, 3, 2, 5, 3, 5, 2, 1, 0, 0, 0, -1, 0, -1, -5, -6, -6, -5, -6, -2, -5, -2, -2, -2, -2, 1, 1, 2, 2, 0, 0, 2, -1, 0, 0, 0, -2, 1, -1, 0, 1, -2, 0, -1, -1, 0, -1, 0, 0, -1, 1, 1, -1, 0, 0, 0, -1, -1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, -2, 0, -1, 0, 2, 2, 0, 1, 0, 0, -2, 1, -1, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -1, 1, 1, 1, 0, -1, 1, 1, 0, 1, 2, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 0, -1, 1, 0, 0, 1, -2, 1, -1, 0, 0, -1, 2, 0, -1, 2, 0, 0, 0, 2, -1, 0, -1, 0, 1, -1, -1, -1, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 1, 0, 1, -2, -1, 1, 0, 0, -1, -1, 2, 1, -1, -2, -1, 1, -2, 0, 0, 1, -1, 0, -1, 0, 1, 2, 1, -1, 1, 0, -1, 0, -2, 0, 0, 1, 0, 1, -1, 0, 0, 0, -1, 1, 1, 0, 0, 1, -1, 1, -1, -1, 0, 0, 1, 0, 0, 1, -1, 0, 1, -1, -1, 1, 1, 0, -1, -1, -1, -1, 0, 1, -2, 1, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 0, 0, -2, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, -2, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 1, 0, -2, 0, -1, -1, 0, 1, 0, 0, -1, 0, -2, 2, -2, 1, -1, 0, 2, -1, 0, 0, 1, 0, -2, -2, 1, -1, 0, -1, 1, 0, -1, 0, 1, -1, -1, 0, 0, 0, 1, -2, 1, -1, 1, 0, -1, -2, 1, 1, 0, -1, 0, 2, 0, 0, 0, 0, -1, -2, 0, 0, -2, 0, -1, 0, -1, 2, 0, 1, 1, -1, 0, 0, 0, -1, 0, 0, 1, 1, -1, 0, -1, -1, 0, 0, 0, 0, -2, -1, 1, -2, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, 0, -1, 1, 1, 0, 1, -2, 0, -1, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, -1, 1, -1, 0, -1, -1, 0, -1, 1, 1, 1, 0, 1, -1, -2, 1, -1, 1, 0, -1, -1, -1, 0, -1, 1, -1, -1, -2, 0, 0, 0, -2, 0, -1, 1, -1, -1, 0, 0, -1, 1, 0, 1, 1, -1, 1, 0, 1, 0, -2, -1, -1, -1, 0, -1, 0, -1, 0, 1, 0, -1, 0, 1, -1, -1, 0, 0, -1, 0, -1, -1, 0, 1, -1, 0, 1, -1, 0, 1, 0, -2, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, -1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, -1, -1, -1, -1, -1, -1, -1, -1, 0, -1, 0, -2, 0, 1, 1, 1, 0, -1, 2, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, -2, 1, 1, 1, -1, 0, 0, 0, -2, -1, 1, 1, 0, -1, 0, 0, 1, 1, 1, -1, 1, -1, 1, 0, 0, 1, 1, -1, 1, -1, 0, 0, -1, 0, -2, 1, 1, -1, 1, -1, -1, -1, 0, -1, 1, -1, -2, 0, 2, 1, 1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, -2, 0, 0, -2, 0, 0, -1, 0, 1, 1, -1, 0, 0, 0, -1, 1, 1, -1, 1, -2, 0, -1, 1, 0, 1, -1, 1, 1, -2, 0, -1, 2, -1, 1, -1, -2, -1, 1, 1, 0, 0, -1, 0, -2, 1, 0, 0, 0, 1, -2, 0, 2, 0, 0, 0, -2, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 1, 0, 0, -1, -1, -1, -1, -1, 0, -1, 1, 0, 1, 0, -1, 1, -1, 0, 0, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, 1, -1, 0, -1, -1, 0, 0, 1, -1, 0, 1, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, 1, -1, 1, 0, 1, 0, 1, -1, 0, 1, 0, 0, 1, -1, 0, -1, 1, -1, 0, -1, 1, 2, 0, 0, 1, 0, 1, 0, 0, -1, 1, -1, 0, -2, 1, 1, -1, 0, 0, -1, 0, 0, 0, 1, 1, -1, -1, 0, -1, 1, -1, 1, -2, -2, -1, 0, -1, 2, 1, 1, 0, 1, -1, 1, 1, -2, 0, 0, -1, 0, 1, 0, 1, 0, 0, 1, 0, -1, 0, -1, 0, 1, 0, 0, -1, 1, 1, 1, -1, -1, 0, 1, -1, 1, -1, 0, 1, 0, -1, 0, 0, -1, 1, -2, 0, 2, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, 0, 1, 1, -1, 0, -1, 0, -1, 0, -1, 0, 1, -1, -1, -1, 1, 0, 0, 0, -1, 1, 1, 0, -1, -1, 2, -2, 0, 0, 0, 0, -1, 0, 0, -1, 1, 1, -1, -1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, -1, 0, 1, 0, -1, 1, -1, -2, -1, -1, 0, 0, 0, 0, 1, -1, 0, 1, 0, -1, 0, -1, -1, -1, 1, 0, 0, 1, -1, 1, 0, 2, 1, 1, 0, -1, 0, 0, 2, 0, 1, -2, 0, -1, 1, -1, 0, 0, 0, 0, 0, 1, 2, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, 2, 0, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, -1, -2, 0, -1, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 1, -1, -1, -1, -1, 1, -1, 0, 1, -2, 0, 0, 1, 2, 1, 0, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 2, -1, 1, -1, 1, 0, 0, 1, -1, -1, 0, 0, 1, 1, 0, -2, 0, 0, 0, 0, -1, 0, 1, 1, 1, -1, -1, 0, 0, -2, 2, 0, 0, -1, 0, 0, -1, 1, 1, 0, -1, -1, -1, 1, -1, 1, -1, 1, 0, 0, 0, 1, 0, -1, 2, -1, 1, 0, 0, 1, -1, 0, -1, 0, 0, -1, 0, 1, 1, 0, -2, 0, 1, 0, -1, -1, 2, 1, 1, -1, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, -2, 0, -1, 0, 0, 0, -1, 0, 1, -2, 0, -1, -1, 1, 0, 0, 1, 1, -1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, -2, 0, 1, 0, -1, -1, 1, -1, 1, 1, 1, 1, 2, 0, -1, -1, 1, -1, 0, -1, 1, 0, 0, 0, -1, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, -1, 0, 0, -2, 1, 0, 1, -1, 0, 0, 1, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, -1, -1, 0, 1, 0, 0, 1, 1, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, 1, 1, 0, 1, 1, -1, -1, 0, 0, 2, 0, -1, 1, 2, -1, 1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 1, 0, 0, 1, 0, -1, 1, 1, -1, 0, 1, 0, 0, -1, 0, -1, 0, 1, 0, -1, 0, -1, -2, -1, 1, 1, -1, 0, 0, -1, 1, 1, 0, 0, -2, 0, 0, 1, 1, -1, 1, -1, 0, 0, 1, 1, -2, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, -1, -1, 1, 0, -1, 1, 0, 1, 0, -1, -1, 0, 1, 0, 1, 0, 2, -1, -1, 0, 0, 0, 0, 1, -2, 2, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, -1, 1, 0, 0, 0, 1, 0, -1, 0, -1, -1, 0, -1, -2, -1, 2, 1, -1, 0, 0, -1, 1, -1, 0, 0, 1, 1, 0, 0, -2, 0, -1, 1, -1, 0, 1, 1, 0, 0, -2, -1, 1, 0, 0, 1, -1, -2, -2, 0, 1, -1, 2, -1, 0, 0, 1, -1, 0, 0, 0, 1, -2, 1, -1, -1, -1, -1, 1, 0, -1, -1, 0, -1, 1, 0, -1, 0, -2, 0, 1, 0, 1, 1, 1, 0, 1, 0, 0, -1, -1, 0, 1, -1, -1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 2, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, -2, -2, 1, 0, 1, 0, 0, -1, 0, -1, 0, -2, 0, 0, 0, 1, 0, 1, 2, -1, 0, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 1, 1, 2, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, -2, 0, -2, 2, -1, 1, -1, 0, 1, 1, 0, 0, 0, 1, -1, -1, -1, 0, 1, 1, 0, 1, 1, 1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 1, -1, -1, 0, -1, -1, 0, -1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 1, -2, 2, -2, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 1, 2, 1, -1, 1, 0, -1, 0, -1, 0, -1, -1, 2, 0, 1, -1, -1, 0, 1, 0, 0, 1, 1, 0, 1, 0, 0, -1, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 1, 1, -1, -1, 1, 1, -1, 0, 0, 0, -1, -1, 1, -1, 1, 1, 0, 0, 0, 1, -1, 1, 0, -1, 0, 0, 0, -1, 1, 1, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 1, 2, -1, -2, 0, 0, 0, 0, -1, 1, 0, -1, -1, 1, -1, 0, 1, 0, 0, 1, -1, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 0, 1, -1, -1, 2, 0, 2, 1, 1, 1, 0, 1, 1, 1, 1, 0, -1, 0, 0, 1, 0, -1, -1, 1, 0, 0, 0, 0, 4, 3, 5, 4, 3, 3, 4, 1, 4, 2, 5, 2, 7, 3, 5, 1, 3, 1, 3, 0, 1, 1, 4, 3, 2, 2, 2, 1, 0, 0, 0, 3, 1, 2, 1, 3, 1, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 3, 1, 3, 3, 3, 4, 0, 2, 1, 0, 0, 0, 3, 0, 1, 0, -2, 1, -2, -2, -3, -4, -4, -3, -2, -1, -1, 0, -1, 1, 1, 2, -1, 3, 2, 3, 3, 2, 1, -3, 0, 4, 1, 2, 0, 0, -1, 0, 1, -3, -1, -3, -3, -3, -4, -4, -3, -1, -2, 0, 0, 0, -1, 0, 3, 0, 1, 1, 3, -2, 0, 3, 2, 0, -1, 1, 0, 0, -2, -2, -2, -2, -2, -4, -2, -4, -3, -2, 0, 0, 0, -1, 0, -1, 1, 3, 1, 0, 1, 0, 0, 2, 2, 0, -1, -2, -2, -3, -1, 0, -2, -2, -3, -1, -1, -4, 0, 0, 0, 0, -2, 0, 0, -1, 0, 3, 0, 1, -2, -2, -1, -2, 0, -1, 0, 0, -1, 0, -1, 0, -4, -2, -3, -2, -2, -3, -3, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, -2, -3, 0, 0, 0, 0, 2, 1, -2, -2, 0, 0, -3, -4, 0, -3, -4, -5, -2, -4, -1, -2, 0, -1, -1, -3, -2, -2, -1, -3, -1, -3, 0, -1, -2, 0, 0, 1, 1, 0, -3, 0, 0, 0, 0, 0, 1, 0, -2, 0, 0, -1, 0, -1, 0, -2, -1, -3, -5, -2, -2, -4, 3, 1, 0, 0, 1, -1, -1, -1, -1, -2, -1, -1, 4, 4, 2, 3, 0, 1, 0, -2, -3, -2, 0, 0, -2, 0, -2, -1, -1, -2, 2, 0, -1, 0, -2, 0, -3, -2, 0, -2, -2, 2, 5, 5, 6, 4, 1, 1, -1, -1, -4, -2, -3, 1, 0, -2, -2, -3, -5, -3, 0, 1, 0, -3, 0, -1, -2, -1, -1, -1, 0, 4, 5, 8, 6, 6, 6, 6, 2, 2, -1, -3, -1, -1, -1, -3, -1, -3, -4, -3, -2, -1, 0, -1, -3, -2, -2, 0, -1, 1, 2, 6, 6, 6, 9, 11, 10, 8, 4, 3, -3, -5, -2, -5, -3, -2, -5, -3, -5, -4, 0, -1, 0, -3, -4, -3, -1, -2, 0, 2, 2, 7, 8, 11, 12, 11, 8, 6, 6, 4, 0, -2, -5, -3, -5, -2, -6, -4, -3, -6, -3, 0, -2, 0, 0, -3, -2, 0, 0, 3, 4, 3, 9, 10, 8, 8, 9, 7, 6, 3, 2, -1, -3, -7, -3, -4, -4, -3, -6, -2, 0, 0, 0, -2, -2, -1, -5, -3, 2, 2, 2, 7, 9, 5, 6, 7, 9, 9, 7, 6, 6, 0, -5, -5, -6, -5, -4, -5, -6, -5, -2, 1, -1, -2, -1, -3, -3, 0, 0, 2, 4, 4, 7, 6, 7, 9, 8, 11, 7, 7, 2, 0, -6, -6, -5, -3, -2, -1, -2, -1, 0, -2, -1, -4, -3, -5, -2, -2, 1, 1, 3, 3, 8, 7, 10, 10, 12, 11, 7, 6, 1, -5, -4, -6, -3, -5, -1, -2, 0, -2, -1, 0, -1, -4, -1, -5, -1, 0, 1, 1, 3, 6, 6, 8, 9, 11, 11, 9, 4, 1, 0, -4, -7, -5, -3, -4, -2, 0, 0, -3, -1, -3, -4, -3, 0, -1, -2, -1, 0, 1, 2, 5, 5, 9, 6, 8, 6, 4, 1, 1, 0, -5, -5, -2, -4, -3, -1, -1, 0, -4, -1, -1, -2, -1, 0, -2, 0, 0, -1, 0, 1, 2, 3, 6, 5, 5, 5, 2, -1, -1, -2, -2, -3, -3, 0, 0, 0, -3, -2, -4, 0, -1, -1, 1, 0, 0, 0, -3, 0, 0, 2, 0, 0, 3, 2, 1, 0, 0, -3, -1, -2, 0, -2, -1, -1, 0, -3, -5, -3, -4, 0, -1, -1, -2, 0, 0, -3, -4, 0, 0, 0, 1, -1, 0, 0, -3, -4, -1, 0, 0, 0, -2, -2, 0, -3, -1, -3, -3, 0, -2, 0, -1, -1, 0, 0, -2, -1, -1, 0, -2, 0, -1, -1, -1, -4, -5, -3, -3, -2, 0, -2, 0, 1, 0, -1, 0, 0, -1, 0, 3, 0, -1, 0, -1, 0, -2, 0, -2, -2, -3, -3, -3, -4, -6, -7, -4, -3, -2, -2, 0, -1, -1, 0, -1, -1, 0, 2, 4, 2, 4, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, -3, -3, -1, -6, -5, -7, -3, -5, 0, 2, 0, 0, 0, 1, 0, 1, 3, 5, 5, 3, 1, 0, 0, -1, 0, -2, 0, -2, 0, -3, -1, -1, -1, -1, -2, -4, -4, -3, 0, 0, 2, 2, 0, 2, 3, 4, 6, 6, 2, 0, 0, 2, -1, -1, -1, -1, 0, 0, -1, -1, 1, 0, -2, -2, -2, -5, -4, -3, -2, 0, -2, 0, 0, 0, 4, 4, 2, 3, 0, 0, 0, 0, -2, -1, 0, -2, 1, 0, 1, 0, 0, 2, 2, -2, -3, -5, -1, -3, -1, -1, 0, -1, 1, 0, 1, 4, 1, 0, 0, 1, 1, 0, -1, 1, 0, 1, 2, 2, 0, 0, 4, 3, 2, 0, -1, -1, -2, -2, -1, 0, -1, 1, 2, 0, 2, 4, 1, 1, 1, 3, -2, 1, 0, 2, 2, 1, 0, 0, 0, 0, 1, 3, 0, 0, 4, 3, 0, 1, 3, 2, 1, 2, 2, 1, 1, 2, 1, 3, 0, 0, -1, 0, 0, 2, 0, -1, 1, 1, 2, 2, 0, 2, 0, 1, 0, 0, 0, 0, 2, 2, 0, 2, 1, 2, 1, 3, 2, 2, 0, 3, 0, 0, 0, 0, 1, 1, -1, 1, 1, 0, 0, 0, -1, 0, 0, 2, 1, -1, 0, 1, 1, 2, 0, 0, 2, 1, 2, 3, 1, 2, -2, 0, 0, 0, 2, 0, 1, 1, 0, 0, 0, -2, 0, 0, -1, 0, -2, 0, 0, 0, 1, 1, 0, 1, 2, 0, 0, 0, 3, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, -2, -1, 1, -1, 0, -2, 0, -1, 0, -2, 0, 0, -1, 0, 0, 0, 0, 2, 2, 0, 1, 1, 1, 1, -2, 0, 1, 1, 1, 0, 0, -1, 0, 0, -2, -2, 0, -1, -2, -2, 0, -2, 0, -1, 0, 1, 2, 1, 1, 1, 1, 0, 0, 1, -1, -2, -2, -1, 1, -1, 0, 0, -3, -1, -1, -2, -2, -3, -1, 0, -1, 0, 0, 1, 0, -1, 1, 1, 1, 0, 1, 0, 1, -1, 0, 0, -1, -1, -2, 0, 0, -3, 0, -3, 0, -2, -2, -2, -1, 0, 0, 0, -2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, -2, -1, -3, 0, -1, 0, -2, -1, 0, 0, -2, 0, -2, 0, 0, 1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, -2, -1, -2, 0, -2, -1, -3, 0, 0, -2, -1, -1, -2, -1, -1, -2, 0, 0, -2, 1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -2, 0, -3, 0, 0, -3, -2, -3, 0, 0, -1, 0, -2, -1, -2, 0, -1, -3, -1, 0, -1, -2, 0, 1, -2, -2, 0, 1, 0, -2, 0, 0, -1, -2, -3, -2, -1, 0, -2, -2, -1, -1, -2, -2, 0, 0, -2, -1, 0, -2, 0, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, -3, -3, -3, -1, -1, -2, 0, -1, -1, -1, 0, -3, -1, -1, -3, 0, -3, 0, -2, 1, 0, 0, 2, 2, -2, 0, 0, -1, 0, -1, -2, -2, -1, -1, -1, 0, 0, -2, -2, -2, -1, 0, -2, -1, -2, 0, -2, 0, 1, 0, 0, 1, -1, 1, 1, 0, -3, -2, -2, 0, -2, 0, -2, -1, -1, 0, 0, 0, -2, -1, 0, -2, 0, -2, -2, -1, 0, -1, -1, 0, -2, 1, 0, -1, 0, 0, -2, -1, -2, -3, -2, -2, -1, -1, 0, -1, -1, -2, -1, 0, 0, 0, -1, -3, -2, -2, 0, -2, 0, -1, 0, -1, 0, 1, -2, 0, -3, -2, -4, -2, -1, -1, -1, 1, 0, -2, 0, 0, -2, -1, -1, -1, -3, -4, -2, 0, 0, 0, 0, -1, 0, 2, 1, -1, 0, -3, -3, 0, -4, -2, -3, -2, 0, -1, 0, -2, 1, 0, 1, 0, 1, -2, -2, -2, -3, -1, -3, 0, 0, -1, 1, 1, 1, -1, -1, -3, -2, -3, -3, -3, 0, -2, -3, -1, 0, -2, 0, 1, 0, -1, -2, -2, -2, -2, -2, -2, 0, 0, -1, 0, -1, 0, -1, 1, -2, -2, 0, 0, -1, -1, -1, 0, 0, -3, 0, -1, -1, 0, 0, -1, -1, -1, -2, 0, -2, 0, -3, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, -3, -3, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, -2, 0, -3, -1, -1, 0, 0, 1, 0, -1, 1, 1, -1, 2, -1, 1, 0, 0, -3, -1, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, -3, 0, -1, 0, 0, -2, 0, 0, 1, 0, 1, 0, -1, -1, 0, -1, 0, -2, 0, -1, -2, 0, 0, -3, 0, -1, -2, -2, 0, -2, -1, -1, 0, -1, 0, 1, 0, -1, -1, 0, 0, 2, 0, 2, -1, 1, 0, -2, 0, -1, 0, 0, -2, -2, 0, 0, -2, 0, 0, -2, -1, 1, 0, 1, -1, 0, -1, 0, 1, 2, 2, 2, -2, 0, 1, 0, 2, 0, -2, 0, 0, -1, 0, 0, 0, 0, -1, -2, -2, 0, 0, 0, 0, 1, 0, 1, -1, -1, 0, 1, 3, 3, 1, 1, 0, -1, 1, 0, -1, 1, 0, 0, 1, -1, 0, 0, 0, -2, 0, 0, -2, 0, 0, 1, 1, -1, 0, 1, 0, 2, 1, 2, -1, 1, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, -2, 0, -2, -1, -1, 1, 0, 0, 2, 2, 3, 1, 0, 0, 2, 0, -1, 0, 0, 0, 1, 1, 2, -1, 0, -1, 0, 1, 2, 0, -2, 0, -1, 1, 1, 0, 0, 0, 1, 2, 1, 0, 2, 1, 2, 0, 1, -1, 1, 1, 0, -1, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, -1, 1, 1, 3, 0, 2, 2, 1, 1, 2, 1, 0, 0, 2, 0, 2, 2, 1, 3, 2, 2, 0, 2, 2, 1, -1, 2, 2, 3, 0, 2, 0, 2, 3, 0, 0, 2, -3, -1, 3, 3, 7, 6, 3, 5, 3, 3, 6, 4, 4, 5, 8, 7, 6, 3, 5, 3, 8, 7, 8, 7, 6, 8, 8, 6, 8, 7, -3, 0, 2, 2, 3, 6, 2, 2, 3, 4, 3, 1, 0, 0, 0, 2, 2, 2, 4, 4, 4, 5, 3, 7, 7, 7, 6, 6, 8, 5, -3, 0, 3, 2, 1, 0, 3, 2, 3, 3, 2, 0, -2, -1, -4, -1, -3, 0, 2, 1, 4, 5, 3, 3, 5, 6, 7, 5, 6, 6, -3, 0, 4, 3, 2, 2, 2, 0, 1, 4, 2, -2, -2, -4, -4, -3, -2, 0, 0, 4, 1, 4, 3, 2, 2, 6, 5, 4, 7, 6, -1, 1, 3, 2, 3, 0, 0, -2, 0, -2, 0, -4, -6, -4, -5, -4, 0, -2, 0, 1, 2, 4, 4, 4, 3, 3, 6, 3, 6, 1, -4, 0, 0, 0, -1, 0, -1, -2, -5, -2, -3, -4, -4, -8, -9, -5, -4, -6, -5, 0, -1, 0, -1, 1, 2, 1, 4, 5, 1, 0, -2, 0, 0, -2, 0, 0, -2, -1, -2, -2, -5, -4, -5, -10, -9, -10, -10, -6, -5, -2, -3, 0, 1, 0, 2, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, -2, -6, -6, -3, -4, -7, -7, -9, -5, -8, -7, -4, -1, 0, -1, 0, 2, 3, 0, 0, -1, 0, 1, 0, 2, 0, -4, -3, -4, -4, -4, -8, -9, -6, -5, -4, -6, -4, -5, -4, -7, -7, -5, -5, -2, 1, 2, 2, 1, -2, -2, -2, 0, 0, 1, -3, -1, -2, -3, -7, -8, -8, -7, -9, -6, -3, -1, -1, -5, -4, -3, -4, -8, -5, -4, -1, 1, 0, -1, 2, 0, -1, 1, 0, 0, -1, -3, -3, -6, -3, -6, -6, -5, -7, -1, -3, -2, 0, 0, -2, -2, -3, -5, -7, -3, -1, -2, 0, -2, 0, 0, -2, 0, 0, -2, -2, -4, -7, -3, -3, -5, -5, -4, -3, -4, -2, 1, 2, 3, 0, 0, -3, -3, -7, -7, -4, -3, -2, -3, -1, -2, -1, 0, -1, -1, -2, -5, -6, -9, -6, -10, -6, -6, -6, -2, -2, 0, 0, 0, 0, 0, -1, -4, -8, -6, -8, -5, -5, -1, -2, -5, -4, -1, 0, -2, -3, -7, -6, -10, -8, -10, -7, -6, -6, -2, -1, -2, 0, -2, 0, 0, 0, 0, -4, -7, -8, -6, -5, -2, -5, -3, -2, -5, -1, 0, -2, -4, -5, -10, -11, -9, -9, -9, -5, -5, -6, -5, -3, 0, 0, 1, 0, 2, -4, -3, -8, -6, -3, -2, -4, 0, 0, -2, 0, 0, 0, -4, -9, -11, -7, -6, -6, -7, -6, -5, -6, -4, -1, 0, 2, 0, 3, 3, -2, -4, -9, -6, -3, -1, -3, 0, 0, -3, 0, -3, -4, -5, -9, -12, -9, -6, -8, -7, -6, -2, -3, -1, 0, 3, 2, 3, 2, -1, -4, -7, -7, -5, -4, -5, -3, 1, 0, 0, -3, -1, -3, -5, -8, -10, -8, -9, -7, -7, -6, -4, 0, 0, 0, 1, 3, 3, -1, -4, -8, -9, -9, -7, -7, -3, -1, 0, 0, 0, 0, -2, -4, -5, -5, -7, -9, -9, -6, -8, -5, -2, -2, -2, 0, 0, 0, 0, -4, -6, -8, -7, -5, -5, -4, -1, 1, 1, 0, 1, 0, -2, -1, 0, -4, -6, -8, -6, -5, -5, -7, -4, -3, -1, -3, -3, -5, -5, -6, -7, -9, -6, -6, -1, -3, -1, 0, -1, 0, -1, 1, -3, 0, -2, -1, -5, -6, -7, -9, -6, -9, -7, -8, -7, -9, -9, -9, -8, -6, -6, -4, -4, -3, -2, -2, 0, 0, -1, 0, 0, 0, 0, 0, -2, 0, -2, -7, -7, -9, -6, -6, -5, -8, -7, -9, -8, -10, -9, -7, -5, -4, -3, -4, 0, 0, -1, -1, 1, 0, -2, 0, -1, 1, -1, 0, -3, -4, -8, -8, -5, -5, -10, -8, -10, -10, -10, -7, -6, -4, -3, -4, -1, -1, -2, -2, 0, 1, 1, 3, 1, 1, 1, -1, 0, -1, 0, -3, -2, -4, -7, -6, -9, -10, -9, -9, -10, -6, -4, -1, -3, 0, -1, 1, -1, 0, 4, 4, 3, 6, 2, 4, 0, -1, -2, 0, 0, 0, -3, -3, -4, -6, -4, -8, -9, -8, -8, -6, -3, -1, 0, 3, 0, 1, 0, 5, 4, 9, 8, 10, 4, 3, 4, 1, 1, 0, 0, -2, 0, -3, -2, -3, -5, -5, -8, -9, -4, -6, -4, 0, 0, 1, 0, 0, 2, 7, 7, 8, 8, 6, 0, 3, 1, 3, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, -6, -4, -6, -2, -1, 0, 0, 0, 0, 2, 3, 6, 8, 7, 7, 7, 1, 2, 2, 0, 0, -1, 0, 0, 0, 4, 3, 3, 3, 0, 0, -3, -3, -4, -1, 0, -2, 2, 4, 4, 6, 5, 6, 5, 4, 6, -1, 0, 0, 2, 0, 0, 4, 4, 5, 3, 6, 6, 6, 5, 4, 2, 1, 0, -2, 0, 0, 1, 1, 3, 6, 9, 4, 4, 5, 4, 1, 1, 4, 5, 7, 6, 8, 7, 6, 7, 8, 7, 10, 8, 6, 3, 6, 4, 3, 2, 5, 4, 4, 7, 7, 8, 6, 5, 6, 7, 2, 0, 3, 4, 2, 1, 2, 3, 4, 3, 5, 4, 7, 8, 8, 6, 3, 3, 2, 6, 6, 4, 2, 4, 2, 4, 4, 2, 1, 0, 1, 1, 2, 2, 2, 0, 1, 1, 4, 2, 3, 2, 1, 6, 6, 2, 5, 2, 3, 3, 1, 4, 1, 3, 3, 3, 3, 2, 2, 0, 0, -1, -1, 2, 0, 1, 1, 0, 1, 2, 3, 0, 2, 0, 4, 4, 3, 0, 1, 2, 4, 2, 3, 4, 4, 3, 2, 4, 4, 0, -2, -1, 2, 0, 0, 2, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 2, 0, 1, 0, 0, 0, 1, 3, 2, 2, 3, 2, 0, 1, 0, 1, 0, 1, 1, 2, 1, 0, 1, -1, -2, 2, 0, 0, -1, 0, 0, 2, 1, 2, 3, 3, 2, 4, 2, 3, 1, 2, 1, -1, 2, 0, 1, -1, 0, -2, -1, 1, 2, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 2, 1, 1, 3, 2, 1, 4, 1, 2, 2, 0, -1, 1, 0, 0, 1, 0, -1, -1, 1, 2, 0, 0, -2, 0, 0, 0, 0, -1, 2, 3, 0, 2, 3, 1, 3, 4, 0, 2, 3, -1, 0, 0, -1, -1, -2, -2, 0, -2, -2, 0, -3, 0, 0, -1, -2, -2, 0, 0, 1, 0, 1, 2, 1, 0, 0, 1, 2, 1, 0, 1, -1, -1, -1, 0, 0, -1, -1, 0, -1, -2, -2, -2, 0, -3, -1, -1, -1, 1, 1, 1, 0, 0, 0, 1, 2, 2, 2, 2, 1, -1, -2, -2, -1, 0, -1, -1, -3, -1, -3, 0, 0, -1, -1, 0, -1, -3, 0, 0, -1, 3, 2, 1, 3, 0, 0, 1, 1, -1, 0, 0, 1, -2, 0, 0, -3, -4, -2, -2, -5, -2, -3, -1, -2, -3, -3, 0, -3, -1, 0, 0, 1, 2, 4, 1, 0, 2, 0, 0, 1, 0, 0, -2, -1, 0, 0, -1, -4, -2, -2, -2, -2, 0, -3, -4, -3, -3, -2, -2, -1, 0, 0, 1, 1, 0, 2, 1, 0, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, -1, -2, -4, 0, -2, -2, 0, 0, 0, -1, -2, 0, -4, 0, 2, 1, 0, -1, 0, 1, 1, 0, 0, -1, 0, -2, -2, -4, -4, -3, -2, -4, -5, -4, -4, -1, -3, -1, -1, 0, 0, -1, -2, 0, 1, 1, 3, 0, 0, -2, 1, 0, 1, -1, 0, -3, -1, -2, -3, -3, -6, -3, -5, -1, -1, -2, -4, -1, 0, -1, 0, -2, -2, -2, 0, -1, 1, 0, 2, 0, -1, 0, 1, 0, 0, -4, -1, -2, -4, -4, -6, -7, -5, -4, -1, -2, -4, 0, -3, 0, -1, -1, -2, -1, -2, 0, -1, 0, -1, 1, 2, 1, -1, -1, 1, -3, -3, -2, -3, -3, -5, -6, -2, -2, -3, -5, -5, -2, 0, -3, -1, 1, 0, -2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, -1, -3, -3, -4, -3, -1, -3, -3, -4, -3, -2, -2, -5, 0, 1, 0, 0, 2, -3, -3, -1, -1, 0, 1, 2, 0, -1, 0, 0, -3, -1, -2, -5, -4, -5, 0, -3, -6, -4, -1, -3, -2, -3, 1, 1, 0, 1, 1, -3, -3, -1, 0, -2, -1, 0, 1, 0, 1, 0, -4, 0, -2, -1, -5, -1, 0, -2, -3, -4, -3, 0, 0, -2, 0, 2, 1, -2, 0, 0, -1, 1, -2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -4, 0, 0, -4, -3, -4, 0, 0, 0, 0, 1, -1, 0, -1, -3, -2, 2, 0, -1, 3, 1, -1, 0, 2, -1, 0, 0, 0, -1, -1, -2, -1, -1, -2, -1, -2, -2, 0, -1, -3, -1, -1, 0, 0, -1, -2, -1, 0, 1, 0, -1, 1, 2, 0, 1, -1, 0, 0, 0, 0, 0, -2, 1, -1, 0, 0, 0, -2, 0, -2, -2, -1, -1, -2, -1, -1, 0, -1, 1, 0, 0, 0, 2, 0, 0, 0, -2, 2, 2, 0, -1, 0, -2, 0, 1, 0, 0, -1, -2, 0, 0, 0, 1, 2, -1, 1, 0, 0, 0, -1, 0, 0, 3, 1, -1, 1, 1, 1, 0, 1, 1, -1, 0, 0, -2, 0, -3, 0, -1, -4, 0, 1, 0, 1, 0, 0, 1, 0, 2, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 2, 2, 0, -1, -1, 1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 1, 1, 1, 3, 0, 3, 2, 4, 0, -1, 0, -1, -1, 0, 0, 1, 2, 2, 1, 2, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, -1, 2, 2, 3, 4, 2, 1, 0, 1, -1, -1, 0, 1, 2, 1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 3, 0, 0, 2, 1, 1, 1, 4, -1, 0, 0, -1, 2, 2, 2, 2, 3, 2, 0, 1, 0, -1, -1, 0, -1, 0, 0, 1, 3, 3, 3, 2, 3, 3, 0, 0, 1, 1, -2, 2, 1, 1, -1, -1, 0, 0, 0, 3, 0, 0, 1, 2, -2, 1, -1, -2, 0, -1, 0, 0, 2, 2, 3, 0, 1, 0, 4, 4, 1, 0, -1, 0, 0, 0, -1, 0, -1, -1, -2, 1, -2, 1, 0, 0, 0, 1, -1, 0, 1, 2, 1, 1, 0, 1, -1, -1, 1, 1, -1, 1, -1, 1, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 0, 0, 1, 0, 1, 0, -1, -1, 0, -2, 0, -1, 0, 1, 0, 1, 0, -1, 1, 0, 0, 1, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, 0, -1, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, 1, 1, -1, 0, 1, 1, 0, 0, 0, -1, -2, -1, 0, 1, 1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 0, 2, -1, 1, -1, 1, 0, 1, 2, 0, 0, 2, 1, -2, 1, -1, -1, -1, 0, -2, 0, 0, -1, 0, -1, -1, 0, -1, 0, -1, -2, -1, -1, -1, 1, 1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, 1, 0, -1, 0, 1, 0, -1, -1, -1, 1, -1, 0, 0, -2, -2, -1, 1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, 1, 2, 0, 0, -1, -1, 1, -1, 1, 0, 1, -1, 0, 1, 0, -1, -1, 0, 0, -1, 1, 1, 1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, 1, 0, 0, 1, 0, -1, 0, -1, 1, 0, 0, 1, 1, 0, -1, 0, -1, -1, 0, 0, 0, -1, 1, 0, 0, -2, 0, 2, -1, -1, -1, -1, 2, -1, -1, -1, 1, 0, -1, -1, 2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, -1, -1, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 2, 0, 1, -1, -1, 0, 1, 0, 1, 1, 0, -2, 0, 1, 1, 0, 1, -1, -1, -1, 0, 1, 2, 0, -2, -1, -1, -2, 1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 1, 1, 0, 0, 1, 0, 1, -1, 0, -1, -1, 1, -1, -1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, 1, 1, -1, -1, 1, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -1, 1, 1, 0, -1, -1, -1, 0, 0, 2, 1, 0, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 1, -2, 0, 0, -1, -2, 1, 1, 1, 0, 0, 2, -1, -1, 1, -2, 1, 1, 1, 0, 0, 0, 0, 1, -1, 1, 1, 1, 0, 0, -1, 1, -1, 1, 0, 1, 2, -1, 1, 0, 1, -2, 1, 0, 0, -2, -1, -2, 1, 0, -1, 1, 1, -1, 1, 0, 0, 0, -1, 0, -2, 0, 0, -1, 1, 0, -1, -1, 0, 0, 0, 1, -1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 2, -1, -1, 1, 1, 0, 0, 0, 0, -1, 1, 1, 0, -1, 1, -1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, -1, 1, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -2, 2, -1, -1, -1, -1, 0, 2, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, -1, -1, 1, -1, -2, 0, 2, -1, 1, 0, -1, 0, 1, 1, 1, -1, -1, 1, -1, -1, -2, 1, -1, 0, 1, 1, 0, -2, 0, 0, -1, 0, -1, 1, -1, 1, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, -1, -1, 1, 0, -1, -2, 1, 1, -1, 0, 1, 0, -1, 0, -2, 1, 0, -1, -1, 1, 0, 0, -2, -1, 0, -1, -2, -1, 0, 0, 0, 0, -1, 0, 0, -1, 1, -1, -1, 0, -1, -1, -1, 0, 0, 0, 0, 1, -1, -1, 0, -1, -1, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 2, 0, 0, -1, 0, 0, 1, 0, 1, -1, 2, 1, 0, 0, 1, 0, -1, 2, 0, -1, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, 0, 0, -1, 0, 1, 0, -1, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -1, 0, 1, -1, 1, 0, -1, 1, 0, 1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 1, -2, -1, -2, 0, 0, -1, 1, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 0, 2, 0, -1, 0, 2, 1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, 1, 1, 1, 0, 1, 0, 1, -1, -1, 0,
    -- filter=0 channel=7
    0, 1, -2, -1, 0, -2, 0, -1, -1, -1, 1, 1, 0, -2, 0, -2, -1, -1, 0, -2, -2, 0, 0, -1, 0, -1, -2, -2, 0, -3, 0, -1, 0, 0, -1, 0, -1, 2, 1, 0, -2, 0, -1, -1, 0, -1, -1, 0, -1, -2, -1, 0, 0, 0, -1, 0, -3, -1, 0, -4, -1, 0, 0, 0, -1, -1, 0, 2, 1, -1, -1, -1, 0, 1, 0, -1, -3, -1, 0, 0, -2, -1, -2, 0, 0, -3, -2, -3, -2, -2, 0, 0, 0, 0, 2, 0, 2, 1, 2, 0, 0, 1, 0, 1, 0, 0, 1, 1, 0, -2, 0, -1, -1, 0, -3, 0, -3, -2, 0, -3, 0, 1, 2, 1, 1, 2, 1, 0, 0, 0, 0, -1, 1, -1, 0, 0, -2, -1, -2, -1, 0, -2, -2, 0, 0, 0, 0, -1, -2, 0, 3, 0, 0, 2, 0, 0, 2, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -3, -1, 0, -1, -2, 0, 0, -2, -1, 0, -1, 1, 1, 2, 0, 0, 3, 2, 1, 0, 2, 0, 1, 0, 1, -1, 0, 0, 0, -3, 0, 0, 0, -3, 0, -3, -2, 0, -3, -2, -2, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, -2, -1, 0, -2, -3, -3, -1, -2, -2, 1, 1, 2, 0, 0, -1, 0, 1, 2, 0, 2, -1, 1, 0, 0, 0, 0, 0, -1, -1, 0, -2, -1, -2, 0, 0, -1, -3, 0, -1, -1, 2, 0, -1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 1, 0, 1, 0, -1, 0, -2, 0, 0, -2, -1, -1, 0, -1, -2, 0, -1, 2, 0, 2, 0, 0, 2, 0, -1, 0, 2, 0, 0, 2, 0, 1, 1, 2, 0, 0, -3, 0, -2, -1, 0, -2, -1, 0, -3, -2, -1, -1, 2, 0, 0, 0, 1, 0, 0, 2, 2, 2, 1, 2, 0, 3, 0, 0, -1, -1, -3, 0, -3, -2, 0, -2, 0, -1, 0, 0, -1, 2, 1, 0, 2, -1, 1, -1, 0, 0, 0, 0, 0, 2, 0, 2, 4, 0, 1, -2, -4, -4, -3, -2, 0, -1, 0, -1, 0, -1, -1, 1, 0, 1, -1, -2, -2, 0, 2, 0, 0, 0, 0, 1, 0, 0, 4, 1, -2, 0, -2, -4, 0, 0, 0, -1, -4, -1, -1, -4, -4, 2, 0, 0, 0, 0, -2, 1, 0, 2, 0, 0, 0, -1, 2, 3, 3, 3, 0, -2, -2, -3, -3, -3, 0, 0, -3, -3, -2, -1, -2, 0, 1, -1, 2, 0, 0, 1, 0, 2, 0, -1, 2, 1, 3, 1, 2, 4, 2, -3, -1, -3, -2, -1, -2, -2, -1, -2, 0, -3, -3, 0, 2, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, 2, 2, 4, 5, 1, 0, 0, -2, -3, -2, -1, -1, 0, 0, -2, -2, -3, -5, 0, 0, 0, 1, -1, -1, 0, 0, 0, 0, 0, -1, 2, 1, 4, 5, 2, 1, -2, -1, -2, -2, -1, -1, -1, -2, -1, 0, -1, -2, 0, -1, 2, 0, 0, 0, -1, 0, 1, 0, 0, 0, 3, 3, 4, 1, 0, 1, -1, -1, -2, -2, -2, 0, 0, -3, -2, -2, -2, -3, 1, 0, 0, 0, 1, 0, 1, 0, 0, 2, 0, 0, 3, 0, 1, 3, 2, 0, 0, -1, -3, -3, 0, -1, 0, 0, 0, -2, -2, -4, 1, -1, 1, 1, 2, -1, 0, 0, 1, -1, 1, 1, 0, 1, 0, 3, 0, 0, 0, -1, -4, -2, -2, -3, 0, -3, -3, -1, -3, -2, -1, 1, 0, 0, -1, 1, 2, 3, -1, 0, 2, 2, 1, -1, 1, -1, -1, 0, 0, 0, -1, -2, -2, -3, 0, -1, -2, -2, 0, -3, 0, 0, 1, 2, 0, 1, 0, 2, 0, -1, 0, 1, -1, 0, 0, 0, 0, -2, -3, -2, 0, -3, 0, 0, -2, 0, -3, 0, -1, -2, 0, 0, 1, 1, 2, 0, 0, -1, 1, -1, -1, 2, -2, -1, -2, 0, 0, -1, -2, -2, 0, 0, -3, -3, -3, -1, -2, -3, -2, -3, 1, 1, 1, -1, 2, 1, 1, 0, 0, 1, 1, -1, -2, -2, 0, 0, 0, 0, -1, 0, 0, -3, 0, 0, -1, -1, -1, -2, -2, -1, 0, 0, 0, -1, 1, 2, -1, 1, 0, -2, -2, 0, -2, 0, 0, 0, -1, 0, 0, -2, 0, -2, -2, 0, -1, -1, -3, -2, 0, -3, 1, 1, 1, 0, -2, 1, 0, 0, -2, 0, 0, 0, -1, 0, -1, -2, -2, 0, -1, -1, -1, 0, -1, 0, -1, -1, -3, 0, -1, -2, -1, 1, -1, 0, 0, -1, 0, -1, -2, -1, 1, -2, -1, -2, -2, 0, 0, -2, -1, 0, -2, 0, -2, 0, -2, -2, -2, 0, -3, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, 0, 0, -1, -2, -1, -2, -1, -3, 0, -3, -2, -3, 0, -2, -2, 0, -1, -1, -1, -2, -2, 0, 0, -3, 0, -1, 0, -2, 0, 0, -1, 0, 0, -3, -2, -5, -4, -1, -1, -2, -3, 0, -4, -4, -1, -3, -2, -4, 0, 0, -4, 11, 8, 6, 7, 4, 3, 5, 2, 2, 1, 2, 1, 4, 4, 4, 3, 4, 3, 5, 2, 3, 0, 2, 1, -3, -3, -1, -2, -3, -2, 7, 9, 5, 5, 2, 4, 3, 2, 0, 0, 2, 2, 1, 2, 1, 1, 0, 1, 1, 3, 0, -1, 1, 0, -3, -4, -2, -3, -5, -6, 8, 7, 6, 1, 3, 1, 1, 1, -1, -1, -1, 1, 1, 0, 0, 2, 0, 3, 0, 0, -1, 0, 0, -3, -4, -2, -6, -5, -5, -4, 9, 6, 5, 0, 0, -1, 0, -2, -3, -4, -2, 0, 0, 0, 1, 4, 2, 4, 0, 2, -1, 1, 0, 0, -2, -2, -2, -4, -3, -3, 9, 4, 2, 2, -2, 0, 0, -3, -3, -4, -3, -1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 1, 1, 0, 0, -1, -2, -4, -6, 11, 5, 4, -1, -1, -4, -4, -4, -5, -4, 0, -2, 1, 0, 0, 1, 1, 0, -1, 0, 2, 0, 0, 0, 2, 0, 0, 0, -2, -3, 10, 7, 0, 0, -4, -4, -4, -5, -7, -6, -5, -2, -2, -1, -3, 0, -1, 0, 0, 2, 1, 3, 1, 3, 0, 0, 2, -2, -2, -3, 7, 5, 2, 0, -1, -3, -6, -7, -10, -10, -6, -7, -3, -3, -4, -3, 0, 1, 3, 2, 2, 3, 3, 2, 4, 2, 0, -1, -2, -3, 7, 5, 1, 0, 0, -2, -2, -5, -10, -7, -10, -10, -6, -7, -3, -3, -1, -1, 1, 7, 6, 5, 5, 3, 4, 2, 1, 1, -1, -3, 11, 7, 5, 3, 0, -1, -1, -5, -6, -8, -8, -9, -8, -6, -5, -5, -2, -2, 0, 4, 4, 2, 2, 4, 4, 3, 0, 2, 0, 0, 8, 8, 4, 3, 2, 0, 0, -4, -7, -7, -6, -7, -7, -6, -8, -9, -8, -5, -2, 3, 2, 2, 4, 3, 1, 3, 3, 3, -1, -2, 7, 7, 3, 1, 1, 0, -1, -2, -5, -7, -7, -7, -7, -6, -10, -7, -8, -7, -3, 2, 5, 3, 2, 2, 3, 2, 0, 1, -2, -2, 8, 4, 1, 1, 0, 2, -2, -3, -3, -8, -8, -5, -8, -5, -8, -9, -9, -9, -3, 0, 5, 6, 5, 2, 0, -1, 2, 0, 0, -1, 7, 4, 2, -1, 0, 2, 1, 0, -5, -7, -6, -6, -5, -8, -7, -11, -8, -5, -2, 1, 7, 5, 4, 3, 1, 1, 0, 0, 0, -1, 7, 4, 1, 2, 1, 1, 0, -2, -3, -8, -5, -6, -8, -9, -7, -7, -10, -4, 0, 3, 9, 10, 6, 3, 3, 2, 0, 1, -1, 0, 6, 3, 0, 1, 1, 0, 2, 1, -4, -6, -6, -7, -5, -8, -6, -8, -8, -6, 0, 4, 11, 12, 10, 8, 2, 4, 1, 0, -1, 0, 8, 6, 1, -1, 0, 0, 1, -1, -5, -3, -6, -8, -6, -8, -7, -10, -5, -5, -2, 5, 6, 10, 9, 5, 3, 3, 3, 1, -1, -2, 5, 3, 1, 2, 1, 0, -2, -4, -6, -6, -6, -7, -5, -5, -8, -9, -8, -8, -2, 4, 6, 9, 7, 7, 3, 3, 0, 0, -1, -4, 9, 3, 2, 2, 2, 1, -1, -2, -4, -4, -7, -5, -6, -5, -7, -10, -7, -8, -3, 1, 6, 7, 7, 5, 1, 1, 2, 0, -1, -1, 5, 5, 1, 3, 2, -1, -1, -2, -4, -9, -9, -10, -9, -9, -8, -7, -7, -4, -1, 0, 2, 4, 2, 2, 2, 1, 0, 1, -1, -4, 5, 5, 5, 0, 1, -3, -2, -5, -6, -9, -9, -8, -6, -7, -9, -5, -5, -3, -1, 0, 4, 2, 6, 4, 4, 2, 0, 2, 0, -4, 7, 5, 3, 1, -2, -2, -3, -4, -8, -9, -7, -10, -8, -7, -8, -8, -6, -3, 2, 2, 3, 5, 5, 5, 2, 1, 3, 1, 0, -3, 9, 3, 3, 0, 0, -3, -2, -3, -5, -3, -7, -7, -9, -8, -7, -5, -2, -1, 1, 2, 5, 4, 6, 4, 2, 4, 1, -2, 0, -4, 7, 6, 2, 0, -2, -5, -5, -4, -6, -5, -3, -5, -8, -7, -6, -4, -3, 0, 2, 0, 5, 3, 5, 1, 1, 3, 0, -1, -1, -3, 7, 7, 3, 0, 0, -3, -4, -4, -3, -2, -4, -3, -2, -2, -1, -2, 0, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, -3, -1, -6, 9, 6, 3, -1, -3, -2, -4, -1, -3, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -2, -3, 0, -1, -3, -6, 9, 7, 2, 0, 0, -1, -4, 0, -1, -2, 0, -1, 2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, -1, -1, -2, -3, -2, -4, -4, 9, 6, 2, 1, 0, 0, -3, 0, -2, -2, -1, 0, -1, 2, 1, 0, 2, 0, 1, 1, 1, -3, -1, -4, -3, -5, -5, -6, -6, -6, 11, 8, 4, 1, 0, 1, 1, -1, -4, -2, 0, 1, 0, 1, 0, 4, 1, 1, 0, 2, 0, -1, -1, -6, -6, -5, -3, -4, -5, -3, 10, 6, 5, 3, 3, 3, 1, 1, 0, 1, 1, 1, 0, 3, 2, 0, 2, 0, 0, 0, -2, -3, -3, -4, -5, -4, -4, -5, -3, -2, 6, 2, 4, 3, 1, 4, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -2, -2, -1, -3, -1, -4, -3, -2, -4, -3, 5, 2, 4, 0, 1, 0, -1, 1, 1, 1, -3, 0, 0, 0, -1, -1, -2, 0, -1, -1, -3, 0, -3, -3, -3, -1, -2, -4, -4, -1, 6, 2, 2, 2, 0, 1, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, 0, 0, -2, -1, -3, -2, 0, -1, -3, -1, -2, -4, -4, -3, 2, 3, 2, 0, 2, -1, 0, -1, 0, 0, -3, -3, 0, 0, 0, 0, 1, -1, 0, -2, -2, 0, -1, -3, -2, -1, -2, -5, -2, -6, 3, 3, 0, 0, 1, -1, 0, -2, 0, -2, -2, -3, -2, 0, 1, -1, -1, 0, 0, 1, 0, -1, 0, -1, -1, -1, -2, -3, -3, -1, 6, 3, 1, 0, 0, -1, 0, 0, -3, -2, -3, 0, -1, -2, -1, -1, -2, 0, 0, -2, -2, -2, 1, -2, -2, 0, -3, 0, -2, -2, 3, 4, 2, 1, -1, -2, 0, -2, -2, -2, -2, -2, -3, -1, -1, -2, -2, 0, 0, 1, 0, 0, 0, -1, -3, 0, -2, -1, -3, -4, 4, 2, 3, 0, -1, 0, -2, -3, -2, -3, -1, -2, -2, -4, -2, -3, -2, -1, 1, 0, 0, 1, 2, 0, 1, 1, 0, -3, -2, -4, 5, 2, 1, 0, 0, -1, -1, 0, -5, -6, -4, -4, -2, -3, -2, -2, -2, 1, 2, 2, 2, 0, 2, 2, 0, 0, -1, -2, -2, -1, 5, 5, 2, 0, 0, 1, -1, 0, -2, -4, -2, -6, -4, -3, -4, -1, -2, -3, -1, 1, 0, 2, 2, 0, 0, -1, 1, -2, 0, -4, 3, 4, 2, 2, 2, 2, 0, 0, 0, -1, -4, -5, -4, -4, -4, -5, -2, -3, 0, -1, 2, 1, 0, 0, -1, -1, 0, 1, -2, 0, 3, 4, 1, 2, 3, 0, 1, -1, -3, -4, -1, -5, -2, -2, -5, -5, -5, -2, -3, -1, 2, 0, 0, 0, -2, -1, -1, 0, -1, -3, 3, 2, 3, 2, 2, 2, -1, -1, 0, 0, -3, -3, 0, -4, -3, -4, -1, -4, -2, -1, 0, 1, 0, 1, 1, 0, 0, 0, -1, -3, 3, 2, 0, 0, 0, 0, 1, 0, 0, -2, -2, -4, -2, -4, -2, -1, -2, -1, -2, 0, 0, 2, 2, 1, 0, -2, -1, -1, -3, -1, 4, 3, 0, 1, 1, 0, 0, -2, -1, 0, -4, -4, -3, -1, -1, -2, -4, -1, 0, 0, 0, 3, 2, 3, 0, -1, 0, -2, -2, -2, 2, 1, 0, 0, -1, 1, 2, -1, 0, -4, -4, -3, -4, -2, -3, -3, 0, 0, 0, 1, 0, 2, 0, 3, 0, -2, 0, -1, 0, -2, 1, 0, 0, 0, 0, -1, 0, 1, -2, -1, -1, -4, 0, -4, -2, -1, -4, -2, -2, -2, 0, 0, 4, 0, 0, 0, 0, -2, -3, 0, 5, 4, 0, 2, 2, -1, 1, -1, -3, -3, 0, -3, -3, -1, -2, 0, -3, -2, -2, 1, 2, 3, 2, 1, 0, 1, -2, 0, -3, -2, 2, 3, 2, 1, 0, -1, 0, 1, 0, -1, -1, -3, -1, -3, -3, -5, -4, -4, -4, 0, 0, 0, 0, 1, 0, -1, 0, -2, 0, -2, 3, 3, 3, 1, 0, 1, 0, 0, 0, -2, -4, -2, -4, -1, -3, -1, -3, -1, -2, 0, 0, 0, 1, 1, 0, 0, 0, 0, -2, -3, 4, 1, 0, 1, 2, 0, -2, -2, -3, -5, -4, -2, -3, -3, -4, -2, -1, -1, 0, -1, 1, 2, 1, 0, -2, 0, -2, -2, -3, -2, 2, 0, 2, 2, 0, 0, -3, -3, -1, -4, -5, -1, -1, -5, -1, -4, -3, -3, -2, 1, 0, 0, 2, -1, -1, -1, 0, 0, -3, -1, 2, 2, 0, 1, 0, -2, 0, -3, -1, -1, -4, -3, -3, -5, -4, -5, -1, 0, -2, 0, 1, 0, 0, 0, 1, -1, -1, -3, -3, -1, 2, 3, 4, -1, 0, 0, -1, 0, -1, -4, -1, -3, -4, -3, -2, -2, -2, -2, -1, 0, -1, 0, 1, 1, 0, -1, -1, -1, -3, -4, 3, 2, 3, 0, 0, 1, 0, 0, 0, -2, -1, -2, 0, -3, -2, -2, -3, -2, 0, -1, 1, -1, 0, 0, 0, -1, -3, 0, -1, -4, 3, 3, 2, 0, 0, -2, -1, -2, -3, 0, -1, 0, -2, -3, -1, -1, -2, -1, 0, 0, -3, -2, -2, -3, 0, -2, 0, -2, -2, -5, 3, 1, 0, 1, 0, -2, -1, 0, -2, -2, 1, -1, 0, -1, -2, -1, 0, 0, -1, -2, 0, -2, 0, -4, 0, -2, -3, -4, -2, -1, 5, 1, 1, 1, 0, -3, 0, 0, -2, 0, 0, -2, -1, 0, -1, 0, -1, 0, 0, -1, -1, -2, 0, -3, -1, -5, -2, -1, -4, -3, 4, 3, 2, 0, 1, 1, -2, -1, 0, 0, -2, -1, -1, -1, 0, -1, 0, -3, -3, -1, -3, 0, -4, -5, -4, -4, -2, -5, -3, -4, 6, 3, 1, 2, 1, 1, -1, -2, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, -2, -3, -1, -4, -2, -1, -2, -3, -4, -5, -6, -6, -1, 0, -2, -1, 0, 1, 1, 0, 1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 1, -1, -1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, -2, 2, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 1, 1, 0, 0, 0, -1, -2, -1, -1, -1, 0, 0, 1, 0, 0, -1, 1, 0, 0, -1, 0, -1, -1, 0, 1, 1, 1, 0, 1, 0, 1, -1, -1, 1, 2, 0, -1, 0, 0, -1, 0, -1, 0, -1, -1, 0, 1, -1, -1, -1, -1, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 1, 0, 0, 1, 0, -1, 0, -1, 2, 0, 0, 0, -1, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 1, -1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 1, 0, 1, 0, 2, 0, 1, 0, 1, 0, -1, 1, -1, -1, 1, -1, 0, 0, 0, -1, -1, 0, 1, 0, 0, 1, 2, 0, 1, 2, -1, 1, -1, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 0, 0, -1, 0, 0, 0, -2, 0, 0, 1, 1, 1, -1, 1, 0, -1, -2, 0, -1, 0, 0, 0, 0, 1, 1, -1, 0, 1, 0, -1, 0, 1, 1, 0, 0, -1, 0, 1, -1, -1, 1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 1, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, 1, -1, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 1, -1, 0, 1, -1, -1, 0, 0, -1, 1, 0, 0, 0, -1, 2, 0, 0, 0, 0, 0, 0, -1, 1, -1, 1, -1, 0, 0, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 0, 2, 0, -1, 0, 0, 0, 1, 1, 1, 1, 0, -1, 0, 1, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, -1, 1, 0, -1, -1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, -1, 1, 1, -1, 1, 1, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 1, 2, 0, -1, 0, -1, 1, -1, -1, -1, 1, -2, 1, -2, -1, 0, -1, 1, 0, 1, 0, 0, 1, 1, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, -1, -1, -1, -1, 0, -1, 0, 0, 1, -1, 1, 0, -1, 0, 0, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, -1, 2, -1, -1, 0, 0, 1, 0, -1, -1, 1, 1, -1, 1, 0, 1, 1, -1, 1, 0, 0, -1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 2, 1, -1, 0, 1, -1, -1, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 0, -1, 1, 0, 0, 0, 1, 1, 1, 1, -1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 1, -1, 0, -1, -1, -1, 0, 1, 0, 1, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, 1, 0, 0, -1, 0, -1, 0, 0, 1, -1, 0, 0, 0, -1, 1, 0, -1, 0, 1, 2, 0, 1, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 1, 0, -1, -2, 2, 0, 0, 1, 0, -2, -2, -1, -1, -1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, -1, -1, -1, 0, -1, 1, -1, 1, -1, 1, -1, 1, -1, 1, -1, 1, -1, 0, 0, 0, 0, 1, -1, -1, 1, 0, 2, 0, 0, 1, 0, -2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, -1, 2, 0, 1, -1, 0, -1, 0, 0, 0, -2, 1, 0, 0, 1, 0, 0, 1, 0, 0, 1, -1, 1, 1, 1, -1, 0, 1, 1, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, -2, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, -1, -2, 0, -1, -1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 1, -1, 1, -1, -1, 2, 1, 0, 2, 2, 0, 1, 0, 0, 1, 1, 0, 1, -1, 0, 1, 0, 1, -2, -1, -1, -2, 0, 1, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, -1, 1, -1, 1, 0, 0, 0, 1, 1, 0, -1, 2, -1, 1, -1, 0, -1, -1, -1, 1, 0, 0, -1, 2, -1, 0, 1, -1, -1, 2, 0, 0, 0, 2, 0, 0, 0, -1, 2, 1, 1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, 0, -1, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 2, 1, -1, -1, 1, -1, -1, 1, 0, 2, -1, 0, -1, 0, 2, -1, -1, 0, 0, 1, -1, -1, 1, 0, -1, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, -1, 1, 0, 1, 1, 1, 0, 2, 3, 2, 2, 1, 0, 1, 3, 5, 5, 6, 3, 3, 4, 6, 6, 3, 5, 3, 3, 5, 4, 2, 2, 3, 2, 1, 2, 0, 0, 0, 1, 2, -1, 0, 1, 0, 0, 2, 5, 2, 4, 2, 4, 4, 4, 4, 3, 0, 2, 2, 0, 3, 4, 2, 1, 0, 1, 0, -1, -1, 0, -2, 0, 0, 0, 1, 1, 2, 1, 0, 3, 2, 1, 3, 2, 3, 2, 1, 0, 1, 0, 2, 1, 1, 0, 0, -2, -1, 0, -2, 0, 0, 0, 0, 1, -1, 0, 1, 0, 1, 3, 4, 1, 3, 2, 2, -1, 0, 2, 0, 1, 0, 0, 0, 1, 0, -1, -2, 0, -2, 0, 0, 0, -1, 2, 0, 1, -1, 0, 0, 1, 0, 2, 1, 0, -1, -1, 0, 1, 2, 2, 0, 1, 0, 2, 0, -2, -2, -3, 0, -3, 0, -2, 0, 1, 0, 3, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, -1, -3, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, 1, -2, -1, 1, 1, -1, -1, 1, 1, 2, 1, 1, 0, 3, 1, 0, -1, 1, 0, -3, -3, 0, -3, -2, -3, -1, -1, 0, 1, 0, 0, -1, -1, 1, -1, 0, 1, 1, 0, 1, 1, 0, 2, 3, 2, -1, 1, 1, -1, -1, -2, -1, -2, -1, -1, -2, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 3, 0, 2, 2, 3, 0, 1, 2, 1, 0, 0, -1, 0, 0, 1, -2, -2, -1, -1, -1, -1, 0, -3, 0, -2, -1, -1, 0, 0, -1, 0, 2, 1, 0, 0, 1, 1, 2, 0, 0, 0, -1, 0, 1, -1, -1, 0, 1, 2, 3, 1, 0, -1, -3, -4, -4, -3, -1, 0, 0, -1, 0, -1, 0, 3, 1, 1, 1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 3, 2, 4, 0, 0, 0, -3, -6, -5, -1, 0, -1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 2, 1, 1, 2, 3, 1, -1, -1, -3, -7, -7, -5, -2, 0, 0, 0, 2, 1, 0, 0, 2, -1, 1, 1, -1, -3, 0, 2, 0, 0, 2, 0, 2, 1, 3, 1, 0, -1, -3, -5, -5, -1, 1, 1, 2, 3, 3, 0, 1, -1, 1, 0, 0, 2, 0, 0, -3, -2, 2, 3, 2, 2, 1, 1, 2, 0, 0, 0, -5, -5, -4, 0, 3, 4, 7, 2, 2, 0, 0, 1, 2, 1, 1, 1, 0, 0, -3, 0, 1, 0, 3, 1, 1, 0, 2, 0, 0, -1, -2, -5, -4, 0, 2, 6, 4, 6, 4, 3, 0, 3, 2, 1, 1, 2, 0, 0, 0, 0, 0, 1, 0, 3, 3, 2, 3, 1, 0, 0, -3, -7, -5, -4, 1, 4, 4, 3, 2, 4, 2, 2, 1, -1, 2, 0, -1, 1, 0, -1, 2, 2, 2, 2, 0, 1, 1, 0, 2, 0, -2, -7, -9, -5, -1, 1, 4, 3, 2, 3, 2, 2, 0, 2, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 3, 3, 3, 2, 0, -3, -6, -7, -9, -2, 0, 1, 2, 4, 3, 0, 2, 1, 1, 1, 1, 2, 0, -1, 0, -2, 1, 0, 0, 3, 2, 1, 3, 1, 0, -3, -2, -7, -5, -2, -2, 1, 0, 1, 3, 0, 0, 0, 1, 1, 0, 2, 0, -1, -3, -3, -1, 0, 0, -1, 1, 0, 0, 1, 0, -3, -5, -6, -6, -3, -1, 2, 2, 2, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, -2, 0, 1, 2, 0, 1, 0, -1, 0, -3, -5, -4, -3, -1, 1, 1, 1, 2, 1, 3, 3, 1, 0, 3, 1, 0, 0, 2, 0, 0, -1, 0, 0, 1, 0, 1, 0, -2, 0, -3, -3, -3, 0, -2, 1, 0, 1, 4, 1, 2, 4, 2, 0, 0, 0, 0, 3, 0, 1, -2, 0, 0, -3, 0, -1, 1, 1, -2, -2, 0, 0, 0, -3, 0, 0, 1, 1, 2, 0, 3, 4, 3, 1, 2, 2, 0, 1, 0, 0, -1, -2, -2, 0, -2, -2, 1, 1, 0, 0, 0, 0, 0, -1, -1, 0, 0, -2, 1, 2, 2, 2, 0, 0, 2, 0, 0, 2, 0, 0, -2, 0, -2, 0, -2, 0, 0, 0, 1, -1, 2, 0, -2, -2, -2, -1, -3, 0, 0, 0, 2, 0, 2, 3, 1, 0, 0, 0, -1, -3, 0, 0, -2, -2, -1, -1, 0, 1, 1, 0, 1, 2, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 0, 1, 1, 1, 0, 0, -1, 0, 0, 0, -2, 0, -1, -1, 1, 0, 0, 0, 3, 2, 1, 2, 1, 0, -1, 0, -1, 0, 0, 2, 1, 2, 0, 0, 2, 0, -1, -1, 0, 2, 0, -2, -1, 1, 0, 2, 2, 0, 2, 2, 4, 1, 0, 1, 1, 0, -1, -1, 0, 0, 1, 0, 1, 3, 4, 0, -1, -1, 0, 0, 1, 2, 0, -1, 1, 0, 1, 2, 5, 3, 4, 4, 2, 3, 0, 0, 1, 1, 3, 0, 3, 2, 1, 2, -1, 2, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 2, 0, 0, 1, -1, 1, 2, 1, 1, -1, 2, 0, 0, 1, 1, 2, 1, 0, 2, 0, 0, 2, 0, 1, 0, 0, 0, -1, 1, -1, -1, 0, 0, -1, 0, 0, 0, 1, 1, 0, 0, 1, 0, 1, -1, -1, 0, 0, 2, -1, -1, 2, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 1, -1, 2, 2, 0, 3, 3, 1, 1, 2, -1, 1, 0, -1, -1, 0, -1, -1, -1, 1, 1, 0, 1, 0, 2, 0, 0, 1, 2, 0, -1, 0, 0, 0, 3, 2, 2, 2, 0, -1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 1, 2, 1, 1, 2, 0, 0, 0, 0, 1, 2, -1, 1, 2, 0, 1, 0, 0, 2, 2, 0, 0, -1, -1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 1, 0, -1, 0, -1, 1, -1, 1, 0, 1, 0, 0, 0, 2, 0, -2, 0, 0, 1, 1, 1, 0, -1, -1, 1, 1, -1, 1, -1, 0, -1, 0, -1, 2, 1, -1, 1, 2, 0, 0, -1, -1, 1, 2, 0, 2, 2, 2, 1, -1, 2, -2, 2, 0, 0, 0, -1, 1, 0, 1, 1, 0, -1, 1, -1, 2, 0, 0, -1, 0, 2, 1, 1, 0, 0, -1, 1, 1, -1, 0, 0, 0, 0, -1, 0, -1, -2, 2, 2, 2, 2, -1, 0, 0, 0, 2, 2, 0, 1, 0, 1, 1, 0, 2, 2, 0, 0, -1, 0, -1, 0, 1, 0, 1, 1, 0, -1, 0, 0, -1, 0, 2, -1, 0, -1, 0, 1, 2, 0, 1, 0, 0, 1, 0, -1, 1, -1, 0, -1, 1, 1, 2, -1, -1, 0, 1, 1, 2, 0, 1, 1, -1, 0, 0, 1, 2, 0, 0, 2, 0, 1, 2, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, -1, 2, 1, 0, 0, 0, 2, 0, -1, 0, 0, -1, 0, 2, 1, 1, 0, -1, 0, 0, 1, 0, 0, 0, -2, 0, 1, 1, 1, -2, -1, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 3, 0, 0, 1, -1, 1, 0, 1, 2, 1, 0, 1, -2, 0, 0, 0, -1, 1, 0, 0, 0, -1, 1, -1, 0, 0, 1, 0, 0, 2, 0, 0, 0, 0, 0, 2, 0, 1, 0, 0, -1, 1, 0, -1, -1, 1, -2, 0, 0, 0, 1, -1, 0, 2, 2, 1, 0, 2, 2, 0, 0, 0, 2, 0, 0, 0, 0, 1, 1, 1, 0, -1, -1, 1, -2, -1, -1, -1, 0, 0, 0, 0, 2, -1, 1, 0, 1, 0, 2, 2, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, -1, 1, -2, -1, 0, 1, -1, 1, 0, 0, 1, 0, 2, 0, 1, 0, 0, -1, 1, 2, 3, 1, 1, 0, 2, 3, 0, 0, 1, 1, 1, -2, 0, -1, 1, -1, 1, 0, 0, 0, 2, 0, 1, 2, 0, 1, 0, 3, 2, 0, 0, 1, 0, 2, 0, 0, 1, 2, -1, -1, -1, -2, -2, 0, -2, 1, 0, 0, -1, 1, -1, -1, 0, 1, 2, 1, 1, 1, 3, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, -2, 0, -2, -2, 1, 0, 1, -2, 0, 0, 0, 1, 0, 2, 0, 1, 1, 2, -1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 1, 0, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, -1, -1, 2, 0, 0, 0, 3, 2, 0, 1, 0, 0, 0, 1, 1, 2, -1, 0, 0, -1, 0, 0, 0, -1, -2, 1, 0, 0, 2, 2, 1, 2, 0, -1, 0, 2, 0, 0, 2, 0, -1, 2, 1, 0, 1, 0, 0, 2, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, -1, -1, 1, 0, 0, -2, 0, 1, -1, -2, -1, -1, 0, 0, -1, -1, 1, 2, 0, 2, 1, 0, -1, -1, 0, -1, 0, 2, 1, 1, 1, 1, 1, 0, 1, -1, 1, -2, -2, -1, 0, 1, -1, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, 1, 1, 0, 3, 1, 1, 0, 1, 0, 0, 1, 0, -2, 1, -1, 0, 0, -1, -1, 1, 0, 2, 1, 0, 0, 0, 2, -1, 0, 0, 2, 1, 1, 0, 0, -1, -1, 0, 0, 0, -1, -1, -1, -2, -1, 1, -1, -1, 0, 0, 1, -1, 0, 2, 0, 1, 0, 1, 0, 0, -1, 1, 0, 1, 1, -1, 0, 0, -1, 1, 1, 0, 1, 0, 0, 0, 0, 1, -1, 1, -1, 1, 1, -1, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 1, -1, 0, -1, 0, -1, 0, 0, -1, -1, 1, 0, 1, 1, -1, 0, 0, -1, 0, 0, 0, 1, 1, -1, 0, 1, 0, 1, 0, -1, -1, 2, -1, -2, 0, 1, -1, -1, 1, 0, 0, 0, -2, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, -2, 1, 1, -1, -1, 0, 0, -1, 0, 1, 0, -1, 2, 0, 0, 2, 2, 1, 1, 0, 0, 0, -2, 0, -2, -2, 1, -1, 0, 1, 0, -2, -1, -1, 1, 0, 1, 1, 2, 2, -1, 0, 0, 1, 1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, 0, -2, 1, -1, 0, 0, 0, 0, 2, 0, 0, 0, 2, 1, 1, 0, 1, 1, -1, -1, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 2, 0, 0, -2, -1, -2, -1, 1, 2, -1, 2, 2, 1, 2, 0, 2, 1, -1, 0, 0, 1, 0, 1, -1, -2, 0, -1, 1, 1, 1, -1, 0, 0, -2, 0, 0, -1, -1, 1, 0, 2, 0, 0, 0, -1, 2, -1, 1, 0, 0, 1, -1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, -1, -1, 0, 2, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, -2, -2, 0, 1, 1, 0, -1, 0, 1, 0, -1, 0, 0, 2, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, 0, -1, 0, -2, 0, -1, 1, 0, 1, -1, 2, 2, 2, 2, -1, 0, -1, -1, 1, 0, 0, -1, 0, -1, 1, 0, 0, 1, 0, 0, 0, 1, -2, 0, -1, 0, 0, 0, 0, 1, 1, 0, 1, -1, 0, 1, 1, 0, 0, 2, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 1, 1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 1, 1, 3, 1, 2, 1, 0, 0, -1, 2, 1, 0, 2, 2, 1, -1, -2, 0, 1, -2, 1, 0, -1, 0, -1, 0, 0, 2, 0, 2, 0, 2, 3, 3, 0, 2, 0, 0, 0, -1, 2, 0, 0, 2, -1, -2, 0, 0, 0, 0, 0, 1, 0, -2, 1, 0, 0, 0, 1, 0, 0, 3, 1, 1, 1, -1, -1, 0, 1, 0, -1, 0, 2, 2, 2, -2, 1, 0, -1, 0, -1, 0, 0, 0, 0, 1, 2, 1, 0, 0, 0, 1, 1, -1, 0, 0, 0, -1, 2, 1, 1, 0, 1, 0, 0, 0, 1, -1, 1, -1, -1, 0, 0, 0, -1, 1, 1, 0, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -2, 1, -1, 0, 1, 0, 0, -1, 0, 0, -1, -2, -2, 0, 2, 0, 0, 0, 3, 0, 1, 1, 1, 0, -2, 0, 0, 1, -1, -1, 0, 0, 0, -1, -1, -1, 0, -1, 1, 0, -1, -2, 1, 1, 1, 0, 1, 0, 2, 1, 1, 0, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 2, 0, 2, 0, 2, 1, 1, 0, 0, 0, 2, 0, 2, 0, 0, -2, -2, 1, -2, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, -1, 1, 0, 0, -1, 0, 0, 0, 1, 0, 2, 0, -1, 0, -2, -2, -1, 1, -1, 0, -1, 0, -2, 0, 1, 1, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 2, -2, 0, 0, 1, 1, 1, 0, -1, -1, 1, 1, 1, 0, 0, 0, 2, 2, 0, -1, 1, 1, 0, 0, 2, 0, 0, 0, -1, -1, 1, 1, 0, -1, 1, 1, -2, 0, -1, -1, -1, 2, 1, 0, 2, 0, 2, 1, 1, 0, 0, -1, -1, -1, 1, 0, -1, 1, 0, 0, -1, 0, 1, -2, 0, -2, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, 0, -1, 0, -1, 1, 0, -1, 0, 2, 0, 0, -1, 0, -2, 0, -2, 1, 1, -1, 1, -1, 0, 1, -1, 1, 1, -1, 1, 0, 2, 2, 0, 2, 1, 1, 1, 1, 1, 1, 2, 2, 1, -1, 1, -1, -1, -1, -2, -2, 0, -2, 0, -1, -1, -1, -1, 0, -1, 1, 2, 0, 0, 2, 2, 0, 1, 0, 0, 0, 2, 1, 1, 0, -2, -2, -2, -2, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 2, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 1, 0, -2, 0, 0, -1, 0, -2, -1, 0, -2, 1, 0, 0, -1, 0, 1, 1, 2, 0, 1, 0, 0, 1, -1, -1, 0, 1, 0, 1, -2, -1, -1, -2, 0, 0, -2, 1, 0, 0, -1, 1, 1, 1, 0, -1, -1, 1, 1, 0, 1, 0, 2, 0, 0, 0, -1, 1, 0, -1, -1, -1, -1, 0, -2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 2, 0, 0, 0, -1, 0, 0, -2, -2, 0, -2, 1, -1, -1, -2, -1, 0, -1, -2, -2, 0, 0, -1, 0, 0, -1, -2, 0, -2, -2, 0, 0, -2, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, -2, 0, 0, -2, -1, -1, 0, 0, 0, 0, -1, 0, -1, -1, 1, -1, 1, 0, 1, 2, 0, 0, 1, 0, 0, 1, 1, 0, 3, 1, 0, 3, 5, 3, 1, 1, 2, 4, 2, 0, 0, 2, 2, 1, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, -2, 0, 0, 2, 0, 2, 2, 1, 4, 3, 2, 2, 1, 1, 4, 0, 2, 1, 3, 0, 1, 3, -1, 0, 0, -1, 0, -2, -3, 0, 0, 0, 1, 2, 0, 1, 2, 2, 3, 2, 4, 3, 3, 1, 2, 1, 3, 0, 3, 3, 1, 4, -1, 0, -1, -1, -1, 0, 0, -2, -1, -1, 1, 1, 0, 1, 2, 0, 0, 1, 3, 3, 1, 3, 3, 3, 3, 3, 0, 2, 0, 4, 0, -2, -1, -1, 0, -1, -3, -1, -2, 0, -1, 0, -1, -1, 1, 1, 1, 0, 0, 0, 1, 2, 2, 2, 3, 1, 0, 3, 0, 4, 0, 0, 0, -2, 0, -1, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, 0, 2, 3, 1, 3, 0, 3, 2, 3, 1, 0, 0, 0, 4, 0, 0, -1, 0, -2, -3, -4, -4, -3, -5, -3, -4, -3, -3, -1, 0, -1, 1, 1, 1, 1, 4, 1, 3, 2, 2, 0, 0, 0, 3, -1, -1, 1, 0, -3, -3, -2, -2, -2, -5, -2, -4, -3, -3, -2, -2, 0, 2, 1, 0, 1, 3, 1, 1, 1, 1, 0, 1, 0, 2, 1, 0, -2, 0, 0, -3, -2, -4, -5, -5, -2, -3, -4, -2, -5, -1, 0, 0, 0, 1, 2, 0, 3, 0, 0, 0, 0, 1, 3, 0, 0, 2, 1, -2, -2, -1, -1, -3, -4, -5, -1, -2, -4, -4, -5, -2, -1, 0, 2, 1, 2, 1, 1, 2, 1, 4, 0, 3, 1, 4, 0, 0, 0, -1, -2, 0, -3, -2, -3, -4, -2, -5, -3, -6, -4, -5, 0, -1, 0, 0, 1, 1, 0, 3, 2, 0, 0, 0, 2, 2, 0, -2, 0, 1, 0, -3, -2, -3, -3, -4, -3, -5, -5, -5, -3, -5, 0, 1, 0, 3, 2, 3, 4, 3, 2, 1, 4, 2, 3, 2, 0, 0, 0, 1, -1, 0, -1, -4, -3, -4, -4, -5, -4, -4, -4, -2, -3, 0, 2, 5, 2, 5, 4, 5, 2, 3, 3, 2, 4, 5, 2, -1, 1, 1, -1, -2, -1, -4, -4, -3, -5, -6, -4, -5, -2, -3, -1, 1, 5, 4, 6, 4, 3, 3, 4, 5, 2, 3, 4, 2, 0, -1, -1, 0, 1, -1, -1, -1, -5, -5, -5, -3, -3, -3, -3, -3, 0, 0, 2, 5, 7, 6, 3, 1, 4, 1, 1, 1, 2, 4, -1, 0, 0, 1, 0, 0, -2, -2, -3, -3, -3, -2, -3, -3, -2, -3, -3, 0, 1, 2, 2, 4, 2, 5, 4, 4, 2, 4, 3, 5, 2, 0, 1, -1, 0, 0, -2, -2, -4, -6, -3, -6, -3, -7, -3, -5, 0, 3, 2, 1, 3, 3, 2, 1, 2, 2, 4, 3, 3, 2, -1, 0, 0, 0, 0, -2, 0, -1, -5, -4, -6, -3, -6, -4, -5, -5, -2, 3, 1, 0, 4, 5, 4, 3, 3, 4, 4, 2, 1, 4, 2, 1, 0, -2, -2, -2, -3, -4, -3, -5, -4, -6, -4, -6, -3, -5, -2, 0, 1, 3, 1, 3, 1, 1, 3, 3, 4, 0, 1, 5, 1, 2, 0, -1, -2, -1, -3, -2, -4, -3, -5, -5, -4, -5, -3, -4, 0, 1, 2, 1, 4, 2, 2, 1, 1, 2, 3, 4, 3, 3, 2, 2, -1, -1, -2, -2, -2, -5, -4, -5, -3, -7, -3, -4, -2, -3, 1, 3, 1, 3, 2, 2, 3, 4, 1, 2, 1, 3, 1, 5, 2, 1, 0, 0, -2, -1, -3, -5, -4, -6, -5, -4, -1, -1, -1, 0, 1, 2, 2, 2, 1, 1, 2, 3, 2, 2, 3, 0, 2, 1, 1, 0, -1, -2, 0, 0, -1, -1, -4, -1, -4, -4, -2, -1, -3, 0, -1, 2, 2, 1, 2, 1, 3, 0, 0, 3, 1, 0, 3, 4, 1, 0, 0, 0, -1, 0, 0, -2, -2, 0, -3, -1, 0, 0, -1, 0, -1, 0, 0, 1, 0, 3, 1, 3, 2, 2, 3, 2, 0, 3, 1, 0, -1, -2, 0, -1, 0, -2, -2, 0, 0, -1, 1, 0, 0, -1, 0, 0, 0, 1, 2, 0, 1, 0, 0, 0, 3, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, -2, -3, 0, 0, -1, -1, -1, 2, 0, 1, 0, 0, 0, 3, 2, 0, 0, 1, 0, 1, 1, 4, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, -2, -1, 1, 0, 0, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 3, 0, 0, 1, 1, 1, 1, 0, -2, -2, -1, 0, 0, 0, 2, 2, 0, 1, 2, 0, 2, 0, 0, 1, 1, 0, 3, 1, 0, 2, 2, 2, 0, 2, 0, 0, 0, -1, 0, -1, 0, 1, 0, 1, 1, 0, 4, 3, 4, 2, 0, 1, 0, 2, 2, 0, 0, 1, 3, 3, 3, 2, 0, 0, 2, 2, 1, 0, 0, 1, 1, 1, 3, 2, 3, 5, 3, 3, 3, 4, 3, 3, 3, 5, 5, 1, 4, 4, 1, 1, 5, -7, -8, -6, -3, -3, 0, 1, -2, 1, 1, 1, 3, 6, 8, 12, 12, 12, 11, 11, 12, 13, 13, 14, 13, 14, 13, 13, 13, 14, 15, -5, -6, -7, -2, -2, -2, -2, 0, -2, 0, 2, 1, 2, 4, 8, 5, 8, 7, 9, 8, 10, 10, 10, 8, 8, 11, 9, 10, 12, 14, -5, -5, -3, -2, -1, -3, -1, -2, -3, 0, 1, 1, 3, 3, 3, 4, 6, 4, 4, 6, 7, 7, 7, 5, 7, 9, 7, 9, 11, 13, -6, -8, -4, -4, -1, -3, -2, -4, -5, -3, -1, 2, 2, 4, 2, 5, 3, 2, 3, 3, 5, 2, 3, 5, 6, 5, 8, 9, 7, 13, -7, -8, -4, -6, -4, -1, -4, -4, -2, -2, 0, 2, 0, 0, 2, 3, 2, 0, 3, 1, 2, 1, 1, 1, 6, 6, 7, 4, 9, 9, -7, -8, -5, -5, -4, -3, -2, -2, -2, -1, 0, 2, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 2, 5, 8, 7, 7, 6, 8, -5, -7, -9, -6, -4, -3, -2, -2, -1, 1, 2, 0, 1, -1, 1, -1, 0, -1, 1, 0, 1, -1, 0, 0, 4, 4, 6, 7, 6, 10, -7, -10, -10, -7, -5, -2, -3, 0, 0, 1, 1, 2, 1, 1, 0, -3, -3, -3, -3, 0, -2, 2, 0, 3, 4, 5, 4, 5, 5, 11, -8, -9, -7, -9, -8, -4, -3, 0, 1, 2, 1, 3, 1, 0, 0, 0, -1, -2, 0, 0, 0, 0, 1, 2, 4, 6, 5, 3, 7, 8, -9, -9, -8, -6, -5, -4, -5, -3, 1, 1, 0, 1, 0, 0, -3, 0, -4, -4, -1, 0, -3, 0, 0, 0, 3, 4, 2, 4, 5, 7, -8, -7, -5, -6, -4, -5, -1, -1, 1, 2, 3, 3, 2, 1, -2, -2, -4, -3, -5, -2, 0, 0, 0, 3, 1, 6, 3, 4, 5, 9, -7, -7, -7, -5, -4, -2, -2, 0, 1, 4, 4, 4, 1, 1, 1, -1, -6, -4, -3, -2, 0, 0, 0, 2, 4, 3, 4, 4, 4, 6, -6, -4, -5, -3, -2, 0, -3, -1, 2, 1, 4, 4, 4, 2, 1, -4, -7, -3, -4, -1, 0, 2, 1, 3, 4, 4, 4, 4, 4, 9, -8, -6, -5, -4, -2, 0, -2, 0, 0, 1, 3, 5, 3, 4, 0, -3, -4, -6, 0, 1, 2, 4, 3, 3, 6, 3, 6, 5, 7, 8, -8, -8, -3, -5, 0, -2, -1, 0, 2, 4, 3, 4, 1, 1, 0, 0, -6, -1, 0, 3, 6, 6, 2, 5, 6, 5, 6, 7, 5, 11, -5, -6, -6, -4, -1, -1, 0, 0, 1, 3, 3, 0, 3, 0, 0, -3, -4, -2, -2, 1, 7, 5, 6, 4, 7, 6, 6, 7, 9, 11, -6, -7, -6, -5, -1, -1, -1, 1, 1, 2, 4, 3, 4, 2, 0, -3, -5, -6, -1, 1, 4, 7, 5, 5, 6, 5, 4, 4, 8, 11, -4, -7, -4, -4, -5, -3, -2, 1, 2, 3, 3, 4, 5, 2, 0, -6, -7, -6, -4, 0, 4, 6, 8, 7, 6, 6, 6, 5, 4, 9, -5, -5, -6, -4, -4, -3, -2, 1, 1, 5, 6, 4, 2, 0, -3, -6, -9, -4, -2, 0, 3, 4, 6, 6, 3, 6, 5, 3, 7, 8, -4, -3, -6, -3, -3, -3, -1, 0, 4, 3, 6, 4, 1, 0, 0, -4, -8, -3, -4, -2, 0, 5, 7, 4, 6, 2, 3, 6, 4, 10, -5, -3, -4, -6, -4, -2, -2, 0, 3, 5, 5, 4, 2, 0, -1, -2, -4, -2, -2, 0, 3, 5, 6, 6, 5, 4, 4, 3, 7, 8, -4, -3, -4, -8, -4, -1, 0, 0, 3, 5, 1, 3, 3, -1, -2, -2, 0, -2, -2, 0, 3, 4, 6, 3, 4, 4, 5, 5, 8, 11, -4, -7, -4, -4, -5, -4, -3, 0, 1, 0, 0, 0, 0, 1, 0, 0, -3, 1, 0, 2, 2, 5, 3, 6, 3, 3, 6, 7, 6, 8, -3, -5, -7, -3, -3, -1, 0, 0, -1, 0, 2, -2, 0, 0, 1, 0, 0, -2, 0, 1, 3, 1, 5, 5, 4, 4, 3, 3, 6, 8, -5, -7, -4, -4, -5, -4, -3, -1, 0, -2, 0, 0, 1, 2, 0, 0, -1, -2, 0, 0, 1, 0, 2, 5, 7, 4, 7, 7, 5, 9, -4, -5, -5, -2, -2, -2, -1, -3, -3, -1, 0, 0, 1, 0, 2, 0, -2, -3, 0, -1, 0, 2, 3, 6, 6, 5, 5, 5, 9, 10, -3, -4, -4, -2, -2, -1, -3, -2, -2, 0, -1, 0, 3, 0, 0, 0, -1, 1, 1, 2, 2, 4, 4, 7, 7, 5, 9, 7, 9, 9, -7, -5, -5, -4, -1, -3, -2, 0, 0, -1, 2, 3, 4, 4, 3, 3, 4, 1, 3, 1, 1, 3, 7, 8, 9, 8, 9, 9, 8, 12, -4, -6, -5, -1, -2, -2, -3, -2, 0, -2, 2, 5, 4, 3, 5, 6, 6, 4, 4, 6, 6, 8, 8, 9, 10, 9, 10, 10, 12, 10, -6, -5, -5, -2, 0, 0, 0, 1, 0, 0, 1, 2, 7, 7, 8, 9, 7, 7, 10, 9, 8, 10, 10, 11, 12, 13, 10, 12, 11, 10, 1, 0, 0, 0, 0, 1, -1, 0, -1, 1, 0, 0, 0, -1, 2, 0, 0, 1, 1, 1, -1, 2, 1, -2, -1, 1, 0, -1, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, -1, -1, 0, 0, 1, -1, -1, 0, 0, 0, 0, -1, -2, 1, 1, 0, 1, 0, 0, 0, 2, 1, 0, 1, 1, 1, 0, 0, -1, 1, 0, 2, 0, -1, 0, 1, -1, 0, 0, -1, 0, -1, -2, -1, -1, 0, -1, -1, 1, 0, 0, 1, -1, 0, -1, 0, 0, 0, -1, 1, 0, 1, -1, 0, -1, -1, 1, 0, 0, 1, 0, 1, 1, -1, 0, 0, 2, 0, -1, 1, 0, -1, 1, 0, 0, -1, 1, -1, 1, 1, -1, 0, 0, 1, 1, -1, 1, 0, 0, 0, -1, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, -1, -1, 0, 0, -1, 1, 0, 0, -1, 2, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, -1, -1, 0, 1, 1, -1, -2, -1, 0, 2, 0, 1, 1, 1, 0, 2, 0, 0, 0, -2, -1, 0, 0, 2, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, 1, 0, 1, -1, 0, 0, -1, 0, -1, 1, -1, 1, 0, 0, -1, 0, 1, -1, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, 2, -1, -2, -1, 0, 0, -1, 1, -1, 0, -1, 0, 0, -2, 1, -1, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 2, 1, 1, -1, -1, -2, 1, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, 0, -2, 1, -1, 1, -1, 0, 0, 2, 0, 1, 0, 1, 1, -1, 1, 0, 1, -1, -2, 0, -1, 0, 1, 1, -1, 1, -1, -1, -1, 0, -1, 0, 0, 0, -1, -1, -1, 0, -1, -1, 1, -1, 0, 1, 0, 0, -1, 0, 1, -1, -1, 0, 1, 0, 1, 2, -1, 0, 0, 1, -1, 1, 1, 1, 0, 1, -1, 0, -1, 2, 0, 0, 0, 0, -1, 0, -1, 1, 0, -1, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, 1, 0, 0, -1, 1, 1, -2, -1, 0, 1, 1, 2, 0, 0, -2, 0, -1, 0, 0, 0, 0, -1, -1, 1, 0, -1, 0, 0, 1, 2, 0, 0, 0, 1, -1, -1, 0, 2, 0, 1, 0, 0, 0, 0, -1, 0, 0, 2, 1, -1, 0, 0, 0, 0, 0, -1, 1, 1, -1, 0, -1, 2, 1, 0, 1, -1, 0, 1, 0, -2, 1, 1, 0, -1, 0, 0, -1, 0, 0, 0, 2, 0, 0, 1, 0, -1, -1, 1, -1, 0, 0, 2, 0, 2, 1, 0, 0, 0, 2, 0, 1, -1, 0, 0, -1, 0, -2, 1, 0, 1, 0, -1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 1, -1, 0, 0, -1, -1, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 1, -1, 1, 1, 1, 0, 1, 1, 0, 1, -1, 0, 0, -1, -1, 1, 1, -1, 0, 0, 0, -1, 2, 0, 0, -1, -1, 0, 0, 1, 0, 1, 1, 0, -1, 1, -1, 0, 1, 0, 1, 1, -1, -2, -1, 1, 0, 0, 0, 1, 1, 0, 2, 1, 0, 1, 0, 0, 1, 1, -1, 0, 0, 1, -2, -1, 0, -1, -1, 0, 1, -1, 0, 1, -1, 1, 0, 2, 0, 0, 0, 1, 1, 1, 0, -1, 0, -1, 0, 2, -1, 0, 0, -1, 1, -1, 0, -1, 0, -2, 1, 0, 0, 1, 0, -1, -1, 1, 2, 0, 0, -1, 0, -1, 2, -2, 1, 0, -1, 0, 1, -1, 0, 0, 1, 0, -1, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, -1, -1, 2, 2, 2, -1, 1, 0, 0, 0, 0, 0, 0, 2, -1, 1, 0, -1, 0, -1, 1, 0, 0, 1, -1, 0, 0, -1, 0, -1, -1, 0, -1, 2, -1, -1, 0, 0, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, -2, 1, -1, -1, 1, -1, 0, 1, -1, 0, 1, 1, 0, 0, 0, 2, 2, 0, 1, 0, -1, 0, 2, 1, -1, 0, -1, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 2, 0, 1, 0, 0, 0, -1, 1, 0, 1, -1, 0, 0, 0, 1, 1, -1, 0, -1, 0, 1, 1, -1, 2, 2, 1, 1, 0, 0, 1, -1, -1, 0, 0, -1, 1, 1, 1, -1, -1, 1, -1, 0, 1, 0, -1, 0, 0, 0, -1, 2, 0, 1, 0, 0, 0, 1, -1, 2, 0, -1, 2, 0, 1, 1, 2, -1, 0, 0, 0, 1, 1, 0, 1, -1, -1, 2, 0, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 1, 1, 0, 1, 0, 0, 0, 0, -1, 1, 0, -2, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0, 0, 1, 0, -1, -1, 1, -1, 1, 1, 0, 1, 0, 1, 0, -1, 0, 0, -1, 1, 2, 0, 0, 0, 0, -1, 1, 0, 1, 0, 1, 0, 1, 0, -1, 1, 0, 0, 2, 0, 0, -2, 1, 0, 1, 2, 0, 0, 1, -1, -1, -1, 1, 2, 1, 0, -1, -1, -1, -1, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, 0, 0, -1, -1, 0, -1, 1, 1, -1, -1, 1, 0, 0, -1, 0, 1, 0, -1, 1, 1, -1, 0, 0, 0, 0, 1, 1, -1, 0, 1, 0, 0, 0, -1, 1, -1, 0, 2, 0, 1, 0, -1, 1, 1, -1, 0, 0, 0, 0, -1, 1, -1, 0, -1, 0, 1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, -1, -1, 1, 0, 1, 1, -1, 0, -1, 1, -1, -1, -1, 0, -1, 1, 1, 0, 0, -1, 2, 0, 0, -1, -1, -1, 1, 0, -1, 0, 0, -1, 0, -1, -1, 0, 1, 0, 1, 0, -2, 1, 1, -1, -2, -1, 0, 1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 0, 0, -1, -1, 0, 1, -1, 1, 1, 0, -1, -1, 0, 0, 0, 1, 2, 2, -1, 0, -1, 0, -1, 1, 2, 0, 0, 0, 1, -1, -1, -1, 1, 1, 1, -2, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 1, -1, 0, 1, -1, -1, 1, 0, -1, 0, 0, -1, 1, 0, 0, -1, -1, -1, 1, 0, 0, -1, 0, 0, 0, 0, -1, -1, 0, 0, -1, 0, 1, 0, 1, 2, 0, -1, 0, -1, 1, -1, -1, 0, 0, 1, -2, -2, 0, 1, 0, 1, 1, 1, 0, 0, -1, 1, 0, -1, -1, 0, 0, 2, 0, -1, 1, 1, 0, 0, 0, 1, -1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 2, 1, 0, 0, 0, -1, 1, 1, 0, 0, -1, -1, 1, 1, 0, 1, -2, 0, -2, 0, 0, 0, -1, 0, 1, 0, 1, 0, 2, 0, 0, 1, -1, -1, -1, -1, 0, 0, -1, 1, 1, 0, 0, -1, 0, 0, 0, -1, -1, 0, -2, 1, 0, 0, 0, -1, -1, 1, -1, -1, 0, 0, 0, 0, 1, 0, -2, -1, 1, 1, 1, 0, 0, 0, 2, -1, 0, 0, 1, 0, -1, -1, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -2, 1, -1, -1, 0, 0, 0, 1, 0, -2, 1, -1, 0, 1, 2, 2, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 0, 0, 1, -1, 0, 1, -1, -1, -1, 0, 1, -1, -1, 0, 0, 1, 1, -1, 1, 0, 0, 2, 0, 0, -1, 0, 0, 1, 1, -1, -2, -2, 0, 1, 1, 0, -1, -2, -1, 0, 0, 0, -1, 1, -2, 1, 2, 0, 0, 1, -1, 1, 0, 1, 0, 0, 0, 2, 0, -1, 1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, -2, 0, 0, -1, 0, 0, 1, 0, 1, 0, -1, -1, 2, 1, 0, 0, -1, 2, 0, 0, 0, -2, 1, -2, 0, 0, -1, 0, 1, 1, 0, 1, 0, 1, -1, -1, 0, 0, -1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 2, 0, -1, -1, 2, -1, 0, 1, 1, 1, 0, 0, 0, 1, -1, 0, 0, 2, -1, 0, 0, -1, -1, 0, -1, 0, 1, 0, 1, 0, 1, -2, -1, 0, 0, -1, 2, 2, -1, 0, -1, 0, -1, 1, 1, -1, -1, 1, -1, -1, 1, 0, 0, 0, -1, 1, 1, 0, 0, 1, 1, -1, 2, 0, 1, 0, 1, 0, 0, -2, 0, 1, 0, 1, 0, 0, -1, 0, 1, -1, 0, 0, 1, 0, 1, 1, 0, 0, -1, -1, 0, -2, 1, 1, -1, -1, -1, -1, 1, -1, -2, 0, 1, 1, 1, -1, 1, 0, 0, 1, -2, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, -1, 0, -1, 1, 1, 0, -1, 2, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 1, 0, 0, 0, -1, -1, 0, 2, -2, -2, -1, -1, 1, 0, -1, -1, -1, 1, 1, 1, -1, -1, 1, 0, 1, 1, 1, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, -1, 1, -1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 0, 1, 0, 1, 0, -1, 1, -1, 1, -1, 1, -2, 1, 0, -1, -1, 9, 4, 4, 4, 2, 3, 3, 1, 1, 3, 4, 3, 7, 7, 8, 10, 8, 8, 7, 9, 5, 5, 5, 2, 2, 0, 0, 2, 2, 2, 6, 3, 2, 1, 1, 3, 2, 0, -1, 0, 0, 3, 2, 7, 4, 8, 6, 4, 5, 2, 3, 2, 0, 1, 1, -2, 0, 1, 0, 1, 6, 3, 0, 1, 0, 2, -2, -3, -3, -2, 0, 4, 3, 4, 5, 5, 4, 6, 5, 2, 0, 0, -1, 1, -1, -3, -2, -2, -2, -2, 4, 3, 0, -2, 0, -3, -4, -4, -2, 0, 0, 3, 1, 2, 4, 6, 6, 2, 3, 2, 3, 0, 0, -1, -1, 0, 0, -3, 0, 0, 6, 2, -2, -1, -2, -4, -3, -5, -2, 0, 2, 2, 2, 1, 4, 3, 4, 3, 2, 0, 0, 2, 2, 0, 1, 3, -1, -2, -1, 2, 3, -2, -1, -5, -3, -4, -6, -7, -3, -2, 0, 1, 1, 1, 0, 0, 2, 2, 1, 2, 0, 2, 1, 2, 3, 2, 0, 0, 0, 2, 2, 1, -4, -2, -4, -6, -8, -5, -5, -3, -1, -1, -1, 0, -1, 0, 1, 0, 0, 2, 3, 4, 2, 1, 5, 2, 2, 0, -2, 2, 4, 0, -3, -2, -4, -5, -5, -6, -4, -6, -4, -6, -5, -4, -2, -1, -1, 0, 4, 5, 6, 7, 2, 6, 6, 4, 5, 1, 1, 0, 3, -1, -2, -2, -1, -3, -6, -7, -6, -8, -8, -8, -6, -3, -5, -5, -2, 2, 1, 5, 6, 4, 6, 3, 5, 3, 5, 3, 0, 1, 5, 0, 0, -1, -3, -1, -3, -3, -4, -6, -4, -6, -5, -6, -7, -5, -5, -3, 0, 4, 1, 3, 3, 2, 1, 2, 4, 3, 0, 0, 2, 2, -1, -2, -1, 1, 0, 0, -3, -4, -4, -4, -5, -6, -9, -8, -9, -7, -1, 1, 2, 4, 0, 2, 1, 3, 2, 0, 0, 2, 2, 0, -3, 0, 0, 1, 0, 1, 1, -1, -3, -1, 0, -5, -7, -12, -13, -10, -4, 2, 2, 3, 2, 2, 0, 3, 1, -1, -1, 2, 3, 0, -3, -1, 0, 0, 3, 1, 0, -4, -1, -2, 0, -8, -10, -15, -12, -7, -2, 1, 6, 8, 2, 2, 0, 0, 1, 0, 0, 0, 2, 0, -2, -3, 0, 4, 3, 2, 0, -2, -2, 0, -2, -6, -10, -13, -14, -9, 0, 7, 11, 9, 9, 5, 3, 0, 0, 1, -1, 2, 1, -2, -3, -2, 0, 4, 1, 0, -1, -1, 0, -1, -2, -6, -9, -12, -10, -5, 2, 11, 13, 15, 9, 4, 2, 1, 4, 0, 2, 0, 0, -3, -2, -1, 1, 1, 4, 0, 0, 0, 0, 0, -3, -3, -10, -11, -13, -6, 4, 11, 16, 15, 12, 8, 4, 3, 1, 1, 0, 3, 1, 0, -3, -3, 0, 1, 1, 0, 0, 1, 0, 0, -2, -5, -10, -12, -12, -8, 0, 7, 15, 13, 10, 8, 3, 2, 0, 0, -1, 0, 2, 0, -2, -1, 2, 3, 0, 0, 0, 1, 0, -3, -1, -6, -11, -12, -14, -11, 1, 7, 8, 12, 10, 7, 2, 1, 1, 0, 0, 2, 4, 1, 0, 1, 2, 2, 0, 0, 0, -3, 0, -3, -5, -7, -8, -11, -13, -7, -1, 2, 5, 7, 5, 5, 2, 0, 0, -2, 0, 2, 6, 1, 0, 0, 0, 0, 0, -2, -2, -1, -2, -4, -7, -7, -11, -11, -13, -7, -2, 2, 5, 5, 3, 4, 2, 0, 0, 1, -1, 1, 2, 2, 0, -4, -1, -4, -4, -3, -2, -2, -4, -4, -6, -8, -8, -11, -8, -2, -1, 5, 5, 4, 4, 6, 1, 2, 1, 0, 0, 0, 4, 4, -1, -3, -1, -4, -1, -1, -5, -3, -5, -7, -7, -9, -8, -8, -3, -1, 4, 3, 6, 6, 7, 6, 5, 2, 0, 2, 0, 0, 7, 3, 0, -2, -2, -3, -5, -5, -4, -4, -7, -7, -10, -5, -4, -2, -2, -1, 1, 5, 6, 8, 8, 5, 5, 1, 0, 0, 0, 1, 5, 0, -4, -5, -2, -5, -5, -4, -3, -3, -1, -5, -3, -2, -4, 0, -3, 0, 0, 1, 1, 4, 4, 3, 3, 2, 0, 1, 0, 0, 4, 1, -3, -2, -5, -4, -4, -2, -3, -2, -1, 0, -1, -2, -2, -1, 0, -3, -1, -2, 1, 0, 4, 2, 3, 1, -1, -1, -1, 1, 5, 0, -1, 0, -3, -2, -4, -2, -4, 1, 1, 1, 2, 3, 0, 0, -3, -3, -2, 0, -1, 1, 2, -1, 1, 0, 0, -1, 0, -1, 5, 0, -2, -1, -1, -4, -5, -3, -2, 0, 0, 0, 1, 2, 3, 0, 0, 0, -1, -2, 0, -1, 0, -3, -3, -1, 0, -3, -1, 0, 3, 1, 0, 0, 0, -2, -4, -2, -3, 0, 0, 0, 1, 3, 4, 3, 1, 3, 1, 0, 0, -1, -2, -4, -2, -3, -2, -3, 0, 1, 6, 5, 1, 0, 3, 0, 0, -3, -4, 0, 0, 0, 3, 5, 7, 5, 2, 2, 2, 2, 0, -3, -3, -1, 0, 0, 0, -1, 1, 1, 10, 7, 4, 3, 2, 2, 2, 2, 0, -1, 0, 2, 3, 7, 8, 8, 7, 5, 6, 5, 1, 3, 1, 1, 0, 0, 0, 2, 2, 2, 2, 3, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -2, -3, -3, -1, -1, 4, 1, 1, 0, -1, 0, -1, -2, 0, -3, -2, 0, 0, 0, 2, 2, 1, 0, 0, 0, 1, 0, -3, 0, -1, -2, -2, -2, 0, -1, 2, 1, 0, 1, -1, 1, -1, -1, 0, -1, 0, -1, -1, 1, 0, 0, 1, 1, -1, 1, -1, -1, 0, 0, -3, -3, -2, -1, -3, -4, 0, 2, 0, 1, 0, -3, 0, -2, 0, -1, 0, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, -2, 0, -2, 0, -1, 0, -3, 2, -1, 1, -2, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, 1, -1, -1, -1, -1, 0, -2, -1, -1, 0, 0, -2, -3, -2, -3, 3, 0, -2, -1, 0, -1, 0, -1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 0, -1, 1, 1, 0, -1, -2, -1, -2, -1, -1, 3, 2, 0, 0, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, -1, -1, 1, -1, -1, -1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 0, 3, 1, 0, -1, -1, -2, 0, 0, -2, -1, -1, -2, 0, 0, 0, -1, 0, 2, -1, 0, 1, 1, 2, -1, -1, -1, 0, 0, 0, -2, 1, 3, -1, -1, 1, 0, 0, 0, 0, -3, -2, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 1, -2, 1, 0, -3, 1, 1, 0, 1, -1, -1, 0, -1, -2, 0, -1, 0, 1, 0, -1, -2, 0, -1, -1, 2, 0, -1, -2, -1, -1, 1, 1, -2, -1, 0, 3, 1, 0, 0, 2, 1, 0, -1, -1, 0, -2, 0, 0, 0, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, -1, 0, 0, 0, -2, 0, 0, 0, 0, 1, -1, 1, -1, 0, -1, 1, 0, 0, 1, -2, -1, -2, -2, -1, 0, 1, 1, 1, -1, 0, 0, 0, 0, 0, -2, -3, 2, 0, 0, 0, 0, 0, 0, 1, -2, -1, -2, 0, 0, 0, 0, -1, -2, -2, -1, 1, 0, 0, 0, -1, 0, -2, -1, 0, -1, -2, 2, -2, 0, -2, 0, -1, 0, 1, -1, 1, 1, 1, 0, 0, -2, -4, -3, -4, -2, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, -2, 1, 0, -1, 0, 0, -3, -3, -3, 0, 0, 0, 3, 0, 0, 2, -2, 0, -1, -1, 0, -1, 1, 0, 0, 0, 2, 1, 0, -1, -1, 0, 0, 0, 0, -2, -2, 0, 0, -2, 0, 1, 3, 0, 0, 2, -1, 0, -2, 0, -2, 0, 0, 1, 1, -1, 0, 0, 1, 1, 0, -1, 0, 0, -1, 0, -2, -1, 0, -1, 1, 1, 3, 1, 3, -1, -2, 0, 0, 0, -2, -3, 1, 0, -1, 1, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, 0, 0, 0, 1, -2, -2, 0, 0, -3, 0, 1, 1, 0, 1, 0, -1, -1, 0, 1, 0, -2, -1, -2, 0, -2, -1, -1, -1, 2, 0, 0, 0, 0, 1, 0, -1, 0, -1, 0, 3, 0, 0, -1, 1, 0, -2, 0, 0, -1, -1, 0, 0, 0, 0, -1, -3, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, -1, 0, -1, 3, 2, 1, 1, -2, 1, -1, -3, -1, 0, 0, 0, -2, -3, 0, -4, 0, 0, 1, 1, 0, 0, 0, 2, -2, -1, 0, 0, -1, -2, 0, 1, 1, 0, -1, -1, -1, 0, 0, -2, 0, -3, 0, 0, 0, 0, -2, 1, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -3, 0, 0, 0, -2, 0, 0, 0, -1, -1, -2, 0, -3, 0, -2, -1, -2, 0, 0, 0, 0, -1, 2, 0, 0, 1, 0, 0, 0, -1, -1, 1, 0, 0, 0, -1, 0, -1, 0, -1, 0, -2, 0, -2, -2, -2, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 1, 1, -1, -1, -2, -2, -2, -2, 0, -1, -1, 0, -2, -2, -1, 0, -2, -1, 0, 0, 0, -2, 0, 0, 1, 0, -2, -3, -2, -3, 0, 0, -2, 0, -1, -1, 0, -2, -2, 1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, -2, -1, 0, -3, -1, -2, -1, -2, -2, 1, 2, 0, -2, 0, 0, -2, 0, 0, 1, -1, -1, 1, 2, 1, 0, 0, 0, -1, 0, -1, -2, -2, -3, -2, -2, -1, -2, -2, -2, 4, 1, 1, 0, 0, -1, -1, -1, 0, 0, -2, 1, 0, 1, 0, -1, 0, 1, -2, -1, 0, -2, 0, 0, -4, -3, -2, -4, -4, -3, 3, 1, 0, -1, 0, 0, 0, -1, 0, 0, -2, 0, 0, 0, -1, 0, 0, -1, -1, 1, 0, -1, -1, -1, -2, 0, -3, -1, -4, -3, 5, 4, 0, 0, -1, 0, 0, 0, 0, -1, -1, -2, 0, 2, 1, 2, 1, 0, 0, 0, -2, -2, 0, -3, -1, -3, -3, -1, -1, 0, 11, 8, 5, 2, 4, 1, 0, -2, -2, -5, 0, 0, 0, 3, 4, 3, 2, 4, 4, 0, 1, -3, -3, -5, -4, -6, -6, -5, -6, -3, 11, 7, 1, 1, 1, 2, -2, 0, -4, -3, -1, 0, 0, 4, 1, 6, 2, 1, 0, 0, -3, 0, -2, -3, -6, -7, -8, -8, -5, -4, 11, 3, -1, -1, 0, 0, 0, -4, -4, -3, -2, 0, 2, 3, 2, 2, 3, 1, 2, -1, -1, -2, -2, -5, -5, -4, -5, -8, -5, -4, 8, 3, -3, -3, -3, -5, -3, -4, -2, -3, 2, 2, 2, 2, 3, 4, 3, 0, -2, 0, -1, 0, -2, -2, -3, -3, -2, -3, -8, -5, 7, 2, -4, -4, -6, -5, -6, -5, -3, 0, 2, 1, 4, 2, -1, 1, 1, 0, -3, -1, 0, -2, 0, 0, -1, -1, 0, -6, -7, -5, 7, 0, -2, -4, -3, -4, -2, -5, -5, -5, -2, 0, -1, 0, 0, 0, 0, -2, 0, 0, 2, 1, 0, 1, 2, 0, -1, -2, -4, -4, 9, 0, -4, -5, -4, 0, -2, -7, -6, -7, -5, -1, -3, -2, -2, -1, 0, 1, 2, 4, 2, 2, 3, 1, 0, 1, 0, -3, -2, -1, 8, 1, 1, 0, -3, -1, -3, -2, -5, -4, -4, -4, -3, -4, -4, -5, -4, 0, 3, 2, 4, 3, 1, 4, 1, 0, 0, -2, 0, -1, 10, 4, 1, 1, -1, 0, 0, 0, -1, -1, -3, -4, -3, -2, -4, -5, -6, -3, -2, 0, 2, 3, 0, 2, -2, 1, 0, 0, -4, 0, 9, 2, 1, 1, 0, 2, 4, 2, 3, 0, 1, 1, 1, -1, -4, -10, -9, -6, -4, -3, 1, 0, 0, -1, -1, 0, -1, -1, -4, -1, 6, 3, 1, 2, 0, 5, 4, 3, 3, 3, 2, 3, 3, -1, -5, -13, -14, -14, -10, -2, 0, 0, -1, -2, -3, -1, -2, -5, -4, -2, 4, 1, -4, 0, 2, 4, 8, 7, 8, 6, 6, 3, 3, -1, -9, -14, -17, -16, -8, 0, 0, 2, -1, -1, -2, -2, -5, -3, -4, -3, 4, -2, -2, -1, 1, 6, 10, 9, 4, 2, 2, 2, 2, -3, -7, -14, -15, -13, -4, 1, 5, 8, 5, 0, 0, -1, -3, -5, -5, -2, 3, -2, -6, -4, 1, 7, 9, 7, 4, 5, 5, 4, 3, 0, -7, -13, -13, -9, -4, 6, 12, 12, 8, 0, 0, -1, 0, -2, -2, -1, 3, -3, -5, -3, 0, 2, 7, 8, 6, 5, 5, 3, 4, -2, -6, -13, -15, -13, -6, 5, 11, 15, 11, 3, -1, 0, -3, -2, -6, -3, 5, 0, -5, -3, -1, 2, 5, 6, 7, 6, 5, 6, 5, 0, -5, -13, -20, -17, -8, 4, 9, 11, 9, 5, -1, 0, -4, -2, -7, -2, 3, -1, 0, -2, 1, 3, 6, 8, 5, 6, 6, 3, 2, -2, -8, -15, -17, -15, -6, 2, 5, 7, 7, 5, -1, 0, -3, -4, -5, -1, 7, 3, -1, 0, 0, 1, 4, 4, 3, 3, 3, 1, 2, -3, -8, -12, -17, -16, -8, 0, 4, 2, 4, 2, -2, -2, -4, -7, -6, -4, 8, 3, 1, 0, -1, 0, 1, 1, 0, 3, 0, 1, 0, -5, -9, -10, -16, -12, -7, 0, 2, 1, 3, 0, 0, 0, -4, -5, -4, -5, 6, 2, 2, 0, -3, 1, 0, 0, 2, 0, 0, -3, -5, -5, -9, -12, -11, -8, -3, 0, 3, 2, 4, 0, 0, -1, 0, -3, -5, -4, 5, 5, 0, 0, -3, 0, -1, 0, 0, 2, -2, -5, -8, -10, -9, -9, -6, -5, 0, 2, 3, 7, 4, 6, 4, 0, 0, -3, -5, -1, 7, 3, -1, 0, -4, -4, -2, 0, 0, -1, 0, -7, -10, -10, -7, -8, -5, 0, -1, 4, 7, 6, 6, 3, 3, 2, -1, -3, -4, -4, 10, 1, 0, -3, -2, -5, -4, -2, -1, -1, 1, -3, -5, -7, -3, -3, -2, -2, -1, 0, 0, 3, 3, 4, 0, 1, 0, -4, -5, -4, 10, 4, -1, -1, -4, -4, -6, -4, -2, 0, 1, 0, 1, 0, 0, -3, -5, -6, -4, -5, -2, -1, 1, -2, -2, 0, -1, -2, -3, -3, 6, 0, -1, -4, -3, -3, -4, -1, -1, 1, 2, 0, 2, 3, 0, 0, -3, -3, -6, -5, -2, -3, -2, -1, -1, -5, -4, -6, -6, -6, 6, 0, 0, -2, -1, -1, -4, -3, -3, 0, 1, 0, 3, 2, 1, -1, -1, -1, -2, -2, -1, -4, -2, -5, -3, -4, -4, -6, -6, -4, 9, 0, 0, -2, -1, -2, -3, -3, -2, -1, 1, 0, 2, 3, 4, 3, 3, 0, -1, -1, -2, -4, -7, -9, -7, -7, -7, -7, -7, -5, 12, 4, 1, 0, 2, 2, 0, -4, -6, -4, -2, 1, 0, 2, 4, 7, 1, 2, 0, 0, -4, -4, -6, -7, -8, -7, -7, -3, -4, -5, 14, 8, 5, 4, 0, 1, 0, 0, -2, -3, -2, 0, 1, 4, 7, 8, 7, 2, 1, 0, -3, -1, -2, -5, -5, -6, -4, -5, -4, -2, 14, 9, 6, 5, 4, 3, 2, 1, 2, 2, 0, 3, 3, 8, 12, 12, 8, 9, 5, 5, 5, 0, 0, 1, -1, -2, 0, -2, -4, -1, 4, 3, 3, 1, 2, 1, 1, 3, 1, 2, 3, 4, 2, 2, 0, 3, 1, 0, 3, 2, 0, 1, -1, -1, -1, 0, 0, 0, 0, -1, 1, 2, 2, 4, 1, 2, 0, 1, 3, 2, 3, 0, 3, 0, 0, 2, 1, -1, -1, -2, -2, 0, -4, -1, -3, -3, -4, 0, -2, -4, 2, 2, 1, 3, 4, 0, 2, -1, 2, 1, 0, 0, 0, 2, 1, 0, 0, 0, -3, 0, -2, -2, -2, 0, -3, -4, -5, -4, -2, 0, 0, 0, 0, 1, 0, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, -1, -1, -1, -1, -3, -3, 0, -3, -1, -2, -5, -3, -1, 1, 0, -1, 1, -1, 1, 0, 0, 3, 1, 2, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, -2, 0, -1, -1, -3, -3, -2, -3, -1, 1, 0, 1, 2, -1, 0, -1, -1, 1, 1, 1, 2, 2, 1, -1, 0, 0, 0, 0, -3, -1, 0, 0, -3, 0, 0, 0, 0, -4, 0, 0, 1, 0, -1, 2, 0, -1, 0, 2, 2, 0, 1, 0, 2, 0, 0, 0, 1, -2, 0, 0, -2, -2, 0, -1, -2, -2, -2, -4, 0, 0, 0, -1, 0, 0, 0, -2, 0, 0, 1, 1, 3, 0, -1, 2, -1, 1, 1, 0, -1, 0, 0, -2, 1, -1, -2, -2, -3, -5, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -2, -2, -1, 0, 0, 0, 1, 1, 4, 4, 1, 0, 2, 1, 1, 0, 0, -2, -2, -3, -2, 3, 0, 2, 1, 2, 2, 0, -2, -2, 0, 0, -3, -2, -1, 0, 2, 2, 4, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, -3, 3, 1, 2, 0, 3, 1, 1, 0, 0, 1, -1, -1, -2, -4, -1, -2, 0, 1, 3, 0, -1, 0, 0, -2, 0, 0, 0, 0, -2, 0, 3, 2, 2, 3, 4, 2, 2, 2, 1, 0, 3, 0, -1, -3, -2, -4, -1, 3, 3, 2, -1, 0, 0, -3, 0, 0, 0, -1, -2, 0, 3, 1, 0, 3, 2, 1, 2, 2, 0, 1, 1, 0, 0, 0, -3, -4, -1, -1, 0, 0, 0, -1, -3, -1, -2, -3, -2, 0, -2, -2, -1, 0, 1, 2, 2, 3, 4, 2, 2, 2, 0, 0, -1, -5, -5, -2, -2, 0, 4, 0, -1, -3, -2, -4, -3, -1, -1, -1, -3, -2, -1, -1, 2, 4, 5, 3, 2, 0, 0, 0, 2, -1, -2, -4, -3, -5, -1, 1, 6, 5, 1, -2, -1, -1, -2, -1, -3, -2, 0, -1, 1, 0, 0, 0, 3, 5, 3, 1, 0, -1, -1, 0, -1, -2, -2, -2, -2, 3, 5, 4, 5, 1, -3, -2, 0, -1, -3, -1, 0, -2, -1, 0, 0, 1, 4, 4, 3, 1, 0, 0, 0, 0, 0, -3, -6, -4, -3, 1, 6, 6, 4, 1, 1, 0, 0, -1, -1, 0, -3, -2, -1, -1, 0, 2, 0, 2, 4, 4, 3, 3, 2, 0, -2, -1, -6, -6, -3, 3, 4, 5, 1, 3, -1, -2, 0, 0, 0, -1, -3, 1, 2, -1, 0, 0, 1, 3, 2, 0, 0, 3, 2, 0, -2, -4, -3, -5, -2, 1, 1, 4, 1, 0, -1, 0, -1, 0, -2, -4, -3, 0, 2, 3, 3, -1, 1, 3, 0, 1, 1, 0, -1, -1, 0, -4, -3, -6, -3, 0, 0, 3, 3, 0, -1, -1, -2, -1, 0, -4, -3, -1, 0, 0, 2, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, -2, -2, -5, -3, -1, 2, 0, 0, 0, 0, -1, -2, -2, -2, -2, 0, 0, 1, 0, -1, 1, 1, 0, 3, 1, -1, 0, -3, 0, 0, -4, -3, -3, 0, -1, 2, 3, 3, 0, 0, -1, -2, 0, -2, -3, -4, -3, -1, 0, 1, -1, 2, 0, 1, 2, 1, 0, 0, -4, 0, 0, -2, 0, -1, 1, 3, 5, 4, 2, 2, 3, -1, -2, 0, -3, -3, -2, -1, 0, 1, -1, 0, 1, -2, 0, 0, 1, -1, -1, 0, 0, -1, 0, -1, 1, 3, 1, 1, 0, 1, 1, 2, 0, 0, -2, -4, -3, 0, 0, 0, -2, -2, 0, -1, -2, 0, 0, 0, 0, -2, 0, 0, 0, 1, -1, 2, 1, 2, 0, -1, 1, 0, 0, -2, -3, -4, -2, 0, 1, 1, 0, 0, -1, 0, 1, 0, 3, 2, -1, 1, -1, 0, 0, -3, 1, 0, -2, 1, -1, 1, -1, 0, -2, 0, 0, -3, 0, -1, 0, 1, 0, 0, 0, 0, 0, 3, 4, 3, 2, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, -4, -2, 0, 1, -1, -1, 0, -1, -1, -2, 1, 1, 3, 1, 0, 2, 1, 0, 0, -1, -1, -1, 0, -1, -3, -2, -2, -2, 0, 0, -1, -2, -3, 2, 0, 0, 0, 2, -1, 0, -1, -1, 0, 2, 2, 0, 0, 0, -1, -3, -1, -3, 0, -4, -3, -4, -2, -2, -4, -3, -5, -5, -1, 2, 0, 1, -1, 2, 0, 0, 0, -1, 1, 1, 0, 2, 0, 0, 0, -2, 0, -2, -3, -2, -4, -2, -5, -5, -3, -5, -3, -2, 0, 0, 0, 1, 0, 0, -1, -2, -1, 0, -1, -1, 2, -1, 1, 0, 0, 2, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 1, 0, 1, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, -1, 1, 0, 1, 1, 0, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, -1, 0, 0, -1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, 1, -1, -1, -1, 1, -1, -1, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, -1, -1, 1, 0, 0, -1, 0, 0, 1, -1, 0, -1, 0, -1, 1, 0, -1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 0, 2, 2, 0, 0, 1, 0, -2, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -1, -1, 1, 1, 2, 1, 0, 0, -1, 0, -1, 0, 1, -1, 0, 0, -2, 1, 0, -1, 1, 1, -1, -1, -1, 0, 0, 0, 1, 1, 1, 0, 0, -1, 1, 1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, -1, 0, 0, 1, 0, 0, -1, 0, 0, -1, 1, 0, -2, 1, 1, -2, 1, 0, 0, -2, 0, 1, 0, 0, 0, -1, 0, 0, -1, 1, -1, 0, 1, 1, -2, 0, -1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 1, -1, -1, -1, 1, 0, 1, 0, 0, 1, 0, 0, -2, -1, 0, 0, 0, 1, -1, -2, -1, 0, 1, 0, -1, -1, -1, 0, 0, 1, 0, 0, 0, -1, 1, 1, -2, 0, 0, 1, -1, 0, 0, 1, -1, 0, -2, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, -1, 0, -1, -1, 0, 0, 0, -1, 1, 2, 1, -1, -1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, 1, 1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 1, 0, 1, 0, 1, -1, 1, 1, 1, 2, 0, 1, 0, 1, -1, 0, -2, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, -2, 0, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, -1, 1, 1, -1, 1, -2, 1, 0, -1, 1, 0, 1, 0, 0, -1, -1, 0, -1, 1, 1, 0, -2, 1, -1, 1, -1, 0, 1, 0, 1, 1, 0, 1, -1, -1, 0, 1, 1, -2, 0, -2, 0, 1, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 1, 1, 1, -1, 0, 0, 1, 1, 2, 0, 1, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 0, 0, 0, -1, -1, -1, -1, 2, 1, 0, 1, 0, 0, 0, -1, -1, 0, 0, 0, -1, 0, -1, -1, 1, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, -2, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 0, 0, 1, 1, -1, 1, -1, 0, 2, -1, -1, 0, 1, -1, -1, -1, -1, -1, 0, 1, 0, 0, 2, 1, 0, 0, -2, 1, -1, -1, 0, 0, 0, 1, 2, 0, 0, -1, 1, 1, 0, 0, 1, 2, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, 0, -2, -1, -1, 1, 2, 0, 0, 1, 0, 1, 1, 0, 0, -1, 0, -1, 1, -1, -1, 0, 1, 1, 1, -2, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 1, -1, 2, -2, -1, -1, 1, 1, 0, -1, 1, 1, 1, 0, -2, 0, 1, -1, 2, 1, 0, -1, 0, -1, 0, 0, -1, 1, -1, -2, 0, 1, 0, -2, 0, -2, 0, 0, 1, -1, 0, 1, -1, -1, 1, 0, 0, -1, 0, 0, -1, 0, 1, -1, 1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 0, 1, -1, 1, -1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 1, 2, 1, 0, 1, -1, 1, -1, -1, 0, 1, 1, 2, -1, 0, -1, 0, 1, 0, 1, 0, -1, 0, -1, -1, 0, 2, 0, -1, 0, -1, 1, 0, -1, -1, 0, 0, 1, 0, 1, 0, 0, 1, -1, 1, 1, 1, 0, 1, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 0, -1, 1, 1, 0, 1, -1, 0, 0, 1, -1, -1, 1, -2, 0, 0, 1, 1, 0, 0, 1, -2, 1, 0, 0, 0, 0, 1, -1, 1, 1, 0, -1, 0, 1, 1, 0, 0, -1, -1, 2, 0, 0, 0, 2, 0,
    -- filter=0 channel=8
    -3, 0, -1, -1, 0, 0, -1, -2, 0, 0, 0, -1, 0, -1, -1, 1, -1, 0, 0, -1, 0, -1, 1, 0, 2, 3, 0, 0, 0, 2, 0, 0, -1, -1, 0, -2, 0, 0, -1, 0, 1, 1, 0, -1, 0, 1, 0, 0, 0, 1, -1, 0, 1, 1, 0, 0, 0, -1, 0, 2, 0, 0, 0, -1, -1, -2, -2, 0, 0, 1, 0, 1, 1, 0, -1, 1, 0, 0, -2, 0, 0, 0, -2, -2, -2, 0, 0, 0, 1, 3, -3, 0, 0, -1, 0, 0, -1, 0, -2, 0, -1, -1, 0, -2, 0, -2, 1, -1, 1, 0, 2, 1, 0, -2, 0, -2, -1, 1, 2, 3, -2, -3, -3, 0, -2, -3, -1, 0, 0, 0, -2, 0, 0, 0, -1, 1, 0, 0, -1, 0, 2, -2, -2, 0, -1, -2, 0, 1, 1, 3, -1, -1, 0, 0, -1, -2, 0, 0, 0, 0, -3, -3, 0, -1, -2, 1, 1, 0, 1, 1, 1, 0, -2, -1, 0, -1, 1, -1, 2, 1, 0, 0, 1, -2, -3, -2, -3, 0, -3, -1, -2, 0, -3, -3, -1, 1, 1, 0, -1, 1, 0, -1, -1, -1, 0, 0, 0, 0, 1, 1, -2, 0, 0, 0, -1, 0, -2, 0, -2, -1, -1, -2, 0, 0, 0, 0, -2, 0, -1, 1, -1, 1, -1, 1, 1, -1, -2, -1, 1, 3, -2, 0, 0, -2, -1, -1, 0, 0, 0, -1, -1, -2, 0, 0, 0, 1, -1, -1, 0, 1, 0, -1, 1, -2, 0, 2, 0, -1, 0, 2, 0, 0, -2, -1, 0, 0, 0, -1, -1, -4, -1, -4, -3, -1, 0, 1, -1, 1, 2, 2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, -2, 0, 0, -1, -1, 0, -1, -3, -2, -4, -1, -1, -2, -3, -1, 0, -1, 2, 2, -1, 0, -2, -1, 0, -1, 0, -1, -1, 0, 2, -2, -2, -1, 0, -3, 0, -1, -3, -4, -1, -3, -4, 0, -2, 0, 1, 0, 0, 0, 0, 2, 1, 1, -2, 0, 1, 0, 0, 1, 2, -1, 0, -2, 0, -1, -3, 0, -1, -3, -3, -3, 0, 0, -1, 0, -2, 0, 1, 1, 0, -1, 1, 0, 0, -1, -1, -1, 0, 2, 0, -2, -2, 0, -2, -2, -1, -2, -4, -3, -1, -3, -2, -2, 0, -1, -2, 1, 0, 1, 0, 2, 1, 0, 0, -2, -1, 0, 0, 0, 3, -2, 0, -2, -1, 0, -3, -2, -1, -1, -1, 0, -1, 0, 1, 0, -1, 0, 0, -1, 0, -1, 3, 0, 0, 0, -3, 0, 1, 1, 0, -1, 0, 0, 0, 0, -3, 0, -1, -2, -2, -2, 0, -1, -1, -1, -2, 0, -2, -1, 0, 0, 0, 1, 1, -1, -2, 0, 0, 0, 0, -2, -3, 0, 0, -1, -1, -3, -2, -4, -2, -1, -3, -2, 0, -1, -1, -1, 1, -1, 0, 2, 2, 1, 1, -2, 0, 1, 0, 0, 1, -2, -3, 0, -1, 0, -2, -4, -3, -3, 0, -2, -2, -2, 0, -2, -1, -2, 0, -1, 0, 0, 1, 1, 1, 0, -1, 1, 0, -1, 1, 0, -2, -2, -1, -1, -2, 0, -4, -1, -1, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 1, 2, -1, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, 0, 0, -2, 0, -1, -1, -1, -2, -1, -2, -2, -3, -1, -1, 0, 1, 0, 1, 0, -3, 0, 0, 1, 1, 1, -1, 0, 0, 0, -3, -2, -2, 0, -2, 0, -2, 0, 0, 0, 0, -1, 0, 1, 0, 0, -1, 2, 0, 0, 0, -3, -1, 0, 0, 3, 0, 0, 0, 0, 0, -2, -1, 0, -3, -1, 0, -1, -1, -3, 0, 0, -2, 0, -1, -1, 0, 2, 0, -2, 0, -1, -2, 1, 0, 2, 0, 0, 1, 0, -2, 0, -1, -1, 0, -1, -3, -2, -2, -1, -3, -2, -1, 1, 0, 0, -1, 0, 1, 0, -2, -2, -1, 0, 1, 2, -3, -1, 0, 0, -1, -2, -2, -1, 0, 0, 1, 0, -2, -1, -2, 0, 2, 0, 0, 0, 0, 0, 1, -2, 0, -1, -1, 2, 2, 4, -1, -2, -1, 0, -2, -2, 0, -1, -2, 0, -3, -1, -1, -1, 1, 0, 1, -1, 1, 1, -1, 0, 0, 0, 0, -1, 1, 2, 0, 3, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -2, -2, 1, 0, 0, 0, 0, -2, 1, 0, 1, -1, 0, -2, 0, 1, 2, 2, 4, 0, 0, -1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 0, -1, -1, -2, 1, 0, 0, 4, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, -2, -1, 0, 0, 1, 1, 2, 2, 0, 4, 3, -1, -2, -2, -1, 0, -2, -1, -1, -1, -2, 0, 1, 0, 2, 0, 0, 2, -2, -1, 0, 1, 2, 2, 2, 0, 0, 0, 3, 3, 3, -2, -1, -2, 0, 0, 0, -2, 0, 0, -3, -1, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 3, 3, 1, 2, 3, 5, 2, 0, 2, 0, 0, 0, 0, 0, 2, 0, 1, 2, 1, 2, 5, 6, 6, 6, 8, 6, 9, 8, 6, 9, 8, 6, 6, 8, 7, 4, 4, 3, 0, 1, 0, 1, 1, 0, 3, 2, 1, 1, 4, 4, 5, 0, 0, 3, 5, 5, 4, 6, 6, 7, 9, 7, 6, 7, 8, 2, 3, 3, 1, 2, 2, 1, 1, 4, 1, 1, 0, 0, 4, 0, 0, 0, -1, 2, 1, 3, 3, 5, 3, 5, 5, 5, 8, 8, 7, 3, 4, 4, 3, 3, 4, 3, 1, 2, 3, 2, 1, 2, 1, 2, -1, -2, 0, 0, 0, -2, -1, 1, 1, 4, 6, 8, 7, 8, 7, 5, 4, 2, 3, 3, 0, 1, 2, 1, 1, 0, 2, 0, 3, 0, 0, -1, 0, -3, 0, -3, -1, -2, 0, 0, 3, 6, 6, 6, 5, 2, 1, 3, 3, 3, 1, 2, 1, 1, 2, 1, 0, 3, 2, -2, -2, 0, -4, -2, -2, -5, -6, -2, -2, 1, 1, 6, 5, 5, 3, 0, 4, 3, 1, 3, 2, 1, 2, 2, 1, 1, 0, 2, -1, -2, -1, -3, -1, -1, -6, -4, -7, -4, -3, 0, 2, 1, 4, 5, 2, 1, 2, 4, 3, 1, 2, 2, 4, 2, 3, 2, 1, -1, 0, 0, -1, -3, -1, -2, -5, -7, -5, -6, -1, -1, -2, 2, 3, 3, 1, 2, 1, 2, 2, 2, 1, 3, 4, 2, 3, 0, 1, 2, 2, -1, -2, 0, -3, 0, -2, -3, -3, -2, -4, -2, -2, 1, 0, 0, 4, 1, 2, 2, 1, 1, 2, 1, 2, 3, 1, 1, 1, 0, 2, -1, -3, -2, -1, -3, -4, -1, -4, -6, -4, -4, -2, 1, 2, 2, 1, 1, 1, 3, 1, 0, 0, 1, 0, 0, 1, 3, 2, 1, 0, 1, 0, 0, 0, -3, -2, 0, -2, -4, -3, -1, -3, 0, 1, 2, 3, 4, 3, 3, 2, 1, 1, 0, 1, 2, 3, 1, 3, 0, 1, 0, 0, -2, 0, 0, -2, -1, -1, -1, 0, 0, -2, 0, -1, 1, 1, 3, 2, 2, 3, 0, 0, 0, 1, 3, 3, 3, 0, 2, 0, 2, 1, -1, 0, -3, -2, -1, 0, -2, 0, 0, -2, 0, 2, 3, 2, 2, 0, 3, 3, 2, 3, 2, 2, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, 0, -4, -3, -4, 0, -1, 0, 0, 2, 3, 2, 0, 2, 3, 0, 0, 0, 1, 3, 3, 0, 2, 0, 1, 1, -3, 0, 0, 0, 1, 0, -1, -3, -3, -2, -3, -1, 2, 0, 1, 0, 2, 2, 3, 3, 2, 1, 0, 2, 3, 0, 3, 2, 1, 0, 0, 0, 0, 2, -1, -1, 0, -2, -4, -1, 0, -1, 0, 0, 4, 3, 1, 2, 2, 2, 0, 0, 1, 0, 2, 0, 0, 3, -1, 0, -2, 0, 1, 0, 2, 0, -2, 0, -4, -5, 0, 0, 0, 4, 2, 2, 2, 2, 1, 3, 0, 0, 2, 2, 1, 3, 3, 2, 1, 0, -1, -3, 0, 0, 2, 1, 0, -3, -3, -3, -3, 0, 0, 2, 4, 2, 0, 3, 2, 0, 0, 0, 1, 3, 0, 2, 1, 3, 3, 2, 0, 0, 0, -1, 0, -1, -3, -1, -4, -5, -3, 0, 2, 0, 4, 0, 3, 3, 2, 1, 0, 2, 0, 3, 4, 3, 1, 0, 1, 0, -2, -3, -2, -1, -1, -2, -2, -2, -6, -6, -5, 0, 0, 1, 3, 4, 2, 2, 3, 2, 0, 0, 2, 4, 0, 2, 1, 2, 0, 0, -2, -2, 0, 0, 0, -3, -1, -3, -4, -3, -5, -2, 3, 1, 2, 4, 2, 3, 1, 1, 1, 0, 2, 1, 1, 3, 3, 3, 1, 0, 0, 1, -2, -1, 0, -2, -6, -3, -1, -3, -3, -1, 2, 4, 2, 4, 1, 2, 1, 1, 2, -1, 1, 2, 3, 2, 2, 2, 3, 2, 0, 0, -1, 0, -2, -3, -4, -4, -4, -4, -4, 0, 3, 4, 3, 3, 0, 2, 2, 0, 0, 0, 1, 3, 1, 2, 1, 2, 3, 3, 3, 0, -1, 0, -1, -2, -2, -3, -1, -3, 0, 0, 3, 5, 5, 3, 1, 2, 0, 1, 2, 3, 2, 2, 4, 3, 1, 2, 2, 3, 0, 1, 0, -1, -3, -5, -3, -4, -3, -4, 0, 1, 3, 2, 2, 4, 1, 1, 0, 0, 2, 0, -1, 2, 2, 4, 0, 1, 2, 4, 0, 0, 0, -2, -1, -3, -1, 0, -1, 0, 0, 3, 5, 4, 5, 3, 4, 0, 2, 3, 1, 2, 0, 3, 2, 3, 1, 2, 1, 3, 3, 1, -1, 0, 0, -1, -1, 0, 2, 2, 1, 4, 8, 6, 6, 3, 5, 3, 2, 3, 3, 2, 0, 2, 1, 3, 2, 3, 1, 0, 2, 2, 0, 0, -1, 0, 2, 3, 5, 3, 3, 6, 7, 8, 7, 7, 2, 4, 2, 0, 1, 0, 1, 0, 3, 3, 2, 1, 2, 2, 2, 3, 0, 3, 2, 3, 2, 6, 5, 7, 6, 7, 10, 8, 8, 8, 2, 3, 3, 3, 0, 1, 1, 0, 0, 3, 5, 4, 3, 4, 4, 4, 5, 4, 7, 7, 8, 6, 6, 7, 10, 8, 8, 10, 9, 9, 1, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 3, 2, 4, 3, 2, 6, 3, 5, 6, 4, 7, 6, 6, 4, 8, 7, 6, 2, 2, 1, 0, 0, 0, 0, 1, -1, 1, -1, 1, 0, 3, 3, 2, 2, 2, 0, 3, 4, 5, 2, 2, 6, 6, 5, 6, 8, 6, 2, 0, -1, 0, 0, 2, 0, 1, 1, 3, 0, 0, 0, 2, 0, 3, 0, 1, 1, 2, 1, 1, 2, 5, 4, 7, 3, 8, 8, 8, 0, 0, 0, 3, 2, 1, 0, 1, 0, 2, 1, 2, 0, 0, 2, 0, 0, 0, 0, 0, 1, 1, 0, 2, 3, 2, 5, 4, 8, 7, 3, 3, 2, 0, 0, 0, 0, -1, 3, 3, 2, 1, 0, 0, 1, 1, -1, -1, 0, 0, 1, 1, -1, 1, 3, 4, 2, 7, 4, 6, 2, 0, 0, 1, 0, 1, 0, 1, 2, 0, 2, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, -2, -1, -2, 2, 1, 4, 3, 7, 4, 1, 2, 0, 1, 0, 0, 0, 3, 1, 1, 0, 0, -3, 0, -1, -2, -2, -4, -3, -3, -4, -3, -1, -1, 0, 0, 1, 2, 4, 3, 2, 1, 2, 1, 1, 0, 2, 1, 0, 0, 0, 1, -2, 0, -1, -2, -1, -3, -4, -4, -4, -3, -1, -1, 0, 2, 0, 4, 2, 5, 1, 0, 0, 0, 2, 1, 0, 2, 2, 1, 0, -1, -1, 0, 0, -3, 0, -2, -3, -4, -1, -1, 0, 0, 0, 0, 0, 1, 4, 4, 0, 2, 2, 2, 0, 0, 0, 0, -1, 1, 0, -2, -1, 0, -3, -1, 0, -3, -2, -1, -3, -3, 0, -2, -2, 1, 1, 0, 1, 4, 3, 3, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, -2, 0, -1, 0, -2, -1, -1, -3, -2, -2, 0, -1, 0, 0, 1, 0, 2, 5, 1, 0, 1, 1, 2, 1, 0, 2, 2, 1, 2, -1, -2, -2, 0, -2, -1, 0, -1, 0, -3, 1, 0, 0, 0, 2, 0, 3, 3, 3, 0, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -2, -1, 0, -2, -1, 0, -1, -1, 1, 0, -1, 2, 1, 4, 4, 0, 2, 2, 1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, -1, 1, 1, -1, -2, 0, 0, -1, 0, -1, 2, 2, 0, 2, 4, 1, 0, 0, 0, 0, 0, 0, 1, 1, -2, 0, -1, -1, -1, 0, -3, -1, -2, -3, -2, 0, 0, 0, 1, -1, 1, 2, 0, 3, 2, 0, 1, 2, 2, 2, 2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, -2, -1, -2, 0, -1, 0, 1, 0, 2, 4, 1, 1, 2, 1, 0, 1, 2, 0, 1, 0, -1, 0, -2, -2, -1, 0, -1, 0, 0, -1, -1, 0, -2, 1, -1, 0, 1, 2, 1, 4, 0, 0, 1, 0, 2, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, -2, -2, -1, -3, 0, 1, 0, -2, 0, -1, 0, 0, 1, 1, 2, 2, 0, 0, 0, 2, 0, 0, -1, 0, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, -1, -2, 0, -3, 0, 0, -1, 1, 2, 2, 3, 1, 2, 0, 1, 1, 2, -1, -1, 0, 1, 0, 0, 0, -1, 1, -2, 0, -3, 0, -2, -2, -3, -3, 0, -1, 0, 0, 0, 1, 1, 1, 2, 1, 3, 2, -1, 0, -1, 0, 0, 0, 0, -1, 0, -2, -1, 0, -1, -1, -1, -1, -1, -1, 0, -3, -2, -1, 0, 4, 2, 1, 0, 2, 0, 2, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, -1, -2, -3, -1, -2, -3, -2, -4, -3, -2, 0, 1, 0, 3, 4, 2, 0, 1, -1, 1, 0, 0, 2, 0, 2, 1, 0, 2, -1, 0, 1, -2, 0, -2, -3, 0, -3, -3, -3, 0, 1, 1, 0, 4, 3, 3, -1, -1, 2, 2, -1, 0, 0, -1, 0, 0, 0, 2, 0, -1, 0, -1, 0, -1, -1, -3, -1, -3, 0, 1, 1, -1, 3, 1, 3, 5, 0, 2, 2, 1, 0, 2, 0, 1, 1, 0, 2, 1, 1, 0, 2, -1, 0, 0, -1, -2, -1, 0, 0, 0, 0, 1, 1, 4, 5, 4, 0, 0, 1, 0, 2, 0, 0, -1, 3, 0, 1, 3, 2, 2, 1, 1, 1, -2, 0, -3, -2, 0, 0, 1, 1, 3, 4, 2, 4, 6, 2, 0, 0, 0, -1, 0, 2, 0, 0, 3, 1, 0, 3, 2, 0, -1, 0, -2, 0, -3, 1, 0, 1, 2, 0, 2, 6, 4, 4, 5, 2, 0, 0, 3, 1, 1, 1, -1, 1, 1, 0, 0, 0, 0, 3, 0, 2, 0, 0, 0, 2, 2, 4, 2, 4, 5, 4, 7, 7, 6, 1, 2, 1, -1, 2, 1, 0, -1, 1, -1, 1, 0, 3, 1, 3, 1, 1, 2, 1, 3, 3, 2, 2, 6, 7, 7, 8, 6, 6, 5, 2, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 3, 4, 2, 2, 3, 3, 6, 5, 6, 5, 8, 7, 6, 10, 9, 6, 0, -1, 0, -1, 1, 0, 1, 1, 0, 0, 1, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, -1, 0, 1, 1, 1, 0, -2, -1, 0, 0, 2, 0, -1, 0, 0, -2, 0, -1, 1, 1, 1, 0, 0, 0, -1, -1, 1, 0, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 1, 1, 1, -1, -1, 0, -1, 1, 1, -1, 1, 0, 0, 0, -2, -1, 0, -1, -1, 0, 1, -1, -1, 2, 1, 1, 1, -1, -1, 0, -1, 0, -1, -1, 1, -2, 0, -1, 1, 1, -1, 0, 1, -1, -1, 0, -1, 0, 0, 1, -2, 1, 1, 1, 0, 0, -1, 1, 1, -1, 2, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 1, -2, 0, 1, -1, 2, 0, 0, 1, 1, 0, -1, 0, -1, -1, -1, 0, 0, -1, 1, 1, 0, -1, 1, -2, 0, 1, 0, 0, -1, 1, 2, 0, 0, 0, -1, 1, 1, 1, 1, 0, -2, 0, -1, -1, 0, 2, 0, 1, 0, 1, 0, -1, -1, 0, -1, 2, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -2, 0, -1, 0, 0, 1, 0, -1, -1, -1, -1, 1, 1, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 0, 0, 0, 0, 2, -1, 1, 0, 2, -1, 0, 0, 2, -1, -1, 0, 1, 0, 1, 1, 0, 0, 0, -1, 0, 1, -1, -1, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 1, 1, -1, 1, 1, 0, -1, 0, 0, -2, 0, 1, -2, -1, 0, -1, 0, -1, 1, 0, -1, 0, -1, -2, -1, 1, 1, 0, 1, 1, -1, 1, 0, -1, 0, 0, 2, 2, -1, 0, -1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 2, 2, 0, -2, 0, 1, 0, 1, 0, 2, 1, 1, 1, -1, 0, -1, -1, 1, 1, -1, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, 0, -1, 1, -1, 0, 0, 0, 0, -1, -1, -1, 1, 0, 0, 0, 0, 2, 1, -1, 1, -1, -1, 0, 2, 0, -1, -1, 0, 2, 1, 0, 1, -1, 1, 0, -2, -1, 1, 0, 1, -1, 2, 0, 0, 1, 1, 1, -1, 0, -1, 1, 0, 1, 0, -1, 0, 0, 0, 1, 1, -1, -1, 0, 1, 0, 0, 1, 0, 0, 1, -2, -1, 0, 0, 0, 1, 0, 0, 2, 1, 1, -1, 0, 1, 0, 0, 0, -2, 0, 0, -1, 0, -2, 0, 0, 0, 1, 0, -1, 0, 0, -2, -1, 0, 1, 0, 1, -1, -1, 0, 0, 0, 1, -1, 0, -1, 0, 1, 0, -1, 0, 1, 1, 1, 0, 1, 0, 0, -1, 1, 2, 0, 2, -1, -1, 1, -1, 0, -1, 1, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 2, 0, -1, -1, 1, 1, -1, 1, -1, 0, -1, 1, 0, 1, -2, 1, 0, -1, 1, 0, 0, 1, 0, 1, -1, -1, 0, -1, 0, 1, 0, 1, 0, -1, -1, 0, -2, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, -1, 0, -1, 1, 1, 1, -1, 0, 1, 0, 1, 1, 0, -2, -1, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, -1, 1, 1, -1, 0, 0, -1, 0, 0, 0, 0, -1, 2, 0, 0, 0, -1, 0, -1, 1, -1, 1, 1, -1, 1, -1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 1, 0, 1, 1, 1, 1, -1, 0, 1, 1, -1, -1, 0, 0, -2, -1, 0, -1, 0, 0, 1, 0, 0, -1, -1, -2, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, -1, 1, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, -1, 0, 1, 0, 2, 0, -1, -1, -1, 0, 0, -2, 1, 1, -1, 0, -1, 1, 0, 0, 1, 0, -2, 0, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, -1, 0, 1, 0, 0, 1, -1, 0, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 0, -1, -1, 1, 2, -1, -1, -1, 0, -1, 1, -1, 0, 0, 0, -1, 1, 1, 0, 0, 1, -1, -1, 0, 0, 1, 1, -1, 0, -1, 0, -1, -2, 1, -1, 0, 0, 0, 2, 1, -1, -1, -2, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 0, -1, 1, 2, 1, 0, -1, 0, 2, -1, 1, -1, 2, 0, -1, -1, 0, 1, -1, 0, 2, 0, -1, 2, 0, 1, 1, 0, 2, 1, 0, 0, 0, -1, 0, 1, -1, -2, 0, 0, 0, 0, 1, 1, -2, 0, -1, -2, 0, 0, 0, 1, 0, -1, -1, -2, 0, 1, 0, 0, 0, 3, 0, 2, 0, 0, 0, 0, -4, -4, -2, -2, -4, -2, -2, 0, -3, 0, 0, -2, 0, 0, -3, -4, -4, -6, -6, -7, -9, -11, -12, 3, 2, 0, 0, -1, 0, -1, -3, -2, -3, -2, -3, -1, 0, 0, -3, -1, -2, -2, 0, -1, 2, -1, 0, 0, -4, -6, -5, -5, -10, 0, 1, -1, 0, 1, -2, 0, 1, 0, 0, -1, -2, -3, -2, -2, -3, -4, -2, -2, -1, 0, 0, 0, 0, -1, -3, -4, -3, -6, -8, 4, 0, 1, 1, 0, 0, -2, 0, 0, 0, 0, -3, 0, 0, -1, -1, -1, -2, -2, 0, -1, -1, 3, 3, 1, 0, -1, -1, -5, -5, 0, 2, 1, 0, -1, 0, 1, 1, -1, 0, 0, 0, 1, -2, 0, 0, -1, 0, 0, -1, 0, 0, 2, 0, 0, 0, 1, -1, -2, -7, 0, 0, 2, 0, 0, 0, 0, 0, 2, 0, 0, -1, 0, -3, -2, 0, 0, 0, 0, 0, -1, 0, 1, 0, 1, 2, 0, -3, -2, -6, 2, 0, 1, -1, 1, 0, 1, -1, -1, -1, 1, -1, 0, 0, -1, 1, 0, -1, 1, -1, 0, 0, -1, 0, 0, 2, 0, 0, -2, -6, 2, 1, 1, 1, -1, 1, 0, -1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 3, 3, 1, 0, -2, 0, -5, -4, 0, 1, 1, 1, -1, -1, 1, 1, 2, 1, 1, 2, 1, 4, 2, 2, 0, 0, 1, 2, 1, 0, 1, 0, 0, 0, 0, -1, -3, -5, 0, -1, -2, 0, -2, -2, -1, -2, 1, 1, 2, 0, 1, 0, 2, 0, 2, 4, 2, 2, 3, 0, 1, 0, 0, -2, -2, -3, -3, -7, 2, 0, 0, -1, -2, -2, -2, 0, 0, 0, 2, 0, 1, 3, 0, 2, 2, 3, 0, 2, 4, 3, 2, 3, 1, 0, -1, -1, -3, -8, 1, 0, 0, -2, -1, -3, 0, -1, 0, 0, 5, 5, 3, 4, 1, 1, 0, 0, 1, 2, 1, 2, 0, 1, 1, 2, 0, -4, -2, -6, -1, 0, -1, -2, 0, -1, 1, 2, 2, 0, 4, 5, 2, 3, 2, 2, 0, 0, 0, 0, 2, 3, 1, 0, 1, 2, -2, -2, -4, -5, -2, 0, 1, -2, -2, -2, 0, 0, 0, 0, 2, 1, 0, 0, 1, 1, 3, 1, 1, 1, 3, 2, 0, 0, 2, 0, 0, -2, -2, -6, 0, 0, 0, 1, -2, 0, 1, 1, 1, 2, 2, 0, 2, 0, 0, 0, 2, 1, 1, 1, 0, 0, 2, 0, 0, 0, -1, -3, -4, -8, 0, 1, -1, -1, 1, -1, 0, 0, 1, 0, 2, 0, 0, 0, -2, 0, 1, 2, 0, 1, 4, 1, 2, -1, -1, 0, -1, -1, -2, -5, 1, -1, 1, 0, 1, -1, 0, 2, 0, 1, 2, 3, 3, 1, -2, 0, 1, 2, 1, 3, 1, 1, 2, 1, 1, -1, -1, 0, -3, -4, 2, -1, 1, -1, 0, -2, 0, 0, 0, 3, 0, 2, 2, 1, -1, 1, 0, 4, 4, 1, 3, 1, -1, -1, 0, 0, -2, -3, -1, -3, 0, 0, 0, 0, 1, 0, 0, 0, 1, 2, 0, 0, 3, 0, -1, 0, 3, 3, 4, 1, 4, 4, -1, 1, 0, 0, 0, -1, -2, -4, 1, 0, -1, 0, 0, 1, 1, 0, 1, 0, -1, 0, 0, -1, 0, 0, 1, 1, 5, 1, 5, 0, -1, 1, -1, -1, 1, 0, -1, -5, -1, -1, -2, 0, -1, 0, -1, 0, 1, 1, 2, 2, 1, 0, -1, 0, 0, 2, 4, 0, 4, 0, -1, -1, -1, 0, -1, -2, -5, -5, -1, 0, -1, 0, -1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, -1, 2, 0, 3, 0, 2, 4, 0, -1, 0, 0, 0, -2, -2, -6, 0, -1, 0, 0, -2, 0, 0, 1, 1, -1, 1, -1, -1, 0, 0, 2, 2, 0, 1, 1, 2, 1, -1, -1, -2, -1, 0, -1, -4, -5, 0, 0, -2, -2, -2, 0, -1, 0, 3, 0, -1, -1, 0, 1, 0, 1, 0, 3, 0, 2, 1, 0, 1, 0, 0, -1, -1, -3, -3, -4, 1, 1, 0, 1, 0, -1, -1, 0, 1, -1, -1, -1, 0, 1, 2, 0, 2, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, -4, -4, -8, 1, 0, 0, 0, 0, 0, -1, -2, -2, 1, -1, -2, -1, 0, 0, -2, 0, 0, 3, 0, 2, -2, -1, 0, -3, -2, -2, -2, -7, -6, 0, 0, 0, 0, -2, 1, -2, -2, 0, -1, -1, -1, 0, -2, -1, -2, -1, 0, -2, 1, 0, 0, 0, -3, -3, -2, -4, -5, -6, -10, 1, 2, 1, 0, -1, -1, -1, -2, 1, -1, 0, -2, -2, -4, 0, -2, -4, -3, -2, 0, 0, 1, -2, 0, -3, -2, -1, -3, -6, -7, 2, 0, 0, 0, 1, 0, -1, 0, -1, -2, 0, -2, -3, -3, -2, -1, -2, -4, -3, -1, -1, -1, 0, -2, -2, -5, -2, -6, -4, -9, 2, 2, 0, 0, -2, -1, 0, -1, -2, 0, 0, 0, -2, -4, -1, -4, -1, -4, -2, -2, -3, -4, -2, -4, -3, -5, -7, -8, -7, -7, -2, 1, -1, 0, 0, 0, 0, -2, -1, 0, -1, 0, -1, -3, 0, -1, 0, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 0, 0, 1, -2, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, -2, 0, -2, 0, 0, -2, 0, 1, -1, 0, 1, -1, -1, 1, -1, 0, 0, -1, 0, 1, 0, -2, -2, 0, -1, -1, 0, -1, 0, -2, -2, -2, 0, -2, 0, 0, -1, -1, 1, 1, 0, 0, 1, 0, -1, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, -1, -3, -1, -2, -2, 0, -1, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, 1, 1, -1, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, -3, 0, -1, -1, -2, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, -1, -2, -1, 0, -2, 0, -1, 0, 0, 0, 0, 0, -3, 0, 0, -1, 0, -2, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -3, 0, 1, 0, 0, 0, 0, 0, -1, 1, -1, -2, -2, -1, 0, 1, -1, 1, 0, 0, 0, 1, 0, -2, 0, 0, 0, 0, -2, 0, 0, -1, 0, -2, 0, 1, 1, 0, 1, 0, 0, 1, 0, -1, 0, 0, -1, 1, 0, 1, -2, 0, 1, 0, -2, -1, -1, -2, -2, -1, 0, -2, -2, 0, 0, -2, 0, 1, 1, 1, -1, 0, 0, -1, -1, 1, -2, 0, 0, 0, -1, 1, 1, -1, -2, -3, 0, 0, -1, -1, 0, 0, -2, 0, -1, -1, 1, 0, 1, 1, 1, -1, -1, 0, -2, 1, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -2, 0, 0, 0, 1, 1, -1, -2, -1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, 0, 1, 0, -3, -2, -2, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, -1, 0, -1, -1, 1, -2, -1, 0, 0, -2, -2, -1, -2, -1, 1, 0, 0, 0, -2, -3, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -1, 0, 1, -2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 1, -2, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 1, -2, 0, 0, 0, 0, 1, -1, -1, 1, 0, 0, 0, -1, 0, 0, -2, -1, 1, 0, -2, -1, 0, 0, -1, 1, 1, -2, -2, 0, 0, -2, -2, -1, 1, 0, -1, 0, 1, -1, -2, 0, 0, -1, -2, 1, -2, -1, -1, 0, -2, 1, -1, 0, -2, 0, 1, -1, -1, 0, 1, -2, -1, 0, 0, -2, 0, -1, -2, 0, -1, -1, -1, -2, 0, -1, 0, -1, 0, -1, -1, 0, -1, -2, 1, 0, 1, 0, 0, -2, -1, -1, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, 0, -2, -1, -1, 0, 1, 0, -1, 0, 1, 1, -1, 0, 0, -1, 0, -1, 0, -2, 0, -1, -2, 0, 1, 0, 0, 0, -2, -2, -3, 0, 0, -1, 0, -2, 0, -1, -1, 0, -2, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, -2, -3, 0, -2, -1, 0, 0, -1, -3, -1, 0, 0, 0, -2, -1, -2, -1, -1, 0, 0, 0, 2, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, -2, 0, -2, -1, -2, 0, 0, 0, 0, -1, -1, 0, 2, 1, -1, 1, -1, 0, -1, 0, 0, 1, -1, -2, -2, -1, 0, 0, 0, -3, -1, -1, -1, 0, 0, -2, 0, -2, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, -2, -1, -1, 0, -1, 0, 0, -1, 0, -2, -2, 0, 0, -1, -1, -2, 0, 0, 0, -1, 0, -1, -1, 0, -1, 0, 1, 0, -1, 0, 0, 0, 0, -2, -2, -2, -2, -1, 0, -2, 0, 0, -1, 0, -1, 0, 1, 1, -1, -1, 0, -1, -1, 1, 0, -1, -1, -2, -2, -1, 0, -1, -1, -2, 0, -1, -2, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, 1, -1, 0, -2, -1, 1, 0, 1, 0, 0, -2, 1, 0, 0, 0, 0, 0, -2, -2, 0, -2, -1, 0, -1, -2, -2, -1, 0, -1, 0, 1, -1, 1, 1, 0, 1, 1, 0, -1, -2, 0, -1, -2, 0, -2, 0, 0, 0, 0, -2, 0, 0, 0, -1, 0, -2, -2, 0, 0, 1, 1, 1, -1, 0, 0, -1, 0, 0, 1, -1, -1, 0, 0, 0, 0, -1, -1, 0, 1, -1, 0, -2, -2, -1, -2, -2, -2, -1, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 0, -1, 1, 0, 0, 0, -1, -2, 0, 0, -1, 1, 0, 0, -1, -1, -2, -1, -1, 0, 0, -2, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, -2, 0, 0, 1, 0, -2, 0, -1, -1, 0, 0, 0, 0, -2, 1, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -2, 0, 0, -1, 0, -2, -1, 0, 0, 0, 0, 0, -2, 0, -2, -2, 0, -2, 0, 0, -1, -2, -1, 0, -1, -1, -2, 0, -3, 0, -2, 0, 0, 0, 1, -2, 0, 0, 0, -1, 0, -1, -1, 0, -2, -1, -1, 0, 0, 0, 0, -1, -2, 0, -1, -1, -1, 0, -3, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1, -1, -1, -2, -1, -1, -2, 0, 0, 0, -2, -2, 0, 0, 0, -1, -1, -3, -2, 0, -2, -2, 0, -1, 1, 1, 0, 0, 0, 0, -2, 0, -1, 0, 0, 0, 1, 0, 0, 1, -2, 0, 0, -1, -2, -2, -2, 0, 0, -2, 0, 0, 0, 0, -2, 0, 0, -1, -2, -2, -2, 1, 0, -1, 1, 0, 0, 1, -2, -2, 1, -1, -1, -1, -2, -1, 1, -1, 0, 0, -2, 0, -1, -1, -1, -1, 1, 0, 0, -1, 1, -1, 0, -1, 0, 0, -2, -1, 1, -1, -2, 0, 0, -1, 1, -1, -1, -1, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -1, -1, 1, -1, 0, 1, -2, 0, 1, 1, -1, 0, 2, 1, 1, 0, 0, -1, 0, 0, -1, -1, 1, 1, -2, -1, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, -2, -1, -1, 0, 0, -1, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 1, -1, -1, 0, 1, 0, 0, 0, 0, 0, 0, -3, -1, 0, 0, 0, -3, 0, -2, 1, 0, 1, 1, 0, -1, 1, -1, -2, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -2, -1, -2, -1, 0, -1, 0, -1, -1, 0, 0, 1, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, -2, 1, 0, -1, -1, 0, 0, -1, 0, -2, 1, -1, -1, 0, -2, 0, 0, -2, -1, 1, 0, 2, 0, 1, 1, 0, 0, 0, 0, -1, 1, -1, 0, -1, 1, 1, -1, -1, 0, 0, -2, 0, 0, 0, 0, -2, 0, 0, 0, 1, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, -2, -2, 1, 0, -1, 0, 1, -2, 0, 0, -1, 0, -2, 0, 0, -2, 0, 0, -1, -2, 0, -1, 0, 0, 0, 0, -2, 0, 0, 0, 0, 0, -2, 1, 0, 0, -2, 0, 1, -1, 0, -1, 0, 0, -2, 0, -1, -2, -1, -2, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 1, -1, -1, 0, 1, -1, -1, 0, 0, -2, -1, -2, -2, 1, -2, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -2, -1, 1, 0, 0, -1, 0, -1, -1, -2, 0, 0, -1, -1, 0, -3, -2, -2, 0, -2, -2, -1, 1, -1, -1, 0, 1, 1, -2, -2, 0, 0, 1, -2, 0, -1, 0, 1, -1, 1, -1, 0, -1, 0, 0, 0, -2, 0, 0, 0, -1, 0, -1, 0, 0, -2, -1, -1, 0, -1, 0, 0, -1, 0, 1, 0, 1, -2, -2, -1, -1, -1, 0, 0, -2, -3, -2, -2, 1, 0, 0, 0, -1, 0, 0, -1, 1, -2, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 1, 0, 0, -2, 0, -2, -2, -1, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, -2, 0, 0, -1, 0, -1, 0, -1, -2, 1, -1, 0, -2, -1, -1, -2, -2, 0, -1, -2, 0, -1, -1, 0, 0, -2, 0, 0, 0, 0, -2, 0, -2, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, -2, -2, 0, -2, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 1, -2, -2, -1, 0, -1, 0, 1, 0, -2, 1, -1, -2, 0, -2, -1, 1, -1, 0, -2, -1, -2, 0, -1, -2, 0, 1, -1, -1, 0, 1, 0, -1, -1, -2, 0, -1, -1, 0, -1, 0, 0, -2, 0, -1, -1, -2, 0, 0, -2, -1, 0, -1, -1, 0, 0, 0, -2, -1, 0, -2, 0, 0, -2, -2, -1, -2, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -1, -2, -1, 0, 0, -1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -2, 0, 0, -2, -1, 1, 0, 0, -2, -2, 0, -2, 0, 0, -2, 0, -2, -2, 0, 0, -2, 0, 0, -2, 0, 0, -2, 0, 0, -2, 0, 1, -2, 0, -2, 0, -2, -1, -2, 1, 0, 0, 0, 1, 1, -1, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, -3, -2, -1, 0, -2, 0, -2, -1, -1, -1, 1, -2, 0, 1, -2, 0, 0, 1, -1, -1, 0, 0, 1, -1, 0, -1, -2, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, -2, 0, 0, -2, -2, 0, 0, -1, 0, 0, -1, -1, -1, 0, 1, 1, 0, 0, -2, -1, -1, 0, -1, 0, 0, -2, -1, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, -2, -2, 0, 0, 0, 1, 0, -2, 0, -1, -3, 0, -1, 0, -2, -1, 0, -1, 0, 0, -1, 0, 1, -2, 0, 0, -3, -2, 0, -3, 0, -2, 0, -2, 0, -2, 0, -3, 0, 0, -1, -1, -2, -1, 0, 0, -1, 0, -2, 0, 0, -1, 1, 0, -2, 1, 0, 0, -3, 0, 1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 2, -1, -1, 0, -2, 0, 0, -1, -1, 0, 1, 0, -1, -1, 0, 0, 0, -1, 0, -1, 0, -1, 1, -2, -1, -1, -2, 1, 0, 0, 0, 0, -2, -1, 0, 0, 1, 1, 0, -1, 0, 2, 0, 1, 0, 0, -1, -2, 0, -1, 0, -2, 0, 1, -1, -2, 0, 0, 1, 2, -1, -1, 1, -2, 0, 1, 1, -1, 1, -1, 0, 1, -1, 2, 0, 0, 0, 0, 1, -2, 0, 0, 0, 0, -2, 1, 1, 0, 0, 2, 0, 0, -1, -1, 1, -1, -1, 0, 1, 0, -1, 0, 0, 0, -1, 1, 0, 1, 0, 0, 0, 0, -2, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, 1, -1, -2, 0, 0, 1, -2, 1, 2, 1, -1, 1, 1, 1, -1, 1, -1, 1, -1, -2, 0, 0, 1, 1, 2, 0, -1, 2, 1, 1, 2, 0, 1, 1, 0, -1, 0, -1, 0, -1, 0, 2, 0, 0, 0, -1, 0, -1, 0, 0, -1, 0, 1, 0, 2, 0, -1, 0, 1, 0, -1, 0, 0, 2, 0, 0, 0, 1, 1, 2, 1, 0, 0, 2, 1, 1, -2, -1, -1, 0, -2, -1, -1, 1, 2, -1, 2, 1, 1, 1, 0, -1, -1, 1, 0, -1, -1, -1, -1, 2, -1, 1, -1, 1, 1, 1, -2, -1, -1, 0, -1, 1, 0, -1, 1, 1, 0, 1, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 1, 1, -1, 0, 0, 1, 0, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 2, 1, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, -1, 0, -1, 0, -1, 0, 0, 0, 0, 0, -2, 1, -1, -1, 0, 0, -2, 0, 1, 2, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 0, 1, 0, 1, 2, 1, -1, 0, 0, 0, 0, 1, -1, -1, 0, -1, -1, 1, -1, -1, 0, 2, 1, -1, 0, 0, 1, 0, -1, -1, 1, 1, 1, 0, 0, -1, -2, -2, 0, 0, -1, 0, 0, 1, -1, 0, -2, -1, 0, 0, 1, -1, 1, 0, -1, 1, 0, 0, 0, 0, 1, -1, 1, 2, 1, 1, 0, 1, 1, 0, 0, 2, 0, 1, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, 1, 0, 0, 0, -1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 2, -1, 0, -2, 1, -2, -2, -1, 2, 1, 2, 2, 0, 1, 0, 1, 1, 0, 1, 0, -1, -1, 0, 1, 0, 2, 1, 1, 0, -1, 1, 0, -1, 0, 0, -2, -1, 1, 2, 2, 0, -1, 0, 0, -1, 0, 2, 0, 2, 0, 2, 0, 0, 1, -1, 0, 1, -2, 0, 2, -1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 0, 2, 0, 1, 1, -1, 1, 1, 0, 0, 0, -1, 0, 0, -2, -2, 0, 0, 0, -2, -1, -2, -2, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, -1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 0, 0, 1, 2, -1, 0, 0, 0, 1, 0, 0, 1, 3, 0, 0, 0, 0, -1, -1, 1, 1, 0, 1, 1, 1, 1, 0, -1, -1, 0, 0, 1, 0, 2, 0, -1, 0, 0, -1, 0, 2, -1, 0, 1, 0, 1, 0, 0, -1, -1, 0, -1, 0, 1, 0, 1, 0, 0, 0, 0, 0, 2, 1, 0, 2, 0, 2, 0, 1, 0, 0, 0, 2, 0, 1, 2, 1, -1, 1, 0, 1, 1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, 2, 0, -2, 1, 2, -1, -1, 0, 0, 2, 1, 1, 1, -1, -2, 1, 1, 1, 0, 0, 0, 2, 0, 0, -1, -2, 1, 0, 0, -1, -1, 0, 0, -1, 1, 0, 0, 2, 0, 1, 2, 0, -1, 0, 0, -1, 1, -2, -2, -2, 0, 0, 0, 1, 0, -1, 0, -1, 1, 0, 1, 1, 0, 2, 0, -1, 1, 0, 0, 1, 1, 2, 0, -1, -2, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, 1, 1, 1, 2, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, -1, 0, -1, 0, 0, 0, 1, -1, 0, 1, -1, 0, 1, 1, 0, -1, 0, -1, 1, 2, 0, 2, 0, 0, 1, 1, 2, 1, 2, 0, -2, 0, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, 1, 2, -1, 1, 2, 0, 3, 1, 2, 3, 0, 1, 1, 0, 0, 0, 1, -2, 0, 0, 0, 0, 1, 0, -1, -2, -2, 0, 0, -1, 1, 0, 2, 0, 0, 1, 0, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 1, 2, -1, -1, 0, 0, 0, 0, -3, -3, -6, -3, -3, -4, -9, -8, -9, -9, -9, -7, -7, -9, -8, -10, -8, -8, -8, -11, -12, -15, -18, -18, -20, -23, -24, -26, -26, -31, -3, -7, -5, -6, -7, -7, -7, -7, -5, -5, -6, -9, -5, -7, -8, -9, -6, -7, -4, -5, -7, -7, -9, -12, -13, -19, -21, -23, -25, -26, -6, -5, -6, -3, -4, -3, -3, -5, -3, -7, -6, -7, -7, -4, -5, -3, -4, -2, -4, 0, -3, -3, -3, -8, -9, -13, -14, -18, -22, -26, -3, -4, -3, -6, -4, -5, -4, -2, -5, -5, -6, -6, -4, -3, -3, -5, -1, 0, 0, -2, -1, 1, 0, -3, -4, -6, -13, -18, -18, -22, -3, -5, -5, -5, -4, -3, -1, -2, -2, -3, -2, -3, -3, -4, -2, -1, 1, 0, 0, 2, 3, 2, 1, 2, -2, -3, -8, -14, -16, -22, -4, -3, -6, -2, -2, -3, -2, -4, -3, -3, -1, 1, 0, -1, 1, 0, 0, 1, 3, 3, 2, 2, 5, 1, -2, -3, -8, -12, -15, -21, -4, -4, -5, -2, -4, -3, -2, -4, 0, -4, -2, -1, 0, 0, 1, 1, 1, 4, 2, 2, 6, 5, 4, 3, 0, -1, -4, -8, -14, -18, -6, -2, -6, -4, -2, -4, -3, -2, -1, 0, 0, 0, 2, 2, 1, 3, 4, 3, 2, 3, 7, 7, 4, 1, -1, -5, -6, -7, -16, -17, -3, -3, -6, -4, -6, -3, -5, -4, -3, 0, 0, 3, 1, 5, 3, 1, 5, 7, 7, 5, 6, 7, 5, 2, 0, -2, -3, -8, -14, -17, -4, -4, -3, -4, -5, -6, -2, -1, 0, 0, 0, 3, 3, 1, 4, 5, 3, 6, 5, 6, 6, 5, 3, 3, 0, -3, -4, -10, -11, -15, -3, -3, -6, -6, -4, -7, -2, -1, -2, -2, 0, 2, 4, 1, 2, 2, 5, 7, 4, 5, 8, 4, 4, 5, 0, -2, -2, -9, -12, -16, -4, -6, -3, -5, -5, -3, -1, 0, 0, 1, 0, 2, 2, 1, 2, 3, 3, 3, 4, 6, 6, 5, 7, 3, 2, 0, -4, -6, -11, -18, -4, -7, -4, -3, -3, -5, -3, -2, 1, 0, 3, 5, 3, 3, 0, 1, 3, 3, 1, 2, 4, 4, 4, 2, 3, -1, -3, -5, -12, -16, -5, -3, -4, -5, -4, -3, -4, -3, 1, 2, 5, 4, 1, 1, 2, 2, 0, 4, 1, 2, 6, 5, 4, 5, 2, -2, -3, -7, -13, -18, -4, -2, -4, -3, -5, -3, 0, 1, 0, 2, 4, 4, 2, 0, 0, 1, 0, 4, 3, 1, 6, 6, 4, 1, 3, 0, -5, -9, -10, -16, -3, -2, -5, -6, -2, -3, -1, -1, 0, 1, 3, 3, 0, -1, 0, 0, 4, 2, 4, 2, 5, 5, 3, 4, 2, -1, -1, -9, -10, -17, -2, -4, -3, -4, -2, -2, 0, 1, -1, 3, 4, 3, 3, 0, 0, 3, 3, 6, 5, 6, 5, 5, 2, 4, 2, -2, -2, -9, -12, -14, -2, -4, -6, -6, -3, -2, -2, -1, 1, 2, 3, 2, 3, 1, 0, 0, 5, 4, 7, 5, 3, 3, 2, 2, 1, 0, -4, -9, -13, -15, -4, -2, -2, -3, -5, -3, -1, 1, 0, 0, 1, 0, 2, 0, 0, 1, 6, 7, 5, 7, 6, 5, 2, 3, 0, 0, -5, -8, -11, -15, -4, -5, -4, -5, -3, -1, 0, -1, -1, 0, 1, 1, -1, 2, 0, 1, 6, 4, 6, 6, 8, 7, 2, 2, 3, 0, -5, -9, -12, -18, -6, -7, -4, -4, -2, -1, 0, 0, -2, 0, 0, -1, -1, 0, 0, 3, 4, 5, 6, 5, 5, 4, 4, 2, 0, 0, -4, -8, -12, -16, -3, -6, -3, -4, -4, -4, -1, -1, -2, 0, 0, -1, 1, 1, 0, 2, 4, 4, 6, 6, 5, 3, 2, 3, 0, -4, -7, -11, -14, -17, -3, -2, -6, -5, -2, -3, -3, 0, 0, -4, -2, 0, 0, 1, 0, 1, 2, 2, 3, 6, 7, 2, 4, 0, 0, -4, -7, -12, -14, -19, -3, -5, -4, -3, -4, -4, -2, 0, -1, -2, -1, -3, 0, 0, 1, 2, 3, 4, 2, 5, 3, 2, 2, 1, -2, -4, -7, -14, -15, -22, -6, -2, -4, -6, -3, -5, -3, -4, -2, -4, -2, -2, 0, 0, 0, 0, 0, 2, 3, 2, 2, 1, 2, 0, -4, -4, -11, -11, -16, -23, -4, -6, -7, -4, -3, -4, -4, -3, -3, -5, -5, -5, -3, -2, -2, -1, 1, 2, 2, 0, 3, 0, 0, -4, -3, -6, -11, -17, -21, -22, -3, -6, -3, -3, -4, -6, -3, -4, -4, -2, -3, -3, -3, -5, -5, -2, 0, -1, 1, 1, 0, -2, -4, -5, -7, -9, -14, -18, -20, -23, -3, -2, -5, -5, -7, -5, -7, -2, -6, -5, -3, -6, -7, -7, -7, -8, -5, -3, -4, -2, -4, -4, -9, -9, -9, -12, -18, -21, -24, -26, -3, -6, -3, -5, -3, -3, -6, -5, -2, -6, -6, -6, -9, -9, -7, -8, -7, -6, -10, -9, -10, -10, -12, -11, -14, -19, -18, -21, -25, -29, -5, -5, -3, -4, -5, -3, -4, -4, -3, -6, -7, -7, -9, -7, -10, -10, -11, -12, -11, -14, -12, -13, -15, -17, -17, -20, -24, -25, -26, -31, -2, 0, 0, 0, -1, -1, -2, 0, 0, 1, 0, -2, -2, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, -1, -1, -2, 0, 1, 1, 0, 0, -2, 0, 0, -1, -1, 0, 0, -2, 1, 0, 1, -1, 0, -2, 1, 0, -1, 0, 1, 0, 1, 0, 0, 0, -1, 0, -1, 0, -1, -1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 1, -2, -1, -1, -1, 1, 0, 0, 0, -1, 0, 1, 0, -1, 1, -1, -1, -2, -1, 0, 0, 1, 0, -2, -2, 0, 1, 1, 0, 1, -2, 0, 1, 0, 1, 0, 0, 0, 0, -2, 0, 0, 1, 0, -1, -2, -1, 0, 0, -1, 0, 0, 1, 0, -1, 1, 1, -1, 0, -2, -1, -1, 0, 0, 0, -1, 1, 0, -1, -1, -2, 0, -1, -1, 0, -2, 0, 0, -1, 0, -2, 0, 0, -1, -2, 1, 0, -2, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, -2, 0, -2, -1, 0, -1, 1, 1, 1, 1, -2, 1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -2, 0, 0, 1, 0, 0, -2, -1, 1, -2, -1, -1, -1, 0, -2, -2, -1, 0, -1, -2, 0, -1, 0, -2, 0, -1, 0, -2, 0, 0, 0, 0, -2, -2, -1, 1, -1, 0, 0, 1, 0, -2, 0, 0, 0, 0, 0, -2, -1, 1, 0, 0, 0, 0, -1, 0, 0, -2, -1, 1, 0, 0, 0, 0, 0, -1, 0, 1, -2, -2, 0, 0, 1, 0, 0, 0, -2, 0, -2, -1, -2, 0, -2, -1, -2, -2, -1, 0, 0, 1, 0, 0, -2, 0, 0, -1, -2, 1, 0, 0, 1, 0, -2, -2, -2, 0, 0, -1, -1, 0, -1, 1, 0, 0, -1, 0, -1, 0, 0, -1, 1, -2, 0, 0, -1, 0, 0, 0, -1, 1, -2, 0, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, -2, 0, 0, 0, 0, -1, 1, -2, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 0, 1, -1, -1, 0, -2, -2, 1, 0, -1, 0, 1, -2, -1, 1, 0, -1, -1, -1, 0, 1, 0, 0, 1, -2, -1, 0, -1, 0, 0, -1, 1, -1, 1, 1, 0, 0, -1, 1, 0, -1, -1, -2, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, -2, 0, -1, -1, 0, 1, 0, 0, 0, 1, -2, -1, -2, -1, 1, 1, 0, 0, -1, -2, 0, 0, -2, 0, 0, -2, 0, 0, -1, -1, -1, 1, 0, 0, -1, 0, 0, -2, 0, -1, 0, 0, 0, -2, 0, -1, -1, 0, -1, 0, -1, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, -1, -2, 0, 0, -2, 0, 0, -1, 0, 0, -1, -2, 0, -1, -1, -1, -2, -1, 0, 0, 0, 0, -2, 0, 1, 1, 0, 0, 1, 0, -1, -1, 0, 0, -1, 1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, -2, 0, 1, 1, 0, 0, 0, 0, -1, 0, -2, 0, -1, 1, -2, -1, 0, -2, 1, 1, 0, 1, 0, 0, 0, -1, 0, -2, 0, 1, -1, 0, 1, 1, 0, 1, 0, -1, -1, 0, -2, 0, -1, -1, 0, -1, -1, 1, -1, 0, -1, 0, 0, -2, -1, -2, 0, 1, 0, -1, 1, 0, -1, -1, 0, 0, -2, 0, 0, -2, 1, 0, 0, 0, -2, -2, 0, 0, 0, -2, 1, 0, 0, 0, -2, -1, 0, 0, 0, 0, 1, -1, -1, -1, 1, 0, 1, 1, -2, -1, -1, -2, 0, 0, 1, 1, -1, 1, 0, -1, -2, 0, -2, -1, 1, 0, 0, 0, 0, -2, 0, -2, 1, 0, -1, -1, 0, 1, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, -2, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, -2, 1, -1, -2, -2, 0, 0, 1, -1, 1, -1, -1, -2, 1, 0, 1, -1, 0, -2, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 1, 0, -2, 1, -2, -1, -1, -1, 0, 0, -2, 1, 1, 0, -2, -2, 0, -1, -1, 0, 0, -2, 0, -1, 0, 1, -1, -1, 0, 0, 0, 1, 0, 0, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 1, 1, -2, -2, -1, 1, 0, 1, 1, 0, -1, 0, -1, 1, 0, -1, -1, 1, 1, -2, -1, 0, 0, -1, -2, -1, 1, -1, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0, 0, -1, 0, 1, -1, 0, -1, 1, 0, 1, 0, 0, -1, -1, -1, 0, 0, 1, -2, -1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 0, -1, -2, 1, -1, 1, 0, 1, 0, 0, 0, 0, 0, -2, -2, 0, -1, -2, 0, 0, -2, 1, -1, 0, 1, -1, 0, 0, -1, 0, 1, 0, 0, 2, 0, 0, -1, 0, 0, -2, 0, -1, 1, -1, 1, -1, -1, 0, -1, 0, 0, 0, -1, 0, -2, 0, 2, -1, -2, 0, 0, -1, -1, 0, 0, -1, 0, -1, 1, 1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 2, 2, 1, 0, 1, 0, 1, 0, -1, 0, 1, 1, 1, 0, 0, 1, 0, -1, -1, 1, 2, 0, 1, 1, 1, -1, 1, 1, -1, -1, 1, 0, 1, -1, 1, 2, 0, 0, -1, 0, -1, -1, 1, 1, -1, -1, -1, -1, 0, 0, 1, -2, 2, 0, 0, -2, -1, -1, -1, 0, 2, 0, 1, 1, 0, -1, 0, 1, 2, 0, 0, 1, 0, 1, -1, 0, -1, 0, 0, 1, 0, -1, 0, 0, 1, 0, -1, 2, -1, 0, 0, 1, -1, 0, 1, 0, 0, 1, 2, -1, -1, -1, 1, 0, -1, -2, -1, 0, 0, 1, 0, 1, 1, 0, -1, 1, 0, 0, 0, 0, -1, 1, 1, 0, 0, 2, 0, 1, 1, -1, 0, 2, 0, 0, 0, 1, 0, 2, 0, 1, 1, 1, 0, -1, 1, -1, 0, -1, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 0, -1, -2, 1, 1, 0, 0, 0, -2, -1, -1, 0, 0, -1, 0, -1, 1, 1, -1, 0, 1, 0, -1, 2, 0, 0, 0, 1, -2, -1, 0, -1, 1, 1, -1, 0, 1, 0, 1, -1, 0, 0, 0, 1, 0, -1, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 0, 1, 0, 0, 1, -2, 0, -1, -1, -1, 1, -1, 0, 0, 1, -1, -1, 0, 0, 0, 1, 0, -1, 1, 1, -1, 1, 1, 2, -1, 2, 0, 1, -1, 0, 1, -1, 0, 0, 1, 1, -2, 0, -1, 0, 1, 0, 1, -2, 0, -1, 1, 0, 2, -1, 0, -1, 0, 0, 0, 0, -1, -1, 0, 1, 2, 0, -1, -1, -1, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 2, -1, 1, 0, 1, -1, -1, -1, 0, 0, 0, 0, 1, 0, -2, -1, 0, 0, 0, -1, -1, -1, -1, -1, 0, 1, 1, -1, 0, 0, 0, -1, 1, 1, -1, 0, 0, -1, 1, -1, -1, -1, 0, 0, 0, -1, 0, 1, -1, 1, 0, 0, 1, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 1, -1, -1, -1, 1, 0, 1, 1, 0, 0, 0, 2, 0, 1, 1, 0, 1, -1, 1, -1, 0, 0, -1, 0, 1, 0, -1, -1, 0, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, -1, 1, 0, -1, -1, 0, 0, -2, 1, 0, 0, -1, 0, 1, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 2, 1, -1, 2, 1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -2, 1, -1, 0, -2, -1, 0, -1, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, -1, -1, -1, 1, -1, 1, 0, 0, -1, 2, -1, 0, 0, -1, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, -1, 1, 0, 0, 1, -1, 0, 0, 0, 0, -1, -1, 1, -1, -1, 0, -1, 1, 1, -1, -1, 0, 0, -2, 0, 0, 0, 0, -1, 0, -1, 0, 0, 1, -2, 1, 1, -1, -1, 0, 0, -2, 0, -2, 0, -1, 0, 1, 0, 0, -2, 0, 1, -2, -1, 0, 1, -1, -2, 1, 0, 1, 0, 0, -1, 0, 1, 1, 0, 0, -1, -1, 0, 1, 0, 0, 0, 0, -1, 0, -1, -1, -1, 1, 1, 0, -1, 0, 1, -1, -1, 0, 0, -1, -1, 0, 1, -1, 1, 0, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, -1, 0, 0, 0, -1, 1, 0, -1, 0, 1, 0, 0, -1, 2, 0, -1, 0, -1, -1, -2, 0, 0, 0, -1, -1, 0, -1, 1, 0, -2, 0, -1, -1, 0, -2, 0, 0, -1, 1, -1, -1, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 2, 1, -1, 0, -1, -1, 1, 1, 0, 0, -1, 0, 1, 1, 0, 2, 1, 0, 2, -1, 0, 0, -1, 0, 1, 1, -2, 2, 2, 1, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, 0, -1, 1, 0, 0, 0, -2, 0, 1, 1, 0, -1, -1, -1, -1, -2, 0, -2, 1, 0, 0, 0, 0, 0, -1, 1, 0, 0, 0, -2, 1, -2, 0, -1, 0, 0, 1, -1, 1, 0, 2, 1, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 0, -1, 1, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, -1, -1, -2, 0, -2, 0, 0, -1, -1, 0, 0, -1, 1, -1, 0, 0, 0, 0, 0, 0, 2, 0, -1, 1, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 1, 0, 0, 0, 4, 3, 2, 1, -1, 0, -1, -2, -2, -6, -5, -5, 0, -1, 2, -1, -1, 2, 4, 2, 3, 4, 1, 2, -1, -2, -4, -5, -4, -7, 4, 0, 0, 1, 0, 0, 1, 0, 0, -4, -5, 0, -1, -1, 0, -1, -1, 0, 3, 2, 2, 5, 3, 5, 3, 0, 2, -1, -3, -6, 2, 2, 3, 2, 3, 0, 0, 1, -1, -2, -3, 0, -1, -1, 0, -2, -3, -2, 1, 0, 3, 4, 4, 2, 4, 3, 5, 0, -3, -8, 5, 1, 3, 0, 1, 1, 2, 1, 1, 2, 1, 1, 0, 2, -2, -2, 0, -3, -2, 0, -2, 0, 0, 2, 2, 3, 5, 0, 0, -5, 4, 5, 2, 1, 3, 1, 1, 0, 3, 0, 1, 0, 0, 0, 2, 0, 0, -3, 0, -2, -2, -1, 0, 3, 4, 2, 3, 0, -3, -7, 5, 4, 2, 3, 2, 4, 3, 0, 3, 2, 2, 2, 3, 0, 0, 0, 0, -2, -2, -5, -4, -2, 0, 0, 3, 2, 2, 0, -2, -11, 5, 1, 2, 0, 1, 2, 2, 1, 2, 1, 0, 3, 2, 3, 2, 0, 0, 0, -4, -2, -4, -3, 0, 1, 0, 0, 0, -1, -5, -8, 1, 4, 1, 2, -1, 2, 1, 2, 2, 2, 4, 5, 2, 3, 0, 1, -1, 0, -2, -1, -3, -2, 0, 0, 0, -1, -1, -2, -5, -7, 0, 3, 2, 1, 0, 2, 1, 1, 4, 3, 2, 2, 4, 2, 2, 0, 1, 2, 0, 1, -1, 0, 0, -1, 0, -2, 0, -1, -5, -7, 0, 2, 2, 1, -1, 0, 0, 1, 5, 6, 5, 6, 3, 3, 1, 3, 1, 1, 3, 1, 0, 0, 1, 0, -2, 0, -2, -1, -6, -8, 1, 1, 2, 0, 0, 0, 2, 1, 3, 7, 6, 4, 6, 5, 1, 0, 4, 2, 2, 1, 1, 0, 1, 0, 0, 0, -2, -2, -4, -8, 0, 2, 0, 0, -1, -1, 3, 4, 6, 8, 5, 7, 5, 4, 1, 2, 3, 0, 1, 1, 3, 0, 2, 0, 1, -3, 0, -3, -7, -8, 1, 0, 1, 0, 0, 0, 1, 4, 6, 5, 5, 7, 3, 0, 1, 0, 3, 1, 0, 2, 3, 0, 0, 0, 1, 1, -2, -3, -6, -9, 0, 2, 1, 2, 1, 1, 1, 3, 5, 6, 6, 5, 1, 1, 0, 2, 2, 1, 3, 4, 3, 1, 2, -1, -1, 0, -1, -2, -4, -11, 2, 1, 3, 0, 0, 3, 3, 3, 7, 4, 5, 4, 0, 0, -1, 2, 1, 2, 5, 4, 4, 2, 1, 1, 1, 0, 0, -2, -4, -9, 3, 1, 0, 0, 4, 3, 4, 5, 4, 5, 7, 2, 0, -1, 0, 1, 5, 7, 5, 5, 1, 3, -1, -2, 0, 0, -1, -1, -4, -8, 0, 4, 1, 1, 0, 2, 3, 3, 6, 4, 4, 5, 1, 0, 1, 2, 6, 6, 5, 5, 1, 0, 0, -2, 0, 1, 0, -3, -5, -8, 3, 1, 3, 0, 0, 3, 5, 5, 6, 5, 4, 2, 2, 0, 1, 1, 5, 9, 8, 2, 3, 0, -2, -3, 0, 0, -1, -2, -4, -10, 3, 1, 2, 0, 0, 3, 5, 3, 5, 5, 2, 1, 0, -1, 1, 2, 4, 5, 3, 5, 3, 0, -1, -1, 0, 1, -1, -1, -1, -11, 2, 3, 0, 2, 2, 0, 3, 7, 2, 3, 2, 3, 0, 0, 0, 1, 3, 3, 2, 1, 2, -3, -4, -3, 1, 0, 2, 0, -3, -8, 2, 0, 1, 0, 1, 4, 4, 3, 4, 2, 3, 0, 1, 1, 1, 0, 4, 5, 2, 1, 0, 0, -3, -3, -1, 0, 2, -1, -3, -8, 0, 0, 0, 0, 1, 1, 5, 6, 1, 3, 2, 4, 1, 1, 2, 0, 5, 3, 0, 0, 0, 1, -1, -3, -1, 0, 1, 0, -5, -10, 1, 1, -1, 0, 1, 0, 2, 1, 1, 2, 4, 0, 3, 4, 1, 5, 2, 0, 0, -1, 1, -3, -1, 0, -3, -1, -1, -1, -5, -8, 3, 0, 1, -1, 1, 0, 2, 3, 3, 3, 2, 2, 3, 1, 3, 4, 0, 0, -1, 0, 0, -1, -2, -3, 0, 1, -2, 0, -7, -8, 2, 0, 0, 0, -1, 0, 1, 3, 4, 4, 2, 1, 2, 4, 4, 0, -1, 2, -1, 2, 0, 0, -1, -1, -3, 1, -1, -4, -4, -12, 2, 0, 0, 0, 0, 0, -1, 0, 3, 3, 1, 2, 0, 1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1, 2, 1, -1, -3, -8, 3, 2, 0, 0, 0, -1, -2, 1, 2, 1, 2, -1, -1, -2, -1, 0, -3, -3, 0, 3, 2, 1, 2, 3, 3, 0, 2, 0, -4, -10, 4, 3, 1, 3, 0, 1, -1, 1, 0, 3, 0, -1, -2, 0, -1, -3, -3, -2, 1, 2, 2, 1, 0, 2, 2, 3, 2, 1, -6, -10, 5, 4, 1, 2, 0, -2, 0, 0, 2, 3, 0, -1, 0, -2, -2, -2, 0, -1, 0, 3, 5, 5, 3, 4, 2, 3, 1, 0, -6, -8, 5, 5, 4, 0, -1, -1, 0, -1, 0, 1, -2, -1, -2, 1, -1, -1, 1, 1, 5, 4, 3, 4, 4, 1, 1, 0, 0, -1, -3, -9, 0, 0, 1, 0, 1, -1, -2, 0, 1, 1, 1, 0, 1, 0, 1, 0, 0, 1, 1, 2, 0, 3, 4, 1, 1, 0, 2, 2, 0, -2, 0, 1, 0, 2, 1, 0, 1, 0, -1, -1, 1, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 2, 2, 3, 1, 3, 1, 3, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, -1, -1, 0, -1, -2, -1, 0, -1, 0, 0, 0, 2, 3, 0, 3, 2, 2, -2, 0, 0, 3, 3, 0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, -1, 1, 2, 2, 1, 0, 0, -1, 0, 2, 0, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 2, 2, 2, -2, 3, 1, 2, 1, 1, 0, -1, 0, 0, 2, -1, 0, -1, -1, -1, -1, -1, 0, 0, -3, -2, 0, 0, 0, 0, 1, 3, 2, 0, 0, 2, 2, 0, 0, 0, 0, 0, 2, 0, -1, 0, 1, 0, 0, 0, 0, 0, -1, -1, -3, -2, -3, 0, -1, 1, 1, 0, 0, 0, -3, 0, 2, 1, 0, 1, 1, 0, 2, 0, 1, 0, 0, -1, 1, 1, -1, 1, 0, 0, -1, -1, -2, -2, -1, 1, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 1, 0, 0, -2, 0, -1, 0, 0, -2, 0, -1, -1, 1, -1, 2, 0, -1, -2, 1, 0, 0, 0, 1, -1, -1, 0, 2, 2, 2, 1, 0, 2, 1, 1, -1, -2, -1, -1, 1, -1, 2, 0, -1, 0, 0, 0, -1, -1, 2, 2, 1, 2, 1, -2, 0, 0, 0, 3, 2, 1, 2, -1, 1, 0, 2, 1, 1, -1, 0, -2, 1, 0, 1, 0, 0, -2, 1, -1, 0, 1, 1, 0, 1, 1, -1, 1, -1, 0, 2, 0, 0, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, 1, 1, 1, -1, -1, -2, 0, 0, 2, 2, 1, 0, 0, 2, 2, -1, 0, 1, 0, 0, -1, -1, 1, 0, 0, 1, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 0, 0, 0, 2, 0, 0, -2, -1, 1, 1, 1, -1, 2, 0, 1, -1, 0, -1, -1, 1, 0, 0, 0, -1, 0, 2, 1, 1, 2, 2, 2, 1, 0, 0, 0, 0, 1, -1, 1, 0, 0, 0, 3, 0, -1, 0, 0, 0, 0, -1, 0, 0, -2, -1, -1, 1, 0, 1, 0, 2, 0, 1, -1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 0, 0, 0, -2, -2, -1, 2, 0, 1, 2, 2, 0, 1, 0, 2, -1, -1, 0, 0, -1, 1, -1, 2, 2, 2, 1, 0, 0, 0, 0, -1, 1, 2, 0, 0, 0, 2, 0, 1, 0, 1, 1, -1, 0, 1, 2, 2, 0, 0, 0, -2, 1, 0, 1, 2, 0, 0, 0, 0, -1, -1, 0, 0, 2, 0, 0, 0, 0, 0, 2, -1, -1, 0, 0, 0, 0, 2, 2, 0, 1, -1, -1, 0, 2, 1, 1, 1, 0, 0, 0, -1, 1, 0, -1, 1, 0, 0, 0, 1, 0, 0, 1, 0, 3, 1, 0, 0, -1, 1, 2, -2, 0, -1, 0, 0, 0, -1, -2, 0, -2, -1, 0, 0, 1, 0, 0, 2, 2, 1, 0, -1, 2, 0, 0, 1, 2, 0, 0, 0, 1, 0, -2, 1, 0, 1, 0, -1, 0, 0, 1, -1, 2, 0, 0, 0, -3, 1, 1, 1, 0, 0, 1, 0, 2, 1, 1, -1, 0, 1, 0, -2, 1, 0, 1, -2, -2, -2, 0, 0, 0, 0, 2, 0, 1, 0, 0, 2, 0, 2, -1, 1, 0, -1, 1, 0, 0, 1, -1, -1, -1, -1, 2, 0, -2, -2, -1, 0, 0, -2, -1, -2, 0, 0, 0, -2, -1, 0, 0, -1, 2, 0, 0, -1, 0, 2, 1, 0, 1, 1, 0, 0, -1, 0, 0, -2, 1, -2, 0, 0, -1, -1, 0, 1, -1, 0, -2, 1, 0, 2, -1, 0, -1, -1, 2, 1, 0, 2, 0, 2, 1, 1, 0, -2, -1, -1, -1, -2, 0, 0, -1, 0, 1, 0, 0, 0, -1, 2, 2, 1, 0, 0, 1, 0, 0, 3, 2, 0, 1, 1, -1, 0, 0, -3, -2, -1, 0, 0, 2, 1, 2, 0, 0, 0, 0, -1, -2, 0, 0, -1, 1, -1, 0, -1, 2, 1, 1, 0, -1, 0, 0, 0, 0, -2, -2, 0, 1, 0, 0, 0, 2, 0, 0, 0, 1, 1, -1, 3, 1, 2, -1, 0, 0, -1, 1, 2, 0, 1, 0, -1, 1, 0, 1, 0, -2, 0, 0, 2, 0, 2, 2, 0, 2, 2, 0, 0, -2, 2, 0, 0, 2, 0, 0, -1, 0, 0, 0, 2, -1, -1, 2, 0, 0, 1, 0, 0, 1, 1, 3, 1, 0, 4, 0, 3, 2, -1, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 0, 2, 1, 0, 2, 0, 3, 2, 4, 4, 4, 2, 4, 3, 0, 0, 0, 0, 0, 0, 8, 5, 2, 0, 1, -2, 0, -3, -1, -6, -6, -5, 0, 0, 2, 0, 0, 2, 2, 6, 8, 7, 7, 5, 4, 2, 0, 0, -4, -10, 8, 4, 3, 2, 0, 2, 0, 0, 0, -2, -4, -3, 1, 2, 2, -1, -3, 0, 1, 0, 3, 8, 8, 8, 7, 3, 4, 2, -4, -7, 6, 5, 3, 2, 3, 1, 1, 2, 2, 3, 1, -1, 0, 0, 2, 0, -2, -3, -3, 0, 1, 0, 4, 5, 5, 6, 3, 0, -1, -10, 7, 6, 4, 3, 5, 3, 0, 1, 4, 1, 2, 1, 2, 2, 2, -1, 0, -3, -3, -4, -3, -2, 1, 4, 5, 7, 5, 0, -1, -12, 4, 3, 5, 2, 2, 2, 3, 3, 3, 3, 0, 2, 3, 1, 2, -1, 0, -3, -5, -8, -6, -7, 0, 2, 3, 2, 1, 0, -6, -9, 7, 5, 2, 1, 1, 2, 4, 5, 2, 3, 4, 5, 4, 1, 1, 0, -1, -4, -1, -4, -7, -6, -5, -3, 0, -1, 0, -1, -5, -12, 4, 5, 3, 2, 0, 0, 3, 5, 1, 4, 1, 5, 4, 4, 1, 0, 1, -2, -1, -2, -6, -4, -3, -3, -2, 0, 0, -1, -8, -15, 4, 2, 1, 2, 1, 0, 0, 3, 1, 3, 6, 4, 6, 6, 2, 3, 3, 0, 3, 0, -3, 0, -1, -4, 0, 0, -2, -2, -6, -13, 4, 0, 3, 0, -2, -3, 0, 1, 2, 5, 4, 7, 3, 6, 2, 2, 1, 0, 1, 3, 3, -1, -1, -3, -2, -2, -4, -6, -8, -13, 3, 0, -1, 0, 0, 0, -2, 3, 4, 7, 10, 9, 7, 4, 3, 0, 3, 2, 1, 4, 2, 0, 0, 0, -2, -2, -3, -5, -10, -14, 3, 3, 0, 1, 0, 1, 0, 2, 6, 7, 10, 8, 9, 6, 4, 2, 3, 2, 2, 0, 1, 2, 2, 2, 0, -1, -2, -4, -7, -14, 4, 3, 0, 1, 0, 0, 1, 4, 5, 8, 8, 6, 4, 3, 3, 1, 4, 4, 1, 1, 0, 0, 0, 1, -1, 0, -2, -6, -7, -15, 4, 1, 0, 3, 0, 3, 3, 7, 8, 5, 7, 4, 3, 1, 1, 0, 2, 5, 1, 4, 0, 1, 1, 0, -2, -3, -3, -6, -9, -15, 4, 4, 3, 1, 2, 3, 5, 6, 7, 5, 4, 4, 2, 0, 0, 1, 2, 6, 3, 6, 2, 1, 0, -3, -1, 0, -2, -3, -6, -14, 4, 2, 3, 2, 1, 5, 4, 6, 5, 5, 7, 2, 1, 0, 1, 2, 6, 5, 7, 9, 6, 2, -1, -1, -1, -1, -3, -2, -8, -16, 3, 4, 5, 1, 1, 2, 3, 6, 7, 7, 8, 5, 2, 0, 0, 3, 8, 10, 9, 8, 3, 0, 0, -3, -2, -3, -4, -5, -9, -15, 2, 1, 3, 2, 1, 4, 2, 6, 5, 4, 6, 6, 3, 0, 0, 3, 5, 8, 9, 8, 2, 1, -1, -5, -2, -2, -2, -3, -9, -13, 1, 3, 3, 2, 2, 0, 4, 8, 5, 3, 2, 4, 4, 0, 2, 2, 3, 8, 9, 6, 3, -1, -5, -5, -4, -3, -2, -3, -8, -13, 2, 1, 2, 3, 1, 4, 6, 8, 6, 3, 3, 1, -1, 0, 0, 2, 3, 6, 4, 3, 1, 0, -2, -4, -3, -2, 0, 0, -4, -14, 2, 2, 2, 0, 0, 4, 3, 8, 5, 4, 2, 2, 0, 1, 0, 0, 4, 2, 2, 2, -1, -3, -5, -6, -4, -3, 0, -1, -4, -14, 3, 3, 1, -2, 0, 1, 5, 3, 5, 2, 1, 2, 0, 2, 0, 3, 3, 2, 0, 0, -1, -1, -2, -4, -3, -3, -1, -2, -5, -14, 3, 1, 0, 0, 1, 0, 1, 4, 3, 2, 3, 0, 0, 3, 2, 2, 1, 2, 0, -2, 0, -1, -5, -5, -3, -2, -3, -3, -8, -16, 4, 2, 1, -1, 1, 0, 3, 4, 4, 4, 4, 2, 0, 1, 2, 2, 3, 0, -2, 0, 0, -4, -4, -7, -6, -2, -3, -3, -7, -16, 1, 0, 2, -1, 1, 0, 0, 1, 2, 2, 2, 2, 3, 3, 1, 2, 0, -1, 0, -2, -3, -4, -7, -3, -5, -1, -2, -5, -8, -17, 3, 4, 0, 2, 0, -1, -1, 1, 4, 3, 0, 0, -1, 1, 1, -2, -4, -1, -2, 0, -2, -3, -1, -1, 0, -1, -2, -3, -11, -14, 3, 1, 1, 2, 0, 0, -1, 1, 3, 3, -1, 0, -2, 0, -1, -5, -3, -3, -1, 0, 2, 0, 0, 0, 0, 0, 0, -5, -9, -16, 4, 4, 2, 3, 2, 0, 2, 0, 4, 0, 0, -2, -3, -3, -1, -5, -4, -4, -2, 0, 1, 0, 2, 2, 0, 3, 2, -2, -6, -11, 4, 4, 3, 1, 0, 0, 0, 0, 3, 1, 0, -1, -4, -4, -2, -3, -2, -1, -1, 3, 2, 2, 2, 1, 1, 3, 0, 0, -7, -13, 6, 6, 2, 0, 0, 0, -1, 0, 2, 0, -2, -2, -2, -1, 0, -2, 1, 1, 0, 3, 2, 5, 0, 2, 0, 0, -2, -1, -5, -12, 10, 8, 5, 2, 1, 0, 0, -1, 0, 1, 0, 0, -1, -1, 1, 1, 3, 2, 4, 5, 4, 4, 2, 3, -2, 0, -5, -4, -8, -9, 0, 1, 2, -1, 0, 0, 0, 0, -3, 0, 0, 2, 0, 0, 0, 0, 2, 2, 4, 4, 1, 0, -1, 0, 0, 0, 0, 1, -3, -2, 0, -2, 0, 0, 0, -2, 0, -2, -3, -1, -3, 0, 2, 0, 0, 1, 2, 4, 5, 4, 1, 1, 1, 0, 0, 1, 0, -1, -1, -4, -1, 0, -1, 2, 0, 1, 0, 0, -2, -3, -2, 1, -1, -1, -1, -2, -1, 0, 0, 3, 4, 4, 2, 1, 0, 0, 1, 0, 1, -3, 1, 1, 2, -1, 1, 0, 3, 0, -1, -2, -1, -2, -1, 2, 0, 0, -1, 0, 1, 0, 2, 2, 3, 1, 2, 3, 0, -1, -2, -1, 2, 0, 0, 3, 0, 1, 0, 3, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, 0, 1, 0, 4, 4, 3, 1, 0, -4, 2, -1, 0, 0, 1, -1, 0, 1, 0, 0, 0, 0, -2, -2, 0, -2, 0, -1, -1, -2, -2, 1, 0, 1, 2, 0, 0, -1, -1, -6, 0, 0, 1, -1, 0, 1, 2, 1, 0, -2, 0, -1, -2, -2, 0, -1, -1, -1, -3, -3, -3, 0, -2, 0, -1, 0, 0, -1, -4, -6, 2, 0, 0, 1, 0, 0, 0, 3, 0, 1, 0, 0, 0, 1, 0, 0, -1, 0, -4, -2, -4, -1, -1, -2, 0, -1, 1, 0, -3, -6, -1, 1, 2, 0, 1, 2, 2, 0, 0, 0, 0, 1, 2, -2, 0, 0, 1, 1, -2, -3, -1, -2, -3, -3, -3, 0, 0, -1, -1, -5, 2, 2, 2, 1, -2, 1, 2, 2, 0, 1, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, -2, -1, -1, 0, -2, -3, -2, -1, -3, -5, 0, 0, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, -2, 1, 0, 0, 1, 0, -1, 1, 0, -3, -3, -1, -3, -1, -2, -2, -3, -6, 0, -1, 0, 0, -1, 0, 0, 3, 0, 2, 1, 0, 1, 0, 0, 2, -2, 0, 0, -2, -1, -1, -3, -2, -3, -3, -4, -1, -2, -7, 2, 1, -1, -1, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 2, 0, 0, 0, -1, -1, -3, -3, -1, 0, -1, 0, -3, 0, -3, -6, 1, -1, 0, 1, 2, 0, 1, 0, 2, 0, -1, 0, -2, 0, 2, 0, 0, -1, -1, 0, -3, -1, -3, -2, 0, -2, -1, 0, -2, -4, 0, 1, -2, 0, 1, 0, 1, 2, 0, 1, 0, 0, 0, -2, -1, 1, -1, 0, 0, 0, 0, -4, -1, -1, 0, -3, 0, -1, -2, -7, 0, 2, 0, 1, 2, 0, 0, 1, 0, 2, -1, -1, 0, 0, 1, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0, -1, -3, -1, -7, 2, 2, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, -3, -3, 0, 2, 2, 0, -1, 0, 0, -4, -4, -2, -2, 0, -3, 0, -3, -4, 0, 2, 1, 1, 1, 0, 0, 0, 2, 0, 2, 2, -1, 0, 2, 1, 4, 4, -1, 0, -3, -4, -2, 0, 0, -3, -1, -1, -4, -5, 2, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 0, 0, 1, 2, 1, 0, 0, -2, -1, -4, -3, 0, -2, -3, -1, -1, -7, 2, 1, 0, -1, 0, 1, 0, 2, 0, 0, 0, -1, 0, 1, 0, 2, 1, 0, 0, 0, -2, -4, -2, -1, -1, -1, 0, -3, -2, -6, 0, -1, 1, 0, 0, 0, 3, 0, -2, 1, -1, -1, -2, -1, 0, 0, 0, -2, 0, 0, -3, -3, -5, -1, 0, 1, -1, -1, -1, -6, 1, -1, 0, 2, 0, 2, 0, 0, 0, -1, 1, 1, 0, 0, -2, 0, 0, 0, -3, -2, 0, -1, -3, 0, 1, 1, -2, -1, -4, -4, 0, -2, 0, 0, 0, 2, 3, 0, -2, 0, -2, 0, 0, 0, 1, 0, 0, -1, -2, -3, -3, -4, -3, 0, -1, -1, 1, -2, -4, -5, 0, 0, 0, 0, 0, 0, 3, 1, 1, 2, -2, -1, 0, 0, 0, 0, 0, -2, -3, 0, -2, -3, -1, -2, 0, 2, 1, 0, -2, -3, -1, 0, 1, 2, 0, 1, 3, 3, 0, 0, 0, 0, 0, 0, 2, 1, -1, 0, -1, -3, -4, -1, -4, -2, -1, 1, -2, -2, -1, -5, -1, -1, 0, 0, -1, 1, 0, 1, 0, 2, 0, 0, 0, 1, 0, -1, -2, -1, -2, -3, -3, -1, 0, -2, 0, 1, 0, -3, -4, -2, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, -1, 0, 1, 0, -2, 0, -1, 0, 0, -3, -1, 0, -1, -1, 0, 0, -4, -1, 0, 0, 0, 1, 0, 1, 2, 1, 0, -1, 1, 0, 0, 0, 0, -3, 0, 0, -1, 0, 0, -2, -1, 1, -1, 0, -2, -2, -4, 2, 1, 0, 0, 0, 1, 3, 0, 0, 0, 0, -2, 1, -1, 0, 1, 0, -1, 0, 1, 2, 2, -1, 0, 3, 2, 1, 0, -1, -4, -1, -1, 1, -1, 0, 1, 1, 2, 1, 2, 0, -1, 0, 0, 0, 2, 0, 1, 1, 1, 1, 0, 1, 3, 0, 1, 2, 3, 0, -1, 1, -1, 0, 1, -1, -1, 1, 0, -1, 0, -1, 1, -1, -1, -1, -1, 1, 1, -1, 1, -1, 0, 0, -1, 1, 0, -1, 0, -1, -1, 1, 1, 0, -1, -2, 0, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 0, 1, 0, 0, -2, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 1, 0, -1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, -1, 0, 1, -2, 0, 0, 1, 1, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, -1, -1, 0, 0, -1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, -1, 2, 0, -1, -1, 1, -1, 0, 0, 0, -1, 0, 0, -1, 0, -2, 0, 0, -1, -2, 0, -1, 0, 0, 0, 1, 1, -1, -1, 0, 0, 0, -1, -1, 0, 0, 0, 1, 2, -1, 1, -1, 0, 1, 1, 0, -1, 0, 1, 0, 1, 0, -1, 0, 2, 0, 1, 0, -1, -1, 1, -1, 0, -2, 0, 0, 0, -2, 1, 0, 1, -1, -1, -1, 0, -1, 0, 0, 0, 1, 0, 0, -1, 0, 1, -1, 0, 0, -1, -1, 0, 0, 0, 1, 1, 0, -1, 0, -1, 0, -1, 0, 1, 0, 0, 0, -1, 0, -1, -2, 0, 1, 0, -2, 0, -1, 0, 2, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 1, 1, -1, 0, 0, -1, 0, 0, 1, 0, -1, 0, 0, -1, 0, 1, 0, -1, 0, 1, -2, 1, -1, 0, -1, 1, 1, 1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -2, 1, 1, -2, -1, -1, 0, 1, 0, -1, -1, -1, -1, 0, 1, 0, 1, 0, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 1, 0, 0, 0, -1, -1, 0, 2, 0, 0, 0, 0, 1, 0, 0, -1, 1, 0, 0, 1, -1, -1, 0, -1, 0, -1, -1, 0, -1, 1, -1, 0, 0, 2, -1, -1, 1, 0, 2, 1, 1, 1, 0, -1, 1, 0, 0, 1, -1, 1, -2, 0, -1, 1, -1, 0, 0, 0, 1, -1, -1, 1, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, -1, -1, -1, 1, -1, -1, -1, 0, 1, 0, 1, 0, -1, -2, 1, 0, 0, 1, 1, 0, 1, -1, 1, -1, 0, 2, 0, 1, 1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, -1, 0, 1, 0, -1, -1, -2, 0, -1, 1, 0, 0, -1, -2, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, -1, 0, -1, -1, 1, 0, 0, 0, 0, -2, 0, -1, 1, -1, 1, 1, -1, 1, 0, 0, 1, 0, 0, -1, 1, 0, 0, -1, -1, -1, 1, 0, 0, -1, -1, -1, 0, 0, 0, -1, 0, 1, -1, 0, -1, 0, 0, -1, -1, 1, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -1, -1, 0, -1, 0, 0, 1, -1, 2, -1, -1, -2, 1, -1, -1, -1, 1, 1, 1, -1, 1, 1, 0, 1, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 2, 1, 1, 0, -1, 0, 0, 0, -1, 1, 0, -1, 0, 0, 0, 0, -1, -1, -1, 0, 1, 0, -1, -1, 0, 0, 1, -1, 1, 1, 0, -1, -1, 1, 1, 1, -2, 0, 0, 0, 0, -1, 0, 0, 0, 2, -1, -1, -1, 0, -1, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, 1, 1, 0, 1, 1, 0, -1, 1, 0, 0, 0, 0, 0, -2, 1, 1, 1, -1, 0, 0, 0, 2, 0, 0, 2, -2, 0, 1, -2, 0, 0, 1, 0, -1, 0, 0, 0, 1, -1, -1, 1, 1, 1, -1, 1, 0, 0, -2, 1, -1, 1, -1, 1, 1, 2, 1, 1, 0, 1, 1, 1, 0, 0, -2, 0, 0, 0, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 1, -1, 0, 1, 0, 0, 0, -1, 0, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -2, 1, -1, 0, 0, -1, -1, -1, 0, 0, -1, 1, -1, 1, 0, -1, -1, 0, -1, 0, -1, -1, -2, -2, -1, -1, -1, 1, 2, -1, -1, 0, -1, 0, -2, 0, 0, -1, -1, -1, 1, 0, -1, 0, 0, -1, -1, 0, 0, 0, -1, -1, 1, 0, 1, 0, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -2, 1, -1, 1, 1, 2, -1, -1, -1, -1, 1, 1, 0, 1, -1, 0, 1, 1, 0, -2, 0, 2, -1, 0, 0, 1, 1, 0, -1, 1, 0, -1, 0, 2, 0, 0, 0, -1, 1, 0, 1, -2, 0, 1, 0, 1, 0, -1, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, -1,
    -- filter=0 channel=9
    4, 1, 2, 2, 4, 3, 1, 0, 0, 2, 0, 0, 0, 0, 1, 1, -1, 2, 3, 3, 1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 4, 1, 1, 3, 2, 4, 0, -1, 0, 1, 3, 0, 1, 1, 0, 0, 0, 1, 2, 1, 0, 1, 0, 0, 1, -1, -1, 0, 0, -1, 2, 2, 0, 1, 4, 2, 1, 0, 0, -1, 2, 0, 1, -1, 0, 2, 0, 3, 2, 0, 0, 1, 0, 0, 0, 1, 3, 2, -1, -1, 0, 2, 0, 1, 3, 0, 2, -1, -1, 0, 1, -1, 0, 1, 1, 0, 0, 0, 0, 1, 3, 1, 0, 1, 0, 1, 4, 0, 0, 0, 3, 1, 0, 1, 4, 0, 2, 0, 0, 0, 2, 0, 0, 1, 2, 2, 2, 2, 1, 1, 3, 3, 3, 0, 3, 3, 3, 0, 2, -2, 0, 1, 3, 3, 2, 1, 1, 1, 0, 0, 2, 0, 0, 2, 0, 3, 1, 1, 3, 4, 2, 1, 2, 2, 4, 4, 4, 2, 3, -1, 3, 2, 2, 2, 2, 0, -1, 1, 0, 2, 4, 2, 0, 1, 2, 2, 3, 2, 3, 0, 1, 1, 1, 1, 1, 1, 2, 3, 0, -1, 3, 3, 2, 0, 0, 1, 1, -1, 2, 1, 3, 2, 3, 0, 3, 0, 0, -1, 2, 1, 3, 2, 2, 2, 1, 2, 4, 3, 1, -2, 5, 2, 3, 1, 0, 0, -1, 0, 0, 2, 0, 3, 1, 2, 2, 3, 0, -1, 2, 1, 2, 0, 0, 2, 3, 2, 1, 3, 3, 2, 2, 4, 3, 1, 0, 2, 0, 0, 1, 1, 1, 3, 1, 0, 2, -1, 0, -1, 3, 1, 1, 1, 0, 2, 1, 1, 2, 4, 0, 0, 4, 2, 0, 1, 0, 0, -1, 0, 0, 0, 2, 0, 1, 0, 1, 0, 2, 0, 1, 1, 2, 3, 1, 0, 1, 1, 4, 2, 2, 0, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 2, 1, 2, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 2, 2, 2, 3, 3, 0, -2, 2, 2, 1, 0, 2, 0, 0, 1, 0, 0, 0, 0, 2, 1, -1, 1, 0, -1, 1, 1, 3, 3, 2, 0, 1, 4, 2, 2, 3, 0, 2, 1, 2, 0, 2, 0, 0, -2, 0, 1, 3, 2, 2, 1, 1, 0, 0, 0, 0, 1, 4, 3, 1, 0, 0, 4, 4, 4, 2, 0, 1, 3, 0, 0, 0, 2, -2, -2, 2, 0, 0, 0, 1, -1, 1, 0, -2, 0, 2, 4, 1, 1, 1, 2, 2, 2, 4, 4, 1, 0, 0, 0, 1, -1, 0, 1, 0, 0, 0, 1, 2, 0, 2, 1, -1, -1, 0, -2, 1, 2, 5, 3, 1, 2, 0, 2, 1, 5, 4, -2, 0, 2, -1, 2, 1, 0, 0, -1, 0, 2, 3, 2, 2, 0, -1, -1, -1, 1, 4, 1, 3, 3, -1, 1, 3, 2, 3, 4, 1, -2, 4, 3, 0, 0, 2, 0, 2, 2, 2, 2, 2, 2, 0, -1, -1, 1, 1, 1, 4, 2, 4, 1, 2, 4, 4, 5, 4, 3, 2, -2, 1, 0, 0, -1, 0, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 1, 0, 1, 2, 0, 1, 0, 0, 3, 4, 5, 4, 4, 3, -3, 3, 2, 2, 1, 0, 0, 0, 2, 0, 0, 0, 2, 2, 1, 1, 0, 0, 0, 3, 0, 0, 3, 2, 0, 5, 4, 2, 2, 0, 0, 4, 2, 1, 1, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 1, 3, 1, 3, 2, 2, 4, 5, 3, 2, 2, 1, 0, 4, 2, 2, 0, 2, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 1, 0, 3, 4, 3, 0, 0, 3, 2, 4, 2, 2, 3, 2, -3, 1, 1, 1, 1, 2, 0, -1, -1, 0, 1, 2, 1, 0, 0, -2, 1, 2, 0, 4, 2, 0, 3, 0, 2, 4, 5, 3, 2, 2, 0, 2, 2, 0, 4, 0, -1, -1, 1, 0, 2, 0, 1, 2, 1, 0, 2, -1, 0, 4, 0, 2, 2, 2, 5, 3, 3, 3, 1, 0, -3, 4, 2, 0, 2, 0, -2, 0, 1, 0, 0, 0, 0, 2, 0, 0, -1, 2, 3, 1, 1, 0, 2, 2, 3, 3, 2, 4, 3, 0, 0, 4, 0, 2, 0, 1, 1, 0, 0, 1, 0, 1, 0, 0, -1, 0, 0, 0, 3, 2, 3, 1, 2, 2, 1, 2, 1, 3, 0, 0, -1, 1, 3, 2, 2, 2, 0, 0, 2, 1, -1, -1, 1, 0, 0, -1, -2, 1, 0, 1, 0, 2, 0, 0, 1, 3, 3, 1, 0, 0, -3, 2, 1, 4, 1, 0, 0, 2, 3, 0, 0, 0, 0, -1, 1, -1, 0, -1, 1, 0, 0, 0, 0, -1, 2, 3, 0, 0, 2, -2, -3, 2, 2, 0, 2, 1, 0, 0, 1, 0, 1, 0, -1, 1, 1, 0, -1, 1, -1, 0, 1, -1, -2, 0, -1, -1, 0, -1, -1, -2, -3, 2, 1, 3, 0, 2, 2, 1, 3, 2, 1, 0, 2, 2, 0, 3, 2, 2, 0, 2, 0, 0, 0, 1, 0, 1, -1, -1, 0, 0, 0, 12, 12, 9, 8, 6, 6, 3, 1, 0, 0, 2, -2, -4, -7, -7, -9, -11, -11, -10, -11, -8, -9, -7, -4, -4, -1, 0, 2, 3, 3, 15, 9, 9, 7, 4, 4, 4, 2, 1, 0, 0, 0, -3, -3, -6, -6, -5, -7, -5, -6, -9, -7, -5, -3, 0, -3, 1, 0, 2, 1, 13, 11, 7, 6, 3, 4, 4, 0, 4, 2, 1, 0, -2, -1, -1, -2, -4, -1, -6, -7, -3, -5, -5, -3, 0, -2, 0, 1, -2, 0, 13, 10, 8, 7, 3, 4, 2, 2, 4, 4, 1, 0, 0, 1, 0, 0, -2, -2, -4, -3, -3, -2, -2, -1, -2, 0, 0, -2, -2, 0, 12, 8, 7, 7, 3, 1, 4, 1, 3, 1, 1, 0, 4, 2, 0, 0, 0, 1, 0, -2, -2, -2, -3, -1, -2, 0, -3, -3, -4, -1, 13, 7, 8, 7, 4, 3, 3, 1, 4, 2, 3, 1, 2, 3, 1, 0, -1, 0, 0, -4, -3, -2, -3, -1, -2, -3, -4, -4, -3, -4, 12, 8, 7, 5, 3, 4, 4, 1, 3, 1, 1, 2, 0, 2, 0, 0, 1, 0, -2, -3, -5, -1, -3, -4, -2, -5, -2, -3, -3, -1, 12, 5, 1, 2, 3, 2, 3, 3, 2, 0, 1, 0, -1, 0, 0, -3, -3, 0, -3, -4, -2, -6, -3, -2, -2, -4, -5, -4, -2, -3, 9, 6, 2, 0, 0, 0, 2, 1, 3, 2, 2, -1, 2, 0, -1, 0, 0, -1, -1, -3, -4, -4, -5, -3, -2, -3, -6, -4, -6, -1, 9, 4, 0, -1, 0, 0, 2, 0, 2, 3, 0, 0, 1, 0, 0, 1, 0, 0, -1, -1, -1, -4, -2, -2, -3, -3, -5, -4, -4, -1, 7, 1, -2, -4, -4, -1, -3, -1, -1, 0, 1, 0, 0, -1, 1, 0, -1, -1, 0, -1, -3, -1, -4, 0, 0, -4, -1, -2, -3, 0, 7, 0, -3, -4, -1, -4, 0, -3, 0, -1, 1, 0, -2, 0, -2, 0, 0, 2, 0, 0, -1, -4, -1, -3, -2, 0, -4, -5, -3, -3, 8, 0, 0, -1, -3, -5, -3, -4, -3, 0, 0, 0, -1, -2, 0, 2, 4, 3, 0, -1, -1, -2, -2, -1, -1, -1, -1, -2, -4, 0, 9, 1, 0, 0, -4, -4, -2, -1, 1, 2, 2, 0, 0, 0, 1, 0, 3, 2, 2, 2, 2, -2, -4, -4, 0, 0, -3, -3, -3, -1, 12, 3, 0, -3, -2, -3, -1, 0, -1, 3, 0, 0, 0, -1, 0, 2, 1, 3, 5, 2, 3, 0, -3, 0, -2, 0, -2, -1, -2, -1, 8, 4, -1, 0, -1, -3, -1, -3, -1, 2, 1, 0, 0, 0, 2, 2, 5, 5, 3, 3, 2, -2, -2, -1, 0, 0, 0, 0, -4, 0, 13, 3, 0, -1, -3, -3, -3, -3, 1, 0, 0, 1, -1, 1, 1, 5, 4, 6, 5, 1, 0, -4, -3, 0, 0, 0, 0, -2, -1, -3, 10, 4, 0, -2, -2, 0, -1, -2, 1, 0, 0, 0, 0, 0, 0, 1, 6, 4, 2, 0, 0, -2, -3, 0, -2, -1, 0, -2, 0, -1, 10, 4, 0, -3, -2, -2, -3, 0, -2, -2, 0, 0, 1, -1, 0, 1, 0, 4, 1, -2, -3, -1, -3, -1, -1, 0, -1, -4, -4, 0, 10, 7, 0, 0, 0, -2, -3, 1, 0, 1, 0, -2, 0, 0, 4, 2, 2, 4, 0, -2, -2, -2, -4, -3, -1, -3, -5, -2, -2, -1, 12, 5, 2, -1, -1, 0, 2, 1, 1, -1, -1, 0, -2, 0, 2, 0, 3, 1, 2, -1, -2, -4, -3, 0, -2, -3, -3, -3, -6, -2, 12, 9, 0, 2, 0, 0, 1, 3, 1, 1, 0, -2, 0, -1, 0, 1, 2, -1, 1, 0, -3, -2, -2, 0, -1, -1, -3, -5, -5, -4, 14, 9, 6, 4, 0, 3, 2, 0, 2, 3, 2, -1, -2, 0, -1, 0, 1, 0, 0, -1, -3, -2, -4, -2, -3, -1, -3, -3, -4, -2, 14, 10, 3, 6, 4, 2, 0, 1, 1, 2, 0, -2, -3, 0, -1, 0, 0, -2, -4, -2, -3, -4, -5, 0, -3, -4, -2, -2, -6, -5, 11, 8, 6, 5, 4, 2, 1, 3, 2, 0, 0, 0, -1, -2, -2, 0, -1, -2, 0, -5, -7, -3, -3, -5, -3, -5, -4, -7, -5, -4, 12, 7, 9, 6, 3, 3, 4, 1, 2, 0, -1, 0, -2, -5, -2, -4, -1, -1, -1, -3, -3, -4, -6, -7, -4, -2, -6, -5, -5, -3, 10, 10, 8, 7, 6, 2, 4, 4, 3, 2, -2, -3, -1, -2, -4, -3, -3, -1, -6, -5, -6, -7, -5, -3, -4, -3, -4, -3, -4, -2, 14, 10, 8, 5, 3, 3, 3, 3, 0, 0, -1, 0, -4, -3, -1, -5, -3, -2, -3, -7, -9, -6, -4, -1, 0, -4, -4, -3, -1, -3, 12, 8, 9, 4, 5, 4, 3, 1, 0, -2, -3, -3, -2, -4, -6, -4, -4, -7, -6, -8, -8, -7, -5, -3, -3, -4, -2, 0, -3, 0, 11, 9, 8, 4, 5, 3, 1, 2, 0, -2, -2, -2, -1, -3, -6, -5, -5, -9, -6, -7, -9, -6, -6, -6, -6, -2, -2, 0, 0, 2, 5, 5, 4, 3, 3, 4, 1, 2, 0, 0, 0, -1, -2, -2, -4, -3, -5, -7, -5, -5, -6, -6, -5, -6, -5, -3, -1, -1, 0, 0, 8, 7, 6, 5, 1, 1, 1, 1, 3, 2, 1, 0, 0, 0, 0, -1, -3, -2, -4, -3, -3, -3, -2, -1, -3, -2, -2, -1, -2, -2, 6, 5, 5, 3, 3, 4, 2, 1, 3, 0, 2, 0, 0, 0, -1, 1, -2, 0, 0, -2, -3, 0, 0, -3, -1, -2, 0, 0, -2, 0, 5, 6, 2, 2, 2, 3, 0, 2, 4, 1, 3, 2, 2, 0, 1, 1, -1, 1, -1, -1, -1, 0, 0, 0, -2, 0, -1, -2, 0, -1, 8, 6, 4, 3, 4, 2, 3, 0, 2, 1, 2, 3, 1, 1, 1, 0, 1, 1, 0, -1, -1, 1, 0, -2, -1, -1, -2, 0, -2, -3, 6, 3, 5, 4, 1, 4, 2, 0, 0, 3, 3, 3, 1, 2, 3, 4, 0, 0, 1, 1, 1, -1, 1, -2, -1, 0, -2, -3, -1, -3, 7, 4, 5, 3, 4, 3, 3, 2, 2, 1, 3, 3, 4, 4, 4, 4, 4, 2, 1, 1, 1, -1, -2, -3, -2, -3, -1, -3, -2, -1, 6, 4, 4, 3, 1, 4, 4, 0, 2, 1, 1, 2, 3, 4, 1, 2, 1, 0, 2, 0, 0, -1, 0, -3, -1, -1, -1, -3, -2, -3, 7, 4, 3, 0, 0, 0, 1, 2, 3, 1, 0, 2, 3, 3, 1, 2, 2, 2, 1, 0, -1, -1, -1, -1, 0, -2, -3, -3, -2, -3, 5, 2, 0, -1, 2, 2, 0, 0, 2, 0, 1, 2, 0, 4, 2, 2, 4, 1, 2, 2, 1, -1, 0, -2, 0, 0, -2, -2, 0, -1, 3, 4, 0, -1, 0, 0, -1, 1, 0, 3, 0, 3, 1, 2, 1, 1, 1, 2, 4, 1, 3, -1, 0, 0, 0, 0, -3, -2, 0, 0, 4, 0, -2, -1, -2, -1, 0, -1, -1, 1, 2, 3, 2, 3, 3, 4, 2, 2, 4, 1, 0, 0, -1, 1, 0, 0, -3, -3, -2, -1, 6, 4, -1, 1, -1, -1, 1, 0, 0, 1, 1, 0, 0, 2, 1, 3, 3, 4, 1, 0, 1, 0, 0, 0, -1, 1, 0, 0, 0, 0, 3, 1, 0, 1, -1, -1, 0, 1, -1, 0, 0, 2, 1, 1, 3, 4, 1, 3, 4, 0, 3, 0, 0, 0, 0, -2, 0, 0, -1, 0, 4, 4, 2, 0, -1, 1, -1, 0, -1, 1, 3, 1, 1, 2, 3, 4, 4, 5, 5, 2, 5, 1, 1, 0, 0, -1, 0, -1, 0, 0, 4, 1, 2, -1, 2, 0, 1, 1, 1, 2, 1, 3, 2, 2, 2, 5, 3, 4, 7, 5, 3, 2, 1, 0, 0, 0, 1, 0, -2, 0, 6, 1, 1, 0, 1, 0, 0, -1, 3, 1, 3, 4, 1, 2, 5, 5, 4, 5, 6, 5, 4, 2, -1, 0, -1, 2, 0, 0, 1, -3, 7, 3, 1, 2, 2, -1, 2, 1, 0, 3, 1, 2, 1, 3, 4, 6, 4, 5, 2, 5, 3, 0, 0, 0, 0, 0, 0, -1, -1, -2, 5, 3, 2, 0, 1, 0, -1, 0, 1, 0, 0, 0, 1, 1, 3, 3, 4, 5, 1, 2, 2, 0, 0, 0, -1, -1, 0, 0, -1, -2, 8, 3, 0, 2, 0, 1, 2, 1, 0, 1, 0, 0, 3, 5, 6, 5, 4, 2, 4, 3, 0, 2, -1, 0, 0, 0, 0, -1, -1, -3, 7, 2, 1, 0, 1, 1, 0, 3, 0, 1, 1, 0, 3, 3, 4, 1, 3, 4, 3, 3, 0, 1, 0, -1, 0, 0, -2, -4, -2, -2, 8, 3, 0, 1, 3, 1, 1, 2, 2, 2, 0, 0, 2, 0, 2, 3, 3, 3, 1, 0, 0, 0, -1, 0, 0, -1, 0, -3, -2, -1, 5, 5, 3, 4, 0, 2, 3, 2, 1, 3, 0, 2, 1, 1, 2, 4, 4, 3, 2, 2, 0, 1, 0, 0, 1, -1, 0, 0, -1, -3, 6, 5, 1, 0, 4, 1, 1, 1, 1, 1, 0, 1, -1, 0, 1, 1, 3, 0, 0, 0, -1, 1, -1, -2, -2, -3, -2, -3, 0, -2, 4, 3, 3, 3, 2, 3, 0, 1, 3, 2, 2, -1, 1, 3, 0, 3, 2, 0, 0, -2, -2, 0, -2, 0, 0, -3, -1, -1, -1, -4, 4, 5, 2, 4, 2, 0, 4, 1, 1, 2, 0, 0, 1, 2, -1, 0, 0, 0, 1, -2, -1, -1, -2, -3, 0, 0, -1, -5, -1, -4, 5, 3, 2, 1, 1, 2, 3, 2, 2, 2, 0, 0, -1, 1, -2, 0, 0, 1, -1, 0, 0, 0, -3, -2, -2, -3, -2, -4, -2, -3, 5, 4, 3, 1, 1, 1, 1, 2, 0, 0, 0, 1, 0, 0, 1, -2, 0, -1, 0, -2, -5, -5, -3, -5, -2, -1, -3, -1, -3, -2, 8, 5, 5, 0, 1, 3, 0, 1, 0, 0, 2, 1, 0, 1, 0, 0, 0, -2, -3, -2, -2, -3, -1, -5, -5, -1, -1, -3, -2, 0, 4, 7, 2, 1, 3, 4, 0, 3, 0, 0, 0, 1, -1, 0, 0, 0, -2, -1, -2, -4, -6, -6, -5, -2, -5, -5, -2, -5, -5, -2, 1, 0, -2, 0, -1, -1, 0, 0, -1, -1, 0, 1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 0, 1, 1, 0, 0, -1, -1, 0, 0, 1, -1, 0, 1, 1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, -1, 0, -1, 1, 1, -1, -1, 0, 1, -1, 1, 0, 1, 0, -1, 2, 0, 0, -1, 1, -1, -1, 0, 0, -1, 1, 0, 0, 0, 1, 1, 0, -1, 0, 0, 1, -1, -1, 0, -1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -2, 2, -1, 0, 0, 1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, 1, 1, 1, 0, 0, -1, 0, -1, 1, 2, -1, 0, 0, 1, 0, 0, 1, 1, 0, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 1, -1, 0, 1, -1, 0, 1, 0, 0, 2, 1, -1, 0, 0, 1, 1, -1, 1, 0, 1, 0, 0, 0, 0, -1, -1, 0, 1, -1, 0, 0, 0, 1, 0, 1, 1, 1, 0, -2, 0, 0, -1, -1, 0, -1, 1, -1, 0, 1, 2, -1, 1, 0, 0, 0, 1, 0, -1, -1, 1, 2, -1, 0, 0, 1, -1, -1, -1, 1, 0, 0, 1, 1, 0, -1, -1, 0, -2, -1, 1, -1, 0, 0, 1, 0, 0, 0, 0, -1, -1, 0, 0, 0, 0, -2, -1, 0, -1, 1, -1, 0, -1, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, 0, 1, -1, -1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, 1, 1, 0, -1, 1, -1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, -1, -2, -1, 0, 0, -1, 0, 2, 0, -1, -1, -1, 0, 1, -1, 0, 0, -1, 0, 0, 1, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, -1, 0, -2, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, -1, 1, 0, 0, 1, 0, 0, -1, 0, -1, 1, -1, 0, -1, 1, 1, 0, -1, 0, -1, 0, 2, 1, 1, -1, 0, 1, 1, -1, -1, -1, -1, 0, -2, 1, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, -2, 0, 0, -2, 0, 1, 1, 2, 0, 1, 0, 1, -1, -1, 0, 0, 0, 0, 1, -1, 0, -1, 0, 1, 1, 1, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, -1, -1, 2, -1, 1, -1, 0, 1, -2, -1, 0, 0, 0, -2, 0, 0, 0, 1, 0, 1, -1, 1, -1, 0, 1, -1, 0, 1, -1, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -1, 0, 0, 0, 1, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, -1, 1, -1, 1, 0, 1, -2, 0, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, -1, -1, -1, 0, 0, 1, 0, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 1, -1, 0, 0, 0, -1, 1, 0, 0, -1, 0, 0, 1, -1, 0, 0, 0, 0, 1, 0, 1, 0, 0, -2, -1, 0, 0, 0, 0, 1, 0, 0, 0, -1, 0, 1, 1, 0, 1, 1, 0, 1, -1, 1, -1, 0, 0, 0, 0, -1, 1, 0, 1, 1, -1, 0, 1, 1, 0, 1, 0, 0, 1, 1, -1, 1, 1, 1, -1, 1, 0, 0, -1, 0, 0, 0, -1, 1, -1, 0, -1, 0, -1, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, -1, 0, -1, -1, 1, -1, -2, 0, 0, 0, 0, -1, 0, 1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 0, -1, 0, 0, -1, -1, -2, 0, -1, 0, -1, 0, 0, 1, -1, -1, 0, 2, 0, 1, 0, 0, 0, -1, 1, 1, -1, 1, 1, 0, 0, -1, 1, 0, -2, 1, 0, 0, 0, 1, 0, 1, 1, -1, 0, 1, 0, 0, 1, -1, 0, 1, -1, 0, -1, 0, 1, 1, 0, -1, 1, 0, 2, -1, -1, 2, 0, -1, 1, 1, 0, -1, 0, -1, 0, -1, 1, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, 0, 1, 0, 1, -1, 0, 1, 1, 0, 1, 0, -1, 1, 0, 0, 0, 0, 1, -1, -1, 0, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -2, 0, -1, 0, 0, -1, -1, 0, 0, 0, 0, 1, -1, 0, 0, 0, 0, 1, 1, -1, -1, -1, 1, -1, 0, 0, 0, 1, 0, 0, 0, -2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, 2, -1, -1, 0, 1, 0, -1, 2, 0, 1, 1, 1, 0, 1, 1, 0, 0, 0, 0, 1, -1, 0, 0, 1, 1, -1, 1, 0, 1, 1, 0, 0, 0, 1, 1, -1, 0, -1, -1, 1, -2, -1, -1, 2, -1, 1, -1, -2, 0, 1, 4, 2, 2, 0, 1, 2, 0, 1, -1, 2, 0, -1, 0, -1, -2, -4, -3, -1, -1, -4, -1, 0, -1, 1, 4, 6, 6, 9, 8, 9, 0, 0, 0, 0, 0, 0, 0, 1, 1, 3, 0, 0, -2, -2, -1, -1, 2, 0, 0, -2, -1, -1, 0, 2, 3, 3, 5, 3, 4, 4, 0, 1, 0, 0, 1, 0, 0, 1, 1, 1, 2, 0, 0, 0, -1, 1, 2, 0, 0, -3, -1, 0, -2, 0, 1, 2, 3, 1, 2, 4, 1, 0, 0, -1, -1, -3, 0, 2, 0, 0, 2, 1, 2, 2, 1, 0, 0, 2, 0, 0, -3, -1, -2, -2, 0, 0, 0, 2, 1, 4, 0, 1, 0, 0, 0, 0, 0, 2, 1, 1, 1, 2, 2, 2, 0, 0, 2, 3, 2, -2, -3, -4, -4, -2, -3, 0, -1, 1, 2, 3, 0, 1, 0, 0, 2, -1, 1, 2, 1, 1, 2, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, -1, -3, -5, -5, -2, 0, 0, -1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, -2, -1, 0, 2, -1, -2, -2, -4, -5, -3, -3, -1, -1, 0, 0, 2, 0, 1, 0, 1, 0, 0, 0, 0, 1, 1, 1, -1, -2, 1, 0, -1, 0, 2, 2, 0, -1, -5, -3, -3, -5, -3, -2, -4, -1, 0, 0, -2, 1, -1, 0, -1, 1, 0, 1, 3, 0, -1, 0, 2, 0, 0, 1, 1, 0, 0, -2, 0, -2, -3, -5, -5, -3, 0, -1, 0, 0, -3, -2, -3, -2, 0, 1, 3, 0, 0, 0, 0, 0, 1, -1, 2, 2, 3, 2, 0, 0, -3, 0, -3, -1, -3, -1, -2, 0, 0, -1, -3, -4, -1, -1, 0, 1, 2, 1, 0, 1, -1, 0, 1, 0, 0, 2, 3, 2, 0, -3, -3, -1, -1, -4, -5, 0, 0, 0, 1, 0, -3, -1, 0, 0, 0, -2, 0, -1, 0, 0, 0, 0, 1, 1, 1, 5, 3, 1, -1, -4, -4, -2, 0, 0, -4, -3, -1, 0, 3, 1, -2, 0, 0, -3, 0, -2, 1, 2, 1, -1, -2, -2, 0, 2, 1, 5, 6, 2, -1, -1, -3, -3, -1, -2, 0, -1, -1, 0, 1, 1, 1, -1, 0, 1, 1, -1, -1, 1, 1, 1, 0, -2, 1, 2, 1, 5, 4, 3, 3, 0, -3, -3, -3, -1, -2, -1, -2, -1, 0, 0, -2, 0, 0, 1, 0, -1, 2, 2, 2, 0, 2, 0, 1, 3, 1, 5, 6, 3, 5, 2, -1, 0, 0, -1, -2, -3, -2, -3, 1, 2, 0, 0, 0, 1, -1, 0, 0, 2, 3, 1, 0, 0, 2, 1, 3, 5, 9, 5, 3, 0, -3, -2, 0, -3, -2, -2, 0, 0, 0, 3, 1, 0, 0, -1, 1, 0, 1, 0, 2, 2, 2, 2, 1, 1, 5, 6, 4, 6, 4, 0, 0, 0, -2, -3, -2, -2, 0, -3, -1, 1, -1, 0, 0, -1, 0, -1, -1, 0, 1, 1, 0, 0, 1, 0, 5, 3, 6, 3, 2, 0, -3, -1, 0, 0, -2, 1, 0, -2, 2, 0, 0, -3, 0, -2, -2, -2, 0, 1, 0, 0, 1, -1, 1, 2, 3, 5, 4, 1, 0, -3, -3, -1, 0, -1, -1, -1, -3, 0, 0, 1, 0, -2, -3, 0, -1, 1, 1, 0, -1, 1, 0, -1, 2, 0, 1, 3, 5, 1, 0, 0, -4, -2, 0, -1, -4, -5, -4, -3, 0, 1, -3, -3, -1, -2, -2, 0, 2, 1, 0, 0, -2, -1, 3, 0, 1, 2, 2, 1, 1, -1, -3, -4, -3, -3, -2, -1, -3, 0, 2, 0, -2, 0, -3, -3, -2, 0, -1, 0, 1, 1, 0, 0, 2, 0, 0, 2, 2, 3, 0, 1, -2, -3, -4, -3, -3, 0, -4, -2, 1, 0, 0, -3, -3, -2, -2, 0, 1, 0, 3, -1, 0, 0, 1, 0, 2, 4, 2, 1, 1, 0, -2, -2, 0, -2, 0, -1, -2, -1, 1, 2, -1, 0, -1, -3, 0, 0, 2, 1, 1, 0, -1, 1, -1, 0, 3, 5, 1, -1, 0, -2, -1, 0, -1, -1, -1, 0, -1, 0, 3, 0, -1, 0, 0, -2, -1, 2, 1, 0, 1, 1, 0, 0, -2, 0, 4, 2, 4, 0, 0, -1, -4, -3, -4, -3, -2, -1, -3, -2, 1, 1, 0, -2, 0, -2, 0, 1, 1, 3, 0, 0, 2, 2, 1, 3, 1, 5, 1, -1, -2, 0, 0, -3, -3, -3, -3, -2, 0, 0, 1, 3, 2, -1, 0, 0, 0, 0, 2, 0, 2, 1, 3, 2, 1, 3, 3, 5, 3, 0, -2, -4, -4, -3, -1, 0, -1, -1, -2, 0, 1, 3, -1, -1, 0, 0, 1, 0, 0, 2, 0, 3, 4, 1, 1, 2, 0, 2, 3, 0, -1, -3, -4, 0, 0, 1, 0, 0, 0, 0, 2, 1, 2, 0, 0, 0, -2, -1, 1, 0, -1, 1, 0, 1, 3, 1, 1, 1, 0, 0, 2, -1, 0, 1, 1, 2, 2, 3, 0, 4, 5, 3, 0, -1, 1, 0, -2, -1, 0, -2, -1, 0, 0, 1, 0, 0, 1, 2, 1, 2, 3, 4, 4, 2, 4, 2, 2, 4, 6, 3, 5, 1, 0, 2, 2, 1, 2, 1, 2, -1, 2, 1, 0, 0, 2, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, 1, 0, 2, 0, 2, 2, 1, 0, 0, 1, 1, 1, 0, 0, 2, -1, 0, 2, 0, 2, 2, 0, 2, 0, 0, 0, -1, 1, 0, 0, -1, -1, 0, 1, 2, 1, 1, 0, 0, 2, 1, 2, 0, 2, 0, 2, 1, 0, 0, 0, 2, 0, 2, 0, 0, 1, 2, 2, 0, 0, 0, 1, 0, 2, 0, 2, 0, 0, 1, 2, 0, 0, -1, 0, 2, 0, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 0, 0, 0, 1, 0, 1, 0, 2, 1, -1, 1, 1, 1, 1, -1, 0, 0, 0, 0, -1, 0, 1, 0, 1, 0, 1, 3, 3, 1, 0, 0, 2, 0, 0, 1, 0, 1, 0, 0, -1, 2, 1, 1, 1, 0, -1, 0, 0, 0, 2, 0, 2, 1, 0, 0, 1, 0, 1, 2, 0, 3, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -1, 0, 1, 1, 0, 0, -1, 1, 0, 0, -1, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, -1, 2, 2, 1, 0, 2, 0, 2, 0, 0, 0, 1, 2, 0, 2, 1, 0, 0, -1, 0, 2, 0, 2, 0, 0, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 2, 2, 1, 0, -1, 2, 2, 0, 0, 1, 0, 1, 0, 2, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 1, 2, 1, 0, 0, 0, 0, 2, -1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 3, 3, 0, 2, 2, 0, 1, 0, 2, 1, 1, 0, 0, -1, 1, 1, 0, 1, 0, 0, 0, -1, 1, 1, 0, 0, -1, 2, 1, 3, 0, 0, 2, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 1, 1, 0, 2, 0, 0, 0, 0, 0, 2, 0, 1, 2, 0, 2, 2, 2, 1, 1, 0, 0, 0, -1, 1, 2, 0, 0, -1, 0, 1, 0, -1, 0, 1, 0, 0, 0, 3, 2, 0, 1, 3, 0, 1, 0, 2, 0, 0, 0, 1, 2, 0, 0, 2, 1, 0, 0, 0, 1, 0, 1, 0, 0, 2, 1, -1, 0, 1, 0, 0, 3, 2, 2, 2, 0, 2, 2, 0, -1, 0, 2, 1, 0, 2, 0, 1, 1, 0, 1, 0, 2, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 2, 2, 0, -1, 0, 0, 2, 0, 0, 0, 0, -1, 2, 1, 3, 2, 0, 0, 1, 2, 0, 0, 3, 1, 3, 0, 0, 2, 0, 1, 1, 2, 0, 2, 2, 0, 1, 0, 1, -1, 2, 0, 0, 2, 0, 0, 1, 0, 0, 1, 0, 1, 1, 2, 0, 0, 0, 1, 0, 3, 0, 0, 0, 0, 1, 1, 0, -1, 1, 0, 2, 0, 0, 1, 0, 0, 2, 0, 1, -1, 0, 1, 3, 1, 1, 2, 0, 2, 1, 0, 1, 2, 2, 1, 0, 0, 0, 2, 0, 0, 1, 2, 0, 1, 0, 0, 1, 1, 0, 1, 2, 1, 0, 2, 2, 0, 2, 2, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 1, 0, 0, -1, 1, 0, -1, -1, 0, 1, 0, 0, -1, 0, 3, 1, -1, 1, 0, 1, 2, 1, 1, 2, -1, 1, 1, 0, 0, -1, 2, 1, 0, 1, 1, -1, 0, 0, 2, -1, 0, 0, -1, 1, 0, -1, 2, 1, 1, 1, 3, 1, 1, 1, -1, 0, 0, 1, -1, 0, 0, 1, 2, 2, 0, 2, 2, 0, -1, 2, 0, 0, -1, 1, 0, 0, 2, 2, 0, 0, 3, 0, 1, 2, 2, -1, 0, 0, 2, -1, 0, 0, -1, 1, 1, 1, 2, 0, -1, 0, -1, 1, 2, -1, 0, 1, 1, 2, 0, 2, 3, 0, 1, 0, 0, 0, -1, 1, 0, 0, 2, 2, 1, 2, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 0, 3, 3, 2, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, -1, 1, 0, -1, -1, 1, 2, 1, 0, 0, 0, 3, 0, 0, 2, 2, 0, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 0, -1, 1, 1, -1, 2, -2, 0, 1, 0, 2, 2, 3, 3, 1, 1, 2, 0, 1, 0, -1, 0, 0, 2, 0, 0, 0, 1, 1, -1, 0, -1, -1, -1, 0, 0, 0, 2, 1, 0, 0, 0, 2, 0, 1, 2, 2, 0, 0, 0, 1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 1, 1, 3, 1, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 2, -1, -1, 1, 2, 2, 1, -1, 0, 2, 2, 0, 1, 2, 0, 2, 0, 1, 2, 2, 0, 0, 3, 0, 0, 0, 1, 2, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 2, 0, -1, -1, 1, 0, 2, 0, 2, 1, 0, 2, 0, 0, 1, 1, -1, -1, 0, -1, -1, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 1, 2, 0, -1, 1, 0, -1, 0, -1, 0, -1, -1, 1, 0, -2, -1, 0, -1, 0, 1, 0, 0, 0, 0, -1, 1, 1, 2, 0, 1, 2, 1, 1, 0, 1, 1, 0, 0, 1, 0, -1, -1, 1, -1, -1, -2, -2, 1, 1, 0, 0, 1, 0, 1, 2, 1, 0, -1, 0, -1, 0, 2, -1, 0, 1, 2, 0, -1, -1, 1, 1, 1, 1, -1, 0, 0, -1, 1, 2, 2, 0, -1, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, 1, 1, 1, 1, 0, 0, -1, -1, 0, -1, 0, 1, 2, 0, 1, 1, 0, 0, -1, 0, 1, 0, 0, 0, 1, 1, 1, -1, 1, 1, -1, 0, -1, 0, 0, -1, 0, 0, 0, -2, 1, 1, 1, -1, -1, -1, 0, 0, -1, 0, -1, 0, -1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 0, 0, 2, 1, -1, -1, 0, 0, -1, 1, 1, -1, -1, 0, 0, 2, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, -1, 1, 0, 0, -1, -1, 0, 2, 2, 1, 0, -1, 0, 1, 1, 0, 1, 0, 1, 0, 2, 0, 0, 1, 0, -1, -2, 0, -2, 0, 1, -2, 1, 0, 0, 0, 0, 1, -1, 2, -1, 0, -1, 0, 0, 1, 2, 0, 2, 1, 3, 0, 0, 0, 0, -2, 0, -1, -1, 0, 0, 0, 0, 0, -1, 0, 0, 2, 1, 0, 0, 1, 0, 1, 1, 0, 1, 3, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, -1, -1, -1, 0, 0, 0, 1, -1, -1, 0, 0, 0, 1, 0, 2, 0, 3, 0, 0, 2, 0, 1, 0, -2, -2, -1, -1, -1, 1, 1, 0, 0, -1, 0, 1, -1, 0, 0, 0, 0, 1, 2, 3, 2, 0, 3, 0, 2, -1, 0, 1, 1, 1, -2, 0, 0, -1, -2, 0, 1, 0, 0, 1, 0, -1, 1, 0, 1, 0, 0, 2, 1, 1, 0, 0, 3, 0, 3, 0, 0, -1, 0, -2, -1, -2, 0, -1, 0, 0, 0, -1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 3, 0, 0, 0, -1, 2, 1, 0, -1, 1, -1, -1, -1, 0, 1, 0, -1, 0, 0, 0, 0, 1, 0, 1, 1, 0, 2, 0, 0, 3, 0, 0, 2, 0, 0, 1, 0, 1, 0, -1, -3, -2, 0, -1, -1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 1, 0, 3, 1, 2, 0, 0, -1, -2, -2, 0, 1, -2, 0, 0, -1, -1, 1, 1, 1, 0, 0, 0, 1, 1, -1, 1, -1, 1, 1, 0, 1, 2, 1, 3, 3, 2, 0, 0, -1, 1, 0, -1, -1, 0, 0, -1, 1, 2, 0, 2, 0, 2, 0, 0, 0, 0, 2, 0, 3, 1, 0, 0, 3, 3, 0, -1, 0, 0, -1, 1, 1, -1, 1, 0, 0, 0, 1, 2, 0, 1, 2, 0, 0, 0, 1, 0, 1, 0, 1, 2, 0, 2, 0, 2, 1, 1, 0, 1, -1, 0, -1, 1, -1, -1, -2, 0, 2, 2, 1, 0, -1, 1, 0, 0, 1, 0, -1, 0, 2, 1, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, -1, 1, 0, 0, 1, -1, 0, 0, 0, 1, 2, 0, 0, 0, 1, 0, 2, 0, 0, 0, 1, 2, 1, 2, 0, 0, -1, -2, -2, 0, 1, 0, -1, 0, 0, -1, 0, 1, 0, 0, 0, -1, 1, -1, 2, 0, 1, -1, 2, 0, 2, 0, 2, 2, 0, 2, 1, 0, 0, -2, 1, 0, 0, -2, 1, 0, -1, 1, -1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 2, 2, 2, 1, 1, 1, 1, 0, 1, 0, -2, -1, 1, -1, 1, 1, 0, -1, 2, -1, 2, 0, -1, 1, 0, 0, 0, 1, 1, 0, 2, 1, 1, 2, 2, 1, 0, 0, 0, 0, 0, -1, 0, -2, 1, 0, 0, -1, 0, 0, 1, 0, -1, -1, 1, 2, 0, 1, 2, 0, 0, 2, 0, 0, 2, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, -1, 2, 1, 1, 2, 0, 0, -1, 1, -1, -1, 2, 2, 1, 0, 0, 2, 0, 0, -2, -1, 0, 0, -1, 0, -1, 0, 1, 0, 0, 0, 2, 1, 2, 1, 2, 0, 2, 1, 1, -1, 0, 0, 1, 2, -1, 2, 0, 0, -1, 0, -1, -2, 0, 0, -1, 0, -1, 0, -1, 2, 1, 1, 2, 0, 0, 1, 0, 1, 0, 2, 0, 0, 1, 2, 0, 0, -1, -2, 1, 0, 0, -1, 0, 0, 0, -1, 2, -1, 2, 2, 0, -1, 2, 1, 2, 0, 0, 0, 0, 3, 2, 0, 0, 2, 0, 0, 1, 1, 0, -1, 0, 0, 1, 0, -2, -1, 0, 0, 0, 1, 0, 2, 0, 2, 1, 2, 0, 2, 3, 2, 1, 3, 0, 2, 0, 1, 2, 0, 1, 0, -1, 0, -2, 0, 0, -2, -1, 1, -2, 0, -1, 0, 0, -1, 1, 0, -1, 0, -1, 0, 0, 1, 0, -2, -1, 0, -2, 0, 0, 0, 0, 0, -1, -3, 1, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -2, 0, 0, 1, 0, -1, -2, -2, -3, -3, -2, 0, -2, -1, 1, -2, 1, -3, 0, -2, 1, 0, 0, 0, 0, -2, 1, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, -3, 0, -1, 0, -2, -1, -3, -1, -3, -1, 0, 0, 1, -1, 1, -1, 0, 2, -2, -1, 0, -1, -1, 0, -2, -1, -1, -1, -3, -4, -2, 0, -3, 0, -1, -2, -1, -3, 0, 0, 2, -1, 0, 0, -1, 0, 0, 0, -1, 1, 0, 0, -2, 0, -2, -3, -2, 0, -4, -1, -2, -2, -3, -3, -4, -3, -3, -2, 0, 0, 1, 0, -3, 0, 0, -1, -2, 0, -1, -1, 0, 0, -2, -1, -1, -2, 0, -1, -2, -3, -2, -5, 0, -2, -3, -1, -4, -2, -2, -1, 1, -2, -2, 0, 1, -1, 1, 0, 0, -2, -2, -1, 0, -1, 0, -2, 0, -3, -2, -3, -3, -3, -1, -2, -1, -4, -1, -2, 0, 1, 0, -2, -2, 0, -1, -1, -1, -1, 0, 0, -1, -2, 0, -1, -1, -1, -1, -1, -1, 0, -2, -1, -2, 0, -3, -3, -1, -3, -2, 1, 1, 0, -2, 0, 0, -1, -2, 1, -1, 0, -2, -1, 0, 0, -2, -2, -2, 0, -2, 0, -3, -4, -1, -2, -2, -2, 0, -2, -1, 0, 0, -2, 0, -1, 1, -2, -2, -2, -1, 0, -2, 0, 0, 0, -1, 1, 0, -1, -2, -2, -2, -1, 0, -3, -1, -1, -2, -4, -2, -1, 0, -2, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -1, -2, -1, -1, -1, 0, -2, -4, -2, -4, 0, -2, 0, -1, -1, -1, -1, 0, 0, -2, 0, -2, -2, 0, 0, 0, -2, 1, 0, 1, -1, -3, -2, -1, 0, -2, 0, -2, 0, -1, 0, -3, 0, -1, -3, -3, -2, 0, 0, -2, -2, -1, -1, -2, -1, -1, -1, 0, 0, 0, 0, -2, 0, 0, 1, -1, -2, -1, -4, -2, -1, 0, -3, 0, -1, 0, -3, 0, 1, -1, 0, -1, 1, 0, 0, 0, 0, -1, 0, 0, 0, 0, 1, 0, 0, 0, -2, -1, -5, -4, -2, -1, 0, -1, -3, 0, -1, -2, 0, 0, -2, 0, 0, 0, -1, 1, -1, 1, -3, 0, -3, -2, -1, 0, 1, -2, 0, -4, -5, -2, -1, -1, -1, 0, 0, -3, -3, 0, 3, 0, 0, 0, -2, -2, -2, 0, 0, -1, -3, 0, -2, -1, 0, 0, 0, -1, -2, -5, -5, -1, -3, -3, 0, 0, -2, -2, -1, -1, 0, -2, 0, 0, 0, -1, 0, -2, -1, -2, 0, 0, -2, -2, -1, -1, 0, 0, -1, -5, -1, -5, 0, 0, -3, -2, 0, -2, -4, -1, 2, -2, 0, 0, 0, 0, 0, 0, -2, 0, -2, -3, -2, 0, 0, 0, 0, 0, -2, -5, -4, -3, 0, 0, -1, -2, -3, -3, 0, -2, 0, 0, -3, -1, -2, -2, 0, 0, -1, -2, -2, 0, 0, -2, 0, 0, -1, 0, -1, -1, -3, -5, -4, 0, -2, -1, -4, -1, -1, -1, 1, -3, -1, 1, 0, -2, 0, 0, 0, 0, -1, 0, -1, -2, 0, 0, 0, -4, -2, -1, -5, -1, 0, -1, -3, 0, -2, -3, -1, 0, 2, 0, 0, 0, 0, -1, 1, -1, -1, 0, -2, -2, 0, -2, -1, -1, -2, 0, -3, 0, -3, -5, -3, -2, -4, -1, -4, -4, 0, -1, 0, -2, 0, -1, 0, 1, 1, 0, -2, -1, -4, -3, 0, -3, -2, -2, -3, -1, -3, -2, -5, -3, -3, 0, -1, -3, -2, 0, 0, -2, 0, 0, -1, -2, -2, 2, 1, 1, 1, 0, -4, 0, 0, 0, 0, -2, -4, -3, -3, -3, -2, -3, -2, -3, -2, -1, -4, -3, -1, -2, 0, -2, 0, 1, 1, 0, 1, 0, -2, -3, -1, -1, -1, -3, 0, 0, 0, -1, -2, -1, -4, -4, 0, -1, -3, -1, 0, -4, -2, 0, 3, 0, 1, -2, -1, -1, 0, 0, -1, 0, 0, 0, 0, -3, -1, -3, -1, -2, -4, -2, -3, -3, 0, -2, 0, -2, -1, -2, -2, 1, 3, 0, 0, 0, -2, 1, 1, 0, 1, 0, -2, 0, -2, 0, -2, -3, 0, -1, -4, -4, -4, -1, -4, -1, -2, -3, 0, -1, 0, -1, 0, 0, -1, -1, -2, 0, 1, 1, 1, -2, -1, 0, -2, 0, -2, -2, 0, -1, -3, -3, -4, 0, 0, 0, -2, -1, 0, 0, 1, -1, 1, 0, 0, -1, -1, 2, 1, 1, 0, 0, 0, 0, 0, 0, -2, -2, -3, -2, 0, -3, -1, -1, -1, -2, 0, 0, -1, -2, 1, 2, 2, 0, 0, -1, 0, -1, 0, -1, 1, 0, -1, -2, -1, -3, -2, -4, -1, -2, -2, 0, -1, -1, -2, 0, 0, -1, 1, 0, 2, 2, 2, 0, -2, 0, 1, 0, 0, -1, 0, 0, 0, -2, 0, -4, -2, -1, -3, -2, -2, -2, -4, -1, -1, 0, -2, -2, 1, 1, 0, 0, 2, -4, -3, -1, -4, 0, -1, -1, 2, 0, 2, 0, -1, -1, 0, 1, 2, 3, 2, 2, 3, 4, 4, 5, 6, 9, 9, 8, 9, 12, 12, -5, -4, -3, -3, -1, -3, -1, 1, 2, 0, 0, 0, 0, 0, 3, 4, 2, 2, 3, 2, 1, 1, 3, 3, 3, 5, 6, 7, 9, 9, -3, -5, -2, -4, -1, 0, -1, -1, -1, -1, 1, 0, 1, 0, 0, 2, 6, 1, 0, 0, -1, -1, 0, 0, 1, 2, 0, 3, 5, 8, -2, -5, -1, -2, -2, -2, 0, 1, -1, 2, 0, -1, -1, 1, 0, 0, 0, 1, 0, -1, -1, -3, -2, -1, -1, 1, 1, 0, 2, 9, -2, -1, -2, -2, -3, 0, -1, 1, 0, 0, -1, 1, 1, 2, 1, 0, 4, 0, -3, -4, -4, -6, -6, -4, -5, -4, -1, 0, 2, 8, -5, -2, 0, -2, 0, -1, 0, 1, 0, 0, -1, 0, 1, 0, 0, 0, 2, 0, 0, -3, -4, -7, -6, -9, -6, -3, -1, -3, 1, 5, -3, -3, 0, 0, -1, 0, -1, -1, -1, 1, -1, 0, 0, 0, 2, 3, 1, 2, -1, -1, -4, -8, -6, -10, -6, -6, -4, -2, 0, 4, -5, -3, 0, 1, 0, 0, -1, 1, -2, -1, -1, -2, -2, 0, 2, 3, 6, 5, 2, 0, -2, -9, -5, -7, -6, -8, -4, -2, 0, 4, -4, -2, -1, 1, 1, 0, -1, 0, 1, 1, 0, 1, 3, 0, 1, 2, 6, 3, 5, 0, -2, -4, -8, -7, -7, -6, -6, -2, -1, 1, -3, -1, -2, 0, 3, 2, 1, 2, 0, 0, 2, 0, 3, 3, 5, 6, 5, 5, 4, 0, -4, -2, -5, -8, -6, -6, -6, -4, -1, 4, -4, -3, -2, 0, 3, 1, 2, 1, 3, 0, 1, 0, 0, 2, 3, 4, 6, 3, 5, 0, -3, -3, -6, -5, -9, -8, -6, -4, 0, 2, -7, -1, 0, 0, 3, 1, 2, 2, 0, 0, 0, 3, 2, 2, 4, 8, 8, 3, 0, -2, -7, -7, -6, -7, -9, -7, -7, -6, 0, 4, -4, -4, 0, 3, 2, 0, 2, 3, 2, 1, 1, 0, 1, 3, 5, 9, 9, 4, 0, 0, -6, -6, -7, -7, -6, -7, -5, -7, 0, 0, -3, 0, 2, 3, 1, 2, 3, 3, 3, 1, 2, 1, 2, 5, 7, 5, 8, 4, 2, 0, -7, -9, -9, -9, -8, -6, -7, -8, -2, 1, -5, 0, 0, 1, 5, 4, 1, 3, 3, 4, 1, 1, 1, 3, 7, 9, 8, 6, 4, 0, -5, -8, -5, -8, -5, -6, -5, -7, -3, 0, -4, 0, 1, 2, 3, 1, 2, 1, 1, 1, 1, 2, 4, 4, 6, 9, 8, 8, 4, 2, -4, -8, -5, -7, -5, -4, -7, -8, -2, 1, -2, 0, 0, 3, 4, 2, 3, 4, 3, 2, 2, 3, 6, 5, 9, 6, 8, 10, 3, 0, -6, -5, -4, -4, -7, -5, -8, -6, -5, 2, -3, 1, -1, 1, 0, 1, 1, 2, 0, 0, 2, 3, 1, 4, 7, 6, 10, 7, 2, -1, -5, -7, -8, -8, -8, -6, -8, -8, -4, 0, -1, -2, 0, -1, 0, 0, 1, 0, 0, 1, 2, 3, 4, 6, 6, 5, 5, 4, 3, -3, -6, -8, -5, -8, -6, -8, -7, -7, -4, 2, -5, -1, 1, 0, 0, -1, 1, -1, 0, 0, 0, 2, 2, 5, 2, 5, 6, 2, 1, -3, -5, -8, -7, -9, -9, -9, -7, -8, -4, 2, -6, -3, -1, -1, 0, 0, 0, -1, -1, -1, 1, 2, 4, 3, 5, 4, 7, 4, 2, 0, -5, -7, -8, -8, -8, -9, -6, -7, 0, 2, -7, -5, -4, -3, -2, -1, 1, 0, 2, 0, 1, 1, 1, 1, 3, 6, 4, 3, 3, 1, -4, -3, -5, -8, -9, -6, -7, -5, 0, 1, -4, -5, -3, -2, -1, 1, 0, -1, 1, 1, 0, 1, 2, 5, 4, 5, 5, 3, 3, 0, -3, -5, -4, -5, -5, -7, -6, -5, 0, 2, -4, -5, -3, -4, -4, -2, 0, 0, 2, 0, 0, 2, 1, 5, 5, 5, 7, 4, 3, 0, -1, -1, -6, -4, -4, -6, -2, -2, 0, 6, -2, -4, -4, -3, -3, 0, -1, 3, 3, 2, 0, 2, 2, 3, 7, 6, 5, 4, -1, 0, -2, -5, -5, -4, -5, -7, -6, -1, 0, 5, -5, -6, -2, -4, -1, -1, 0, 0, 0, 0, 2, 4, 4, 3, 6, 8, 9, 5, 2, -2, -2, -1, -6, -6, -5, -4, -2, 0, 1, 8, -6, -5, -3, -2, -1, 1, 0, 2, 1, 2, 3, 3, 5, 6, 7, 8, 6, 5, 0, -1, -1, 0, -1, -1, -4, -5, -3, 0, 3, 7, -4, -5, -3, -1, 0, 0, 1, 1, 0, 2, 5, 2, 5, 5, 6, 9, 5, 5, 1, 0, -1, 0, 0, 2, 2, 0, -1, 2, 3, 7, -1, -3, -5, -1, -1, 0, 0, 0, -1, 1, 4, 2, 5, 4, 7, 5, 8, 7, 7, 1, 3, 2, 3, 3, 2, 4, 2, 2, 5, 9, -2, -5, -2, -1, -1, 0, -3, -1, -1, 0, 0, 0, 5, 2, 3, 4, 5, 9, 7, 7, 6, 7, 8, 5, 8, 6, 8, 9, 7, 12, 2, 1, 0, 2, 2, 0, 0, -1, 0, -1, 0, 1, 0, -1, 1, 0, -1, -1, 0, 1, -1, -1, 1, 0, 1, -1, -2, -1, -1, 0, 2, 0, 2, 2, 0, 2, 0, 0, 0, 2, 0, 0, 2, 2, 1, -1, 1, 0, 0, 1, 1, -1, 1, -1, 1, 1, 0, 1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 0, 2, 1, 2, 0, 0, 0, 1, 1, -1, 0, 1, 1, -1, 1, 0, 1, -2, 1, -1, 0, 0, 0, -1, 0, 0, -1, 1, -1, -1, 0, 0, 1, 0, 2, 1, 2, 0, 0, 1, -1, 0, -2, 0, 1, 0, -2, 0, 0, 2, 0, 2, 1, -1, 0, 0, 0, 0, 0, 1, 0, 2, 0, 2, 0, 0, 0, 0, 0, -1, 0, 2, 0, -1, -1, 0, -2, 1, 2, 0, 1, 0, 1, -1, 0, 0, 2, 1, 1, 1, 1, 0, -1, 1, 2, 2, 0, 1, 0, 2, 1, 1, -1, 1, 1, 0, 0, -2, 2, 0, 0, -1, 2, 2, 1, 0, 2, 0, 0, 0, -1, 1, 0, 2, 1, 0, 0, 0, 0, 1, 0, 0, 2, -1, 0, -1, 0, 0, 0, 1, -1, 0, 2, 2, -1, 0, 1, 0, 1, 0, 0, 0, 1, 2, 2, 0, -1, 0, -1, -1, 0, -1, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, -1, 0, 1, 1, 0, 0, -1, 0, 0, -1, 1, 1, 2, 2, 0, 1, -1, -1, 1, 2, 1, 0, 1, 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 2, 0, -1, 1, 2, 2, 0, 1, 1, 1, -1, 0, 0, 1, 1, 0, 2, 0, 0, 0, -1, 1, 0, 2, 2, 1, 2, 0, 1, 2, 0, -1, -1, 0, 0, 1, 0, 1, -1, 0, 2, 0, -1, -1, 0, -1, 0, 0, 1, 0, -1, 0, 2, 2, 1, 0, 0, 0, 2, 0, 1, 0, -1, 0, 0, 1, 0, 2, 1, 0, 0, 1, 0, 0, 2, -1, 0, 1, 0, 1, 1, -1, 0, 0, 2, 1, 1, 0, 0, 0, 2, 1, 0, 2, 0, 2, 0, 0, 2, 2, 0, 0, 0, 0, -1, 1, 1, -1, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 0, 0, 2, 0, 0, 0, -1, 1, -1, 2, 1, -1, 0, 1, 0, 0, -1, -1, 0, 0, 0, 0, 0, 1, 0, 0, -1, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, -1, 1, 0, 1, 0, 0, 0, 0, -1, 0, -1, 1, 0, 2, 0, 1, 0, 1, 0, 1, 0, 2, 1, 0, 0, 1, -1, 0, 0, 0, 1, 2, -1, -1, 0, 0, -1, 0, 1, 1, 0, -1, 0, 0, 1, 1, 0, 1, 2, 2, 0, 2, 0, 0, -1, 1, 1, 0, 0, 0, 2, 0, -1, -1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 1, -1, 1, -1, 1, 1, 0, 0, 0, 1, 0, 1, -1, -1, 0, -1, -1, 1, 1, 0, 0, 1, 2, 0, 2, 1, 0, 0, 1, 1, 0, 1, 2, 1, 0, -1, -1, 1, 1, 0, -1, 0, -1, 1, -1, 1, 0, 0, 1, 1, 2, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 2, 2, -1, 0, 0, 1, 1, 0, -1, -2, -1, -1, 0, -1, -1, 1, 0, 1, 1, 2, 0, 2, 0, 0, -1, 1, -1, 2, 0, 1, 2, -1, 0, 0, 1, 1, 1, -1, -1, -2, 2, 1, 2, 0, 1, 2, 2, 1, 0, 0, 0, -1, 0, 1, 2, -1, 1, 1, -1, 1, 2, -1, 1, -1, 0, 1, 0, 1, 0, 1, 0, 1, 2, 2, 0, 0, 0, -1, 2, 0, 1, -1, 2, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, -1, -1, 1, -1, 1, 1, -1, 1, 1, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, -1, 2, 1, 0, -1, 0, 1, 1, -1, 0, 0, -1, 0, 1, 1, 0, 0, 0, 2, 1, 0, -1, 1, 0, 0, -1, 1, 0, 0, 1, 0, 2, 1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, 1, -1, 0, 1, 0, 0, 1, -1, 0, 0, 1, -1, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 1, -1, -1, -1, 1, 0, 2, 1, 0, 2, 0, 2, 0, 0, 0, 1, 0, -1, 1, -1, 0, 0, 1, 0, -1, 0, 1, -1, -1, 0, 0, -1, 0, 0, -2, -2, 0, -1, -1, 2, 0, 2, -1, 0, 0, 0, 1, -1, -1, 1, 0, 0, 0, -1, 0, 1, -1, -1, 0, -1, -2, 0, -1, 0, 0, 1, 0, 0, 2, 0, -1, 1, 2, 2, -1, 0, 0, 2, 0, 0, 0, 0, 0, 0, -1, -1, 1, 0, 0, 0, 0, -1, -1, -1, 0, -1, 0, 1, -1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, -2, -2, -1, 1, 0, 0, 0, -2, 0, 0, -2, -1, 0, 0, 1, -1, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, 1, -1, 1, 1, -1, -1, 1, 0, 1, 0, 0, -1, 1, 0, 2, 1, -1, -1, -1, 0, -1, -1, 2, 0, 0, 0, 1, -1, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1, -1, -1, 0, 1, -1, 0, -1, 1, 0, 1, 1, 0, -1, 0, -1, 1, 0, -1, 0, 0, 1, 0, 0, -1, -1, 0, 1, 1, -1, 0, 1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 1, 0, 0, 0, -1, 0, 0, 0, 0, -2, 1, 0, 1, 0, -1, -1, 0, 1, 0, 1, 0, -1, 0, -1, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, -1, 0, -1, 2, -1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, -1, 0, 1, 0, 1, 1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, -1, 1, -2, 0, 1, 0, 1, 2, 1, 1, 0, -1, 1, 0, 0, -1, 0, 0, 0, 0, 0, 1, -1, 1, 0, 0, -1, -1, -1, 0, 0, 1, 2, 0, -1, 0, -1, 0, -1, -2, 0, 0, 1, 0, -1, 1, 1, -1, 1, 0, -1, 1, -2, -1, 1, 0, 0, 0, 1, 0, 1, 0, 1, 1, 0, -1, -1, 0, 1, 1, 0, -1, 0, 0, 0, 0, 1, -1, -1, 1, 1, 1, 0, -2, -1, 0, 1, 1, 0, 0, 0, -1, 0, 1, 0, -1, 1, -1, 0, 0, 0, 1, 0, -1, 0, 1, 0, 1, 0, 0, 1, -1, 0, -1, 1, 0, 0, -1, 1, 0, 0, 1, 0, 0, 2, -2, 0, -2, 0, -1, -1, 0, -1, 0, 0, 0, 0, -2, 1, 0, 2, 0, -1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 2, 0, 0, 1, -1, -1, -1, -1, 0, 1, 1, 0, -1, 1, 0, 1, 1, -1, -2, 0, -1, 1, 0, 0, 0, -1, -1, 1, 1, -1, 0, 1, 1, 0, -1, 0, 1, 0, 1, 0, 0, -1, 2, 0, -1, -1, 1, 2, 0, -1, -1, 0, -1, 0, 0, 1, -1, 0, 0, -1, 0, 1, -1, -1, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 1, 0, 1, -1, 0, 1, 1, -1, -1, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, -1, 1, 0, 1, -1, 1, -1, 0, 0, 0, -1, -1, -1, 0, 0, -1, 1, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 0, -1, 2, -1, 0, 0, 1, 0, 1, 0, 1, 0, 0, 1, -1, 0, 0, -1, 1, -1, 1, -1, 0, 0, 0, 1, 0, -1, 0, 1, -1, 0, 0, 0, 0, 0, -1, -1, -1, 0, -1, -1, 0, 0, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, -1, -1, 0, -1, 1, -1, -1, -1, -1, 0, 0, 0, 1, 0, -1, 0, 0, 0, 1, 0, 0, -2, 0, 0, 1, 0, 0, 0, 1, 1, 2, -1, 1, 0, 1, 1, 0, 0, 0, 0, -1, -2, 1, -1, 1, 1, 0, 1, 0, 1, 1, -1, 0, 0, 2, -1, 0, -1, 0, -1, 0, -1, -2, 1, -2, 1, 0, -1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 2, -1, 1, 1, 0, -1, 1, 0, 1, -1, -1, -1, -1, 0, -1, 0, -1, 2, 1, -1, 1, 0, 1, 1, 0, 0, -1, -1, 1, 0, 1, 1, 0, 0, 0, 0, -2, 0, -1, 0, 1, 0, 0, 2, 1, 1, 0, 1, 0, 0, 1, -1, 0, -1, 1, 1, 0, -1, 1, 1, 0, 0, 1, -1, -1, 0, -1, 2, -1, -1, 2, 1, 0, -1, 0, -1, 1, 0, 0, -1, 1, 0, 1, -1, 0, 1, 0, -1, -1, 0, -1, 0, 2, 1, 0, 1, -1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 2, 0, 1, 0, 0, 0, -1, -1, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, -1, 0, -1, 0, 0, -1, 1, 0, -1, 0, 0, -1, -1, 0, 1, 0, -2, 0, 1, 0, 1, -1, 1, -1, 1, 0, 0, -2, 0, 0, 2, 0, 1, 0, -1, 1, 1, 1, 0, 0, 2, 0, 0, 0, 0, 1, 2, 0, 0, 2, 0, 2, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, -1, 1, -1, 0, 1, 1, 0, -1, -2, -1, -1, 0, -1, 0, 0, -1, 0, 2, 1, 0, 1, 0, -1, 1, 0, -1, 1, 0, 0, -1, 1, -1, -2, 1, 0, 0, -1, -1, 1, 0, 1, 1, 1, 1, -1, 0, 1, -1, 0, 0, -1, 0, 0, -1, 0, 0, -1, 1, 0, 1, -1, 0, -1, -1, 1, 0, -1, 0, -1, 0, -1, 0, 0, 0, -1, 0, -2, 2, 0, -1, 0, -1, 0, -1, 0, 1, -1, 1, 0, 2, 0, 0, 1, 1, 1, 1, 1, 1, 1, -1, -1, 0, 0, 0, -1, 0, -1, -1, 0, 1, 0, -1, 0, 1, 0, -1, 0, 0, 0, -1, -1, 0, 0, 1, 1, 0, 0, 11, 7, 6, 4, 5, 2, 1, 1, 2, 0, 0, -3, -7, -10, -12, -9, -10, -9, -10, -7, -7, -6, -4, 1, 2, 9, 10, 9, 12, 16, 11, 9, 6, 4, 2, 1, 0, 2, 1, 0, 0, -4, -5, -5, -5, -5, -4, -4, -8, -7, -7, -5, -2, -1, 1, 6, 6, 7, 7, 10, 10, 5, 2, 1, 1, 0, -1, 0, 0, 0, 1, 0, -3, -2, -1, -1, -1, -3, -6, -4, -4, -3, -1, 0, 1, 1, 1, 3, 3, 11, 6, 4, 3, 2, 0, 0, 0, 1, 1, 1, 1, -1, -1, 0, 0, -2, 0, -2, -3, -6, -6, -4, -5, 0, 1, 0, 0, 0, 2, 9, 8, 6, 4, 3, -1, -1, 0, 0, 1, 0, 0, 0, 0, 0, 0, -1, 0, -3, -4, -6, -4, -8, -7, -3, -3, -5, -4, -4, 3, 7, 9, 5, 1, 3, 2, 0, -1, 2, 1, 0, -1, -2, -3, -3, -1, 0, -1, -4, -3, -6, -5, -9, -6, -6, -9, -5, -4, -5, 1, 8, 4, 3, 0, 0, 1, -1, 1, 2, 0, 2, -3, -1, -1, -3, -5, -1, -2, -2, -3, -7, -6, -7, -7, -7, -9, -6, -8, -5, -2, 3, 3, 1, 0, 0, -1, 0, 0, 0, 0, 0, -3, -2, -4, -2, -3, -5, -1, -3, -5, -6, -7, -10, -6, -8, -10, -7, -8, -5, 0, 3, 1, -1, -2, -4, -1, 0, 2, 0, 1, 0, 0, -1, -3, -3, -5, -3, -3, -3, -2, -1, -8, -7, -9, -7, -8, -6, -8, -5, -2, 5, 1, -6, -8, -4, -3, -1, 0, -1, 0, -1, 0, -2, -5, -2, -2, -3, 0, 0, -1, -5, -8, -5, -5, -4, -7, -8, -3, -2, 0, 4, 0, -4, -6, -5, -5, -2, -1, -2, 0, 0, -4, -3, -3, -5, -4, 0, -2, 0, -1, -6, -7, -9, -4, -5, -6, -7, -4, -3, -1, 6, 0, -4, -5, -7, -5, -3, -5, -4, -1, -1, -2, -3, -6, -4, -4, 0, 1, 0, -1, -5, -8, -6, -6, -5, -4, -2, -6, -3, 1, 6, 3, -3, -3, -4, -5, -6, -5, 0, 0, -1, -1, -2, -6, -5, -2, 1, 1, 0, 0, -2, -8, -7, -4, -5, -4, -3, -6, -3, 2, 8, 2, 0, -1, -6, -3, -3, -3, 1, 3, 0, -1, -5, -3, -2, -1, 2, 5, 6, 4, 1, -7, -9, -7, -5, -5, -4, -4, -3, 0, 5, 7, 0, -1, -2, -2, -2, -3, 1, 2, 3, 0, -4, -3, -4, 0, 4, 5, 8, 3, 0, -3, -5, -7, -5, -5, -1, -1, 0, 0, 6, 6, 1, -1, -4, -1, -2, 0, 1, 3, 0, 0, -1, -2, -3, 0, 5, 8, 8, 4, 0, -7, -6, -6, -4, -1, 0, -1, 0, -2, 5, 5, 0, -1, -3, -2, -2, -3, 1, 1, -1, 0, -3, -4, -1, 1, 6, 6, 3, 1, -5, -8, -5, -3, -4, -1, -1, -4, -1, -1, 5, 6, 0, -3, -6, -2, -4, -2, -3, 0, -1, 0, -3, -5, -1, -1, 4, 2, 1, -3, -2, -9, -7, -5, -5, -1, -3, -2, -4, -1, 7, 4, -1, -3, -2, -3, -5, -3, 0, -2, 0, -3, -2, -3, -4, -2, 1, 4, 0, -3, -4, -8, -6, -4, -6, -6, -6, -7, -3, -2, 7, 6, 0, -5, -5, -6, -4, 0, 0, 0, 0, -3, -3, -4, 0, 0, 2, 0, 0, -2, -4, -3, -6, -4, -7, -4, -5, -9, -4, 0, 7, 4, -2, -3, -3, -2, -2, 0, 2, 0, 0, -1, -3, -1, -1, 2, 2, 2, 0, -2, -5, -3, -7, -7, -5, -5, -8, -8, -3, 0, 7, 6, -1, 0, -1, -4, -1, 1, 4, 3, 2, -4, -3, -3, -4, 0, 0, 2, -2, -2, -5, -7, -6, -3, -4, -6, -5, -5, -5, -3, 5, 5, 0, -1, -4, -1, 0, 1, 2, 2, 0, -3, -5, -3, -3, 0, 1, 0, -3, -3, -6, -6, -7, -3, -4, -6, -7, -6, -3, 0, 5, 6, 3, 0, -1, 1, 1, 1, 2, 0, 0, -4, -4, -2, -1, -2, 1, -1, -3, -6, -9, -8, -5, -6, -5, -7, -6, -8, -6, -2, 4, 4, 4, 0, -1, 3, 1, 1, 2, 3, -1, -1, 0, -5, -3, -2, 0, 2, -3, -5, -8, -10, -9, -8, -8, -7, -8, -9, -4, -1, 8, 7, 2, 4, 1, 2, 2, 4, 3, 0, 1, -1, 0, -5, -2, 0, 1, 0, -1, -5, -6, -11, -11, -8, -8, -8, -5, -4, -4, 1, 7, 8, 4, 2, 0, -1, 1, 3, 3, 0, 0, 0, -3, 0, 0, -2, 2, 0, -4, -8, -8, -9, -10, -3, -4, -4, -3, -2, -2, 1, 10, 5, 3, 2, 0, 0, 0, 1, 0, -1, -2, -2, 0, 0, 0, -3, 0, -2, -2, -6, -10, -9, -5, -4, -3, -3, -2, -1, 2, 6, 12, 8, 4, 3, 0, -1, 3, 1, 1, -2, -3, -1, -1, -3, -4, -1, 0, -5, -5, -5, -5, -4, -2, -3, -1, -2, 0, 3, 2, 7, 15, 7, 5, 1, 0, 0, 2, 0, 1, 0, -3, -4, -4, -3, -3, -6, -6, -7, -8, -7, -7, -4, -2, -1, -1, 1, 4, 2, 6, 9, 15, 4, 4, 2, 4, 0, 0, 2, 0, 0, 0, 1, 0, -2, 0, -3, -3, -2, -2, -3, -4, -3, -1, -2, -1, 1, 0, 3, 3, 2, 3, 5, 6, 5, 3, 2, 0, 0, 0, 1, 0, 1, 1, 0, 0, 0, -1, -1, -3, 0, -1, -1, -1, 0, -1, -1, 2, 0, 0, 0, 0, 3, 3, 1, 0, 3, 0, 2, 0, 1, 2, 0, 0, 2, 0, -1, 1, -1, -2, 0, -1, -1, 0, 0, -1, 1, 1, 0, 0, -1, 0, 2, 5, 1, 1, 1, -1, 2, 0, 2, 0, 1, 1, 0, 0, 0, -1, 0, 0, 1, 0, -1, 0, -1, -2, 0, 0, 0, -1, -1, 2, 3, 2, 1, 2, 3, 1, 0, 0, 1, 0, 0, 1, 0, 2, 0, 0, 2, 1, 0, -2, 0, 0, -1, -1, -1, 1, -2, -1, 0, 1, 5, 2, 3, 2, 2, 0, 2, 0, 3, 0, 0, 0, 0, 1, -1, 2, 1, 1, 0, 0, 0, -2, -2, 0, -1, -1, -1, -2, -1, -1, 5, 3, 2, 2, 0, 0, 3, 3, 2, 1, 0, 0, 1, 0, 0, 0, 1, -1, 0, 0, 1, 0, -3, -1, -2, -2, -1, -2, -2, 0, 4, 1, 0, 0, 0, 2, 1, 0, 1, 0, 0, 0, 1, -2, 0, 0, -1, 0, 1, 0, 1, -1, 0, -2, -2, -3, 0, -2, 0, 2, 1, 1, -1, -2, 1, -1, 1, 0, 0, 1, 0, -1, -1, 0, -1, 0, 0, -1, 0, -1, -2, -1, 0, -1, -3, -2, -2, 0, 0, 1, 3, 1, 0, 0, -2, -2, -1, 0, 0, -1, 0, 0, 1, -1, 1, -1, 0, 0, 0, 0, 0, 0, -1, 1, -2, 0, -2, -1, 0, 0, 0, -1, -2, 0, -1, 0, 0, 0, 2, 0, -1, -1, -2, 0, 1, -1, 0, 2, 2, 0, 0, -2, -2, 0, 0, 1, 0, 0, -1, 1, 3, -1, -2, 0, 0, -1, -1, 1, 1, -1, 1, -2, -1, -2, 1, 0, 1, 0, 3, 2, 0, -3, 0, 0, -1, -1, -1, 0, 0, 0, 2, 0, 0, -2, 0, -2, -2, 0, 0, 0, 0, 1, 0, 1, 1, 2, 1, 2, 3, 2, 0, -1, 0, 0, -1, -1, 1, 0, -1, 2, 0, 0, 0, 1, -1, -1, 0, -1, 0, 1, 0, 1, 0, -1, 1, 0, 2, 2, 4, 2, -2, -2, -2, -1, -1, 0, -1, -1, 0, 0, 1, 1, -2, 0, -1, -2, -2, 0, 2, 1, -1, 0, 0, -1, 0, 1, 2, 3, 4, 1, 0, -1, 0, 0, 0, 0, -1, -2, 0, 1, 1, 0, -1, 0, 0, 0, 0, 0, 2, 0, 0, 2, 1, -1, 0, 0, 3, 4, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 1, -1, -1, 0, -2, -2, -1, 0, 0, 1, 0, 1, 1, 1, 0, 2, 3, 0, 2, 1, -2, 0, 0, 1, 0, 1, 0, 0, 1, 3, 2, 1, 0, -1, -1, 0, 1, 0, 1, 2, 1, 0, 1, 2, 0, 3, 1, 2, 0, -2, 0, -1, 0, 0, 1, -1, 0, -1, 1, 1, 1, 1, 0, -3, -2, -1, 1, -1, 0, -1, 0, -2, 0, 2, 1, 0, 3, -1, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 2, 4, 0, -2, -1, -2, 0, -1, -1, 0, -1, 1, 0, 0, 1, 0, 0, 1, 0, 1, 0, 0, 0, -2, 0, -2, -1, -1, -1, 0, 1, 2, 0, 1, 0, 0, 1, 2, 0, 2, 0, 0, 0, -1, 1, 0, 3, 3, 3, 0, 0, 2, -1, -1, 0, 1, -2, 0, -2, -1, 0, 3, 0, 1, 0, -1, -1, 0, 1, 0, 0, 0, 0, -2, 1, 2, 1, 0, 1, 2, 1, -1, -2, 0, 0, -2, 0, -1, 0, -1, 0, 2, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 0, -1, -1, -3, 0, 0, 0, 0, -2, 0, -1, -1, 3, 3, 3, 0, 0, 0, 2, 1, 0, 0, -1, 0, -2, -1, 0, -1, 1, 1, 0, 0, -2, -2, 0, 0, 0, 0, 0, 0, -2, 1, 2, 1, 1, 2, 1, 0, 1, 1, 2, 0, -1, -1, -2, -1, 1, 0, 0, 0, 0, -1, 0, -1, -1, 0, 0, -3, -4, 0, 1, 2, 3, 4, 4, 0, 0, 0, -1, 2, 0, -1, 1, 0, 0, -1, 0, 2, 0, 0, 1, -2, -3, -3, -1, -1, -2, -2, -3, -1, 1, 3, 4, 1, 1, 0, 1, -1, 2, -1, -1, 1, -1, -2, 0, 1, 0, -1, 0, 0, 0, 0, -1, 0, 0, 0, 0, -3, 0, -2, -1, 1, 4, 3, 0, 0, 0, 1, 2, 2, 0, 1, 1, -1, -1, 1, -1, 0, -1, 0, 0, -2, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 4, 4, 2, 2, 0, 1, 1, 0, 0, -1, -1, 1, 0, -1, -1, 0, -1, 0, -3, -3, -2, -3, -2, 0, 0, -1, 1, 2, 3, 3, 2, 4, 4, 0, 3, 0, 0, 1, 0, -1, 0, 0, -2, -2, 0, -3, -3, -1, -3, -2, -4, -1, 0, -2, 1, -1, 2, 0, 1, 4, 20, 16, 12, 7, 7, 3, 4, 2, 1, 4, 1, -1, -3, -5, -6, -4, -4, -8, -12, -8, -11, -8, -5, -2, 2, 7, 10, 11, 13, 18, 17, 11, 10, 4, 3, 0, 1, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, -3, -8, -7, -6, -8, -3, 0, 3, 3, 5, 7, 10, 16, 16, 9, 7, 4, 3, 0, 0, 2, 3, 3, 4, 4, 0, 3, 0, 1, 1, 0, -3, -5, -8, -6, -2, -2, -1, 3, 0, 0, 6, 14, 15, 12, 6, 3, 3, 0, 1, 5, 5, 2, 1, 1, 2, 1, 3, 2, 2, 0, -2, -6, -7, -4, -5, -5, -4, 0, 0, 0, 1, 13, 17, 12, 7, 7, 5, 0, 3, 2, 3, 4, 3, 0, 0, 0, -1, -1, 1, -1, -3, -4, -6, -4, -4, -4, -7, -6, -5, -2, -1, 9, 13, 6, 5, 5, 2, 4, 1, 3, 5, 1, -1, -2, -3, -3, -2, 0, 0, -1, 0, -5, -7, -6, -7, -9, -9, -7, -5, -3, 1, 8, 13, 6, 4, 2, 2, 1, 4, 3, 4, 4, 1, 0, -3, 0, -2, 0, 0, 0, 0, -3, -6, -9, -8, -9, -8, -11, -8, -7, -3, 7, 10, 1, 0, -1, 0, 3, 4, 3, 3, 5, 1, 0, -1, 0, -4, -3, -1, 0, 0, -2, -1, -5, -3, -6, -6, -10, -8, -5, -2, 6, 6, -2, -6, -3, -3, -2, 0, 2, 1, 3, -1, -3, -2, -5, -2, 0, -1, 0, 3, 0, -1, -6, -6, -5, -6, -8, -6, -3, 2, 7, 6, -3, -6, -7, -4, -2, 0, -1, 1, 1, -2, -4, -2, -3, -3, 0, 1, 2, -1, 0, -5, -7, -4, -4, -2, -3, -5, 0, 2, 7, 4, -2, -4, -5, -7, -3, -4, -2, -1, -3, -2, -4, -3, -5, -1, 2, 6, 5, 0, -4, -7, -6, -6, -3, -1, -2, -3, -1, 0, 7, 8, 0, -3, -4, -5, -7, -5, 1, 2, 1, -1, -2, -7, -4, 0, 5, 6, 5, 3, 0, -3, -6, -5, -3, 0, -3, -2, 0, 0, 9, 10, 2, -1, -1, -3, -3, -3, 0, 5, 4, 0, -3, -6, -2, -2, 4, 8, 9, 9, 7, 1, -5, -5, -4, 0, -1, 0, -2, 0, 8, 11, 2, 0, -2, -1, -2, 0, 0, 2, 5, 0, 0, -4, -1, 0, 5, 12, 13, 12, 6, 1, -2, -1, -3, 0, 1, 0, 1, 3, 11, 12, 1, -2, 0, -3, -1, -2, 4, 4, 6, 1, 0, 0, -1, 3, 9, 14, 14, 11, 9, 1, -2, 0, -2, 1, 0, 2, 0, 3, 10, 15, 2, 0, -2, -1, -3, -2, 1, 2, 2, 3, 0, 0, 0, 5, 8, 12, 13, 10, 2, -2, -3, 0, 0, 0, 0, 0, -1, 1, 9, 11, 1, -2, -6, -4, -6, -1, 0, 0, 2, 1, -2, -1, -3, 1, 6, 6, 8, 2, -1, -3, -4, -5, -1, -1, 0, 0, 0, 0, 9, 10, 3, -2, -3, -2, -3, -2, -3, 0, 1, 0, 0, -1, -2, 0, 6, 4, 6, 3, -1, -4, -2, -4, -1, -4, -1, -1, -2, 1, 8, 11, 1, -3, -6, -5, 0, 1, 1, 1, 1, 0, -2, -3, 0, 2, 6, 6, 7, 1, 0, -1, -1, -4, -5, -2, -3, -5, -3, 0, 10, 12, 1, -4, -4, -6, -3, 0, 3, 3, 2, 1, -2, -2, 0, 2, 6, 5, 4, 4, 1, 0, -3, -5, -5, -4, -4, -4, -2, 1, 8, 14, 4, -3, -2, -2, -1, 1, 3, 5, 4, 0, -1, -2, -2, 2, 5, 5, 2, 1, -1, -2, -3, -2, -3, -3, -3, -3, -3, 0, 10, 11, 7, -1, 0, -3, 0, 1, 7, 6, 3, 0, -2, -4, -2, 3, 6, 5, 0, -2, -2, -4, -1, -4, -3, -4, -5, -5, -2, 0, 9, 13, 5, 4, 0, -1, 0, 4, 7, 5, 2, -1, -4, 0, -1, 1, 5, 5, 0, -2, -4, -6, -4, -3, -5, -4, -6, -7, -5, 0, 7, 12, 7, 6, 4, 3, 3, 5, 7, 4, 0, 0, 0, -1, 0, 0, 4, 4, 4, 0, -6, -7, -5, -7, -5, -7, -7, -8, -6, -1, 9, 11, 9, 4, 5, 1, 3, 3, 3, 3, 3, 1, 0, 0, 0, 0, 1, 5, 1, 0, -7, -8, -9, -5, -6, -6, -7, -8, -5, 1, 11, 14, 9, 4, 4, 3, 0, 3, 4, 2, 2, 0, 2, 0, 0, 2, 0, 4, 2, -2, -9, -11, -10, -4, -2, -3, -1, -5, -2, 2, 12, 16, 11, 5, 3, 0, 0, 3, 2, 0, 0, 0, 2, 1, 2, 1, 0, 2, 1, -3, -9, -9, -6, -2, -2, 0, 2, 1, 2, 6, 14, 12, 7, 3, 1, 3, 1, 2, 0, 0, 0, 0, 2, 1, -1, 0, 0, 1, 0, -3, -2, -3, -3, 0, 0, 3, 1, 2, 6, 9, 18, 15, 8, 5, 5, 2, 2, 4, 3, 2, -1, -2, -3, 0, -2, -2, -3, -6, -4, -6, -4, -1, 0, 3, 1, 2, 5, 8, 11, 16, 22, 15, 11, 5, 6, 3, 5, 1, 0, -2, -3, -4, -2, -7, -8, -10, -11, -13, -15, -12, -11, -9, -1, 0, 3, 5, 6, 10, 13, 15, 21, 6, 4, 2, 6, 0, 1, 3, 0, 4, 1, -3, -2, -3, -3, -6, -5, -3, -6, -3, -3, -2, 0, 2, 1, 1, 3, 7, 7, 8, 7, 3, 5, 4, 1, 1, 0, 0, 1, 0, -1, 0, -2, -2, -2, 0, -3, -5, -5, -4, -1, -2, 0, 0, 3, 4, 3, 3, 6, 4, 6, 2, 2, 2, 1, 3, 3, 4, 3, 1, 2, 2, 0, 0, 0, 2, 1, -1, -2, -4, 0, -2, 0, 0, 1, 3, 0, 0, 3, 3, 5, 4, 3, 4, 1, 2, 1, 0, 2, 3, 0, 0, 0, 1, 0, 0, 0, 0, -2, 0, 0, -1, 1, 2, 2, 5, 0, 1, 5, 4, 7, 4, 4, 4, 3, 0, 3, 2, 2, 2, 0, 2, 4, 2, 2, 1, 1, 1, -2, -1, 0, 0, 1, 0, 3, 3, 3, 3, 0, 5, 7, 4, 1, 1, 4, 0, 0, 4, 2, 1, 2, 0, 0, 3, 2, 2, 1, 2, 0, -1, 0, -1, 0, 1, 1, 3, 2, 1, 0, 4, 8, 2, 2, 3, 3, 2, 0, 2, 3, 0, 0, 0, -1, 1, 2, 1, 2, 1, 1, 1, -1, -1, 0, 2, 2, 0, 0, 0, 3, 4, 8, 0, 0, 3, 5, 3, 2, 2, 0, 0, 1, -1, -1, 0, 0, -1, 2, 0, 0, 0, -2, 0, -2, 0, 0, 0, 0, 0, 2, 4, 5, 0, 1, 0, 3, 3, 1, 0, 0, 0, 1, 0, 2, 0, 0, 1, 1, 0, 0, 2, 0, -2, -1, 0, -1, 0, 0, 1, 0, 1, 7, 0, 1, 0, 1, 3, 1, 4, 1, 2, 2, -1, 0, -1, 2, 1, -1, 2, 0, 1, 1, 2, 0, 0, 0, 0, 0, 2, 1, 2, 6, -3, -1, -2, 0, 0, 1, 3, 0, 0, 1, 2, 1, 0, 1, 1, 2, 1, 0, 0, -1, -1, 2, 1, 0, 0, 0, 0, 2, 4, 7, -2, -4, 0, 0, -2, 2, 1, 2, -1, 0, 0, 0, -1, 0, 1, 4, 0, 0, 0, 0, 1, 1, 4, 0, 3, 0, 0, 0, 5, 8, -3, -2, 0, 0, 0, 0, 0, 0, -1, -2, -3, 1, 1, 0, 1, 1, 1, 1, 2, -1, 1, 0, 3, 2, 1, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 1, 1, 2, -1, 0, 0, -1, 0, 3, 2, 2, 2, 3, 0, -1, 0, 1, 2, 0, -1, 1, 1, 4, 9, 0, -2, 0, 2, -1, -1, 1, 4, 2, 1, 1, 0, 1, 0, 2, 5, 3, 3, 3, 0, 0, 3, 0, 1, 1, 1, 0, 0, 3, 7, -2, 0, 0, 0, 0, -1, 3, 2, 2, 1, 1, 1, 1, 3, 3, 3, 4, 5, 1, 3, 0, 2, 1, 0, 0, 2, 0, 0, 4, 7, 0, -1, -1, 1, 0, 1, 0, 4, 3, 1, 1, 2, 3, 4, 2, 6, 6, 6, 4, 2, 2, 1, 4, 4, 3, 2, 0, 2, 2, 7, 1, -2, 0, 1, 0, -1, 1, 3, 0, 0, 0, 0, 0, 1, 3, 5, 3, 2, 2, 1, 3, 1, 2, 2, 4, 1, 2, 3, 2, 6, -2, 0, 0, 2, 0, -2, -1, -1, -1, 0, -1, 0, 0, 2, 0, 5, 2, 0, 0, 0, 0, 3, 2, 0, 1, 1, 3, 1, 2, 8, 1, -1, -2, 2, -1, 1, 0, 0, 1, 0, 1, 2, 1, 0, 3, 5, 4, 0, 0, 2, -1, 1, 2, 1, 2, 1, -1, 1, 2, 7, -2, -2, -2, 1, 0, 1, 0, 1, 0, 0, -1, 0, 0, 4, 4, 3, 2, 3, 4, 0, 0, 0, 2, 0, 1, -1, -1, 3, 2, 8, 0, -1, -1, 0, -1, 0, 1, 0, 0, 1, 0, 1, 0, 1, 5, 3, 3, 3, 3, 3, 3, 2, 0, 3, 1, 1, 0, 0, 1, 7, 0, 1, 2, 1, 0, 0, 2, 1, 0, -1, -2, -1, -1, 2, 4, 0, 0, 0, 1, 0, 1, 3, 4, 0, 0, 2, 0, 0, 4, 5, 0, 0, -1, 1, 1, 2, 1, 0, 2, -2, -2, -2, -1, 0, 1, 3, 2, 0, 0, 1, 1, 2, 5, 3, 1, 0, 0, 0, 2, 7, 0, 2, 1, 3, 3, 4, 0, 0, 0, 0, -2, 0, 0, 1, 2, 2, 2, 1, -1, -1, -1, 0, 2, -1, -1, 0, 0, 0, 4, 8, 1, 3, 4, 2, 2, 3, 1, 2, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 1, 2, -1, 0, 0, -1, -3, 0, 1, 4, 8, 2, 0, 1, 3, 3, 3, 3, 0, 1, 0, 0, 0, 0, 1, 2, 0, 0, -1, -2, -3, -2, 1, 0, 1, -1, -1, -1, 1, 4, 6, 1, 0, 1, 2, 1, 2, 2, 0, 1, 3, 1, -1, -1, 2, 0, 2, -1, 1, -2, -1, -1, 0, 0, 2, 0, 0, 1, 1, 2, 8, 1, 4, 3, 1, 0, 3, 0, 0, -1, 0, 0, 3, 0, 0, 0, -1, 0, 1, -2, 0, 0, 0, 0, 2, -1, 0, 0, 0, 3, 7, 0, 2, 0, 1, 1, 2, 0, -1, -1, 1, -1, 2, 1, -1, 1, 2, 0, 1, 1, 3, 1, 0, 1, 2, 0, 0, 2, 1, 5, 9, -1, 0, -2, 1, 1, -1, 0, 0, -2, -1, 0, 0, 0, 1, 2, -1, 1, -1, -1, 0, -1, -1, -1, 1, 0, 0, 1, 0, -1, 0, 1, 0, 1, 1, -1, -1, 0, 1, 0, 0, 0, 0, 0, -1, 0, 1, 0, 0, 1, 1, -1, 1, -1, 1, 2, -1, -1, 0, 1, 0, -1, 1, 0, 0, 0, 0, -1, -1, 0, -1, 0, 0, 0, 1, -1, 0, 0, 0, 1, 0, -1, 0, 1, 1, 0, -1, -1, 1, 1, 0, -1, -2, 1, 1, 1, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 0, 1, -1, 1, 0, 0, 0, 1, 0, 1, 1, 0, -1, 0, -1, 1, 1, 2, 0, -1, -1, 0, -1, 1, 0, -1, 0, 2, -2, 1, -1, -2, 1, 1, 0, 1, -1, 0, -1, 0, 0, 1, 1, 0, 0, -2, -1, 1, 1, -1, -1, -1, -1, 0, 2, 0, 0, 1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 1, 0, 1, -1, -1, 2, -1, 0, 0, 0, 0, 1, 1, 0, 0, -1, 1, 0, 1, 1, 0, 0, 1, 1, -1, 0, 1, 0, -1, 0, 0, 1, -2, -1, 2, 0, -1, 0, 0, -1, -2, 0, 0, 0, 0, 1, -2, -1, 0, 1, 1, -1, 0, 0, 2, -1, -1, 0, 0, 0, 0, 0, 1, 2, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 1, 1, 0, 0, 1, 0, -1, 0, 0, 0, 1, -1, 1, 0, -1, 2, 0, 1, 1, -1, 1, 2, -1, -1, 1, 1, -1, 1, 0, 0, 1, 0, 1, 0, 1, 1, -1, 0, 1, -1, -1, 0, -1, 0, 1, 0, -1, -1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 1, 0, 1, 0, 0, 0, 1, -1, 0, 0, 1, 2, 1, -1, 0, 1, -1, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 0, 0, 0, -1, 2, 1, -1, 2, 0, 1, -1, 0, 0, 0, 0, 2, 1, 1, 0, -1, 1, -2, -1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0, 1, 0, 0, 0, -1, 0, 0, -1, 0, -1, -1, -1, 0, 0, 0, 0, -1, 2, 0, -1, 0, 0, 1, -2, 0, 1, 1, 1, -1, 1, 0, 0, 1, 0, 0, 1, -1, 0, -1, 0, 0, 1, 0, 1, 1, 1, -1, 0, 0, 1, 0, 0, 0, 0, 1, -1, 1, 0, -1, 1, 0, 2, 0, -1, 0, 0, 0, 0, -2, 1, 1, 0, 1, 0, 0, 1, -1, -1, 0, 0, 1, 0, 0, -1, 0, -1, 0, 0, -2, 0, -1, 0, 0, 1, -1, 2, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, 1, -1, 0, 0, -1, 1, -1, 1, -1, 0, -1, 0, 0, -1, 0, 0, 1, -1, 2, 0, -2, 1, 0, -1, -1, -2, 0, 0, -1, -1, 0, -1, 1, 1, -1, 1, 0, 0, -2, 0, 0, 1, -2, 0, 0, -1, -1, -1, 1, 0, 0, 1, -1, 1, -1, 0, 0, -1, 0, -1, -1, 1, -1, 0, 0, -1, 0, -1, 0, -2, -1, 1, 0, 0, 0, -1, 0, 1, 0, -1, 0, -1, 1, -1, 0, 1, 0, 1, 0, -1, 0, 1, -1, 0, -1, 1, 1, 1, 0, -1, 1, -1, 0, 1, 1, 0, -1, 0, 1, 0, 0, -1, 0, 0, -1, -1, -1, 0, 0, 1, 1, -1, 0, 0, -1, 1, -1, 0, 1, 0, 0, 1, 0, 0, 0, -1, 0, 0, 0, 1, -1, 0, 1, 1, 0, 1, 0, 0, -1, 0, -1, 0, 0, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, -1, 1, 1, 1, 0, 1, 0, 2, 1, 1, -1, 1, -1, -1, -1, 0, 2, 1, 0, -1, 0, -1, 0, 0, 1, 0, 0, -2, -1, 0, 0, 1, 0, -1, 0, 0, 0, 0, -2, 0, 0, -1, 0, 0, 2, 1, -1, 1, -1, 0, 1, 1, 0, 0, 0, -1, 0, -1, 0, 1, 1, -2, -1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 0, 1, 1, 2, 0, -1, 1, -1, 1, 1, 0, 0, 1, 0, 0, 1, 1, 0, -1, 0, -1, 0, 1, 0, 0, 0, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, 0, -1, 0, -1, -1, 2, -2, -1, 0, 0, -2, 0, -1, -1, -1, 0, 0, 1, 0, -1, 0, 0, 1, 1, 0, 0, 0, -1, 1, -1, 1, 0, 0, 1, 0, -1, 1, -1, 1, 0, -2, -1, 0, -1, -1, -1, -1, 0, 0, 1, 1, 0, 0, 0, -1, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 2, -1, 1, 2, 1, -1, -1, 2, 0, 0, 2, 0, 1, 0, 2, -1, -1, -1, -1, 1, 0, 0, 0, -1, -1, -1, 0, 0, 1, 0, 1, 0, 1, 1, -1, 0, 1, -2, 0, -1, 1, 0, 0, 1, 1, -1, 2, 0,

    others => 0);
end iwght_package;
