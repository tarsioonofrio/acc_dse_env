library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    713, 734, 729, 738, 729, 722, 746, 765, 740, 683, 626, 624, 643, 649, 629, 
    714, 737, 746, 753, 748, 784, 751, 707, 618, 531, 487, 453, 489, 592, 630, 
    614, 636, 746, 755, 754, 788, 653, 486, 414, 515, 560, 491, 432, 424, 580, 
    488, 450, 733, 760, 721, 638, 608, 467, 421, 553, 614, 506, 427, 325, 478, 
    646, 620, 745, 784, 853, 737, 679, 490, 383, 476, 667, 521, 426, 358, 344, 
    699, 738, 778, 692, 805, 820, 759, 572, 394, 545, 762, 539, 457, 429, 340, 
    715, 709, 687, 658, 598, 762, 850, 670, 507, 604, 726, 499, 430, 477, 461, 
    784, 743, 600, 634, 609, 819, 743, 619, 522, 624, 700, 508, 444, 511, 551, 
    836, 796, 617, 620, 614, 624, 608, 531, 533, 603, 585, 443, 359, 507, 642, 
    847, 812, 659, 573, 632, 496, 605, 672, 531, 573, 421, 291, 373, 619, 707, 
    740, 819, 670, 717, 853, 611, 657, 742, 554, 368, 281, 291, 352, 462, 470, 
    491, 723, 754, 941, 939, 518, 404, 393, 347, 301, 294, 301, 313, 336, 329, 
    288, 444, 730, 968, 590, 321, 306, 294, 286, 276, 287, 312, 342, 344, 355, 
    294, 277, 529, 761, 410, 327, 318, 294, 291, 298, 298, 315, 298, 311, 347, 
    306, 266, 312, 405, 292, 283, 318, 314, 325, 336, 309, 288, 364, 400, 277, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 40, 0, 0, 3, 86, 179, 112, 30, 0, 0, 
    9, 0, 0, 0, 0, 80, 61, 54, 79, 266, 368, 282, 199, 34, 0, 
    202, 13, 0, 0, 0, 38, 218, 211, 197, 274, 320, 231, 190, 80, 0, 
    445, 348, 46, 62, 427, 396, 385, 240, 177, 164, 366, 262, 193, 146, 17, 
    538, 491, 106, 45, 427, 427, 420, 287, 194, 264, 491, 281, 226, 222, 130, 
    532, 532, 115, 0, 197, 341, 532, 369, 287, 371, 462, 268, 207, 248, 212, 
    587, 584, 307, 122, 172, 517, 499, 333, 232, 294, 388, 272, 230, 257, 91, 
    679, 664, 457, 331, 233, 300, 256, 250, 233, 192, 232, 193, 122, 92, 9, 
    618, 646, 511, 417, 412, 225, 292, 444, 311, 243, 193, 106, 133, 54, 9, 
    569, 611, 515, 524, 689, 498, 564, 632, 447, 247, 250, 325, 394, 379, 349, 
    640, 639, 584, 715, 823, 518, 473, 470, 454, 446, 487, 522, 560, 579, 579, 
    617, 567, 570, 801, 599, 501, 501, 472, 469, 491, 545, 589, 614, 618, 658, 
    657, 562, 609, 735, 493, 524, 516, 491, 505, 548, 592, 616, 603, 660, 705, 
    668, 603, 549, 533, 453, 478, 518, 509, 534, 578, 581, 556, 637, 763, 619, 
    
    -- channel=2
    235, 248, 247, 250, 246, 242, 254, 263, 251, 218, 192, 199, 212, 214, 206, 
    243, 254, 253, 255, 251, 301, 248, 237, 179, 164, 143, 130, 145, 187, 207, 
    196, 199, 255, 259, 254, 256, 210, 134, 104, 152, 157, 134, 110, 104, 191, 
    143, 147, 246, 259, 254, 200, 196, 117, 105, 139, 192, 132, 112, 71, 135, 
    179, 205, 241, 233, 305, 221, 214, 143, 97, 124, 210, 143, 118, 88, 72, 
    175, 247, 257, 208, 269, 243, 267, 167, 116, 164, 232, 146, 119, 108, 80, 
    186, 237, 215, 222, 181, 256, 273, 208, 144, 183, 218, 141, 113, 132, 125, 
    226, 247, 156, 212, 158, 256, 219, 176, 153, 192, 215, 144, 110, 140, 166, 
    255, 249, 172, 199, 180, 166, 185, 167, 150, 184, 170, 110, 86, 155, 207, 
    274, 248, 203, 167, 177, 123, 179, 224, 141, 155, 98, 49, 93, 204, 230, 
    247, 255, 205, 235, 292, 166, 180, 214, 145, 85, 52, 49, 69, 111, 110, 
    98, 212, 218, 313, 277, 122, 84, 80, 61, 38, 36, 38, 46, 51, 49, 
    28, 84, 210, 325, 141, 52, 41, 41, 36, 31, 34, 45, 49, 47, 64, 
    29, 27, 106, 250, 80, 50, 51, 38, 34, 38, 34, 38, 32, 43, 42, 
    36, 23, 41, 83, 32, 29, 39, 44, 50, 60, 39, 31, 66, 78, 22, 
    
    
    others => 0);
end gold_package;
