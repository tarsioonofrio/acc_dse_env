library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -1951, -2797, -14671, 3654, 3015, 1817, 2111, -762, 5167, -2454, -1388, -1390, 2736, -2045, 2488, 1138, -4497, -2030, -1124, 3216, -3699, 2732, 4299, 1974, -6667, 3268, -4680, -5118, 482, 3638, 4848, 1600,

    -- weights
    -- filter=0 channel=0
    -14, 2, 5, 13, 12, 4, -12, -20, -5,
    -- filter=0 channel=1
    -18, -8, 0, 3, -11, 7, 12, -17, 2,
    -- filter=0 channel=2
    17, -7, 15, 16, 12, -13, 5, -19, 18,
    -- filter=0 channel=3
    9, 18, -18, 17, 19, 5, 11, -14, 3,
    -- filter=0 channel=4
    14, -19, -15, -7, -2, -10, -5, -8, -13,
    -- filter=0 channel=5
    -10, -17, 0, 2, 1, 4, 15, 7, 6,
    -- filter=0 channel=6
    -2, -4, 7, 12, 0, 6, 2, 17, -5,
    -- filter=0 channel=7
    -1, 3, 15, -21, -8, 13, 12, -18, 6,
    -- filter=0 channel=8
    -11, 14, 9, -15, 17, 0, -4, 16, 7,
    -- filter=0 channel=9
    -3, 7, 1, -11, -14, -13, 4, -11, -1,
    -- filter=0 channel=10
    -12, -3, 1, -4, -16, 20, -11, 8, -10,
    -- filter=0 channel=11
    6, 8, -5, 19, -8, 11, -19, 5, -10,
    -- filter=0 channel=12
    11, -13, 17, -20, 0, 7, -1, -3, 19,
    -- filter=0 channel=13
    -16, 16, 14, 10, 3, 0, -1, -14, 6,
    -- filter=0 channel=14
    9, 6, -16, 14, -20, 20, -14, 0, -10,
    -- filter=0 channel=15
    -13, 16, 13, -3, 16, -14, -8, -3, 9,
    -- filter=1 channel=0
    -9, 12, 0, 4, -20, -9, -18, -8, -17,
    -- filter=1 channel=1
    18, -11, 19, 6, 7, -5, 0, -19, 11,
    -- filter=1 channel=2
    -6, -5, 12, 0, 20, -16, -19, 13, 0,
    -- filter=1 channel=3
    1, 9, 18, -7, -16, 14, -15, 15, -13,
    -- filter=1 channel=4
    18, -17, -20, 4, 0, 19, -10, 12, 8,
    -- filter=1 channel=5
    13, -2, 8, 7, 13, -18, -6, 13, 12,
    -- filter=1 channel=6
    -1, -6, -7, 8, 2, -19, -16, 11, 0,
    -- filter=1 channel=7
    17, 10, -10, 7, 17, -12, 0, -14, 17,
    -- filter=1 channel=8
    -1, -14, -4, 10, 3, -19, -21, 7, -14,
    -- filter=1 channel=9
    -9, 7, -1, 20, -12, 14, 0, -15, 13,
    -- filter=1 channel=10
    -4, 13, 5, 10, 11, -12, -18, 0, -16,
    -- filter=1 channel=11
    0, 6, -13, 17, -19, -6, 17, 11, 16,
    -- filter=1 channel=12
    20, -9, -3, 9, 3, 1, -19, 0, 4,
    -- filter=1 channel=13
    -16, 3, -1, -19, -20, 10, 4, 0, -2,
    -- filter=1 channel=14
    -17, -6, -13, 18, -16, -11, 9, 11, -6,
    -- filter=1 channel=15
    -16, -9, 18, 10, -2, 1, -19, -2, -11,
    -- filter=2 channel=0
    -53, -50, -8, -39, -53, -51, -39, -26, -41,
    -- filter=2 channel=1
    -6, 0, 18, 23, 15, 27, 17, 34, 28,
    -- filter=2 channel=2
    -22, -20, -1, -29, -16, 1, -10, -18, -9,
    -- filter=2 channel=3
    -8, -38, -27, -47, -43, -43, -21, -33, -23,
    -- filter=2 channel=4
    20, 35, 12, 23, 20, 12, 24, 1, 23,
    -- filter=2 channel=5
    12, 6, 19, 25, 2, 18, 15, 13, 0,
    -- filter=2 channel=6
    -4, -7, -5, -13, -10, -27, 3, -28, -12,
    -- filter=2 channel=7
    3, 2, -36, 0, -11, -12, 14, -31, -32,
    -- filter=2 channel=8
    4, 6, 17, 6, 17, 13, -7, 8, -17,
    -- filter=2 channel=9
    11, 13, 32, 52, 53, 15, 53, 26, 38,
    -- filter=2 channel=10
    32, 23, -11, 35, 30, 23, 27, 24, 16,
    -- filter=2 channel=11
    -17, -29, -38, -35, 0, -14, -12, -25, -18,
    -- filter=2 channel=12
    14, 18, 0, 1, -16, 3, -17, -12, 6,
    -- filter=2 channel=13
    12, 54, 25, 66, 54, 40, 55, 67, 46,
    -- filter=2 channel=14
    -25, 14, 18, 4, 16, -15, -25, -1, 19,
    -- filter=2 channel=15
    2, -29, -5, -4, -28, -13, 0, -30, -24,
    -- filter=3 channel=0
    22, 16, 16, -7, -1, 10, -14, 18, 11,
    -- filter=3 channel=1
    13, -15, -4, -19, 10, 6, -9, -18, 14,
    -- filter=3 channel=2
    1, 17, -12, 21, 11, 15, 16, 16, 12,
    -- filter=3 channel=3
    -8, -18, 4, -6, 12, -5, 0, -10, -2,
    -- filter=3 channel=4
    15, 15, 25, 15, -18, -7, -22, 21, 11,
    -- filter=3 channel=5
    -15, -8, -9, 16, 8, -1, -3, 23, 10,
    -- filter=3 channel=6
    16, 12, -5, 3, 10, 4, 19, -9, -13,
    -- filter=3 channel=7
    2, 9, 7, -11, 7, 12, -2, 16, -2,
    -- filter=3 channel=8
    6, 2, 2, -10, 2, -9, 8, -7, 5,
    -- filter=3 channel=9
    18, 14, 17, -17, 0, -10, -1, -17, 23,
    -- filter=3 channel=10
    -24, 7, 3, -24, 16, 13, 20, -8, -14,
    -- filter=3 channel=11
    1, 1, -18, 20, -9, 20, -13, -18, 14,
    -- filter=3 channel=12
    -19, 8, -15, 12, 8, -12, -20, 7, 15,
    -- filter=3 channel=13
    -14, -4, 17, -14, -18, 8, 0, 0, 13,
    -- filter=3 channel=14
    12, -14, -12, 18, -12, -7, 4, 9, -15,
    -- filter=3 channel=15
    11, -13, 20, 13, 1, 16, 2, 1, -11,
    -- filter=4 channel=0
    8, -9, -13, -15, -3, 29, -5, 14, 9,
    -- filter=4 channel=1
    6, 33, 23, 0, 14, 27, 24, -5, 25,
    -- filter=4 channel=2
    -20, 8, -12, 5, -22, -17, -19, 6, 12,
    -- filter=4 channel=3
    10, 16, 24, 8, 15, 39, 0, 29, 28,
    -- filter=4 channel=4
    -9, -6, 0, -12, -30, -18, -32, -14, -19,
    -- filter=4 channel=5
    29, 23, 42, 26, 19, 14, -5, 20, 33,
    -- filter=4 channel=6
    -10, -4, 31, 7, 18, 15, -9, 15, 5,
    -- filter=4 channel=7
    2, -12, -19, 5, -27, -28, -24, 0, -25,
    -- filter=4 channel=8
    8, -10, 0, 6, 10, 1, 1, -4, 5,
    -- filter=4 channel=9
    -36, -13, -7, -32, -21, -32, -13, -37, -12,
    -- filter=4 channel=10
    30, 25, 24, -7, -9, 11, -20, 16, 17,
    -- filter=4 channel=11
    2, -6, 12, -22, 2, -6, 14, 14, 4,
    -- filter=4 channel=12
    8, 14, 3, 19, -10, 10, 2, -10, 1,
    -- filter=4 channel=13
    34, 28, 40, -10, -2, 5, 8, -8, 9,
    -- filter=4 channel=14
    34, 8, 45, 29, 13, 36, 10, 12, 13,
    -- filter=4 channel=15
    -21, 8, -9, -19, -1, -6, -32, -32, 2,
    -- filter=5 channel=0
    18, 6, -17, -7, -8, 0, 14, -15, -8,
    -- filter=5 channel=1
    6, -17, 18, -2, 21, -13, -24, 13, -1,
    -- filter=5 channel=2
    -8, -8, -17, 28, 0, -2, 14, 4, -7,
    -- filter=5 channel=3
    6, -5, -15, -11, 0, 8, -8, 0, -18,
    -- filter=5 channel=4
    -2, 1, 0, -9, -1, 1, -14, 0, -10,
    -- filter=5 channel=5
    12, 15, 1, -15, 15, 25, -24, 21, 6,
    -- filter=5 channel=6
    16, -7, -4, -17, -19, 4, 9, 2, 11,
    -- filter=5 channel=7
    0, -9, 2, -4, -3, -1, 24, 7, 15,
    -- filter=5 channel=8
    17, -7, -10, -16, 14, 1, 15, 2, -5,
    -- filter=5 channel=9
    17, 0, 8, 20, 0, 10, 0, -12, 18,
    -- filter=5 channel=10
    -15, 1, 12, -10, 11, 26, 19, 7, -15,
    -- filter=5 channel=11
    9, 2, 6, 5, 4, -10, 8, -18, -12,
    -- filter=5 channel=12
    -9, 7, -19, 17, 0, -6, -17, -7, 14,
    -- filter=5 channel=13
    -24, 22, 27, -32, -10, 26, -28, 23, -1,
    -- filter=5 channel=14
    -13, -1, 2, -5, -11, -14, -4, -18, -6,
    -- filter=5 channel=15
    24, 0, -13, 23, -6, -2, 12, 9, -19,
    -- filter=6 channel=0
    -2, 23, -9, 10, 5, -13, 13, 23, -13,
    -- filter=6 channel=1
    20, 12, -11, 14, 8, -15, -3, 20, -25,
    -- filter=6 channel=2
    -4, 8, 23, 1, -13, 25, -10, -17, 1,
    -- filter=6 channel=3
    -2, -7, 0, -17, -8, -17, -10, -17, -19,
    -- filter=6 channel=4
    16, 20, 11, 13, 27, -20, 22, 20, -19,
    -- filter=6 channel=5
    -3, -14, -27, -14, -21, -5, -5, 15, -16,
    -- filter=6 channel=6
    -6, -4, 10, -11, 4, 14, 5, -10, -2,
    -- filter=6 channel=7
    -8, 0, -4, -10, 17, 9, 4, 17, 13,
    -- filter=6 channel=8
    -13, -12, -15, 16, -6, 0, 0, 14, 0,
    -- filter=6 channel=9
    26, 11, 24, 13, 10, -15, 8, 1, -15,
    -- filter=6 channel=10
    5, -12, 5, 28, -17, 4, 29, -7, -9,
    -- filter=6 channel=11
    0, 11, -15, -8, 22, -3, 10, -8, -17,
    -- filter=6 channel=12
    -8, 17, -4, 19, -12, -13, 6, -12, 21,
    -- filter=6 channel=13
    23, -7, -5, 24, 19, -9, 39, 10, -35,
    -- filter=6 channel=14
    -5, -8, -26, 11, 15, -4, -7, 18, 13,
    -- filter=6 channel=15
    22, 14, 10, 6, 8, -3, 20, -11, 0,
    -- filter=7 channel=0
    -13, -16, -14, -31, -28, -27, -25, -5, 14,
    -- filter=7 channel=1
    -6, 20, -3, 14, 28, 15, -16, 15, 18,
    -- filter=7 channel=2
    6, -9, -23, -1, -14, 15, 5, 0, -20,
    -- filter=7 channel=3
    -11, -29, -9, -9, -27, -11, -10, -2, -1,
    -- filter=7 channel=4
    5, 28, 30, 7, 30, 13, 21, 17, 15,
    -- filter=7 channel=5
    -9, -4, -11, -7, 0, -19, 10, -1, -12,
    -- filter=7 channel=6
    10, 0, -10, -17, 13, 8, 3, 6, 15,
    -- filter=7 channel=7
    29, 14, -5, 0, 13, 10, -10, 11, 17,
    -- filter=7 channel=8
    13, -2, 2, 7, 7, 17, -11, 17, 15,
    -- filter=7 channel=9
    46, 36, 41, 25, 50, 42, 44, 45, 37,
    -- filter=7 channel=10
    -2, 20, 9, 15, -6, 4, 17, 31, -7,
    -- filter=7 channel=11
    -24, 12, -12, -3, 3, 8, -1, 1, -10,
    -- filter=7 channel=12
    -1, 10, 7, -11, 20, 1, 11, -14, -2,
    -- filter=7 channel=13
    28, 10, 29, 32, 16, 23, 33, 44, -5,
    -- filter=7 channel=14
    -18, -6, -3, 2, -21, -5, -25, -1, -14,
    -- filter=7 channel=15
    15, 9, 0, 0, 9, 6, 14, 14, -15,
    -- filter=8 channel=0
    -4, -20, 9, 0, 11, 0, -16, -19, 11,
    -- filter=8 channel=1
    24, 20, 11, 20, 25, 3, 29, 10, 19,
    -- filter=8 channel=2
    -5, 3, 5, 0, -11, -19, -20, -15, -12,
    -- filter=8 channel=3
    12, -2, 29, -1, 21, 15, 3, 21, 22,
    -- filter=8 channel=4
    7, -3, -18, -3, -7, -26, -24, 8, 16,
    -- filter=8 channel=5
    21, -6, 20, 6, 28, 18, 14, 4, 17,
    -- filter=8 channel=6
    19, 9, -12, 10, 0, 16, -2, 23, -5,
    -- filter=8 channel=7
    -16, -1, 2, -26, -2, -6, -15, -18, 3,
    -- filter=8 channel=8
    -13, 5, 17, 11, 20, -1, 17, 15, 7,
    -- filter=8 channel=9
    -18, -23, -31, -1, -24, -26, -7, -14, 2,
    -- filter=8 channel=10
    10, 12, 29, 9, -15, 24, -5, 12, 14,
    -- filter=8 channel=11
    -3, 17, -4, -17, 6, -18, -3, 18, 20,
    -- filter=8 channel=12
    -2, 2, -4, -5, 0, -21, 4, -5, -10,
    -- filter=8 channel=13
    17, 14, 16, -11, 6, -3, 21, 6, 2,
    -- filter=8 channel=14
    -3, 21, 33, 13, 2, -4, -1, 28, 13,
    -- filter=8 channel=15
    -28, -19, 2, -29, 0, 4, -20, 9, -13,
    -- filter=9 channel=0
    -28, -30, -13, -21, -25, -31, -22, -35, -37,
    -- filter=9 channel=1
    -10, 3, 8, -5, -1, 11, -10, 25, -7,
    -- filter=9 channel=2
    17, -13, 12, -1, -1, -28, 3, 11, -5,
    -- filter=9 channel=3
    -1, -5, -24, -2, -8, -21, -19, 6, -28,
    -- filter=9 channel=4
    7, 4, -3, -12, 6, 17, -12, 26, 25,
    -- filter=9 channel=5
    0, 2, 6, 2, 3, -8, 22, 9, 0,
    -- filter=9 channel=6
    -14, -19, 6, -3, -14, -10, -11, 0, 3,
    -- filter=9 channel=7
    18, -11, 0, 22, -17, -4, -9, -19, -19,
    -- filter=9 channel=8
    4, -20, -10, 15, -12, 7, 11, -18, -14,
    -- filter=9 channel=9
    19, 29, 0, 15, 30, 4, 12, 25, 13,
    -- filter=9 channel=10
    11, 29, 10, 4, 18, 1, 20, 17, 11,
    -- filter=9 channel=11
    -17, 11, 4, 1, 5, -3, 9, 11, 0,
    -- filter=9 channel=12
    -4, 5, 1, -14, 6, -18, 18, 16, -9,
    -- filter=9 channel=13
    27, 37, 26, 41, 14, 22, 14, 21, 11,
    -- filter=9 channel=14
    -23, -3, -9, -8, -16, -20, -4, 16, -18,
    -- filter=9 channel=15
    -9, 12, 6, -14, -7, 8, 11, 10, -20,
    -- filter=10 channel=0
    1, -22, 11, 0, -17, 12, 13, 3, -12,
    -- filter=10 channel=1
    -8, -15, 7, 17, -5, 8, -3, -15, -21,
    -- filter=10 channel=2
    0, 11, 14, -2, -16, 5, 17, 6, 11,
    -- filter=10 channel=3
    -30, -1, -2, 5, -29, -23, -9, -23, -10,
    -- filter=10 channel=4
    30, 17, 0, 24, 12, 4, -6, -9, -13,
    -- filter=10 channel=5
    8, 15, -20, 8, 12, -6, -13, 7, 12,
    -- filter=10 channel=6
    12, 6, 0, -3, -12, 19, -21, -15, 12,
    -- filter=10 channel=7
    0, 5, -18, 2, -18, -17, 20, 16, -14,
    -- filter=10 channel=8
    -6, -16, -7, 13, 2, -21, -15, -18, -13,
    -- filter=10 channel=9
    27, 36, 4, 30, 4, -8, 5, 14, 23,
    -- filter=10 channel=10
    30, 0, 4, 25, 0, 6, 26, -9, -5,
    -- filter=10 channel=11
    18, -21, 0, 18, -17, 12, 16, -1, 13,
    -- filter=10 channel=12
    0, -10, -18, 3, -20, -17, 17, 4, -18,
    -- filter=10 channel=13
    29, 26, 0, 35, -4, 0, 13, -6, -21,
    -- filter=10 channel=14
    -20, -15, -24, -16, -24, -1, -3, -4, -24,
    -- filter=10 channel=15
    23, 4, 11, 18, -7, 20, -11, -5, 5,
    -- filter=11 channel=0
    -2, -20, -4, 18, 3, -6, -7, 1, -18,
    -- filter=11 channel=1
    19, -12, 7, -4, -4, -14, -14, 5, 13,
    -- filter=11 channel=2
    8, 14, 15, 0, 14, 1, 16, 11, 9,
    -- filter=11 channel=3
    -7, 12, 2, 13, 9, 13, -12, -8, -15,
    -- filter=11 channel=4
    -17, 6, -16, 10, 1, 3, -12, 6, -13,
    -- filter=11 channel=5
    -18, 1, -9, 14, 4, 17, 5, 14, 0,
    -- filter=11 channel=6
    12, -16, 1, -12, -7, 20, -8, -20, -12,
    -- filter=11 channel=7
    5, 0, -17, -19, 6, -5, 3, -6, 20,
    -- filter=11 channel=8
    -18, -20, 7, -4, 9, 4, 9, 10, 1,
    -- filter=11 channel=9
    11, -4, -13, -20, 14, 6, 10, 16, 14,
    -- filter=11 channel=10
    -1, -18, -5, 2, 17, 18, 9, -5, 18,
    -- filter=11 channel=11
    -8, 1, 13, 15, 11, 14, -16, 19, -10,
    -- filter=11 channel=12
    -6, -4, -20, 1, -4, 7, 3, -14, 15,
    -- filter=11 channel=13
    2, -13, -12, 17, 15, 8, -13, -20, -16,
    -- filter=11 channel=14
    -2, -16, -4, -3, 0, 14, 8, 15, 20,
    -- filter=11 channel=15
    -12, 14, -7, -11, -2, 8, 7, -8, -3,
    -- filter=12 channel=0
    -10, 11, 7, -20, 20, 7, -9, 21, -2,
    -- filter=12 channel=1
    25, 11, 14, 11, -1, 5, 22, 31, 24,
    -- filter=12 channel=2
    -8, -2, -20, 5, -18, 13, 0, -2, -20,
    -- filter=12 channel=3
    1, 3, 22, 26, 26, 0, 21, 17, -8,
    -- filter=12 channel=4
    5, 10, -5, 1, -8, -18, 15, -4, 8,
    -- filter=12 channel=5
    -4, 10, -6, -2, 3, 10, 26, 23, 2,
    -- filter=12 channel=6
    -18, 6, 8, -15, 12, 12, 21, -9, -15,
    -- filter=12 channel=7
    0, -28, -26, 8, -26, 1, -25, -18, 2,
    -- filter=12 channel=8
    18, -17, 16, 11, 12, 2, -15, 4, 3,
    -- filter=12 channel=9
    1, -27, -3, -12, -17, -29, -27, 4, -12,
    -- filter=12 channel=10
    -14, 23, -12, 20, 18, 12, 16, 14, -1,
    -- filter=12 channel=11
    2, -12, 0, 12, -15, -8, 8, -10, -11,
    -- filter=12 channel=12
    12, 13, 0, -20, -10, 2, 14, -18, -9,
    -- filter=12 channel=13
    -11, 17, 5, 18, 22, 11, 1, 8, 0,
    -- filter=12 channel=14
    26, 26, 28, 11, 13, 0, 0, 25, 24,
    -- filter=12 channel=15
    13, -9, 0, -24, -26, -5, -6, 11, 9,
    -- filter=13 channel=0
    7, 7, -6, -20, -4, -18, -24, -3, 13,
    -- filter=13 channel=1
    3, 4, -11, -13, -12, 0, 7, 1, 12,
    -- filter=13 channel=2
    -9, 9, -16, -4, -11, 6, -13, 14, 6,
    -- filter=13 channel=3
    -20, -19, -13, -14, 4, 6, 0, -18, -9,
    -- filter=13 channel=4
    -12, 23, 20, 17, -1, -9, 1, 28, 0,
    -- filter=13 channel=5
    14, 7, -13, 2, 16, -24, -8, 16, 2,
    -- filter=13 channel=6
    0, 0, 1, -9, -13, 6, -23, 8, 9,
    -- filter=13 channel=7
    6, -4, -16, 23, -2, 4, 2, -12, -6,
    -- filter=13 channel=8
    -19, -15, -18, 8, -1, 17, 0, 14, 4,
    -- filter=13 channel=9
    29, 14, 10, 36, 22, 24, 20, 35, 20,
    -- filter=13 channel=10
    11, -17, 4, -6, 15, -8, 6, 13, -9,
    -- filter=13 channel=11
    5, 3, 15, 8, -21, -6, -19, -20, 15,
    -- filter=13 channel=12
    19, 5, 6, -15, 7, -16, -18, 16, -7,
    -- filter=13 channel=13
    22, -7, 0, 22, 20, 27, 29, 24, 29,
    -- filter=13 channel=14
    -1, -3, -22, -16, -5, -10, -5, 10, -11,
    -- filter=13 channel=15
    -7, -11, -12, -10, -3, 21, 3, 2, 16,
    -- filter=14 channel=0
    5, 1, 26, 11, 8, 2, 10, 13, 28,
    -- filter=14 channel=1
    2, 25, 1, 9, -2, 20, 10, 3, 34,
    -- filter=14 channel=2
    11, -12, 16, 4, -12, 8, 11, 11, -9,
    -- filter=14 channel=3
    35, 18, 24, 30, 24, -2, 12, 28, 26,
    -- filter=14 channel=4
    -29, -29, 17, -20, 0, -3, -11, -25, 22,
    -- filter=14 channel=5
    5, 27, 3, 0, 23, 30, 22, 38, 4,
    -- filter=14 channel=6
    22, 9, 4, -9, 12, 26, 15, 12, 32,
    -- filter=14 channel=7
    -22, -25, 1, -4, -12, 4, 0, -26, -17,
    -- filter=14 channel=8
    -3, -5, -14, 7, 5, -21, -18, 20, 15,
    -- filter=14 channel=9
    -22, -38, -24, -32, -13, -27, -25, -24, -18,
    -- filter=14 channel=10
    8, 5, 21, 9, 24, 9, 7, 5, -1,
    -- filter=14 channel=11
    -18, -9, 16, -11, -20, -17, 0, -11, -6,
    -- filter=14 channel=12
    4, 18, 11, 5, -7, -15, -8, 17, 2,
    -- filter=14 channel=13
    14, -4, 35, -10, 14, 38, 19, 24, 6,
    -- filter=14 channel=14
    8, 0, 35, 29, 31, 1, 17, 35, 22,
    -- filter=14 channel=15
    8, -26, -12, -13, -23, 0, 1, -19, -11,
    -- filter=15 channel=0
    -4, -10, 20, -19, 18, -4, 4, 2, 17,
    -- filter=15 channel=1
    -15, -11, 13, -3, 0, 9, 18, 0, -15,
    -- filter=15 channel=2
    -20, 14, -13, 5, -21, -20, -6, 16, -18,
    -- filter=15 channel=3
    12, 11, 0, -5, -14, -18, -20, -12, 2,
    -- filter=15 channel=4
    10, -3, 9, 3, 10, 0, -15, 1, 20,
    -- filter=15 channel=5
    -13, 9, 19, -7, 0, -10, -13, 17, 1,
    -- filter=15 channel=6
    3, -9, 3, 17, -16, -11, -13, -20, -19,
    -- filter=15 channel=7
    7, 11, -16, 2, -14, 7, -9, 11, 7,
    -- filter=15 channel=8
    14, 18, 16, 5, -14, -12, 9, 5, 16,
    -- filter=15 channel=9
    6, -2, -3, -7, 9, -3, -15, 13, -10,
    -- filter=15 channel=10
    -6, 0, -2, -19, 12, -4, -14, -12, -17,
    -- filter=15 channel=11
    -10, 11, -21, -3, -19, 12, 20, 0, -9,
    -- filter=15 channel=12
    -18, -13, -3, -21, -20, 6, 1, 12, 6,
    -- filter=15 channel=13
    2, -3, 2, 22, -14, 15, -20, -13, -7,
    -- filter=15 channel=14
    -6, 0, -12, -14, 5, -9, 3, -1, 14,
    -- filter=15 channel=15
    19, -9, 2, 13, 15, 18, 5, -18, -7,
    -- filter=16 channel=0
    -3, -6, 13, -14, -20, -15, 16, 18, -3,
    -- filter=16 channel=1
    -7, -10, -4, -2, 8, -2, -13, 10, 26,
    -- filter=16 channel=2
    13, 4, 15, 19, 22, -9, 4, 9, 1,
    -- filter=16 channel=3
    -8, 8, 15, -8, -7, 19, 14, -4, 13,
    -- filter=16 channel=4
    -11, -18, 26, -13, -2, -3, 13, 24, 31,
    -- filter=16 channel=5
    -17, 14, 25, -7, 8, 20, -15, 20, 13,
    -- filter=16 channel=6
    14, 12, 7, 10, -12, 4, -11, 18, 7,
    -- filter=16 channel=7
    0, 15, 10, -13, 2, 8, -8, 14, -1,
    -- filter=16 channel=8
    -1, 8, -19, -7, 9, -3, -2, 14, -14,
    -- filter=16 channel=9
    -16, 1, -1, 6, -19, 21, -11, 15, 11,
    -- filter=16 channel=10
    12, 24, 8, -4, 0, 24, 21, 19, 20,
    -- filter=16 channel=11
    7, -21, 1, -1, -20, -3, -16, -5, 17,
    -- filter=16 channel=12
    13, 18, -19, 19, -19, -17, -1, -21, -8,
    -- filter=16 channel=13
    -25, 18, 13, -13, 27, 3, -7, 22, 12,
    -- filter=16 channel=14
    8, -10, 0, -10, -13, 4, -8, 4, -5,
    -- filter=16 channel=15
    -2, 19, 10, -5, -16, -11, -5, 1, 12,
    -- filter=17 channel=0
    -5, 8, 0, 17, 5, -3, 16, 16, -6,
    -- filter=17 channel=1
    22, 3, -18, 17, 36, -15, 15, 19, -5,
    -- filter=17 channel=2
    0, -11, 16, 32, 13, 22, 21, 12, 6,
    -- filter=17 channel=3
    3, -11, -18, -23, -3, -10, -11, -6, -15,
    -- filter=17 channel=4
    31, 20, -10, 8, 17, -5, 34, 47, 6,
    -- filter=17 channel=5
    15, -11, -37, 6, 19, -16, 25, -13, -10,
    -- filter=17 channel=6
    15, -12, 15, 25, 19, -9, 19, 27, 17,
    -- filter=17 channel=7
    -3, 11, -9, 18, 6, 7, 31, -12, 19,
    -- filter=17 channel=8
    16, 2, 18, 14, -18, 10, 10, -4, 20,
    -- filter=17 channel=9
    31, 28, 9, 15, 31, -7, 28, 18, 3,
    -- filter=17 channel=10
    36, 2, -27, 24, -3, -3, 17, 7, -22,
    -- filter=17 channel=11
    16, 15, 1, 0, 7, 4, 3, -2, 12,
    -- filter=17 channel=12
    18, -5, -14, 19, -14, -1, 2, 8, 3,
    -- filter=17 channel=13
    33, 24, -48, 41, 29, -26, 52, 39, -4,
    -- filter=17 channel=14
    -18, 1, 4, 11, 10, 1, -9, 9, -21,
    -- filter=17 channel=15
    19, 19, 32, -14, -5, 27, 5, 8, 30,
    -- filter=18 channel=0
    13, 0, 9, 1, 13, -4, 7, 3, 10,
    -- filter=18 channel=1
    3, -15, 9, 14, 19, -9, -15, 0, -2,
    -- filter=18 channel=2
    14, 14, -16, -7, 11, -8, -11, 9, -4,
    -- filter=18 channel=3
    -8, 8, -1, -14, -1, 6, -6, 11, 7,
    -- filter=18 channel=4
    -15, 16, -18, -5, 4, -16, -4, -16, 0,
    -- filter=18 channel=5
    -15, 3, -12, -16, -14, 5, 17, -4, 13,
    -- filter=18 channel=6
    21, 14, 8, 18, 13, -17, 9, 22, 23,
    -- filter=18 channel=7
    -3, 9, -7, -5, -4, -2, 22, -6, -6,
    -- filter=18 channel=8
    15, 0, -2, 11, 0, -16, -8, -4, -2,
    -- filter=18 channel=9
    -11, 16, 21, 16, 2, -16, -19, 9, -15,
    -- filter=18 channel=10
    11, -3, 9, 24, -3, 11, 23, -18, -10,
    -- filter=18 channel=11
    11, -17, 14, 7, -4, 13, 18, 11, -7,
    -- filter=18 channel=12
    -19, 20, 16, -19, 11, -2, -4, -16, -2,
    -- filter=18 channel=13
    -11, 12, -17, -17, 20, 10, -5, 22, -13,
    -- filter=18 channel=14
    0, -14, 8, -7, 8, 20, 5, 1, 17,
    -- filter=18 channel=15
    -13, 0, 0, -13, -6, 16, -18, 19, 23,
    -- filter=19 channel=0
    12, 18, -5, 29, 15, 27, 36, 6, 25,
    -- filter=19 channel=1
    3, -15, -6, -38, -21, 24, -28, 8, 6,
    -- filter=19 channel=2
    17, 17, 4, 0, 19, 36, 25, 32, 35,
    -- filter=19 channel=3
    -9, 16, 15, 16, 4, -6, -16, 18, -11,
    -- filter=19 channel=4
    7, 18, 7, -3, -17, -1, -3, -16, 38,
    -- filter=19 channel=5
    5, 6, -11, -2, -12, 12, -27, 13, 38,
    -- filter=19 channel=6
    6, 4, 18, 5, -9, 2, 16, 19, -10,
    -- filter=19 channel=7
    25, 37, 0, 8, 27, -7, 18, -1, 31,
    -- filter=19 channel=8
    9, -8, -10, -12, 11, 11, 0, 12, -10,
    -- filter=19 channel=9
    -27, -17, 9, -13, -1, 1, -34, -8, 0,
    -- filter=19 channel=10
    10, 19, 4, 0, 10, 26, -12, 32, 36,
    -- filter=19 channel=11
    27, -7, 6, 24, -12, -6, 30, -13, 14,
    -- filter=19 channel=12
    16, 10, 13, 9, 10, -18, -17, 4, -8,
    -- filter=19 channel=13
    -26, 7, 30, -60, -19, 43, -59, -21, 60,
    -- filter=19 channel=14
    -4, -17, 14, -20, 6, 29, 11, 21, 25,
    -- filter=19 channel=15
    -1, 32, 16, 22, 7, 11, 10, 2, 26,
    -- filter=20 channel=0
    1, 16, -12, -17, 7, -17, 16, -4, -6,
    -- filter=20 channel=1
    -17, -18, -2, -26, 6, -9, -16, -2, -11,
    -- filter=20 channel=2
    -1, -10, 11, 12, -12, -8, 30, -5, 10,
    -- filter=20 channel=3
    0, -12, 1, 12, 3, -7, -7, 0, 12,
    -- filter=20 channel=4
    -6, -1, -1, 17, 33, 29, -16, 33, 24,
    -- filter=20 channel=5
    -2, 4, -22, 16, 4, -14, 13, -9, 17,
    -- filter=20 channel=6
    1, 0, 19, 10, 14, 2, 16, -15, -2,
    -- filter=20 channel=7
    16, 2, 3, 0, -6, 22, 21, 2, -18,
    -- filter=20 channel=8
    8, -19, -16, 5, 4, 14, 19, -16, -4,
    -- filter=20 channel=9
    15, 10, 15, 14, 23, 32, 27, 32, 9,
    -- filter=20 channel=10
    20, 22, 6, 8, 24, 0, 22, 13, 2,
    -- filter=20 channel=11
    -6, 6, 11, -16, 14, -9, 10, -4, 7,
    -- filter=20 channel=12
    19, -14, 5, -6, -16, 0, -1, -5, -15,
    -- filter=20 channel=13
    12, -6, 7, 6, 10, 28, -9, 28, -1,
    -- filter=20 channel=14
    -23, -16, 14, -26, 6, 0, -14, -14, 4,
    -- filter=20 channel=15
    2, 12, 14, -8, 17, 2, -16, -13, 8,
    -- filter=21 channel=0
    -16, 3, -3, -29, -4, 7, -30, -23, -7,
    -- filter=21 channel=1
    -4, 9, -10, 8, -6, 8, -9, -5, 21,
    -- filter=21 channel=2
    -5, 5, 2, 23, -8, -19, 3, -3, -5,
    -- filter=21 channel=3
    -12, -22, -30, -17, -28, -16, 4, -9, -27,
    -- filter=21 channel=4
    0, 13, -5, -6, 19, 25, 31, 24, 2,
    -- filter=21 channel=5
    -24, -28, -8, -2, -21, -20, 10, -12, -7,
    -- filter=21 channel=6
    -6, -6, -9, -5, 5, -5, 14, -21, 13,
    -- filter=21 channel=7
    -8, -8, -8, 9, -5, -4, 3, 5, -1,
    -- filter=21 channel=8
    -9, 10, -9, 14, -16, 20, 17, -19, -6,
    -- filter=21 channel=9
    34, 40, 40, 12, 28, 37, 19, 32, 15,
    -- filter=21 channel=10
    9, 20, 9, 4, 19, 14, 2, -4, -21,
    -- filter=21 channel=11
    -20, -10, 4, -7, -14, 16, 0, 3, 11,
    -- filter=21 channel=12
    -3, 9, -15, -12, -4, -20, 20, -8, -15,
    -- filter=21 channel=13
    18, 3, -2, 23, 33, 17, 7, 41, 24,
    -- filter=21 channel=14
    -22, -1, -9, -32, -31, -28, -34, -14, -21,
    -- filter=21 channel=15
    -5, -10, 7, 2, -9, 22, -2, 11, -3,
    -- filter=22 channel=0
    -8, 1, -19, -12, 7, 4, 2, -10, 10,
    -- filter=22 channel=1
    6, 7, -2, -12, 24, -6, 13, -12, -12,
    -- filter=22 channel=2
    -14, -18, -8, -13, 17, -11, 14, -8, -19,
    -- filter=22 channel=3
    0, 2, -10, 26, 17, 19, -13, 13, 5,
    -- filter=22 channel=4
    -16, 16, -18, -15, 2, -2, 8, -10, 6,
    -- filter=22 channel=5
    16, -4, -10, -2, -8, -6, -3, 4, -16,
    -- filter=22 channel=6
    1, -15, 0, 11, 8, 10, -3, 15, 6,
    -- filter=22 channel=7
    -15, -2, -1, -1, 5, 0, 6, 9, 19,
    -- filter=22 channel=8
    -12, -15, 20, -18, 16, 6, 3, -16, -4,
    -- filter=22 channel=9
    -18, -23, -10, -1, 9, -8, 7, -25, -19,
    -- filter=22 channel=10
    0, 26, 17, 8, 4, -8, 2, -16, -20,
    -- filter=22 channel=11
    -18, 20, -17, 18, -15, 15, 21, 0, -15,
    -- filter=22 channel=12
    15, 0, -15, -20, 11, -18, -6, -12, -17,
    -- filter=22 channel=13
    26, 10, -9, -5, 20, 3, 24, -6, -3,
    -- filter=22 channel=14
    -7, 28, 14, 16, 12, -2, 20, -2, -3,
    -- filter=22 channel=15
    -12, -3, 0, 9, -14, 8, -16, 5, -19,
    -- filter=23 channel=0
    -33, -15, -12, -28, -39, -8, -1, -6, -13,
    -- filter=23 channel=1
    49, 27, 36, 20, 7, 35, -11, 9, 22,
    -- filter=23 channel=2
    -45, -37, -11, -47, -22, -28, -26, -24, -27,
    -- filter=23 channel=3
    -2, 17, 26, 30, 24, 6, 44, 34, 32,
    -- filter=23 channel=4
    0, -31, -14, -31, -10, -32, -8, -35, -35,
    -- filter=23 channel=5
    40, 46, 52, 11, 26, 20, 8, 35, 22,
    -- filter=23 channel=6
    0, 8, 14, -15, -8, 13, -16, -17, 19,
    -- filter=23 channel=7
    -20, -25, -43, -28, -45, -45, -8, -19, -12,
    -- filter=23 channel=8
    8, 16, -5, -7, 2, -2, -17, 18, -14,
    -- filter=23 channel=9
    -37, -48, -18, -13, -36, -46, -36, -47, -19,
    -- filter=23 channel=10
    20, 17, 43, 6, 21, 42, 19, -4, 16,
    -- filter=23 channel=11
    -2, -14, -25, -14, -7, 2, 10, 11, -10,
    -- filter=23 channel=12
    -3, -15, -10, -11, 7, -11, 17, -19, -16,
    -- filter=23 channel=13
    46, 39, 42, 6, 39, 34, -11, -8, 28,
    -- filter=23 channel=14
    40, 12, 45, 43, 31, 23, 3, 11, 44,
    -- filter=23 channel=15
    -14, -14, -9, -12, -12, -37, -40, -16, -35,
    -- filter=24 channel=0
    -19, -7, -27, -1, -15, -17, -34, -33, 6,
    -- filter=24 channel=1
    -12, 4, 13, 12, 28, 15, 22, 29, 29,
    -- filter=24 channel=2
    6, 5, -12, 18, 5, -2, 19, -19, -12,
    -- filter=24 channel=3
    -3, -29, -35, -18, -2, -34, -16, -20, -16,
    -- filter=24 channel=4
    17, 13, 1, 9, 26, 17, 28, 43, 4,
    -- filter=24 channel=5
    -23, -11, -31, -5, -21, 7, -18, -7, -23,
    -- filter=24 channel=6
    -10, 6, 6, -9, -13, -11, -21, -25, 0,
    -- filter=24 channel=7
    -1, -14, -22, 26, 9, -15, -4, -15, 13,
    -- filter=24 channel=8
    11, -7, 6, 18, 17, -4, 0, 10, 3,
    -- filter=24 channel=9
    17, 41, 27, 47, 18, 20, 40, 11, 39,
    -- filter=24 channel=10
    10, 14, -13, 25, 12, 10, -5, 21, 19,
    -- filter=24 channel=11
    -8, 11, -15, 6, -7, -6, 8, -20, -24,
    -- filter=24 channel=12
    -2, 4, 15, 13, 12, -13, 14, -11, 10,
    -- filter=24 channel=13
    29, 27, 11, 46, 41, 20, 15, 52, 18,
    -- filter=24 channel=14
    -9, -27, -19, -2, 0, -20, -27, 10, 15,
    -- filter=24 channel=15
    12, 1, 5, 12, -6, 23, 3, -3, 5,
    -- filter=25 channel=0
    20, -2, 10, 12, -4, -11, 13, 18, -19,
    -- filter=25 channel=1
    11, 16, 12, 0, 9, 7, 11, 11, -12,
    -- filter=25 channel=2
    -19, 2, -5, 6, -19, -3, 11, -19, 14,
    -- filter=25 channel=3
    -15, -11, 3, 5, 10, 19, -11, -13, 11,
    -- filter=25 channel=4
    11, 14, 13, -8, 11, -16, -19, -3, -7,
    -- filter=25 channel=5
    17, 12, -13, -20, -15, 16, -3, -16, 7,
    -- filter=25 channel=6
    8, -10, -8, -13, 11, -11, 19, 17, 20,
    -- filter=25 channel=7
    5, 13, 7, -3, -14, -18, 4, 0, -9,
    -- filter=25 channel=8
    20, -12, -18, 1, 3, -17, -20, -16, -17,
    -- filter=25 channel=9
    2, -5, -20, -20, 5, -2, -10, 19, -11,
    -- filter=25 channel=10
    -4, -20, -15, 9, -2, 18, -10, -12, -3,
    -- filter=25 channel=11
    -6, -17, -1, 0, 3, 3, 13, 3, -5,
    -- filter=25 channel=12
    2, 13, -17, 19, 9, 9, -20, 19, -15,
    -- filter=25 channel=13
    -8, 2, -4, -13, -10, -1, 5, -4, -21,
    -- filter=25 channel=14
    -9, -9, -17, -4, -7, 9, -6, 15, -11,
    -- filter=25 channel=15
    18, 14, 6, -4, -12, -4, -15, -4, 10,
    -- filter=26 channel=0
    -8, -21, 19, 7, 18, 6, 9, 13, -14,
    -- filter=26 channel=1
    -12, 16, 10, 7, 21, -27, 3, 2, -10,
    -- filter=26 channel=2
    10, 1, -2, 27, 10, -7, 17, 12, 12,
    -- filter=26 channel=3
    -37, 3, -30, -28, -21, -3, 4, -12, 5,
    -- filter=26 channel=4
    38, 37, 33, 43, 18, 8, 34, 33, 27,
    -- filter=26 channel=5
    8, -19, 0, -5, -9, -10, 10, -24, -6,
    -- filter=26 channel=6
    -1, -17, 9, 5, 20, -2, 12, -5, -2,
    -- filter=26 channel=7
    -6, 7, -2, 12, 24, 22, 2, 4, -10,
    -- filter=26 channel=8
    11, 12, 2, 8, -16, 2, -11, 16, 15,
    -- filter=26 channel=9
    31, 39, 18, 41, 22, -5, 39, 33, -3,
    -- filter=26 channel=10
    -5, -2, 15, 7, 11, -6, 0, 18, -24,
    -- filter=26 channel=11
    15, 1, 14, 8, -5, -14, 19, -14, 13,
    -- filter=26 channel=12
    -10, -7, -12, -3, -11, 16, 14, -12, 3,
    -- filter=26 channel=13
    18, 11, 23, 37, 28, -13, 44, 6, -4,
    -- filter=26 channel=14
    -19, -8, -26, -29, 5, -18, -8, -7, -18,
    -- filter=26 channel=15
    -1, 7, -2, 0, 31, 26, 15, -1, 12,
    -- filter=27 channel=0
    1, 0, -8, 21, -2, 15, 7, 5, 20,
    -- filter=27 channel=1
    -2, 2, 18, 9, 12, 21, -15, 0, 14,
    -- filter=27 channel=2
    12, -17, -5, 12, 19, -5, 19, 10, 21,
    -- filter=27 channel=3
    -3, -7, -8, -5, 8, -18, 19, 18, -5,
    -- filter=27 channel=4
    2, 0, -9, 15, -11, 20, -3, -7, -4,
    -- filter=27 channel=5
    8, -9, -4, 0, 10, 13, 20, -10, 3,
    -- filter=27 channel=6
    -16, 0, -5, -11, 14, -3, 13, -15, -18,
    -- filter=27 channel=7
    -3, -13, -16, -4, 18, -15, -10, -3, 16,
    -- filter=27 channel=8
    10, 12, 15, 3, -15, 10, 16, 11, -10,
    -- filter=27 channel=9
    -14, -2, 15, -15, 0, -10, -14, 8, -11,
    -- filter=27 channel=10
    6, 2, 12, 11, -13, 19, 9, -5, 15,
    -- filter=27 channel=11
    -16, 18, -3, 13, 8, 2, -14, -2, -7,
    -- filter=27 channel=12
    -14, -9, 19, 2, -11, -19, -10, 4, 0,
    -- filter=27 channel=13
    -3, 10, 8, -3, -17, -18, -11, -20, -6,
    -- filter=27 channel=14
    5, 16, 14, -14, -19, 14, -11, -15, 10,
    -- filter=27 channel=15
    -20, -2, -4, 4, 7, 21, 8, 20, -8,
    -- filter=28 channel=0
    -17, 20, 21, -11, -5, -16, 0, 9, 20,
    -- filter=28 channel=1
    -13, 21, -3, 4, 8, 15, 24, 12, -22,
    -- filter=28 channel=2
    -12, -19, 5, -2, -19, -3, -6, 6, -17,
    -- filter=28 channel=3
    -21, 16, 19, 1, 6, 5, 20, 2, 8,
    -- filter=28 channel=4
    0, 5, -8, -3, -3, 7, 15, -4, 9,
    -- filter=28 channel=5
    22, -16, -8, -3, 0, -20, 0, 14, -20,
    -- filter=28 channel=6
    -3, -8, -15, -5, -5, -16, 19, 5, 17,
    -- filter=28 channel=7
    -13, -9, -3, 13, -12, -11, 8, 22, 7,
    -- filter=28 channel=8
    -13, -12, -16, -9, 16, -9, -16, 10, -6,
    -- filter=28 channel=9
    -16, -8, 11, 12, -5, -19, 0, 21, 0,
    -- filter=28 channel=10
    12, -6, 10, 9, -9, -4, 14, 10, -14,
    -- filter=28 channel=11
    8, 6, -11, 0, 20, 0, -4, -15, 8,
    -- filter=28 channel=12
    -7, 10, 19, -6, 17, -3, 7, -12, -15,
    -- filter=28 channel=13
    -3, -3, -20, 29, -2, -34, 7, 15, -21,
    -- filter=28 channel=14
    18, -14, -14, -2, 13, 11, -15, -13, -5,
    -- filter=28 channel=15
    -6, -4, 24, -15, -8, -3, -8, 7, 4,
    -- filter=29 channel=0
    21, -12, -10, -17, 9, -11, -20, -2, -12,
    -- filter=29 channel=1
    -11, -15, -18, 3, -17, -6, -5, -10, -4,
    -- filter=29 channel=2
    19, -10, -16, 8, 2, 8, -21, 20, -11,
    -- filter=29 channel=3
    -17, 12, -2, 20, 2, 1, 11, -11, -4,
    -- filter=29 channel=4
    -16, 19, 5, -10, 9, 6, -15, 13, -20,
    -- filter=29 channel=5
    8, 15, 0, 4, -18, 8, 5, 11, -2,
    -- filter=29 channel=6
    -7, 20, -7, 9, -9, 0, 18, 6, 16,
    -- filter=29 channel=7
    2, -5, 4, 19, 4, 17, -21, 10, 9,
    -- filter=29 channel=8
    -7, 1, 3, 0, -3, 15, -14, -4, -17,
    -- filter=29 channel=9
    4, -6, 15, -20, -7, -7, -21, 6, -16,
    -- filter=29 channel=10
    -20, -16, 9, -15, -4, -13, -6, 13, -12,
    -- filter=29 channel=11
    13, -3, -8, -18, 5, -13, 6, -2, -21,
    -- filter=29 channel=12
    19, 6, -1, -5, -3, -2, -15, -17, -10,
    -- filter=29 channel=13
    2, 3, -9, 7, -10, 4, 16, 13, -9,
    -- filter=29 channel=14
    5, -2, 0, 12, -12, -8, -1, 0, -2,
    -- filter=29 channel=15
    -2, 15, -12, -20, 19, -19, 3, 10, -7,
    -- filter=30 channel=0
    -7, 5, 25, 13, 29, 5, -10, 9, 0,
    -- filter=30 channel=1
    2, 6, -21, 6, -27, 4, 2, 3, -12,
    -- filter=30 channel=2
    18, 5, 10, 1, 21, -6, -7, 2, -4,
    -- filter=30 channel=3
    -1, -18, 8, 9, 2, -8, 8, -17, -2,
    -- filter=30 channel=4
    4, -11, -3, 20, 4, -17, 12, -3, 3,
    -- filter=30 channel=5
    13, -26, -19, 3, -26, -7, -13, 5, 12,
    -- filter=30 channel=6
    25, -2, 6, 5, 16, -15, 10, -3, -3,
    -- filter=30 channel=7
    -13, 11, 3, -17, -8, 0, -1, 23, 25,
    -- filter=30 channel=8
    16, -19, 15, -17, 1, -19, 18, -10, 12,
    -- filter=30 channel=9
    -7, 9, 6, 11, 7, 18, -9, 15, 1,
    -- filter=30 channel=10
    21, 3, 20, 19, -11, 17, 6, 18, -6,
    -- filter=30 channel=11
    8, -8, 8, 1, 17, 6, -5, 10, 0,
    -- filter=30 channel=12
    -13, -20, 10, -5, 7, 13, -3, -8, 17,
    -- filter=30 channel=13
    20, -10, 3, -5, -29, -8, 22, -23, 11,
    -- filter=30 channel=14
    9, 8, 5, 5, -16, 9, -2, -15, -13,
    -- filter=30 channel=15
    -6, -11, 14, 25, -11, 9, 18, 19, 0,
    -- filter=31 channel=0
    10, 12, -17, -6, -14, 5, -9, -16, 20,
    -- filter=31 channel=1
    2, -14, 18, -17, 0, -12, -1, 2, 16,
    -- filter=31 channel=2
    3, -5, 19, 12, -15, 7, 8, 8, 1,
    -- filter=31 channel=3
    15, -6, -13, -16, -18, -17, -9, -12, 22,
    -- filter=31 channel=4
    16, -19, 9, -11, -8, 10, 3, 8, 0,
    -- filter=31 channel=5
    -3, -9, 12, -14, -9, -13, 12, -4, -17,
    -- filter=31 channel=6
    -10, 11, 0, -10, 17, -7, 11, -10, -10,
    -- filter=31 channel=7
    0, -7, 20, 19, -1, -7, 16, -18, 16,
    -- filter=31 channel=8
    -19, 0, -10, 18, 15, 5, -11, 0, -9,
    -- filter=31 channel=9
    6, 19, -15, 1, 3, -14, -7, -11, 6,
    -- filter=31 channel=10
    12, -12, 16, 0, 15, 11, -3, -1, 10,
    -- filter=31 channel=11
    18, 20, -11, -12, 12, -6, -16, -8, 11,
    -- filter=31 channel=12
    7, 10, 18, -9, -12, -20, 3, 15, 0,
    -- filter=31 channel=13
    -18, -7, -19, -15, 14, -4, 24, -6, 3,
    -- filter=31 channel=14
    6, 2, 7, 17, 3, -9, 4, 18, 16,
    -- filter=31 channel=15
    12, -11, 0, 13, 15, -6, -19, -1, -5,

    others => 0);
end iwght_package;
