-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;


-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity ifmap_36k_layer0_entity12 is
    generic (
        DEVICE: string := "7SERIES"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic_vector(2-1 downto 0);;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(11-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
 end ifmap_36k_layer0_entity12;

  architecture a1 of bram is

    begin

    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
       BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
       DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
       DO_REG => 0,                     -- Optional output register (0 or 1)
       INIT => X"000000000000000000",   -- Initial values on output port
       INIT_FILE => "NONE",
       WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
       SRVAL => X"000000000000000000",  -- Set/Reset value for port output
       WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
       -- The following INIT_xx declarations specify the initial contents of the RAM
       INIT_00 => X"001700130015004100a400bc00b700b200aa00ac00ba00ba00b800b700b600b7",
       INIT_01 => X"00b400a4007f005c006b006e009900c200c300c900c500c600c900c800c700c5",
       INIT_02 => X"001700130015002e009900ca00bf00b200a4009e00a900b700ba00b800b400b2",
       INIT_03 => X"00b400ad008a0056004a006a00b400ce00cf00d500d000ce00cf00cd00cc00ca",
       INIT_04 => X"001700140017001f007f00c800b900a8009f009e009a00a200b200b200b300b2",
       INIT_05 => X"00b500be00b6007d0047007200c500d100d500d800d500d300d400d300d000ce",
       INIT_06 => X"0017001500180017006300bd00af00a000a800a800a6009500aa00ba00bf00c3",
       INIT_07 => X"00c300c800bc008d0063009200d200d600d500d400d400d500d900d900d700d6",
       INIT_08 => X"0019001700170015004800aa00a5009700af00b700b9009b0092009d00a900bc",
       INIT_09 => X"00c500c400b2008d007900ac00d300db00dd00d900d900d900d600d400d100ce",
       INIT_0A => X"001a001b001a00170031008f00a4009a00a900c200c800a60082007d00800097",
       INIT_0B => X"00a500a50094008f009300b600bc00c900d400d900d500db00dc00d700d700d3",
       INIT_0C => X"001e001a001b00190025007d00b400ab00a900c500ca00b3008b0071007a0082",
       INIT_0D => X"00770085007a008c00b900cb00bf00c900d700da00d700db00dc00da00dc00e0",
       INIT_0E => X"005e0030001f0024006400af00c100a800a300c000c600c300ae0091008e0084",
       INIT_0F => X"006a0079007a008b00c000d100bd00d500f200ed00ef00e800d000d500de00e5",
       INIT_10 => X"00b4009e0072007a00b100be00be00a0008500ad00c500c800c200b900a70092",
       INIT_11 => X"008100810085008d00b100c900bd00dc00f100eb00e800d500bd00c700e100ea",
       INIT_12 => X"00c500c000b200ba00c100c300c5009d008000a300b900bf00c100c300b20097",
       INIT_13 => X"007200810083008600aa00c200d000ea00ec00f000eb00c900b900bb00d000eb",
       INIT_14 => X"00ca00c400bb00c000c800cd00c50097009500af00b800bd00c100bb00a80088",
       INIT_15 => X"007500800080008100a700b500cd00f000f300f300ee00ce00ba00bb00c100dd",
       INIT_16 => X"00cd00cd00c500c000cb00d000c200a000a800bf00c100bf00c100ac00920077",
       INIT_17 => X"007c008e0085008700a700b000bf00ea00f300f100ec00d700ba00b800b900c4",
       INIT_18 => X"00ce00cc00c800c100c500c700bf00b400ac00b300b700ad00ae00ae00980083",
       INIT_19 => X"008d00a6008e009a00a900ac00bf00e600f000f100ef00e400c800ba00b800c0",
       INIT_1A => X"00d200ca00c600bf00c900b400b100ca00ab009a008e008e00a800a80093009c",
       INIT_1B => X"00af00a9009600a4009e00a000c500e600f100f100f400f200e200bf00c300d7",
       INIT_1C => X"00d300c900c700c000cf00aa00a100d700bd00ba00ad00ac00be00b10089007f",
       INIT_1D => X"00b400ae009600a000af00b000c100ec00f500f200f300fb00ef00c900d400e1",
       INIT_1E => X"00d300c400c500c100d100b5009a00d900ce00c500c300b900aa00ad00a60098",
       INIT_1F => X"00a300b800a6009800c000b500af00cc00ee00f300f400f700df00d500e200e2",
       INIT_20 => X"00d600c200b400b500c500c4009b00c600d600c000ae00b700ad00a100ae00b2",
       INIT_21 => X"008000a400bd009300a700b4009c0076009d00d700ef00eb00ce00d600ea00e4",
       INIT_22 => X"00d700c600a600a300b400ca00be00b900cf00d200cd00d600c100ae00b000ad",
       INIT_23 => X"0081008900bf009900a300c800ab00870074009000b800c100bb00d200ef00eb",
       INIT_24 => X"00d800cd00ae00a400b900cb00d200c200bf00d300da00e200e100cb00be00b3",
       INIT_25 => X"0097007900a8009e00a700c200aa00ac009a0083009900a900a200b800de00ec",
       INIT_26 => X"00d800d000c000b400c500ca00d100d200ba00bd00c500cc00d100d500cf00b5",
       INIT_27 => X"00b20095009200af00b700ae009c00ab00a3009400a900b400a600a000ac00cc",
       INIT_28 => X"00da00d500ca00b600bf00cb00c900ca00ca00c300c100c000b200c600cf00c7",
       INIT_29 => X"00d300cb00a600bb00b1009b009300a600a700ab00b600af009c009c009f00a7",
       INIT_2A => X"00d900d700d100ba00b300c800d000c800d100d700d200ba00a100b600c400c2",
       INIT_2B => X"00cb00cf00be00b9009b008e009b00a600ac00b300ad009f0096009e009e008f",
       INIT_2C => X"00d600d500d600c000a900c500da00d900d700d900d400c300aa00b300c300bf",
       INIT_2D => X"00be00c000c000aa0084008e00a700aa00aa00b300ad009d009d00930086007d",
       INIT_2E => X"00d500d100d300ca00a800c100d800de00df00de00d300cd00c200c200c900c6",
       INIT_2F => X"00c600c400bc00990086009b00ab00a700a600bd00b200a500a3008e00850089",
       INIT_30 => X"00d300ce00ce00ca00af00bf00d300d500d600d800c600ab00c200ce00c900c9",
       INIT_31 => X"00c800c500b100960090009e00a7009d009f00b500b000a80098009600950090",
       INIT_32 => X"00d200cc00c900c100b500bc00d000d200cd00ce00a0007a00b100d000c600c2",
       INIT_33 => X"00c100b800a60096008b009c00a00099009b00a0009f009b00980098008c0083",
       INIT_34 => X"00d200ca00c600bb00ae00b200cd00d600d100cb00a4008300b400ca00bb00b6",
       INIT_35 => X"00b600a9009d008b00860099009a00900097008d0083008d009d009b00960093",
       INIT_36 => X"00d200c800c200b500a800a800c400d700d400c700bd00b800cb00b900ad00ac",
       INIT_37 => X"00a3009b00930076008300940091008d00900084007f0085009500a300a2009c",
       INIT_38 => X"00d000c200bd00b400a2009e00bd00d300d300c500c200c700bf00ac00a300a4",
       INIT_39 => X"009e00930082006d008900900090009100900084007c0086009700a2009f0093",
       INIT_3A => X"00c200b100b000b5009f008f00b300cd00d000c700c200be00b500a5009c00a1",
       INIT_3B => X"009500880070007200890085008a00920092008300830090009600950094008d",
       INIT_3C => X"00ac009d00a500b200a70085009c00c700ce00c700c700c200a000850084008b",
       INIT_3D => X"008c007e006b007e00820081008a0095008d008c0091008e0088008c00950098",
       INIT_3E => X"009700860090009b009e007d008200b700c500bf00b700a500800067005e0069",
       INIT_3F => X"007700700075007c0079007d008b008f008b008c0081007d00840095009b0096",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INIT_40 => X"001300150010002f008300930093008e008700890090008e008d008c008c008f",
       INIT_41 => X"008c007e00600049005f005d008200a4009b009c009b009d009e009b00980097",
       INIT_42 => X"001400140011001f007a00a1009b0092008a0088008b00950098009600920097",
       INIT_43 => X"009f00960075004900410058009c00af00a800a900ab00ad00ac00a800a400a3",
       INIT_44 => X"0014001400140015006600a20097008c008d00950088008b009a00990098009f",
       INIT_45 => X"00a600ab00a1006d003a006100b100b700b300b200b100b200b100ad00a900a6",
       INIT_46 => X"0014001400150011004f0099008c0082009700a4009d0087009900a600a900b0",
       INIT_47 => X"00b000af00a100760052008500c400c300bd00b700b400b300b300b100ad00ab",
       INIT_48 => X"00150014001500130038008900820077009c00b200b300920084008b009400a7",
       INIT_49 => X"00af00a900980078006d00a700ce00d200d100c900c300bf00ba00b600b100ac",
       INIT_4A => X"00160016001700160026007300820078009200b900c3009e0076006c006b0084",
       INIT_4B => X"0092008f00810084008f00b700be00c700cf00d100cc00d100d100ca00c700c2",
       INIT_4C => X"0018001300150014001e007100a10094009700ba00c200aa0080006200690071",
       INIT_4D => X"00680074006b008000b200ca00c000c500ce00cf00d100d700d800d600d700da",
       INIT_4E => X"005800290018001d006000ae00ba009c009500b500bd00ba00a4008400810076",
       INIT_4F => X"005c006b006c007c00b400cc00bb00ce00e600e000e700e400cd00d300dc00e2",
       INIT_50 => X"00b10099006d007500af00bd00b70093007800a100bc00c000b800ad009a0083",
       INIT_51 => X"007300730077007f00a600c500bc00d800e900e200e300d300bc00c600e000e8",
       INIT_52 => X"00c200bc00af00b600bf00c200be00900073009800b100b600b700b600a4008a",
       INIT_53 => X"006600760077007b00a000bd00d000e900e800eb00ea00cb00bb00bd00d100eb",
       INIT_54 => X"00c700c000b700bb00c600cd00bf008a008800a500b000b500b800af009a007c",
       INIT_55 => X"006b007600770078009e00b000cd00f000f300f400f200d400c000c000c600e0",
       INIT_56 => X"00c900c900c100bb00c900d100bc0092009b00b600b900b700b7009f0084006b",
       INIT_57 => X"00730085007c007e009e00aa00bd00eb00f600f600f200de00c200c000c000ca",
       INIT_58 => X"00cb00c900c500bd00c400c600b700a5009f00aa00b000a500a400a2008a0078",
       INIT_59 => X"0085009f0087009200a100a500bd00e700f400f800f700ea00d000c300c100c7",
       INIT_5A => X"00d000ca00c400b900c100a7009c00b900a100910087008700a1009e0089008f",
       INIT_5B => X"00a400a4009500a20099009d00c300e400f200f700f900f500e800c700cc00de",
       INIT_5C => X"00d200cc00c500b600bf008e007d00c100b500b100a600a700b800aa00820072",
       INIT_5D => X"00a500aa0098009e00ab00ae00bd00e700f200f400f500fb00f200cf00dd00e9",
       INIT_5E => X"00d400c800c500b900bd0091007000c000c700be00bd00b400a400a700a00089",
       INIT_5F => X"009200b000a2009100b800b100a800c300e800f100f500f900e400dd00ec00eb",
       INIT_60 => X"00d800c700b600ae00b0009b006e00ad00d000ba00a800b200a8009b00a700a4",
       INIT_61 => X"006e009600b10086009a00ab00900068009100d100ee00ed00d200dd00f300ed",
       INIT_62 => X"00db00ce00a9009e00a300a7009500a200ca00cd00c800d100bc00a800aa00a1",
       INIT_63 => X"0070007800ad0087009300ba009b00730062008400b200bc00b900d400f300ef",
       INIT_64 => X"00dd00d600b300a100af00b500b300b100bd00cf00d400dd00dc00c500b800ab",
       INIT_65 => X"008b00670095008c009700b10094009300830070008a009c009700b100d900ea",
       INIT_66 => X"00df00da00c600b200c200c200be00c800ba00b800bf00c700cb00d000c800b1",
       INIT_67 => X"00ab0087007f009e00a8009b0083008f0089007e0094009f00930090009e00c5",
       INIT_68 => X"00e100dd00d000b700bf00c700be00c200c600bc00be00ba00ab00c100c600bf",
       INIT_69 => X"00cf00bf009400a900a00087007b008d008e0095009f009800870088008c009a",
       INIT_6A => X"00de00dd00d600be00b300c300c800be00c600cd00d100b2009700b300b600b5",
       INIT_6B => X"00c500c400ae00a50086007c00890093009900a10099008b0083008b008b007d",
       INIT_6C => X"00db00da00db00c600aa00bf00d200cf00cb00ce00cf00b4009c00ae00b400b0",
       INIT_6D => X"00b600b500b00096006f007d00960098009800a1009a008a008a00800073006a",
       INIT_6E => X"00da00d600d900cf00aa00bc00d200d500d400d300c700b600ae00ba00ba00b5",
       INIT_6F => X"00ba00b600ab008500720089009a0095009400ab009f00920090007b00730076",
       INIT_70 => X"00d800d400d400d100b300bd00cf00cd00cd00cd00b1008a00a700c300bb00b6",
       INIT_71 => X"00b900b5009e0082007d008d0096008c008d00a3009d0095008500830082007c",
       INIT_72 => X"00d700d200d000c800bb00be00ce00cc00c600c400830050009100c200b800ae",
       INIT_73 => X"00ae00a5009300830078008b008f00880089008e008c00880085008500790070",
       INIT_74 => X"00d700d000cd00c200b500b700cd00d100cc00c200810051008e00ba00ab00a1",
       INIT_75 => X"00a1009500890078007300870089007e0085007b0070007a008a008800830080",
       INIT_76 => X"00d600cd00c800bc00b000af00c600d400d000c000a0008e00aa00a8009b0095",
       INIT_77 => X"008d0085007f0064007100830080007b007e0072006c00720082009000900089",
       INIT_78 => X"00d200c400c000b700a900a600c000d200d100c000b600b400ab0099008d008c",
       INIT_79 => X"0086007d006f005c0078007e007e007f007e00720069007400850090008d0081",
       INIT_7A => X"00c400b300b300b900a6009700b500cc00cd00c200ba00b300a6009200850088",
       INIT_7B => X"007e0072005d00610078007300780080008000710071007e008400830082007b",
       INIT_7C => X"00b100a100aa00b800ae008c009c00c300c900c100bf00b600910071006c0073",
       INIT_7D => X"0076006a0059006e0072007000780083007b007a007f007c0075007a00820086",
       INIT_7E => X"009d008c009700a100a60082008000b100bf00b700af009a0070005300470053",
       INIT_7F => X"0063005e0065006e006c006c0079007e0079007a006f006b0073008400890084",

       -- The next set of INITP_xx are for the parity bits
       INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

       -- The next set of INIT_xx are valid when configured as 36Kb
       INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
       INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
       DO => DO,      -- Output data, width defined by READ_WIDTH parameter
       ADDR => ADDR,  -- Input address, width defined by read/write port depth
       CLK => CLK,    -- 1-bit input clock
       DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
       EN => EN,      -- 1-bit input RAM enable
       REGCE => REGCE, -- 1-bit input output register enable
       RST => RST,    -- 1-bit input reset
       WE => WE       -- Input write enable, width defined by write port depth
    );


-- End of BRAM_SINGLE_MACRO_inst instantiation
