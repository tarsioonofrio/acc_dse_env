library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    -63, 126, 276, 171, 3, 65, -74, -22, -39, 177, 193, 129, -22, 186, -321, 27, 60, 81, -9, -63, 38, -44, -152, -10, 136, 81, 129, -30, 265, 152, 203, 31, 81, -278, -39, 33, 65, 294, 124, 124, 181, -134, -30, 36, 72, 174, -168, -142, 142, 328, -153, 90, -95, -40, 78, -30, 368, -75, -232, -105, -126, -172, 213, -418, -129, 38, 101, 105, -40, 188, -268, 77, -280, 31, 41, -189, 77, 57, -156, 75, -278, 69, -68, 102, -91, 100, -80, -7, -114, 204, 73, 65, 48, 190, 208, -107, 156, 225, -16, -2, -9, -89, -44, -148, -293, -176, 15, 76, -35, 234, -111, -232, -141, -48, -129, 237, -108, 181, 37, 239, 199, 120, -173, -56, 153, 37, 41, -116, 11, -216, 196, 21, 56, -100, 196, 111, 28, -127, 60, 193, -100, 117, -63, 114, 484, 137, 136, 2, -109, 150, 211, -139, 76, 83, -14, -107, -160, -81, -7, 158, 171, -135, -47, 185, 182, -137, -41, 231, -14, -20, 419, -30, -1, -151, -90, -149, 97, -203, -324, 4, -120, -24, 38, 48, -167, 422, 3, -83, 407, 80, -153, 38, 17, 149, 121, -255, -40, 125, 163, 319, 161, -204, 24, 58, -135, 41, 71, 80, -164, 146, -102, 129, -76, 111, 43, -59, 32, -116, 44, -43, -185, -171, -117, 17, 70, 95, -121, 265, 155, -104, -21, -55, 69, 276, 64, 379, 279, -164, -243, -142, -37, 20, 29, 158, 328, -48, -87, 171, -25, 419, -131, 175, -44, -60, 100, -207, -318, 2, 79, -200, -117, -40, -49, -13, 51, -104, -48, -2, 123, 19, -51, 15, 85, 97, -35, -196, 80, 158, 300, -303, 146, -310, 18, 397, -20, -92, 245, -9, 445, -62, 41, -81, -70, 177, -43, 187, 9, -44, -65, -194, -47, -115, 276, -25, 137, 84, 234, 19, 2, 98, 121, 188, 147, 139, 159, 212, -166, 326, -148, 219, 17, -3, -223, 104, 51, -79, -190, 322, -54, 20, -64, 346, 243, -257, -12, -149, -281, -132, -97, 16, -69, -36, -72, 66, -136, 23, -73, 94, -158, 131, -180, -148, 33, 267, 58, 137, -59, 26, -57, 92, -148, -38, -44, -18, 462, 38, 201, -66, -127, 256, -84, -3, 135, 312, -206, -164, -185, -67, -81, 238, 271, -336, -233, 141, -203, 102, -10, 50, 37, 184, 171, 15, -209, -172, -13, 10, 164, -62, 207, 85, -130, 41, 75, 56, -40, -60, -63, -203, -1, 68, 44, 26, 92, 22, 36, 297, -20, 88, 38, -139, -105, 40, 177, 59, 75, -79, 35, 341, -52, 79, 48, 142, 179, 157, 112, -44, 151, 274, -538, 106, 64, 17, -14, 146, 1, -53, 2, 22, -17, 124, -31, 41, -154, -37, -26, 214, 61, 129, 4, 83, -148, -116, 428, -134, -1, -102, 227, -94, -3, -19, -1, -170, -71, 60, 237, 318, 43, 120, -56, 141, 194, 129, 200, 28, 126, -66, 107, 16, -113, -91, -144, -100, 18, -35, -272, 372, 211, 71, 128, -57, -42, -167, 64, 32, -26, -66, -44, 67, -46, -103, -42, -290, 155, 169, 224, -68, 128, 0, -110, 108, -90, 239, 107, -144, -76, -46, 91, 93, 75, -63, 3, 43, 29, 20, 425, -21, 9, -2, 5, -25, -61, 113, 45, -59, 228, -14, 13, 39, -110, -36, 25, -8, 54, 79, 169, 95, -63, 36, 1, 81, -104, 34, 92, 97, -222, 171, -30, 297, 321, 90, 10, -21, 48, -1, -47, 34, 201, 253, -69, 406, -204, 253, 110, -25, -137, 280, 230, -106, -189, -53, 14, 23, -138, -264, -214, -4, -103, 227, 63, 321, 35, -111, -84, -35, -255, -15, 30, 66, 18, -118, -138, 87, 168, 103, -184, -29, -15, 46, -14, -131, -85, 49, -63, 15, -227, 269, 179, 132, 96, 83, 27, -62, 119, 39, 288, 285, 355, -143, -179, -173, -165, -128, 71, -167, 64, -4, -52, 58, 73, 36, 28, -141, 23, 26, -23, 65, 306, -190, 82, 45, 64, 106, 154, 69, -36, -101, 103, -128, 91, 134, 228, -98, 287, -45, -4, 11, 146, 31, 130, -19, 285, -35, 102, 141, 70, -5, -14, 230, 109, -127, -364, 27, -32, -93, -85, 80, 29, -239, -129, 124, -90, -67, 202, 84, -89, 23, -252, -35, 176, 61, 78, -31, 221, -338, 143, 367, 157, -229, -132, 14, 248, -108, -152, 94, -74, -201, 122, 208, -103, 314, 370, 5, 323, 115, 17, 115, 116, 176, -98, -279, 43, -125, 73, -45, 43, -46, 181, -99, 105, 280, 326, 50, -64, 257, 163, 83, -155, 36, 203, 177, 45, -107, 124, 152, -287, -61, 74, 77, 125, -64, -111, 55, 97, -221, 148, 39, 21, 4, -267, 32, 16, 21, -256, 57, 176, -42, 139, 3, -113, 284, -166, -236, 55, 301, -172, -107, -8, 94, 161, -277, -14, 63, -101, 58, -28, -9, -59, -155, -64, -64, -133, 100, 168, -85, 49, -183, 286, -71, 39, 96, -124, -146, -68, 178, 287, -104, 64, 84, 95, -2, -26, -26, 125, 134, 132, -38, -45, -142, 145, -242, 57, 118, 62, -149, -184, -126, 41, -46, 343, -185, -140, -202, 103, -86, -41, -192, -86, 273, -86, 141, -274, -61, 213, -11, 106, 43, 62, 180, 101, -46, -73, 11, 63, 98, -156, -80, 91, 210, 332, -72, 153, 25, 45, 215, -100, -8, 225, 20, 195, 106, 244, 9, 269, 75, 128, 17, 100, 162, 171, -31, -91, 50, 39, -91, -157, 17, -93, 23, 214, -245, 31, 218, 10, -108, 288, -133, 45, 60, 43, 82, 2, 43, -55, -84, 98, 364, -157, -125, -49, -143, -38, 12, -37, -175, 188, -23, 23, 10, -126, -90, -43, -93, 217, -25, 54, 9, 49, 40, -114, 36, -73, 296, -52, -226, -116, 112, 132, -96, 32, -155, 204, 206, -47, -96, 58, 222, -130, 13, 175, 30, 150, 332, -253, 180, 221, -104, -158, -39, -82, -34, 52, 207, 2, -152, -36, 47, 128, -28, -89, -104, 7, -77, 24, -80, -68, -98, 146, -2, 19, 190, 104, 252, 230, 76, 54, -39, 21, 25, -188, -132, -82, 321, 77, 241, -126, 250, 115, -113, 21, 212, -77, 17, -100, 283, -26, 114, -87, -18, 70, 343, 282, 162, 130, -77, -44, 89, 213, 94, 13, 91, -17, 123, 47, 455, 248, 112, 82, -223, -6, 55, -10, 83, 161, -25, 68, -113, -300, 57, -39, 5, 91, 75, -92, 108, -28, -34, 152, -80, -225, -24, -31, 132, -166, 35, -171, 265, -220, -13, 48, 394, -58, -71, -46, 176, -19, 71, 42, -293, 55, -10, 67, 77, 222, 44, 119, 39, 122, -196, 3, -182, 128, 18, -58, -28, -89, 94, 62, 214, 29, -47, -5, 176, 4, -22, -52, 35, 99, 119, -89, 11, -17, 80, 2, 146, 174, -45, 246, 6, 26, 118, 190, -72, -106, 64, -229, -207, -122, 342, -145, 61, 68, -55, 66, -160, -37, 141, -7, -208, -233, 221, -142, 40, -149, 142, 108, 85, -51, 339, -113, 157, 66, 122, 114, 115, 47, 89, 107, -154, -94, 243, 201, -52, 321, 5, 90, 34, 89, 104, 194, -242, -144, 19, 124, 22, -85, -98, 121, 68, -213, -76, -74, 5, 618, 127, -217, -240, 177, 56, 417, -45, 26, -10, -247, 184, 26, 230, 32, 4, 119, -179, 41, -61, -95, -57, 198, 305, -168, 56, 220, 22, -38, 113, 46, -223, 15, -55, 30, 49, 30, 262, 7, -76, -52, 186, 115, -71, -358, -61, -108, -96, -168, 76, -209, -136, 47, 38, 344, -34, -115, 23, -341, 130, 135, -133, -9, -104, -267, 22, -74, 64, 59, -12, 169, 397, -59, 0, -77, 32, -157, 62, -33, 95, 86, -134, -171, -56, -247, 117, 128, 97, 109, 91, 196, 60, 579, -66, -188, -230, -9, 176, 208, 65, 167, -126, 304, 273, 313, -178, -152, -67, 230, 118, -190, -11, -11, -373, 122, -33, -10, -76, 85, -298, 84, 82, -102, -15, -10, -179, 71, -130, 365, 10, 33, 108, 117, -221, 159, 8, 259, 45, -269, -109, -75, 22, 239, 78, 173, 234, 186, -15, -142, -23, -161, 181, 255, -5, -23, 10, -75, -88, 56, -9, 191, -134, -9, 182, -22, 14, 47, 85, 65, 95, -224, 147, 187, -14, -213, -40, -167, 86, 6, -235, 46, -211, -146, -118, -48, -17, -43, 186, -13, -142, -15, 410, -74, 110, -10, 26, -21, -80, 30, -154, -113, -13, -20, 79, -106, -39, -14, -222, 45, -110, -396, 85, 472, 0, 141, -23, 200, -50, 123, 30, -38, -84, 83, 30, 38, 111, -97, -150, -131, 73, -17, 9, -473, 62, 63, -28, 180, 80, 89, 232, -186, -59, 221, 43, 6, -15, 87, 121, -199, 98, 232, 79, 197, 80, -140, 35, 17, 160, -65, 165, -83, 95, -109, 81, -16, -68, -31, -254, 2, -31, -134, -107, -201, 121, 47, -70, 308, 146, -238, -62, -99, 130, 89, -101, -92, 92, 330, 95, 43, 149, -103, -228, -92, -17, 16, -5, -90, -90, -43, 65, -133, 397, 109, -76, 62, -294, 223, 148, 117, -36, 332, 89, -42, 131, 92, -57, 382, 96, -104, -113, 19, 82, 200, 141, -47, -86, -8, 121, -340, 228, 255, 21, -54, 52, -226, 167, 346, 143, 56, -227, 53, -217, -32, -101, 53, -57, 242, 115, 107, 288, -140, 41, -4, 107, 72, 30, -146, -123, -127, 162, 115, 53, -151, -59, -71, 190, -303, 382, -50, 235, -18, -138, -42, 161, 141, 284, -3, 136, -114, 52, 21, 33, 112, -17, -82, 52, -44, 88, -107, -120, 232, 100, 85, -176, -244, 26, -42, 4, -98, -72, -26, 75, -83, 10, -49, 424, 102, -196, 286, -35, -22, -42, -128, 316, 53, 81, 218, 150, -81, 235, 254, -373, -90, 187, 9, 26, 164, 19, -124, -248, 108, -24, -34, -218, 21, 229, -147, -62, 161, -69, 268, 91, -241, 160, -1, 53, -11, -111, -74, -100, -75, -35, -131, -44, 169, -156, -135, 326, -80, -55, -102, -24, -125, 67, 92, -89, -171, -57, -170, -96, -61, -1, -61, -205, 167, -59, -116, -136, -65, -13, -113, 184, 33, 75, 201, -159, 201, -54, -17, 113, -16, -134, 26, 218, 273, 340, 416, 715, 65, 96, -95, -120, -133, -31, 146, 77, -24, -152, 185, 155, 103, -367, -100, 84, 13, -65, 6, 122, 68, 28, -97, -14, -158, -57, -31, 117, -97, 293, -107, -41, 50, -94, -109, 16, -140, -71, -45, 67, 321, -162, 298, -90, 115, 94, -157, 288, 119, 132, -71, -88, 57, -146, -249, 118, -16, -106, -5, 22, 269, 62, 276, 24, -20, -371, -87, -49, 61, 99, -102, 150, 112, 116, 174, 15, -45, 102, 200, 153, 274, -20, 49, -244, 114, 25, -77, -211, -52, 120, -237, 25, 100, -185, 162, 35, 84, 99, 122, 126, 70, 204, 257, -227, 187, -246, 256, 0, -198, 230, -38, 144, 159, 87, 28, 14, 253, -54, 38, -47, -96, 115, 28, 23, 57, 38, 39, 108, 19, -41, 132, -114, 75, 153, -46, -74, 92, -159, -153, -102, 441, 243, 71, -203, 379, -72, -3, -51, -209, -88, -119, 84, -187, 82, -206, 65, -70, -39, 199, 244, -17, -180, 77, -77, 142, 188, 91, -81, 9, 225, -154, -188, -169, -10, 325, 46, 83, -108, -347, -94, 168, -177, -96, -227, 63, -39, -155, 56, -145, 98, 38, -89, -168, -72, -131, 202, -252, 121, 467, 69, 93, 345, 56, 193, 138, 311, -103, 206, 92, 139, 87, 113, -335, -58, 464, 139, -179, 9, 476, 61, -244, -165, -12, 89, -115, 78, 75, 37, -185, -115, -73, 22, 84, 134, -31, 105, -122, 189, 159, -289, -171, -173, 150, -79, 95, 70, 136, 64, 235, 65, 87, -12, 63, -91, 261, -59, 187, 184, -78, -105, -114, -63, 239, 225, -193, 60, -207, -103, 39, -205, -56, 98, 385, 73, -115, -123, 31, 311, -160, 162, -294, 59, 105, 51, -169, -70, 108, 57, -3, 84, -173, -33, 22, 351, -49, 32, 108, -119, 121, 16, -276, 371, -117, 43, -79, 28, -34, -79, 250, 83, 279, -338, -398, 69, 38, -150, 208, 62, -100, 104, 248, 238, -42, 25, 89, -46, -62, -124, -18, -94, 175, 20, -75, -17, 274, 89, 7, -22, -33, -182, 294, 19, 69, 76, -130, -37, 124, -102, -299, -182, 88, -51, -4, 380, 14, 19, 153, -92, -138, -154, -129, -85, 24, 72, 137, -27, 111, 173, -69, 295, 319, -45, -193, 44, 406, 190, -75, 187, -168, -139, -62, 86, -46, 90, 63, 38, 62, -166, 51, -32, -83, -45, 139, 131, -27, 26, -146, 60, 98, -260, -480, 139, -226, -173, -113, 151, 119, -99, -18, 121, 130, -111, 19, 119, -83, 235, -78, -138, 154, 94, 100, 28, -71, 11, -71, 57, 218, 19, 313, 52, -172, 146, 33, 68, -14, -249, -229, 250, -9, -5, -168, -192, 63, 152, 89, 119, -15, 9, -138, 57, 18, 152, 149, -28, 124, 27, 81, -74, -52, 127, -34, 101, 397, -392, 8, -37, -40, 131, -70, 48, -231, 90, -126, 77, 5, 10, -148, 2, -141, -86, -31, 39, -161, 67, -85, 322, 248, 267, 100, -82, -261, -84, -22, 84, 159, 9, -145, -114, -107, -135, -92, 178, -54, -79, -180, -157, -5, -131, -128, 385, 93, 329, 111, 17, 205, -9, -1, -273, 70, 74, -110, 308, 86, -128, -211, 27, -195, 2, -221, -235, -220, 28, 243, -6, 25, -163, 41, 132, -4, 47, 121, 69, -115, -9, -63, 47, 136, -61, 293, -44, -85, 267, -331, -22, 30, 322, -56, 237, 141, -212, -132, 119, -25, -54, 320, 202, -81, -213, 40, 138, -10, 310, -47, 9, 91, 32, -44, -109, -227, -117, 116, -151, -130, -276, 63, -168, 205, 114, 191, -8, 148, 337, 103, 48, -66, 151, -342, 26, -132, -32, 77, -72, -31, 132, -13, 109, -80, 161, -129, -78, -103, 3, -105, 235, 
    
    
    others => 0);
end gold_package;
