library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=2
    -6993, -2941, 264, 3156, 9225, -10518, 12743, -7809, 6545, -5077,

    -- weights
    -- layer=2 filter=0 channel=0
    8, 12, -35, -55, -52, -4, 59, -5, 5, 45, -49, -20, -61, 13, 10, -13, 14, -6, 11, -57, 0, 18, 0, 4, -27, 31, 21, 15, -5, 0, 4, -12, 29, -29, 16, -48, -2, 14, -43, 7, 6, -46, -71, 5, 3, 6, 35, 28, -96, -5, -5, -71, 0, -22, -5, 12, 18, 46, 37, -18, 10, -5, 43, -38, 10, -5, -13, 6, -55, 1, 18, 8, 0, 13, -70, 32, -53, -2, 13, 7, -45, 17, 3, -26, 6, -6, 18, -31, -14, 55, 19, 39, -8, -35, 2, 2, 39, -49, 39, -30, -22, -1, -2, 8, 6, -35, -62, 7, -7, -4, 41, 10, -106, -40, 13, -16, 6, 22, -43, 1, -6, 35, 35, -28, 2, -13, 53, -31, 4, -6, -2, -41, -23, -14, 2, -2, -5, 14, -23, 23, -34, 0, 10, -11, -23, 11, -10, -24, -1, 20, 5, 5, -8, -6, 22, -22, -9, -45, 18, 17, -9, -39, 9, 8, 18, 0, -20, -12, -7, 32, -60, 28, 0, 2, -11, 8, -38, -11, 6, 5, 17, -1, -9, 4, 18, 31, -34, 0, 2, -16, 41, -39, -9, -5, -35, -40, -39, 13, 33, 7, 3, 19, -42, 30, -31, 16, 1, 2, 13, 32, -22, -22, 0, 34, -10, -13, -3, 20, 19, 17, -1, -11, 8, 3, 17, -7, 24, 43, 71, 6, -23, -12, 6, -32, -31, 19, 8, 0, -6, 0, -77, 49, -1, -10, 26, 28, -5, -10, 6, 0, -7, -31, 7, -33, 26, -40, 1, 11, -28, -60, -71, 6, -2, 7, 17, 28, -35, 15, 0, 3, -8, 6, 27, 58, 5, -54, 9, 36, 4, 15, 5, 21, 24, 7, 8, -87, 24, -6, -16, -11, -9, 24, 47, 16, -35, -11, -1, 0, -79, 20, 1, -4, -26, -26, -24, 28, 8, -54, -4, 37, 3, 8, 5, -1, -15, -47, -1, -17, 20, 12, 11, 9, -6, -36, -51, -2, -27, -6, -6, 12, 0, 15, -47, 21, 8, 6, 12, 5, 2, -59, -6, 2, -5, 7, 7, 3, 22, 0, -16, -4, 57, 3, -55, 9, 5, 9, -15, -7, -14, -14, -3, -37, -53, 22, -1, 0, -6, -5, -13, 54, 1, -38, 16, -2, -1, -5, -17, 20, -75, -24, 7, -52, 34, 0, 9, -6, -29, -44, -44, -8, 12, 2, 1, 18, -5, -7, -64, -1, -19, -4, 11, -27, 18, -57, -2, -5, 2, 40, 3, 3, 26, -29, 1, 15, 8, 11, -27, 14, 25, 1, -5, -6, -40, -3, -8, -35, -42, 10, -1, 0, -3, -9, 61, 68, 5, -1, -9, 0, 17, 3, 35, 25, -87, -20, -1, -17, 21, 19, -10, 2, -11, 2, -9, -11, 37, -7, 4, 0, -40, 40, -44, 1, -9, -7, -4, -8, 10, -22, 10, 15, -35, -37, -4, 19, -3, -9, -3, -3, 42, 3, 20, 3, -1, -11, 0, 8, -49, -11, -1, -5, -35, -9, -4, -12, -7, 3, -22, -44, 6, -25, 1, -22, 5, 4, -15, 45, 50, -13, 17, -17, 42, -29, 7, -8, 0, -11, 0, 4, 25, 0, -17, -24, -41, 11, -38, -7, 1, 5, -66, 25, -17, -1, -6, 6, -20, -21, 21, 37, 36, 17, -5, -48, -1, -11, 33, -46, 31, -26, 36, 19, -27, -1, -9, 7, 25, 3, -6, 0, 2, -13, -48, -44, 11, -29, 21, 18, 4, -4, -33, 20, 82, -28, 0, 12, -3, -40, 4, -3, -2, 35, 18, 10, 29, -3, -6, 15, -24, 58, 0, 12, -13, 8, 3, -15, -22, -14, 2, 15, -13, -15, -7, 22, 24, 4, -12, -18, 6, 1, 52, -69, 28, 29, 39, 6, -24, -2, -12, -16, -8, 10, 0, 13, 1, 31, -58, -8, 1, -10, 15, 1, 19, 8, -3, 15, 38, 9, -3, -1, 15, -27, 3, 4, 0, -17, -15, 7, 27, 3, -1, 12, 8, 16, 5, 19, -14, 0, 15, -19, 0, -2, -8, 43, 33, -34, -2, 7, 52, -1, 2, -9, -22, -3, 7, -19, 42, -2, 52, 32, -13, 7, -6, -27, -21, 7, -6, -2, -31, 8, -5, 13, 10, 44, 1, 47, 48, 8, -8, 7, 29, -14, 4, 9, -19, 6, -2, -1, -1, -6, -4, -8, 27, -9, 9, 3, 23, -18, -15, -6, 8, 7, 27, 37, -10, 4, -9, 13, 31, -6, 26, -4, 25, 12, -2, -15, 0, 0, -21, -36, -1, 0, 16, 12, -25, -11, 4, -3, -9, 17, 3, -4, -2, 14, 14, 18, 11, -33, -9, 10, 26, 6, -15, 9, -63, -25, 4, -4, 18, 4, 7, 10, 1, 0, -14, -1, 19, 3, -14, -8, 13, -11, -14, -1, 19, -6, -16, -11, 1, 0, -9, 5, 24, 1, -8, -7, 13, -17, -2, -17, 27, -19, 0, -2, 17, 15, 14, 10, -17, -12, 3, 23, 17, -2, 5, 0, -21, 18, 40, 68, -6, -35, -11, -22, -14, -4, 11, 9, -51, -41, 0, -23, 13, 44, 5, -13, -8, 3, -46, -24, -10, 0, -5, 6, 38, -21, -30, -11, -9, -5, -34, -26, -25, -13, 2, -14, -1, 29, -24, 27, 10, -35, -9, -19, -7, 8, -15, -29, 22, -10, 2, -15, -20, 6, -4, 34, -20, -5, 7, 1, -26, 18, 59, 75, -5, -26, -37, 23, 18, 22, -26, 31, -64, -37, -12, -39, -15, 49, -4, -8, -6, 15, 3, 0, 20, 9, 19, -23, -1, 49, -20, -8, 27, 7, 42, -32, 1, -34, 2, 40, -27, -24, 0, 45, 0, -12, 6, 28, -7, 1, 41, -41, 40, -8, -5, -3, -17, 7, -4, 2, 6, 16, 0, -39, 5, -25, -37, -52, -9, -60, 15, -3, 28, -14, -48, 6, 90, 50, -12, 0, 22, -60, -5, 1, 6, 7, -28, -12, 2, 0, 9, -28, -21, 23, 9, -20, 34, 2, 1, 15, 4, 49, -2, 43, 8, -45, 43, 63, -8, 26, -15, -4, 7, -14, 42, -20, 20, 1, 30, 10, -7, 5, -13, -33, 42, 1, -3, -9, 27, 18, -51, -40, -3, 13, 32, 16, 20, 9, -21, 35, 106, 35, -15, -15, -8, -32, -5, 1, -12, -9, -16, 14, 5, 9, 14, 9, 5, 0, -10, 3, -32, 0, 20, -4, 2, -3, 0, -6, -12, 1, 22, 28, 24, 20, -1, -16, -44, -13, 17, 7, 63, -39, 46, 25, -27, 1, 3, 20, -19, -15, 3, 11, -16, 35, -2, -31, -4, 22, 12, -12, 20, 18, -22, 42, 50, -21, 9, 9, -20, -11, -11, 0, 11, -8, -10, 52, -20, 9, -19, 24, -26, -16, -21, 3, -20, 0, 48, 18, -3, -12, 13, -5, 22, -9, 8, 1, 36, 10, 3, -4, 0, 2, -33, 50, 43, -53, 33, 36, -9, 7, 19, -57, -1, 19, 2, 20, -16, 25, -21, -18, 5, 26, -7, 30, 26, 7, -14, 3, 41, -15, 32, -13, -8, 19, -7, 0, 4, -26, -11, 30, -4, 6, -5, -8, -20, -28, 0, 3, -40, 1, 30, 20, -4, -1, -1, -6, 30, -11, 11, 9, 23, 30, -20, -56, -44, -5, -3, -33, -33, -58, 14, 19, -24, 4, 2, -35, 0, -1, -6, -13, -9, -17, 14, 45, -1, 102, 12, -5, -26, 19, 5, -6, -4, -24, -6, -13, -2, 25, 0, 6, 13, -13, 0, 9, 20, -3, 15, 12, 45, -28, 14, -13, -43, -4, 7, -48, 12, 21, 17, -39, 11, 15, 27, 59, 13, -14, 11, 19, 11, -37, -40, 22, 25, -71, 45, -19, -50, 6, 15, 32, 44, 6, -10, 22, -29, 21, 85, 61, 5, 21, 0, 25, -35, 2, 13, 51, 3, -20, 20, -15, 30, 84, -9, -7, -58, 29, -15, -43, 28, -6, 15, -3, 40, 5, -42, -13, -1, -1, 38, -62, 5, -29, -14, -2, -1, -23, -10, -27, -11, -43, 10, 17, -13, 10, -35, -21, 50, 11, 29, -10, -42, -6, 3, -24, 0, -7, 5, -13, -39, 6, 63, 49, -6, 22, -13, -8, 2, 7, 7, 15, -36, -22, -19, 24, 30, 54, 0, -6, -16, 15, -26, 0, 1, 6, 11, -19, -10, 2, -14, -11, 19, -6, -50, -16, 4, -24, -4, 17, -12, -40, -18, 23, 23, -38, -1, -12, -6, -29, 23, -53, -5, 9, -11, 13, -9, 4, 9, 4, 38, -8, -6, -40, 13, -47, -47, -11, -5, 1, 28, -4, -27, 1, -30, 14, 30, 2, -30, -8, 18, -68, -4, 4, 10, -19, -22, -13, 6, 8, 11, 3, -1, -2, -28, -26, -7, 2, -1, -3, 20, 12, -10, -37, 5, 7, 33, 69, -3, 32, -5, 4, 16, -15, -8, 2, 13, -15, 0, 4, -21, 0, -38, 15, 64, -46, -10, -5, -1, -12, 4, -2, -3, -10, 20, 12, 11, 12, -3, 16, 54, -11, -17, 19, 7, 32, 10, 9, -20, -24, 4, 44, 4, 1, 18, -27, 12, -8, -17, 13, -46, -5, 35, 1, 22, -10, 32, -50, 25, 10, 50, 26, -17, 13, -3, 17, -38, -50, 2, 37, -14, -66, 38, -6, -46, -6, 12, -27, 14, -62, 6, -8, -2, -15, 12, 12, -6, -36, -14, 5, -19, 9, -5, -21, 16, -17, -12, 22, -16, 28, -6, 11, -8, -6, 25, 72, 17, -3, 25, 0, -22, -30, -4, -18, -29, -4, 36, -4, 22, 16, 46, -5, 27, -25, 17, -10, 42, -13, 22, 20, -52, -69, -14, 45, -19, -47, 64, 52, -59, 0, 43, -46, -29, -31, -6, 0, -17, 17, 22, -53, -10, 21, -21, -5, -21, 41, -11, -55, 9, -44, 1, 14, -10, 29, -7, -1, 11, -45, -12, 47, 9, -9, 22, 6, -7, 17, -12, -12, -21, -6, 32, 16, 4, -15, 11, -23, 45, 25, 32, -1, 10, 18, 17, 8, -54, -43, 7, 16, 9, -76, 55, 1, -44, -8, 24, -44, 25, -13, -8, -30, 2, -11, 19, -20, -7, 67, -34, 7, 14, 14, -2, -21, 44, -37, -20, 10, -23, 31, 1, 3, 8, -41, -1, -3, 9, -8, 4, 18, 22, -61, -13, -26, -17, -4, 22, -40, 16, -3, -1, -36, 10, 13, 31, 43, -15, 14, 15, -14, -28, -16, 2, -8, 33, -74, 22, -8, -29, 7, 10, 12, 44, -52, -8, 4, 7, -41, 52, 12, 0, -26, -14, 37, 3, -5, 4, 23, -7, -61, -11, 16, -15, 77, 4, 4, -18, -17, -39, -28, 9, -7, -16, 6, 6, 42, -45, 6, 10, -18, 39, -68, 1, -17, -40, -7, -10, 36, 39, 23, 4, 1, 1, 4, -7, 18, -40, -23, -14, 6, 17, -21, 0, -2, -12, -8, 20, 0, 0, -11, -8, -16, 21, 36, -9, -60, 17, -2, 2, -15, 19, 18, 2, 5, -27, 3, -17, 26, 11, 9, -6, -15, -14, -23, 5, 7, 19, 0, -24, -37, -30, -14, 12, 2, -39, -6, 6, -9, -10, -17, 1, -31, 13, 52, 29, -24, 13, -60, 24, 11, 15, 17, -6, -4, -58, 47, -9, 2, 0, 6, 60, 5, -3, 2, -10, -33, 0, 9, -2, -10, 23, 0, 10, -20, -16, 8, 16, -20, 9, 12, 5, -16, -7, 9, 16, -14, -10, -3, 26, 0, 6, 36, -12, 21, -23, -5, 8, 2, 50, -24, 7, -23, 0, -26, 9, 20, 9, 48, 0, -38, -20, -9, 3, 17, -29, -39, 30, -14, -23, -22, -29, 4, -26, 0, 33, -35, 8, 0, -22, -21, 25, 19, 3, -60, 15, -23, 36, -8, -14, 26, 20, -20, -3, 28, -26, -9, -6, 2, 40, -61, -10, 34, 18, -4, 10, 28, 5, -2, 3, 7, -38, 1, 75, -38, 25, -1, 24, -77, -3, 14, 19, 25, -38, -9, 21, 7, -30, -30, -43, -46, 46, -43, 0, -8, -29, -9, 3, -62, -3, -50, 1, -15, 6, -52, 8, 53, 2, 10, 38, 26, 8, -8, -23, -16, -9, -26, -28, 8, -14, -29, 9, -1, 29, -52, 34, 46, 19, -1, 7, -7, -14, -59, 6, 30, -21, 2, 20, 11, -18, -25, 9, -24, -8, 10, 34, -16, 0, 25, 9, 20, -21, -82, -11, 6, -30, -34, 17, 2, -54, 0, -5, -41, 24, -24, -5, -49, 18, -4, 8, 6, -8, 4, 24, 32, -6, -24, -39, -23, -37, -15, -45, 22, -7, -15, 4, 0, 13, -43, -29, 27, 9, 1, 5, 30, -13, -46, -40, -22, -25, -1, 38, 1, -2, -6, -5, -15, 17, 27, 32, -17, -17, 16, 15, -18, -18, -32, 3, 27, -43, -35, -14, 0, -40, 2, -12, -9, -7, -16, -12, -8, 25, -30, -36, -8, -10, 20, 10, -3, 10, -9, -9, -29, 15, 5, -52, 30, -50, -2, 0, 0, -17, 32, -40, 1, 13, 9, 0, 46, -22, -38, -45, 7, -14, -6, 18, -27, -2, -22, -3, -60, 40, 5, 34, 10, -12, 18, 0, -43, -20, -10, -8, -46, -1, -33, -48, 8, -4, 3, 23, -50, 10, -6, 4, 16, 33, -24, -6, 21, 6, -82, 15, -7, -57, 0, 14, 31, -8, -22, 2, 9, -9, -27, 0, -12, -6, -45, -12, -9, 7, 7, 14, 16, 0, 12, 8, 10, -12, -8, 24, -43, 6, -42, -1, -3, 5, 2, 2, 60, 17, 10, 12, -41, -28, 1, -12, -29, 45, -31, -30, 24, -33, 4, 6, 0, 40, 0, 0, 34, 0, 14, 6, 3, 1, -5, 8, 10, 34, -8, 25, 29, 11, -7, -6, -1, -22, 22, 0, 6, -44, -20, -38, -29, 17, -2, -4, -9, -24, 3, -8, -22, -1, 6, 12, 0, -17, 7, -4, 9, 9, 33, 26, 45, 33, -30, 14, 2, 31, 25, -31, 13, 65, 50, 0, 33, -18, -7, -3, 17, 64, -4, -6, 13, 3, 15, 23, 40, 12, 14, 31, -18, 76, -11, 7, 5, -51, -36, 23, -12, -35, 35, 0, 4, 0, -20, -31, 5, -23, -3, -18, 16, 11, -7, 19, 11, 7, -9, -7, -25, 0, -46, -11, -19, -1, 19, 15, 39, 26, -10, 11, -26, 17, -7, -53, -82, -15, 8, 22, 12, -15, -12, 10, 33, 13, -19, -6, 23, -3, -11, 36, 60, 9, -22, 18, 52, 56, 15, 0, 34, -22, -23, 27, -18, -54, -11, 3, -1, 28, -30, 18, 2, 0, 0, -7, 51, 13, -20, 29, 48, -18, 2, 17, 25, 5, -28, -34, -40, -1, 54, 26, -36, 20, 1, -7, -15, 28, 4, -15, -14, 3, -1, 15, 5, 15, -9, 14, 30, -3, -8, 4, 5, 13, -18, 26, 35, 7, -46, 26, -10, 36, -10, -12, 10, -33, 0, -3, -1, -13, -18, -9, -13, 17, 3, 29, 9, 41, 3, 27, 37, -28, -10, 30, 9, -16, 12, -2, 22, 10, -20, -23, -26, 34, 48, 3, -41, 13, 8, -15, -11, 14, -13, -12, 17, -2, -30, 2, 16, 2, 2, 8, 26, 23, 20, -5, -4, 14, -14, 4, 11, 5, -23, -6, 36, -33, 16, -35, 23, -6, 29, 9, 7, 40, -15, 2, -10, 40, 32, 1, 28, 1, -9, 13, 24, -22, -29, 26, -9, -1, -15, -27, -12, -34, 0, 4, -38, 1, 8, 3, -32, 59, 2, -29, 4, 20, -20, 35, -4, -33, 19, 5, 2, 12, -2, 7, 16, 11, -13, -1, -12, 4, 0, -14, 5, -4, 9, -18, -4, -3, 25, -32, -10, 19, 17, 8, 16, -58, -10, 8, -5, 4, 7, -1, 14, 38, -3, 9, 22, -71, -20, -13, -25, -9, -1, 18, -1, -22, -31, 7, 0, -7, -1, 9, 0, -2, 19, -1, -3, -51, -19, -13, -75, -10, 7, -6, 7, -16, -6, 11, -12, 18, -29, 6, 12, 34, 23, -48, 35, 10, -42, -22, -37, -57, 8, -42, 16, 31, 8, 24, 16, -22, -1, -4, -12, 11, 2, -31, -6, -14, -5, -1, 11, -76, 30, -18, 38, -11, 11, -2, -26, -20, -8, -13, 39, 44, -37, 4, 50, 6, -3, 8, 4, -19, 17, 5, -61, 11, -17, 7, 41, -16, 8, -2, 0, -19, 0, -3, 6, 45, 68, -86, -21, -6, 34, 23, 24, 57, 11, -20, 13, 48, -53, 1, 11, -5, -27, -6, -4, -10, -33, -33, -36, -26, 6, -9, 2, -92, -5, -15, 17, -27, 2, 6, 11, -9, -50, -26, -5, -35, 12, 26, 17, 8, -47, 28, -58, 10, 8, -72, 20, 15, 19, -59, 23, -19, 6, -10, -6, -29, 14, -11, 20, 26, -10, 46, 49, -5, 21, 29, 24, 52, -33, -10, 10, -77, -34, 28, 6, -12, 11, -11, 3, 2, -59, -30, -8, -27, -6, 12, 14, 1, -13, 30, 30, -7, 2, -48, 2, -14, -46, -13, -24, 23, 19, 22, -9, 18, -13, 16, -60, 63, 4, -37, -18, 13, 10, -32, 19, 6, 4, 15, 31, 0, 10, -4, 20, 14, -1, 51, 40, 5, -18, -2, 46, 25, 0, -6, 8, -61, -25, 28, -17, 7, 9, 0, -4, 29, -3, 49, 13, -4, -10, 7, 20, -32, 9, 34, 9, -1, -9, -6, 8, 20, -29, -3, -2, -9, 21, 0, 0, 17, -10, 31, -55, 15, 6, -23, -23, 0, 9, 41, 12, -18, -4, 2, 21, 9, 3, -2, 23, 5, -14, 15, 49, -5, -8, -9, -7, 31, 13, -3, 26, -51, -5, 40, -26, 12, 10, 1, 0, 28, -10, 4, 13, 9, 2, 28, 1, -38, 9, 44, 21, -12, -1, -9, 27, 26, -29, -8, 0, 18, 11, -19, -30, 3, -12, 30, -16, 12, -11, -12, 31, -29, -21, 44, 16, -9, -7, 17, -12, -29, 16, -8, 22, 0, -11, 1, -22, 13, 14, -21, 15, -5, 5, 11, 51, -25, -7, 36, -25, 14, -41, -11, -11, 27, 19, 7, -12, 7, 4, 38, 17, -13, 5, 18, -21, -11, 4, -16, 17, 29, -22, 0, 10, 4, 5, -15, -16, -19, 8, -3, -14, 40, -15, -1, -13, -17, -2, 15, 1, -23, 1, 13, 6, -14, -6, 3, 15, 17, 37, -18, 52, -2, 17, -17, 9, 11, -2, 9, 54, 32, -5, 8, -11, 35, 16, -3, -3, 13, 0, 12, -18, -17, -9, 21, 8, -71, -31, 16, 12, 25, 1, -76, 5, -13, -13, -21, 1, 28, -16, -6, 6, -9, -15, 29, -34, 10, 12, 21, -25, -16, 15, -17, -1, 4, 0, 0, -26, 3, -16, 2, 17, 36, 28, -38, -8, -2, 38, -23, 0, 8, -4, -10, 11, 29, 8, 11, -6, 2, -55, 6, 0, 1, -13, -11, -39, 17, -10, 2, 7, -25, 14, 25, 36, 30, -6, -59, -41, -25, -64, -18, 8, 12, 0, 24, 1, -1, -32, 0, 34, 15, 42, 3, 7, 31, -11, -38, 18, -15, 5, -6, -10, -10, -16, -8, 9, 23, 31, -70, -103, 0, 15, -3, -30, 46, 18, -32, 27, 93, -35, -1, 14, 21, -27,
    -- layer=2 filter=0 channel=1
    -6, 2, -23, 60, 33, -38, 46, 5, -18, 0, -47, 58, -48, -8, 7, 2, -47, 19, -21, -9, -33, 4, 18, -30, 25, 7, -3, 8, -21, 7, 47, -5, 14, -2, -17, 10, 15, 10, 15, 4, -15, 46, -4, 29, 6, -5, 8, -12, 51, -2, 1, 30, 1, 60, 30, -26, 10, 0, 21, 37, 5, 16, -10, 39, -3, 0, 7, 3, 8, -5, 0, 9, -3, 3, 0, -18, -20, 0, 14, -11, -39, -33, -5, 25, -32, 12, -26, -23, -5, -33, -13, -44, -12, -1, -10, 33, -17, -24, 10, -1, -1, 13, 18, 3, -12, 40, 1, 15, -7, -5, -28, 7, 42, 3, -8, -7, 3, 3, 62, -26, 1, -11, -35, 22, 32, 10, -25, -16, -3, -15, -9, 2, 28, 7, 7, -1, -4, 10, 9, 21, -16, 0, 10, 6, -8, -19, -8, -20, -2, 6, -15, 39, 29, 0, -1, 18, 7, 24, 41, -6, -6, -13, -26, 2, -29, 9, -8, 3, 1, 41, -1, -4, -10, 6, -12, 22, 24, 27, -1, -20, 10, 32, 24, -10, -5, 6, -30, 7, 1, -23, 1, 35, 1, -11, -20, 3, 1, 0, 23, 10, -3, 13, 16, 16, -18, -8, -3, -6, 21, 0, 7, -24, 10, -32, 12, 4, -21, -6, -7, 11, -4, 7, 12, 6, -1, -44, -3, 8, 9, -20, -14, 11, 5, -27, 12, 2, 6, -12, -14, -25, 39, 38, -9, 14, 11, 35, -11, -10, -6, -5, -5, 10, -10, 18, -11, 19, 0, -8, -28, 15, 14, 6, -2, 8, -5, 29, -14, 1, 10, 10, 3, 3, -49, 7, 1, 19, 20, 4, 19, -11, 6, 15, -23, 22, -12, -41, 22, -2, 45, -58, -31, 13, 51, 10, 5, 0, -9, 6, 50, -9, 0, -15, 7, 9, -7, -48, -6, 28, 22, 21, 1, -14, -13, -4, 9, 26, -19, 16, 0, 9, -1, -10, -43, 19, 30, -15, -13, 9, -11, 21, 15, -30, -5, -11, -24, -6, -5, -60, 0, 27, 7, 12, -11, -19, 17, 8, -13, -15, -5, -38, -24, 2, -8, -3, 4, 5, 26, 8, -4, -7, -6, 26, -3, 3, -7, 0, -11, 8, 28, -50, -11, 13, 4, -12, 39, -4, -31, -15, 21, 29, -9, -1, -36, 2, 0, 8, -43, 15, -5, -25, 3, -1, -15, -12, 15, 20, 1, -18, -8, -9, 0, 23, 16, 13, -35, 34, -35, -16, 1, 56, -35, -8, -12, 34, 19, 22, -10, -16, -21, 28, 19, 20, 13, 11, -12, 27, 51, 5, 2, 10, 2, 24, 21, 1, 9, -10, 1, 26, 27, -29, -23, -11, 0, 11, 15, -10, -39, 4, -9, 1, -21, -33, -6, -18, 14, 1, -8, 3, -17, 10, -5, -1, 15, 7, -43, 1, -12, -34, -41, -33, -19, -19, 1, 11, 9, -21, -2, -9, -11, 1, -37, -27, 34, -12, -30, 6, 18, 8, -5, -29, 25, 24, 4, 1, 0, -6, 11, -3, 2, -7, -1, 4, 26, -5, 11, 11, 7, -20, 1, -7, -7, 26, -10, -1, 24, -30, 1, -7, 10, -4, 8, 4, -7, -3, -1, 11, 1, -3, 31, -7, 4, -32, -18, 7, -18, 5, 0, 18, -14, -34, 1, 15, -1, 4, -9, -4, 1, 2, -24, -12, -6, -9, 2, 0, 7, 1, 0, -21, 2, -6, 27, -31, -11, 18, -20, 16, 35, 7, -7, 0, -25, 25, -4, -6, 18, -8, 10, 0, 13, -36, -11, 25, 17, -5, 1, 0, 39, 21, -3, 6, -5, -7, 20, 7, 10, -1, 0, -37, -10, 9, -39, 21, -16, 11, 18, -5, -15, -29, -34, -43, 0, -17, -23, -13, -15, 2, -2, -24, 8, -24, 6, 19, -22, 22, 15, 41, -3, 6, -14, -47, 8, 11, -30, -21, -44, -3, 10, -12, -11, 7, -11, -14, -16, -4, 21, 22, 31, -7, 22, 7, 16, 4, -24, -15, -8, 3, -3, -4, 38, -21, 32, -29, 47, 17, -10, 11, -6, 16, 7, -5, 15, -35, -27, -34, -15, -19, -44, -43, -47, 0, 0, 15, 24, -58, -2, -25, 15, 41, 0, -37, -9, -71, -39, -3, -3, 16, -86, -53, -37, -38, -15, -16, 7, -22, 5, -6, 0, -2, 2, 16, 29, 8, 24, 1, 0, 6, -14, -11, -4, 3, 24, 8, 44, 11, 12, 11, 21, -7, 11, 12, -2, 5, 17, 17, -9, -17, 5, -75, 0, -25, 27, -24, -17, 0, -8, -12, -15, -22, -4, -19, 14, -9, -23, -21, 4, -21, 3, -39, 34, 26, -59, 11, -13, 7, 12, 20, 16, -11, -8, 8, 22, 0, 37, 2, -12, -7, 2, 20, 4, -21, 17, 4, -7, -7, -12, -2, 12, -3, 35, -22, 41, -5, 2, -14, 3, 17, -20, 30, -11, 2, -7, -4, -33, -4, -8, -5, 0, 0, -3, -29, -37, -11, -11, 15, 27, 22, 13, -35, 5, 2, 20, -4, 59, 0, -4, 25, 1, 24, 17, 16, -4, -26, 1, -5, 8, -28, 7, -1, 25, -1, 9, -9, 25, 34, -7, 10, 32, -11, -2, -13, 10, 4, -29, 9, -5, -14, 15, -12, -28, 9, -6, 41, 23, 10, -34, -16, -36, 18, -54, -5, 16, -5, -15, -28, 25, 0, 8, -11, -2, 21, 18, -16, -1, -26, 15, -1, -13, -25, -20, -13, 8, 31, 10, 29, -17, 13, 8, -17, 1, -39, -18, 4, 5, -7, -8, -1, -5, 10, 1, 12, 31, 4, 6, 5, -28, -39, -23, -25, -14, 11, -12, -54, -7, -19, 8, -14, 8, 23, -34, -7, -12, 15, -74, -22, -5, 8, -25, -26, 6, 5, 5, -4, 8, -9, 31, 31, -10, 33, 6, -54, -30, 9, 34, 8, 9, 13, 0, 9, 17, 8, 1, -17, 15, -48, 25, 17, 2, -1, 4, -34, -16, -9, 21, 26, 23, 5, -7, 11, 18, -6, 14, -36, -25, -10, -37, 48, -12, 17, 17, -6, 17, -2, 0, -60, 7, -39, -43, -40, -10, -11, -18, -22, 3, 20, 4, 11, 6, -44, 17, -13, -3, -20, 1, 5, -9, 11, 20, 12, -3, 6, 6, 18, 62, 3, -3, -3, 16, -90, 0, 25, 13, -8, 8, -43, -1, -4, -2, -7, -1, 3, 7, 18, 41, -14, 26, -73, 6, -14, 14, 39, -12, 4, 45, 0, -8, -68, -45, -36, 3, -78, -10, -5, -36, -1, 19, -26, 10, -21, 0, 29, -7, -28, -28, -26, 0, 36, -12, -4, 15, 41, -6, -18, 17, -22, -1, -7, 12, 2, 5, -1, 35, -48, -2, 48, -14, -5, 37, -49, 22, -24, -23, 12, -16, 0, 9, 41, 45, -12, 44, -81, 31, -2, -7, 44, -70, 38, 19, 20, -40, -68, 7, -30, -62, -78, -80, -37, -55, -9, 10, -60, -6, -38, -9, 0, -5, -46, -65, 11, 0, 0, -24, -32, 41, 21, -16, -34, 0, -29, 10, -23, 64, 43, -1, 6, -30, -16, -1, 19, 13, -6, 24, -32, -15, -10, 9, 39, -13, 0, 13, 18, 48, -17, 38, -84, 77, 25, -14, 9, -67, 30, -7, 15, -61, -37, -42, -35, 16, -44, -40, -12, -31, 1, -7, -13, 30, -33, -12, 14, 17, -15, -36, -83, 4, -58, -28, 7, 42, 39, -6, -12, 11, -31, 11, 0, 47, 27, 0, -6, 31, -62, 26, -7, 24, -8, 17, -24, 0, 3, 14, 8, 1, 7, 20, 32, 44, -13, 9, -25, 26, 34, -21, -12, -35, 35, -3, 3, -32, 8, -18, -24, -8, 0, -65, -23, 5, -9, -20, 4, -4, -13, 4, 0, 7, -9, -15, 16, 8, -23, 3, -15, -84, 16, 11, 2, 32, 6, -3, 21, -58, 0, -10, 3, -13, -32, 0, -52, 22, -8, -22, 29, -19, -9, -8, 49, 9, -12, -21, 14, -3, -25, -55, -32, -43, -20, -10, -20, -48, -2, -3, 13, -62, 19, -6, -44, -72, 6, -41, -14, -8, 3, -16, -42, 24, 4, -10, 20, 17, 10, -27, -5, -7, -67, 3, -33, -19, -3, 28, -11, 37, 45, 16, 6, -3, -2, 1, -9, -7, -17, 7, -12, -10, -6, -34, -14, 22, -31, 0, -12, 15, 8, 10, 20, -36, 7, -25, 28, -4, 0, 21, -19, -37, -24, -12, -2, 12, 19, -7, -25, -17, 10, -30, -33, 6, -3, -31, -1, -24, -7, 9, -25, 26, 4, 5, 44, -8, -2, -19, -6, -24, -23, -5, 11, 7, -14, -1, 0, -5, 32, 0, -11, -4, -66, -39, 18, 5, 8, 19, 9, -27, -24, -51, 37, -11, 8, 7, -12, -9, -15, 22, -1, 28, -6, 21, 14, -28, 6, 17, -8, -20, 6, -9, 28, 28, -42, -73, -20, -3, 11, -25, -30, -2, -16, 0, 19, 47, -8, -22, 12, 9, 43, -1, -14, 55, 4, 78, 4, 33, -14, 8, -3, 34, -26, 9, -8, 29, -105, -40, 0, 26, 5, 11, -11, -16, -45, -34, 10, -19, 0, 17, 39, 33, -26, 24, -8, 32, 15, 11, 43, -51, 47, 43, 3, -65, -3, -33, 31, -33, -52, -21, 11, -36, 9, 16, -43, -5, -38, 2, 35, 32, -29, 21, 11, -4, 46, 8, -11, 3, 38, 24, -38, 39, -38, 53, 8, 2, 2, 0, 9, 1, -52, -33, 28, 13, -12, 49, -20, 41, -8, -38, 35, -29, -6, 22, 38, 52, 18, 38, -53, 18, 0, 1, 25, -59, 81, 31, -30, -45, -22, 1, -8, 4, -71, -75, -13, -53, -7, 0, -92, 26, -23, -5, 19, 24, 10, -4, 13, -2, -32, 12, -28, -40, 0, 34, -23, 43, -59, -6, 13, 79, 58, -4, -7, 8, -102, -21, 43, -12, -7, 32, -14, 14, -33, -18, 25, -31, -11, 19, 8, 40, -20, 12, -53, 32, 2, 4, 25, -79, 81, 12, -45, -103, -1, -69, 0, 2, -44, -109, -32, -23, 9, -2, -73, -4, -18, 5, 17, 21, 5, -11, -41, 3, -119, -10, -15, -35, 26, 52, -2, 24, -30, -19, -15, -8, 48, -9, 9, 27, -70, -9, -1, 0, 4, 33, 3, -14, 9, 31, 7, 0, -4, 27, -10, 1, -31, 21, -62, 18, 17, -27, -28, -1, 39, 0, -25, -87, 28, -44, 24, -26, -20, -50, -31, -11, -3, 8, -100, 0, -15, -3, 5, 0, 29, -19, -38, 2, -62, -35, -36, -62, 58, 53, 39, -5, 11, 11, -4, 27, 17, 0, -10, -7, 5, 3, -26, 6, -9, -24, 17, 5, 3, 22, 37, -18, -4, -25, 32, -32, 12, -46, -19, -54, 15, 7, -48, -22, 7, -4, 2, -54, 1, 11, -37, -24, -15, -33, -36, 1, -1, -1, -34, -6, 10, 5, 23, 27, 1, 30, 30, 6, -38, -9, -9, -71, 4, -11, 3, 37, 20, 26, 15, -34, 10, 5, 6, 4, -32, 10, -17, 11, -1, -7, -46, -12, -18, 22, -47, -34, -8, 9, 18, -3, -25, -8, 16, -93, -9, 2, -70, -50, -4, -16, 38, -72, 0, -25, -63, -24, 31, -18, -80, -3, 6, -10, 7, -4, 20, -9, -5, 30, -2, 0, 45, -3, -49, -68, -21, -84, -78, -24, -24, 27, 38, 9, -1, -10, -71, 1, 5, -22, -5, -10, -18, 20, 0, 47, -16, -14, -27, -50, -75, -7, -3, 21, 44, 9, -14, 15, 23, 89, -12, 23, 10, -51, 62, 25, -15, -43, -19, 37, -62, -10, -21, -46, -1, -44, 2, 42, -22, 8, -37, 9, -4, 57, 0, -19, -36, 3, -23, -36, -39, 42, 16, 39, -28, 36, -23, 3, 27, -12, 4, -11, -13, -5, -35, 2, 33, -3, -9, 0, 11, -36, -28, -23, -42, -23, 4, -24, 49, 7, -12, 9, 37, 16, 13, -12, -17, -20, 24, 11, 20, -1, -27, -33, 18, -4, 16, 62, -41, -27, 4, 21, -3, -31, -45, -8, 46, 5, 24, 18, 2, 4, -29, -66, -2, 50, 15, 32, 45, 9, -54, 4, 3, -5, -1, -1, -14, 34, 5, -22, 53, 13, 12, 19, 37, 10, 9, 28, -23, -25, 2, 62, 53, 30, -3, 41, 40, -19, 17, -10, 43, -67, 29, 15, 17, -47, -4, 5, -30, -18, 2, 9, -1, -48, 8, -2, -43, -7, -48, -1, 14, 19, 8, 5, 33, 9, -24, -30, -39, -5, 31, 23, 62, 12, -57, -6, -3, 34, 56, -9, 11, 19, -3, -27, 39, 17, -3, 36, 39, 6, 23, 56, 0, -23, -11, -3, 34, 14, 22, 21, 34, 21, 15, -10, 14, -94, 31, 27, 52, -75, -13, -15, -1, -1, -10, 44, -46, -30, 4, 18, -53, 12, -23, -1, 5, 3, 37, 0, -65, 3, -33, -13, -13, 67, 64, 44, 59, 50, -36, -29, 4, 55, 1, 4, 1, 19, -60, -9, 28, -8, -11, 40, 20, 12, -42, 11, -32, -11, -9, -8, 46, 21, -64, 13, -8, -29, 27, 13, 3, -26, 17, 48, 49, -17, -22, -39, 54, -10, -16, 10, -77, -29, -1, 28, 15, 8, -50, -1, 36, 6, -3, 42, -16, -8, -50, -30, -17, 43, 12, 43, 21, 13, -31, 1, -6, 36, 24, 6, -4, -7, -60, 4, -49, 35, 2, 8, -64, 5, -32, -9, -35, -11, 3, 34, -17, -15, 8, -34, -29, -60, 10, 15, -89, -60, -25, -16, -17, 2, -24, -39, -30, -27, -31, -45, -102, -31, -7, -5, -19, 4, -36, -5, 2, -4, -52, 68, 28, -1, -55, -64, -74, -44, 6, -19, -15, 21, -2, -23, 23, -30, 2, 8, -7, -24, -47, -43, -3, 12, -8, -14, 4, 8, -56, 36, 0, -24, 8, -20, 2, -6, -38, -31, 19, -57, -59, -10, -86, -43, -14, 0, -3, -62, -40, -2, -49, -26, 24, -1, -14, 0, 8, -11, -40, -41, -7, -7, -18, 3, -2, 0, -34, 2, -26, 15, -35, -114, -37, -41, -16, 7, 53, -40, 3, 21, -102, 1, 11, 28, 40, 8, 6, 71, -9, 26, -7, -56, 12, -25, -30, -40, -10, 50, 38, 18, -57, 1, 18, -17, -1, 44, -4, -86, 44, -19, 19, -85, -20, 31, -5, 19, -63, -9, 21, -37, -2, -16, -7, -17, -12, 9, -14, 40, 18, 5, -59, -1, -8, -14, 20, -67, -10, 24, -20, 45, 19, -46, 47, -8, -8, 5, -8, 46, 10, 21, 21, 34, 0, 2, 29, -47, 22, -19, -61, -48, -7, 42, 18, 7, 23, -16, 47, -31, -8, 41, 16, -91, 56, 0, 67, -47, -39, 21, 1, -34, -51, 1, -22, -15, 0, -35, -8, -40, -34, -4, -27, 15, 33, -16, -54, -8, -17, -20, 7, -15, -26, 9, 48, 9, -19, -15, 14, 0, -3, 7, -4, 29, 6, 32, 8, 9, 1, 11, 40, -11, 17, 2, 3, -17, -17, 63, 24, 19, -3, -21, 80, -48, 16, 10, 11, -60, 17, -4, 60, -55, -20, -36, -52, -5, 5, 85, -44, -24, -8, -1, 11, -46, -16, 10, -33, 14, -7, 6, -55, -1, -12, 21, -10, 52, -12, 28, 62, -11, -15, -11, 4, 16, 18, 2, 9, 61, -8, 30, -18, 12, -9, 27, 40, 0, 21, -18, -12, -4, -10, 39, 61, 5, -11, -13, 53, -9, 29, 37, 12, -50, 19, 10, 59, -20, -8, -38, -20, 17, -10, -6, -57, -13, 7, 15, -10, -18, 12, -11, 10, 25, -11, 30, 10, 4, -8, -11, 13, 10, -10, 36, 98, -26, -12, -5, 4, 66, 6, 11, -3, 28, -71, 29, -19, 24, 4, 11, -5, 23, -24, -27, 16, -11, 12, 6, 9, -16, -15, -24, 24, -5, 23, 22, -23, -13, 34, 22, 15, 5, -29, -51, -17, 11, -1, -11, -46, -59, 0, 2, 15, -3, 5, -12, 29, 21, -37, 13, 21, -11, -21, -30, 18, -45, -20, 46, 53, -23, -53, -38, 31, 44, 49, -5, -6, 9, -28, 22, -50, 26, -1, 14, -5, 16, -42, -58, -17, -22, 8, -15, -14, -11, -2, -53, -30, -39, -2, 10, -132, 4, -5, -21, 15, 7, -38, -84, -3, -47, 5, -29, -20, -54, -9, 0, -3, 11, 15, -1, -25, -1, -19, 59, 16, 2, 2, -20, -81, -38, -22, -1, -1, -41, -16, -41, 31, 36, 22, 0, -14, -15, -20, -22, -11, 1, 1, -26, 93, 0, -31, 61, 26, 0, 3, -42, 1, -27, -63, -21, 34, -51, -34, -70, -13, 63, 0, -25, 10, -56, -33, 32, -62, 17, 36, -28, 23, -21, -7, -21, -36, -83, 3, 2, 7, -27, 34, -31, -16, -14, -17, 58, 22, -43, -22, -42, -1, 37, 33, -7, -54, 63, -119, -9, -5, -30, -9, -30, -23, 81, -9, 4, 45, 1, 22, -17, 6, -46, 9, 72, -15, 25, -36, -21, -7, -37, -36, -9, 16, 61, 24, -39, 64, -69, -17, 18, -42, 30, -58, -27, 39, -33, 0, -16, -85, 14, -4, -3, -28, 17, -5, -74, 3, 4, 0, 17, 18, -6, 14, -28, 8, 53, 18, -20, 32, 50, -6, -7, 0, 28, -25, 19, -18, 90, -5, 3, 71, -21, -15, -33, 41, -46, -3, 38, -2, 46, -18, -2, 14, -2, -9, 27, 21, 36, 14, -11, 62, -12, -26, 26, -18, -83, -60, -15, 40, -22, -2, -47, -28, 16, -5, 10, -64, 50, -29, -10, -105, -9, -14, 35, 12, -9, 9, -49, 15, 0, 8, -56, 69, 91, 7, 5, -19, -2, 0, 26, -23, 54, -9, 12, 64, -39, 10, -49, 0, -43, 1, 52, -3, 30, -19, -3, -15, -22, 11, 68, 10, 32, 17, -12, 53, 3, -27, 6, 2, 29, -37, 0, 49, -62, -4, -29, -13, 4, -16, 5, -17, 33, -22, -22, -30, -5, 17, 8, -8, 26, 2, -22, 38, -5, 2, -49, 21, 68, 6, -1, 6, 26, -42, 49, -24, 42, 6, 1, 19, -16, -8, -32, -5, -45, 0, 8, 0, 16, -18, -28, 7, -10, 28, 34, 31, -12, 39, -10, 61, -5, -31, -31, 3, -35, -58, -6, -14, -48, -7, -20, -25, 7, -15, 6, -8, -7, -24, 6, -4, 1, 20, 13, -14, 11, 25, -1, 51, -17, -20, -20, 25, 40, 29, -7, 0, -4, -64, -23, -2, 31, 8, -18, 5, 9, 16, -40, 9, -47, -5, 60, 13, 26, -39, -11, -30, -23, 26, 23, 2, 10, 18, -27, 14, 6, -42, -88, 19, -4, -42, -72, 21, -61, 1, -5, -20, 5, 24, -4, -5, -48, 10, 36, 37, -5, -1, 22, -6, 3, 15, 7, 21, -32, -25, -11, 4, 62, 32, -6, -7, -24, 0, 51, -8, 49, -2, 17, 57, -42, -20, -24, -21, -16, -12, -38, 24, -23, -14, -46, -35, -48, -12, -28, -76, 55, 31, -37, -18, 42, -43, -35, 18, 20, -16, -1, 53, -41, -9, 4, 14, -20, 27, -9, -7, -49, -8, 42, 70, 0, -39, 3, 25, -68, 1, -37, -10, -103, -9, -58, -1, 54, 24,
    -- layer=2 filter=0 channel=2
    -4, -21, 28, 9, 30, 11, -17, 5, 6, -13, 4, 9, 18, -29, 15, -6, 44, -33, 8, -3, -6, 17, 9, 0, -2, -23, -3, -40, -1, -23, 14, 15, -13, -34, 5, 25, -20, 0, 22, -11, -11, -22, -23, 0, -9, 3, -32, -31, 45, -10, 3, 34, -1, -51, -14, -4, -29, 0, -49, 32, 3, -14, -25, -47, -2, 3, 2, -40, 17, 3, 1, 3, 2, -3, 21, -13, 19, -22, 27, 6, 18, -37, -12, -7, 9, -24, 32, 32, 22, -14, -22, -4, -26, -66, 29, 12, 0, 2, -43, 31, 6, -6, 15, 1, -13, -19, 40, 1, 2, -12, 0, -15, -9, 0, -6, 0, -2, -58, -11, -9, 15, -9, -27, 23, -8, 10, -27, 0, 8, -18, -9, -25, -1, 19, -16, -7, -15, -8, 17, -20, 19, -26, -3, 8, 19, -2, -22, 0, 16, -39, 1, 35, 4, -23, 35, -7, 7, -38, 18, -9, -9, -21, -14, 10, -6, -17, 16, 1, 5, -14, 47, -9, 9, 13, -29, -4, -9, 29, 0, 5, -16, -48, -10, 0, -9, -22, 3, 15, -17, -13, -8, 14, 10, -12, 5, -16, -26, -8, -9, 7, -19, 30, 39, -13, 1, -7, -19, 5, -10, 4, -28, 0, 0, -31, 23, 0, -20, -25, 46, -5, -2, -91, 9, -8, -31, -30, -13, 11, -15, 3, 9, -6, 14, -4, -1, -1, -7, -13, -32, 12, -1, -2, 1, 14, -6, -14, -2, -4, 6, -25, -6, -12, 0, -1, -24, -11, 7, -7, -1, -48, -14, -2, 4, 2, -8, -6, -26, -7, -1, 0, 14, -1, -22, -11, -27, 0, 6, -18, 27, -46, -9, -21, 18, -12, 22, -75, 13, -21, 2, -28, 7, -7, -39, 11, 8, -10, 2, -47, 47, 6, -8, 4, 26, -1, -71, 10, 2, 84, 4, -47, 1, 10, -45, -31, 19, 34, 2, -9, -16, 0, -7, -21, 19, -25, 10, 5, 14, -10, 12, -3, -18, -50, 22, -17, 22, -5, 45, 4, -19, -1, 1, 6, 22, -32, -29, -5, 6, 12, -9, -21, 0, -14, 9, -10, 2, -18, -41, -9, 27, 8, -4, -10, 8, -8, -7, -32, 6, 1, -51, 25, 10, 46, -5, -35, -21, 21, -50, -6, 22, 59, -8, 0, -19, -29, 11, -15, 34, -5, -2, 7, 11, 1, 12, 11, -9, -39, 27, -34, 30, -5, 39, -4, 3, 8, -16, 3, 18, -27, -27, 0, 0, -36, 12, -31, 56, -1, -22, -23, -21, -10, 13, -23, 31, -11, -13, -37, 0, -3, -8, 2, -41, 0, -41, -45, 7, 4, -14, -28, -37, 3, -12, 0, 27, 17, -16, 2, -1, -20, -7, -13, 7, 36, 11, 2, 11, -7, -4, -14, -39, 8, 18, -38, -14, -4, -43, -54, 1, 12, 1, 2, 55, -2, -44, 4, 14, -31, -6, -51, 33, 19, 20, -4, -30, 10, -25, 0, 15, 7, 15, 37, -11, -12, 7, 11, -32, 7, -21, -16, -6, 32, -20, -23, 25, 24, 0, 3, -38, -21, -5, -28, 11, -27, 3, 3, -25, -1, -8, 5, 37, -5, 28, 30, 5, -7, -4, 6, 0, -9, 16, -23, 37, -6, 11, -27, -21, -24, -32, -3, 0, -40, 8, -18, 9, -9, -5, -13, -37, 12, 8, 7, -8, -4, 2, -9, 43, -21, -7, 0, -18, -13, -16, 43, -12, -22, -5, -18, -3, 9, 5, -6, -14, -4, -2, -15, -7, -16, 8, -12, -16, -20, 13, 11, 39, 6, -20, 18, 63, -26, -7, 25, -13, -10, 3, -22, -7, 5, 3, -31, 28, 13, 14, 22, 32, -28, -5, 3, 38, -4, -23, 7, 7, 9, 36, 42, -4, -5, 1, -21, 15, -2, -6, 30, -2, 4, 14, 37, 6, 27, 21, 0, -3, 5, -8, -18, -8, -28, 4, -17, 37, -13, 7, -12, -15, -16, -16, -13, 1, -4, -29, -20, 28, -26, -5, 9, -30, 7, 18, -18, -26, 32, -12, -10, 15, -1, 2, 42, 19, -21, -22, -35, -25, 9, -4, 12, -33, 1, 12, -3, 0, 4, -25, 2, 21, 1, -9, 1, 8, -8, -13, 21, -6, -3, -31, -5, -13, -3, -1, -15, 15, -12, 8, -18, -21, -3, 0, -3, -18, 15, -13, -1, 13, 0, -14, 0, 40, 22, -11, 14, -27, -6, -1, -23, -11, 21, 6, -42, -15, -17, 4, -11, 11, -61, -9, -46, 6, -12, 16, 15, -13, -12, 23, 36, 7, 2, -21, -6, 19, -4, 1, 27, 4, -8, -3, 10, -5, -5, -17, -20, -18, -9, 0, -40, 49, 3, 15, 2, 29, -17, 2, -6, 16, -5, 15, 0, -2, -5, 19, 7, -1, 48, 11, 14, 1, -9, 22, -26, 16, 34, -21, 18, -4, -14, -21, 19, -10, -5, -4, -28, 33, 4, -10, -5, -2, -12, -8, 12, -4, 6, -25, 24, -2, 10, -2, -16, -11, 0, -21, -6, 1, -12, 6, -6, 0, 5, 30, -4, 10, 31, -26, -22, 24, -27, 0, -3, 9, -1, 3, -7, -3, 3, 5, 6, 3, -25, 7, -8, 30, -9, 6, -31, -9, -1, -25, 3, 15, 13, 3, -8, -10, -29, -1, 10, 44, 12, -25, 8, -16, -7, -2, 6, 31, -1, 8, -22, -32, -2, 0, -12, -29, 11, -5, 0, 4, 15, 8, -13, -27, 12, 7, 24, -24, 0, -9, -31, -8, -8, 8, -2, -9, 13, -7, -6, -35, -3, 32, 49, -27, -7, 13, -10, -7, -10, -2, -37, -14, 31, -7, 1, 59, 7, -36, 48, 23, -66, 15, -78, 28, 21, 29, 9, -10, 15, 32, 14, 15, -12, 0, -23, -19, 3, 7, -3, -17, 23, -25, 12, 0, 38, 6, 20, -3, -2, 4, 34, -32, -42, 15, -60, 15, -52, 2, -16, 7, 44, -1, 29, 21, -5, 39, 35, 24, -13, 11, 12, -29, 7, 2, -18, 6, -15, -6, 17, 12, 29, -1, 33, 31, -31, 9, -12, 5, -18, 16, -13, 8, -6, 51, 31, -13, 5, 17, 13, 2, 6, 0, 10, -13, 8, -20, 31, 9, -24, 17, -29, 33, 20, 5, 12, -7, -25, 9, 0, -3, -43, -7, -9, 13, 30, 0, 24, -16, -2, -41, 47, 51, -26, -7, 24, -12, -8, -4, 0, 0, 42, 11, -5, -17, 35, -1, 13, 45, -42, -33, -54, 44, 22, 0, -14, -24, -1, 41, 16, 9, 8, -22, -13, -26, 9, -10, 16, 10, 12, 25, 35, -5, -36, 37, 21, -54, -34, -10, 4, -17, -39, -19, -17, 21, 20, -12, -6, 5, 40, -32, -23, -7, 0, -35, -31, 69, -17, 24, -26, -4, -1, -9, -15, -21, 70, -16, 0, -6, 15, 21, -13, 9, 10, -22, -59, 11, 8, 36, -27, -6, 31, 32, -28, 5, -3, -59, -18, 30, -4, 3, -2, 22, -5, -12, 62, 5, -78, -7, -37, -76, -22, 4, -18, -10, -24, -8, 14, 21, 11, 8, -19, 31, 57, -29, -6, 35, 3, -10, -18, 24, -21, 13, 37, -28, 4, -34, -23, 9, 69, -5, -3, -10, -55, 9, 48, 22, -32, 4, -44, -18, 1, 29, -28, -2, -4, 6, 22, -12, 7, -25, -39, 2, 32, -3, 10, 48, -42, -18, 12, 4, -26, 11, -31, -86, -7, -17, -3, 35, -17, 25, 9, 21, -17, 10, -4, 14, 17, -26, 22, 5, -2, 14, 19, -12, 27, -1, 29, -13, -8, 1, -38, 10, -18, 10, -19, -8, -18, -26, 13, 26, -15, -4, -8, 2, 8, 12, -35, 7, -6, 20, 35, -7, 5, -13, 2, 8, -1, 5, -26, 2, 7, -12, 33, 0, 10, 18, -49, -48, -18, -47, 7, 1, 4, 9, -20, 55, -20, 1, -2, 21, 34, 13, -1, -70, -6, 15, -1, 21, 6, 26, -2, 21, -8, -30, -72, 1, -1, -31, 25, -8, -18, -23, 33, 7, -35, -25, 38, 38, 17, -32, 52, 12, -4, 13, 11, 9, -7, 0, 24, -31, -9, 8, -9, -54, 26, 0, -17, -10, 8, -6, -5, -52, 25, -9, 19, -14, -31, -1, -68, -2, 14, -4, -17, 2, -31, 8, 10, -7, 7, -14, 25, -37, 10, 29, -2, 0, 1, 29, -18, -29, -51, -10, 18, 57, -12, -11, 55, 38, 0, 10, -24, -6, 20, 6, 2, 29, 28, 30, 26, 13, 3, 7, 15, -49, 18, 4, -2, -53, -1, -15, 0, -11, 25, 28, -4, -12, 3, 14, 19, 19, 14, -3, 15, 15, -57, 1, -16, -6, 11, 11, 27, -42, -10, 24, 40, 10, 24, 13, 0, -7, -9, 50, 8, -9, -29, -6, 5, -24, 0, -15, 22, 53, -33, 29, -18, -12, -10, 8, -34, -30, -4, 50, 16, 9, -1, 10, 22, -33, -6, 3, 3, -44, -4, 23, 8, 5, 47, 20, 8, 17, -1, -38, 0, 2, 18, 4, -41, 12, -16, 4, 4, 13, 30, 1, 32, -17, -2, -12, 13, 59, -8, 5, -32, -6, 0, -23, 11, 13, 28, 6, -32, -55, 25, 6, 37, 14, -7, -6, -37, 7, -2, 44, 7, -10, -10, -25, -18, 1, 7, -40, 10, -8, -22, 0, 14, -12, -7, 21, 19, 11, 25, 5, -17, -22, -26, -28, -12, -4, -19, -31, -17, -15, 15, -9, -14, 23, 41, -18, -27, -16, -12, -35, 4, 54, -35, -1, -18, 1, -13, -26, 9, 25, 46, 8, -29, -17, 34, -15, 24, -33, 32, -42, -45, 37, 21, 78, -32, -34, -20, 24, -49, 21, -5, -33, -27, -14, -1, -3, 41, 36, -3, -3, 63, -4, -27, 9, -52, 11, -38, 1, 12, 9, -32, 42, -13, 21, 4, 11, -11, -10, 33, -3, 0, 19, 1, -8, -19, 35, -39, 9, 28, -2, 0, -3, -11, 5, 45, -3, -6, -19, 13, -10, 2, -46, 8, -44, -41, 21, 7, 38, -7, -6, -2, -23, 6, 1, -1, -28, 7, -16, 19, -1, 21, 17, 31, -40, 40, 1, -9, -9, -38, -42, -9, -1, -6, 40, -1, 20, 23, 22, 0, 5, -7, 17, 48, -3, 13, 0, 2, 13, 45, 37, 0, 21, 27, 5, -10, -2, 0, 23, 39, 4, 21, 17, -14, -28, 13, 20, 2, 15, -44, 16, -3, 6, 24, 0, 14, 2, -1, -4, 4, 29, 3, -23, 11, -6, 18, 13, 43, -46, 42, 1, 37, 13, -21, -64, 14, -47, -3, 25, 0, 29, 3, 24, 5, 4, -5, 0, 4, -2, 13, 8, 0, 16, 24, -9, 22, 10, -10, 8, -1, 8, -73, -5, -20, -1, 15, 25, -28, -56, 35, 29, -40, 2, -17, 39, 10, -50, 26, 0, 1, -17, 9, 4, -9, 7, 13, -56, 23, 8, -2, -63, 24, -19, 13, -11, 58, -3, -10, -44, 2, -10, 22, -10, -14, 28, -8, 33, 26, 5, -19, 29, -41, 10, 12, 22, 4, 19, 29, -18, 18, 24, 21, 25, 5, -26, -7, 10, -45, 11, 16, 20, -11, -18, 38, 16, -33, 19, -28, -9, 31, -12, -19, -6, 12, 31, 43, 20, 7, -5, -3, -19, -5, 0, -9, -29, -17, -24, -26, -3, 17, 24, 34, -35, 30, -3, 19, -5, 19, 5, -24, 10, -48, 6, -20, 21, -27, -21, 31, 20, 8, 3, 24, -16, -9, 15, 16, -13, -1, 19, 20, -7, -37, 0, -8, 30, -19, -47, 32, 28, 0, 23, -51, -56, -13, 11, 3, 0, -9, 60, 35, -3, -2, 7, -28, -13, -29, -12, -3, -34, -18, -5, 40, -11, 39, 27, 21, -4, 29, -71, 16, 32, 25, 0, 5, -13, -12, 7, -5, 20, -12, -43, -8, -5, 11, -35, 2, 17, -27, 20, -10, 5, 8, 30, 8, -14, -17, 16, -55, -7, -26, -23, 55, 4, 4, -15, -72, -11, 0, 27, 6, -51, -5, 4, 25, 14, 7, -28, -49, 3, 1, 10, 2, -12, 22, -31, 49, -8, 30, 9, -28, -34, -47, -14, -22, 18, -10, -9, 13, -34, 26, -9, -7, 27, 11, -24, -22, -13, -5, -38, 30, 28, -29, 3, 9, 29, -2, 39, -6, 22, 29, -18, -41, 19, 8, -2, 12, 25, 5, -54, -69, 38, 8, 35, 66, 25, -10, -4, 5, 3, -10, -43, -1, 17, 10, -7, 54, 0, 5, -28, 53, -7, 14, 0, -11, -24, -33, -18, 4, 28, -16, 29, -32, -21, 13, -2, -18, 15, 10, 6, -24, -9, 0, -21, 16, 15, -42, -16, -2, 0, -7, 14, -33, 12, 18, -14, -17, -9, -21, -21, -17, 16, -18, -13, -49, 1, -5, 8, -6, 61, -9, -55, 1, 0, 5, -7, -5, 41, -5, -9, 22, -24, 8, -12, 63, 2, 25, -28, -56, -52, -8, -37, -22, 26, -5, 20, 0, 34, 23, 9, -16, 3, 5, -4, 5, 16, -3, 13, 20, -8, 40, -8, -2, -29, -2, 34, -37, -20, 12, -36, -5, 24, -36, -54, 11, 2, -14, 15, -22, 5, -38, -57, 0, 0, -13, -23, -6, -22, -2, 10, 15, 7, -8, -11, -1, -25, 55, -23, 13, 9, -56, -4, -8, 27, 18, -50, -36, 30, 10, 1, -11, 40, 38, -8, -14, -7, -11, 0, 18, -25, 1, 4, 42, 38, 6, 8, 22, 35, 0, 22, -22, 25, -19, -4, -6, 30, -22, -24, -1, 15, 0, 32, -20, 9, 2, -54, 40, 35, 2, -35, 0, -1, 2, 6, -28, -30, 11, -6, 7, -39, 35, -26, 42, -3, 38, 40, -7, -50, -8, -8, 15, -14, -21, 0, -25, 42, 5, -11, -9, 0, -3, -7, 11, -25, 9, 13, 2, -19, 8, -9, 12, 11, -3, 43, 24, 1, -23, 1, -24, -23, -17, 37, 14, 12, -7, 24, -20, 17, 25, -23, 36, 28, -2, -15, 20, 10, -4, 27, -9, -15, 10, -10, -1, 13, -19, -24, 1, 3, -49, 0, 5, -26, 10, -20, 16, -29, 9, 39, -29, 18, -9, -4, -3, 31, -37, -4, 26, -24, -2, 9, 43, -44, 0, 28, 19, 19, 4, -38, -16, 18, -55, 0, -24, -1, -12, -14, -13, 52, -22, 45, 1, -23, -10, -40, 35, 35, -14, 15, 23, 1, 3, 29, -23, -3, -12, -5, 9, -49, -15, -43, 39, -3, -20, 9, -1, -5, 32, 6, 30, -13, -29, 31, -48, 21, 6, -6, -12, 35, 7, -35, 17, -8, 10, 6, 5, -9, -18, 31, -11, -7, 3, -2, -38, 28, -30, 33, -26, -9, -22, -25, 42, 17, 14, -15, -38, -30, 0, 0, -20, -14, -12, 29, 0, 0, 5, 13, -16, 33, -21, 5, -5, -3, -11, -34, 41, -3, 25, 18, 0, -12, -3, 7, -10, -6, -22, 34, -30, 8, 3, -3, 0, 27, 2, -25, -7, 0, 8, -35, -7, -4, -5, -18, -28, 2, -9, -18, -12, 16, -15, -16, -40, -21, -30, -19, 25, 11, 24, -1, -83, 30, 1, -4, 6, 8, -8, -10, -7, -10, 0, 15, 12, 27, 12, -4, -19, -7, 2, -13, 36, 11, 77, 17, 17, -35, 20, 12, -12, 17, -16, 32, -38, -14, 11, 5, 1, -1, -6, -21, -3, -11, -7, -19, -17, 1, -21, -11, 13, 9, 3, -3, -36, 12, -4, 3, -41, 10, 17, -20, 15, -7, -5, 7, -64, -3, 6, -3, 1, 38, -14, 5, -19, 14, -9, 0, 11, 38, 16, -7, 38, -37, 24, -29, 0, 2, 1, 2, 9, -63, 3, -26, -12, 8, 4, 34, -24, 8, 17, 3, -20, 28, -12, -12, 28, -1, 9, 6, 13, -21, -44, 4, -17, 23, -14, -76, -6, 2, -17, 30, -11, 4, 9, -31, 3, 3, -27, 35, -12, -1, 7, -26, 25, 1, -3, -32, 13, 1, 4, 13, -14, 38, -4, 6, 6, -48, 22, -33, 45, 4, 5, -8, 15, 12, 12, -28, 19, 22, 8, 38, -35, 28, -23, 8, -6, 35, -47, -14, 22, -4, 2, 44, 23, -43, -26, 0, 21, -2, -12, 9, -10, 22, -17, 4, -5, 1, -15, 7, 26, 2, -10, 35, -19, -20, -1, -55, -7, -2, -21, 14, 26, 3, -10, 15, -20, 23, 6, 11, -10, -8, 49, -84, 33, -1, -17, 32, -27, -31, 14, -35, 13, 42, -27, -1, -12, 9, -38, -3, 2, 28, 2, 10, -7, -27, 0, -3, -17, -20, 36, -13, -30, 9, 2, 36, -9, -7, 31, -18, -14, 16, 31, 43, 21, -50, 4, 10, -9, 4, 28, -43, 59, 0, 5, 16, -42, 5, -10, -5, -26, 27, -25, 9, -28, 4, 6, 48, 30, -3, 23, -18, -16, 1, -17, -36, 4, -5, -11, 5, 21, -44, 54, 1, -16, 4, 10, 15, -9, -50, -4, 0, -18, 29, -28, 6, -33, 16, -11, 9, -21, -2, 10, 2, 39, 14, 37, 20, 6, -9, -19, -5, -55, 11, 0, 2, 69, 32, 4, 47, 4, 19, -5, 20, -15, 14, -11, 2, 12, -37, 29, 15, 20, -6, -28, -10, -30, -1, -24, -39, 7, -37, -14, 0, -34, -40, 25, -7, -2, -32, 24, -17, -30, -73, -1, 5, -44, 22, 31, -1, -63, 13, -5, -58, 14, 1, 37, -1, 49, 0, -2, -48, 11, -29, -16, 4, -29, 6, 25, 16, -36, 29, 34, 76, -30, 10, -6, 9, -2, -26, -1, 4, -15, -35, -4, 17, 29, -6, 62, -6, 20, 20, -12, 47, -2, -10, 3, 33, -27, -51, -17, 3, -10, -49, 21, 0, -50, -31, 0, -16, -60, 11, -6, -22, -53, 38, 0, -44, -24, -16, 38, -40, 60, -47, -5, -8, 23, -45, -19, -15, -6, -9, 11, 12, 34, 11, 38, 34, 0, 24, 8, 28, -4, 4, 7, 3, -23, -19, 4, 4, 6, 1, 6, -28, -43, 18, -29, -6, -19, -35, -30, 33, -10, -69, -23, -7, 2, -31, 28, 20, -20, -34, -8, -25, -42, 10, 13, -1, -17, 36, 10, -31, -27, -41, 33, -17, 77, -9, 0, 4, 7, -12, -31, -6, -31, -10, 9, 30, 2, 23, 46, 59, -40, 34, -4, 7, 18, -7, -7, 6, -25, -14, 0, -8, 4, -3, -17, -9, 6, -24, -8, -29, -31, 1, 10, 11, -19, -66, -66, -4, -5, 17, 38, 7, -12, -4, 0, -9, -22, 13, -11, 1, 9, 5, 1, -47, -28, -16, 7, -21, 42, 24, -28, 11, 16, -14, -2, -1, 14, -41, 15, 58, -34, 4, 22, 2, -37, 11, 3, 2, 8, 4, -13, -11, -8, -15, 6, -36, -9, -13, 1, -14, -5, 16, -6, -24, -1, 52, 38, 25, -19, -34, -35, -7, 3, 32, -11, -13, 0, -4, 10, -2, -19, -8, -14, 5, -5, 23, -11, 1, -36, -8, -28, -13, 8, -33, -28, 34, 46, -25, 10, 13, -10, -82, 13, 29, 13, 15, 3, 0, -26, 9, -4, 11, -9, 16, -30, -6, -47, 9, -15, -26, -15, 3, 0, 13, 4, 5, 6, -31, 13, 81, 24, -2, 16, -37, -18,
    -- layer=2 filter=0 channel=3
    0, 3, -50, 13, 8, -7, 19, -1, -27, 0, -2, 35, -4, -18, 3, -4, 28, -8, 6, 4, 8, 21, -37, -20, -1, -12, 17, -18, -36, -18, -9, 10, 20, 18, 14, -15, 8, -30, 6, -2, -12, 17, 29, 0, -2, -43, 19, -26, -13, -11, 2, -16, -6, 15, -22, -54, -13, 4, 32, 11, -31, -8, 18, -14, 2, 8, -34, 56, -4, 7, -12, -4, -17, -9, 10, -8, -38, -2, -3, -3, 20, -4, -10, 44, 13, 0, -50, -18, -25, 18, -20, -12, -34, 26, -49, -8, 44, -5, 42, -2, 23, -12, 9, -5, 2, 22, -12, -6, -10, -24, 13, -8, 5, 13, -4, -23, 1, 16, 6, 7, -12, 0, 29, 9, -20, -9, 0, -36, -8, -2, 10, 10, -12, 4, 13, 1, -22, 7, -1, 8, -2, -3, 6, -7, 34, -14, -3, 18, 21, -15, -31, 2, -3, 48, 0, -8, -1, 29, -20, 7, -7, -28, -48, -14, 3, 42, 17, 10, -16, 0, -20, 7, 0, -4, 0, 6, 3, -13, -1, -68, -7, 32, -27, -6, -25, 15, 15, -3, -14, 22, 19, -9, 6, 8, 11, 26, 13, 1, -3, -3, -19, -24, 9, 27, -14, 3, 10, -7, 49, -20, 5, 12, 21, 18, -18, -8, 25, 11, 11, -26, -26, -4, -22, 9, 19, -18, -16, -19, -24, 7, -3, 5, 3, 32, 7, 4, -5, 0, 28, -13, 2, -1, 4, 4, 1, -1, -21, -12, 3, 26, -35, -2, -3, -7, -1, -2, -1, 3, -6, 37, 13, 13, 24, -10, -41, -41, -8, 4, -14, -43, 14, -7, -16, 5, 36, 28, 29, 0, -31, -19, 16, 5, 22, -20, -14, 5, 49, -4, 47, 12, -4, -6, -26, 12, 16, -5, -17, 15, 11, 12, 3, 0, 37, -15, 1, -2, -8, -49, -16, 39, -26, -22, 20, -5, -20, 5, -5, 7, 32, -4, 3, -6, -10, 1, -14, -19, 16, 10, -17, -3, 5, 28, -42, -8, 6, -1, 13, -7, -17, 20, -9, -17, -15, -7, -11, 3, -19, -41, -10, 24, 32, 12, 1, 39, 18, 0, -24, -34, 0, -9, 8, 24, -1, 12, 3, -4, 9, 0, 33, -3, -2, -43, -13, 6, -32, -17, 34, -8, -38, -7, 0, 19, 14, 36, 9, 1, -10, 31, 3, -7, 0, -6, -34, -10, 32, 13, -33, 8, -13, -2, 0, -36, -23, 38, 12, -6, -25, -40, -8, -37, -7, -59, -19, -21, 7, 11, 27, 38, 4, -5, -33, -33, -7, -1, -33, 5, -24, 3, -7, -46, 6, -25, 33, 35, 0, -13, 10, 22, -9, -32, 14, 23, -59, -12, -37, 4, -22, 21, 5, -7, -30, 11, -31, -1, 32, -8, -7, 12, 17, 5, -12, -18, 9, -12, -52, 29, 1, -2, 40, 1, -11, 4, -19, -4, 2, 27, -9, -7, 7, -3, 16, -2, 28, 4, -14, -4, -10, -4, 4, 38, 9, 12, -4, 0, 23, 28, 10, -45, -5, -12, -13, 0, -53, 21, 32, -3, 19, 9, -6, 10, 19, 31, 2, 7, -16, 52, 15, -14, 27, 3, -11, 9, -9, 15, -10, -2, 2, 10, -26, -8, -17, 13, 3, -4, -25, 22, 5, 30, -38, 19, -14, 0, 5, -9, 20, -1, 5, 4, -2, -25, 0, 3, -14, 15, -39, -4, 1, -1, -7, 17, -8, 0, -6, -38, 0, -1, 2, -15, 9, -6, 0, -6, -10, -9, -2, 12, 1, 12, 5, 36, -17, -27, -28, 7, -17, 7, 41, 39, 31, -23, 15, 12, 47, -27, 0, 22, 0, 1, 22, 35, 16, -32, -24, -43, -33, 14, 26, 15, 9, 3, 6, 11, 0, 21, 3, -6, -12, -4, -19, 21, 4, 1, -12, 12, -11, 3, -8, 8, 13, -9, -46, -14, 2, 5, 21, 4, -20, -2, -2, 0, 9, 0, -10, 13, 17, -30, -7, -10, -33, -25, -17, 20, 4, 35, -20, -6, 7, 15, 17, -13, 20, -12, -1, 7, 10, -24, -8, 1, -28, -5, 29, -15, 12, -23, 4, 33, -40, -4, 6, -13, 13, 35, -27, 19, -8, 35, -15, -5, -3, -14, -9, 11, 34, 6, -6, 14, 20, -15, -4, 11, 8, -1, -21, -8, 1, 10, -13, -18, 20, -4, 8, 0, -30, 5, -7, -14, -16, 10, -3, 0, 39, -37, 10, 1, 51, -13, 1, 17, -12, 20, 9, -9, -12, 7, 32, 11, 7, 26, 8, 33, -16, 3, -6, 5, 0, 3, -39, 4, 4, 31, -18, 3, 12, -24, 0, -14, 9, 1, 43, -25, -5, -12, -9, -3, 20, -7, -18, -10, 5, 5, -14, 7, -5, 3, 9, 3, -15, 16, 10, 2, -3, 15, -7, 5, 23, -15, -45, 23, 14, -1, -15, -21, 14, -44, -8, -24, 10, -22, 28, 9, 25, -33, 0, 1, -26, 20, 0, -5, 27, 23, 26, 20, 1, 18, 18, -14, 35, -6, -13, -20, 24, 10, -60, 0, -3, -11, -23, -12, 3, -8, 17, -3, -5, 4, -25, 16, -3, 4, 31, -5, -19, -26, 1, 5, -32, 5, -12, -5, 9, 6, 16, 14, 49, -16, -16, -26, -21, -5, 3, -26, 22, 4, -23, -23, 27, -12, 8, 0, 12, 6, -20, -2, 17, -1, 3, 3, -7, 28, 0, -14, 34, 37, -10, 29, 20, 19, 14, -16, 15, 16, -6, -25, 6, 6, 31, -36, -10, -7, -31, 17, -8, 21, 33, 4, -19, -11, 25, -3, -32, 8, 4, -12, -20, 0, -10, 2, 33, 13, 3, 1, 13, -8, -4, -30, -4, 10, 16, -5, -4, -3, -41, -10, -21, 24, -7, -1, 17, 24, -20, -10, -3, 37, 16, 2, 10, -9, -7, -25, 3, 25, -26, 27, 2, -46, -10, 1, 25, 13, 5, -5, -2, -3, 4, 13, -8, 2, 0, 0, -9, 19, 18, 45, 13, 19, -2, 8, -6, -3, -50, 4, -36, 0, -25, 13, -4, -22, 15, -68, -6, -34, 24, 3, -24, -9, 15, 6, 4, 0, 12, 4, 15, 6, -21, 14, -3, -4, -14, 25, 12, -16, -6, 24, -3, 7, -8, -5, -3, 6, -63, -11, -27, -5, 16, 21, 6, -4, 34, 19, 13, 2, -12, -8, -39, -31, 22, 21, 50, 5, -9, -6, -14, -45, -64, 36, -53, -3, -11, 19, -42, 9, -27, -40, 13, -19, 2, 14, -6, 9, -34, -3, 1, -24, 29, 4, -2, -7, -15, 35, -8, -11, -36, 12, 5, 27, -7, 3, -37, -41, 42, 4, -24, 25, -22, 3, -11, -25, -18, -28, -2, 0, -14, 13, 32, -30, 30, -4, -46, -11, 21, -12, 11, 10, -6, 5, 22, -14, -17, 2, -45, -3, 26, 75, 13, 13, -23, -39, -18, -7, 33, 2, -14, 51, -33, 18, 15, -10, 30, 8, 19, 32, -1, 56, -8, 19, -12, -5, 2, 17, 9, 108, 44, -17, 48, -25, -49, -15, 4, 9, 11, 17, -44, -16, 0, -1, 0, 5, 24, -17, 16, -2, -42, 17, -8, -8, 40, -22, 17, 12, 30, 5, -15, 2, -50, -18, 29, -17, -16, 7, 13, -28, 13, -3, 35, 1, 32, 20, -31, 6, 30, 12, 50, 4, -2, -9, -8, 14, -11, 6, -23, -8, -32, -30, -7, 11, 21, 12, 45, -15, -52, 12, -8, 33, 22, -4, 21, -12, 6, 1, -7, 7, 9, 4, -25, -2, -16, 14, -46, 16, 22, -6, 3, -7, 28, -26, -32, -9, -15, -1, 10, -3, 10, -60, -38, -34, 8, -16, 15, 16, 23, 4, 21, -7, 4, -11, 17, 9, -2, 11, -21, 14, -7, 13, 12, 12, -38, 0, 6, 25, 5, 10, 5, 4, -25, 29, -5, 18, -15, -22, -13, 1, -5, 16, -19, 7, -25, 15, 0, -5, 5, -31, -14, 39, -5, -15, 0, -9, 16, -23, 19, 14, 54, -2, 14, 5, 6, -26, -21, -62, 18, -3, -33, -3, 27, -7, -7, 4, 21, -7, 15, 0, 13, 9, -10, 11, -4, 17, -6, 6, 8, -48, -6, -15, 1, 6, -11, 0, -2, -6, 25, 17, 26, 14, 17, -41, -8, 12, -5, 18, 4, 6, 23, 8, 0, -32, 24, 14, -9, -21, -5, 5, 23, -4, -21, 35, 27, -12, -7, 27, 12, -7, 20, -5, -9, -33, 24, -10, 3, -5, -18, 10, 10, 7, 3, 4, 0, 21, 8, 7, 0, 39, 21, 20, 17, -22, -10, -55, -30, 18, -27, 29, 19, -2, -20, 8, 21, 6, -15, 44, -8, 4, 26, -15, 4, 9, -2, 5, -16, -43, 18, -23, 12, 18, 7, 4, -31, 2, -19, 14, 1, -16, -17, 13, -3, -33, -11, -47, 19, -28, 17, -14, -12, 2, -13, 0, 14, 0, 10, 0, 1, -1, -9, 9, -4, 18, -49, -11, 17, -5, 2, -20, -3, -46, 21, -17, -33, 8, -11, 10, 12, 5, -30, -32, 10, 7, 24, -18, 3, -13, -24, 4, 5, -18, 18, -10, 29, -1, 6, -11, 2, 0, -40, 21, -95, 0, -7, 42, -44, -65, -44, -5, 2, -14, 25, -16, -8, 39, 5, 7, 19, -23, 7, 1, 0, -18, 11, 28, 0, -24, -54, 16, -24, -2, 3, 46, 0, 19, 24, -13, -53, 30, -15, 15, 2, -35, -16, -8, 13, -5, -43, -5, 33, -39, -41, -7, -7, -36, -20, 0, 37, -6, 14, 7, 8, -20, -60, 5, -94, 9, 65, 31, -17, -28, -46, -41, 12, -25, 23, -15, -19, 30, -52, 32, -11, 1, 16, 2, -4, 9, -30, 22, -1, 12, -38, -22, -46, -11, 9, 52, -1, 27, 9, 1, -82, -17, -7, 23, 1, -7, -66, -18, -7, -6, -8, 18, 31, 0, -54, -1, 27, 15, -4, -30, 30, -19, 30, 4, 75, -29, -44, 24, -37, 21, 21, -14, 3, -98, 10, -39, 18, -14, 21, -5, 26, 2, 24, 17, 0, 13, 22, 6, 4, 6, -30, 15, 5, 4, -9, 5, -11, -19, 6, 40, 8, -10, 74, 19, -81, 2, -3, 32, 4, -27, -34, -33, -2, -5, -17, 0, 3, -8, -23, 4, -20, 1, 1, 14, 16, -14, -4, 7, 9, 11, -41, 6, -22, -9, 29, 22, 1, -22, -1, -8, 0, -48, 25, -4, 0, -9, -24, 9, 29, -4, 26, 0, -9, -4, -24, 29, -6, -9, -16, -2, -12, 13, -4, 21, 10, 10, 53, -19, -23, 41, -15, 31, -5, 5, 0, -64, 0, -3, -17, 1, -27, -11, -3, 6, -6, -30, -1, -1, 24, 10, -7, 0, -27, -19, 1, 15, 33, 27, 5, 1, 30, -2, -3, -47, -5, -25, 15, 10, -3, -12, -8, 41, 13, -21, 4, 0, -5, 23, -14, -4, -3, -1, -5, -37, -10, -32, -2, 19, -15, -25, -52, -12, 18, 15, 13, 14, 27, 14, -4, -12, 0, 2, -11, 19, 10, 16, -27, 8, 0, -25, 13, -17, -25, 23, 10, -1, 0, -15, -8, 28, 19, -18, -3, -14, -23, -17, 21, -22, 15, -20, 28, -6, -29, 20, -12, -1, 0, 7, -16, -3, 20, -4, -22, -9, 4, -1, -34, 8, -37, -2, 3, 1, 5, 6, -21, -28, 16, -6, 4, -49, 14, -4, -13, -7, 0, 0, -21, -13, -19, -21, -52, 1, -11, -42, -27, -3, -15, 8, 6, 6, -30, -27, -31, 16, -14, 5, 5, -38, -33, -10, 11, -1, 0, -58, 12, -22, 9, 34, -67, 3, 20, 4, 0, 0, 10, 12, -20, -15, 4, 24, -40, 41, -42, -30, -7, 3, -19, 3, -16, -4, 5, -12, -18, -26, 0, -19, -14, -18, 1, 5, -7, 38, 14, -11, -62, -9, -4, 14, -8, -4, 8, 23, 4, 8, 17, -23, -22, 3, -43, 14, 46, 5, -47, -45, 4, -14, 14, -39, 2, -4, -1, -9, -7, 14, 1, 11, 7, 2, 25, 17, 6, -11, 5, -1, -11, 12, -17, -9, 0, -9, -7, -8, 23, 20, -25, -4, -13, -8, -1, -45, -18, -3, -6, 2, -44, 0, 0, -47, -39, 5, 11, -8, -1, 15, 10, 1, -9, 4, 0, 0, -41, 0, -68, 5, 64, -11, -15, -49, -25, -2, 24, -51, 14, -23, 2, -2, 61, 28, 19, 27, 7, -9, 30, 16, -13, 0, -5, 3, -8, 4, -16, -23, -3, 40, 41, 3, 11, 13, -16, -7, 9, 30, -6, -11, -37, -3, 2, 0, -33, -14, -14, -5, -54, -3, 6, -7, 7, 1, 18, -5, 11, 2, 38, -10, 0, 41, -12, 0, 45, -30, -27, 11, -27, 10, 28, -62, 29, -27, -6, -5, 9, 4, 31, -1, 4, -4, 27, -28, -26, -6, 5, -13, -43, 14, -10, -50, 3, 44, 23, -5, -36, -9, -28, 1, -14, 9, -4, -22, -13, -2, 6, 10, -21, 0, -6, 0, -54, -6, -11, -11, 7, -37, 18, 45, 10, -11, -37, -30, 6, 13, -3, 5, 6, -17, -35, 1, -15, -15, -9, -17, 7, 15, -6, -20, 2, 9, 11, -39, 12, 11, 1, -8, 21, -14, 5, -8, -35, 29, -5, -12, 8, -6, 14, -4, 1, 3, -25, 13, -15, -27, 7, -36, 0, -10, -10, 0, -5, 18, -29, -2, -13, 0, 9, -15, 24, 23, 16, -4, -8, -6, 36, 0, 11, -2, 17, -2, -36, 12, -4, -11, -5, -31, 3, -30, -11, 16, 9, 6, -8, 17, 14, 11, 11, 0, 3, 14, 4, -6, 10, -5, -7, 33, 7, 18, -3, 5, -16, 30, -36, 7, 5, 10, -10, 0, 12, -16, 16, -14, 9, -6, 17, 27, 8, 12, -11, -3, 12, -17, 1, 3, -13, 5, 1, 0, -91, 15, 5, 5, 23, -10, 2, 9, -11, -19, 11, -21, 20, -26, 27, -1, 25, 37, -36, -26, 4, 7, 7, 10, 23, 3, 30, 0, 0, 24, -29, -5, -10, -22, -2, 6, -4, 10, 26, 22, 25, 8, 21, -9, 14, 12, 14, 37, -13, 2, 0, 29, 13, 9, -58, -8, 1, -15, 10, -4, -20, -5, -19, 0, -17, -24, -32, 46, -30, 10, 1, 9, -34, 49, -3, -24, -3, -16, 14, -1, 26, -9, -25, 14, 6, 1, 7, 4, -15, 3, -1, 4, -4, 10, -7, 5, -24, -11, -9, 13, 5, 2, 22, -8, -3, 8, 5, -12, -16, -17, 12, 4, -3, 0, -42, 17, -14, -28, -25, 1, 8, -19, -8, 8, -4, -1, 11, 0, -20, 1, -38, 42, -14, -2, 39, -34, -19, -26, -31, -25, -3, -47, 22, 0, 17, -20, -33, 7, 10, 16, 5, 3, -3, 20, 4, -5, 3, 7, -8, 14, -30, -31, -4, -2, 8, 49, 49, 2, -23, -1, 35, 20, -32, -18, -3, 7, 4, -7, -19, 3, 3, -28, -61, -11, 32, -2, 3, -24, 0, 14, 6, -6, 24, -10, -7, 19, -10, 0, 63, 2, -1, 12, -12, -1, 18, -5, 14, -12, 5, -5, 25, 8, -55, 4, 14, -6, 4, 1, 8, -20, 5, 52, -19, 21, 3, -12, -8, -18, -2, -7, -6, 10, -9, -24, 20, 0, 15, -41, -43, 30, 2, -10, -24, 4, -22, 11, -35, 6, 22, 15, 1, -29, 1, 2, -9, -12, 41, -3, 10, 8, -15, 2, -6, -9, 14, -21, -1, 16, 42, -59, 13, 5, 0, -33, -51, -21, 7, 26, -9, 9, 19, -26, -26, -10, 1, 10, -18, 0, 7, 15, 10, -15, 5, -11, 1, -3, -34, 10, -18, -2, 12, -39, 23, -1, 3, 5, -2, 21, -4, -5, -35, 6, -8, 20, 7, -11, 15, 34, -15, -12, 25, -21, -9, 34, -27, -6, -6, -45, -20, 21, 5, -35, 12, -26, 9, 11, 4, -7, 19, 3, 29, 25, 4, 7, 20, 15, 0, -6, 5, -2, -57, 7, 0, -26, -13, 4, 12, 5, 17, -13, -20, -1, -18, -20, 1, -43, -32, -9, 0, -4, -8, -3, -15, 8, -15, 0, 7, 10, 8, -3, 11, 25, 0, 4, 8, 1, 6, 30, 42, -19, -3, -10, -53, 11, -8, 2, 22, -37, -14, 8, 9, -2, -25, 10, 3, -1, 4, 0, -4, -16, -15, -19, -5, -26, -7, -8, -2, 21, -7, 5, -2, -17, 20, 2, 36, 1, -19, 0, 20, -29, 10, 10, 10, 7, -4, 0, 9, 27, 4, 3, 13, -27, 24, 19, -24, -3, -9, 1, 2, 25, 11, 72, 46, -44, 8, 6, 17, 5, 19, 1, 7, -6, -23, -8, -2, 48, 21, -26, 18, -4, -4, -2, 6, -6, 17, 0, 5, 12, -17, -51, 5, -15, 5, 12, -19, 18, 2, 12, 20, -20, 47, 6, 5, 10, 9, 49, 6, 0, -11, 11, 6, -3, 9, 11, -11, -17, -11, 16, -16, 11, 22, -2, 1, 0, 4, 43, 5, 15, -28, -17, -1, -6, -13, 9, 9, -23, 4, 4, 38, 37, -24, 0, -16, 27, 18, -11, -1, -9, 3, -17, -6, -13, 20, -26, 0, -4, -4, -28, 16, -15, 20, 12, 15, 5, 22, 9, 1, -4, -5, 6, 6, 6, -21, 17, 1, -14, -50, -6, -23, 9, -12, -40, -19, 2, 16, 3, 20, 2, -8, 29, 31, -32, 7, -3, -30, 0, -16, 0, -10, -6, 25, 7, 17, 25, -50, 15, -64, 8, 12, -7, -5, 19, 14, -21, 5, 6, -17, 32, -57, 7, -14, 17, 19, -2, 14, 17, -13, 5, 53, -5, -20, -22, 8, -8, -11, -2, -6, -30, 10, 5, -38, -5, 2, -5, -28, 20, -37, 11, -12, -8, 2, 9, 15, 3, 24, -30, 41, -16, -19, -12, 9, -20, -12, -15, -29, 4, -32, -19, -13, 13, 7, 16, 7, 2, -9, -11, 12, -18, 3, 20, -8, 9, -16, -7, -12, 51, 9, 15, 19, 12, -11, 21, 34, 36, -40, -8, 9, 26, -11, 12, -12, -25, 0, -4, -41, -8, -13, 24, 15, -2, -4, 3, -1, -6, 19, 1, -5, 0, -5, -22, -19, 36, 17, -47, 1, -11, -13, -29, -22, -5, 17, 30, -58, -13, 10, 34, 13, 10, -7, -9, 45, -2, 2, 17, 3, 7, 1, -3, 7, -37, -3, -14, -14, -7, -15, -6, -8, 19, -35, -34, -1, -1, 6, -4, -18, -8, 3, -12, -28, 3, 36, 11, 38, -3, -1, 2, 1, -6, 46, 6, 12, 34, 18, -7, -22, 1, -3, -12, 6, -21, 21, -45, -5, 7, -38, -16, 9, -14, 12, 1, 9, -1, 4, 0, 21, -12, 7, -16, -10, -2, 13, 25, -12, 16, -5, 9, 6, 27, -3, 5, -13, -38, -13, -20, 16, 11, 8, -7, -5, 39, -51, 14, -16, -11, 6, -19, 60, -1, 2, 12, -31, 9, 25, 3, -2, 52, 40, -19, 0, 8, 1, -7, -59, -12, -2, 20, -26, -10, 49, 22, -13, 2, 0, 4, 0, 3, 14, -18, 3, -22, 7, -17, 56, 1, -3, 46, -2, 9, -28, -16, -1, -5, 6, 22, -12, -19, 13, 14, 6, 16,
    -- layer=2 filter=0 channel=4
    -9, -5, 11, -58, 22, -21, -9, -6, -13, -30, -15, -8, 1, 6, 9, 2, 56, -33, 12, 26, -13, -39, -16, 26, -20, 40, -25, 27, -7, -7, -17, -9, -45, 11, -56, -6, -5, -65, 6, 2, -33, -44, 37, -3, -6, -23, 9, -27, 0, -88, -1, 44, 1, -28, 11, 15, -30, 2, 0, 24, -23, 17, -9, 35, 0, 1, 9, 6, 6, -4, -1, -4, 15, -29, -65, 30, -8, -49, 6, 8, 24, -9, 30, -11, -3, -7, 13, -4, -10, -21, -13, -1, 18, 27, 10, -13, -32, -3, 0, -8, 0, -29, 14, -12, -10, -15, 6, -4, -5, -5, -25, -43, -39, -88, -9, -22, -6, -5, 12, 0, -21, -7, 11, 5, 0, 8, 0, -8, 3, -11, -9, -24, 2, 2, -37, -7, 19, -40, -45, 28, 6, -45, 5, -8, -3, -4, 36, -2, 4, 17, 26, -39, -21, -37, -24, -11, -1, 28, -5, -9, 4, 2, -28, 8, -9, -19, 11, -1, 10, -29, -11, 5, 11, -36, -2, -32, -3, -85, 0, -25, -7, -5, 20, -11, -31, 0, -12, -3, 10, -15, 0, -32, -2, -11, 14, 13, 14, 13, -24, -4, 41, -37, -48, 32, 14, -4, -1, -12, 15, -13, 30, -23, -11, 32, 3, 35, -26, 7, -25, -12, 8, 45, 6, 0, -56, 16, 19, 22, 51, -22, 17, 6, 12, 27, -32, 28, 4, 0, -26, -25, -13, -74, -6, -33, -16, -17, 12, 18, -27, 0, -23, 4, -8, -8, -23, -54, -12, -7, 13, 6, 11, 8, -35, -5, 40, 2, -19, -31, 24, -32, -14, -13, 61, -29, 43, -57, 13, 12, 24, 23, -6, -22, -7, 3, 3, 38, -21, 10, -67, -4, -5, -8, -5, -27, 5, -5, 15, 21, -29, -3, -11, -1, -3, -25, 36, -8, -12, -13, -15, -17, 31, -5, -14, 24, -53, 12, 8, -5, -1, -7, 9, -1, 8, 27, 15, -13, -49, 10, 19, -42, 8, 0, 41, -15, 2, 2, 17, 2, 25, -72, 14, 9, -8, 24, -26, -17, -33, -4, 5, 26, 8, 2, -43, 30, -15, 4, -9, -10, 6, 0, 13, -27, 48, 2, 2, -21, -34, -30, 66, -17, -5, -58, -29, -6, -10, -15, -31, 0, -37, 0, 0, -8, -18, 10, -6, -5, 3, 8, 41, -19, -26, -10, 12, -43, 29, -32, 32, -5, 4, 2, 39, 49, 10, -40, -6, 5, -5, 21, -38, -22, -29, 40, -20, 1, -51, -22, -6, 9, -38, 0, -5, -26, 11, 0, -4, 8, 51, 17, -7, -51, -2, -27, 66, -98, -1, -39, -10, -34, -37, -22, -16, -18, -43, 2, 3, -5, -19, 48, 2, 0, 7, 4, 29, -9, -30, -5, -6, -21, -16, 16, 3, 1, 32, -7, -11, 38, -4, -4, -16, 20, 15, 24, 7, 31, 2, 41, -1, 17, 12, -8, 8, 43, 13, 10, 43, -20, 12, 9, 0, 27, 8, 2, -3, -15, 16, -18, -61, -66, -3, 6, 6, -18, 14, -18, -26, -7, 3, -5, -7, 13, -27, 4, 10, -2, 5, -5, 1, -9, -45, -10, 15, -15, -40, 5, -1, -22, 18, 0, -11, 49, 6, -12, -28, 29, 0, 30, 1, -5, -18, 21, 4, 11, -21, 5, 17, -27, -50, -4, -12, -17, 10, 1, 17, -2, -14, 12, -5, -29, -1, -17, -44, -77, -13, -35, -4, -32, -4, -8, 8, -17, 25, 8, 12, -5, -15, -58, 0, -6, 18, -34, 11, 2, -22, 6, 23, -7, -73, -3, -8, -45, -2, 6, -41, 33, 14, -54, -16, 59, -1, -5, 13, -24, -5, 6, -1, 31, 2, 19, -14, -12, 2, -6, -17, 8, 13, -8, 32, 31, -67, 10, -4, -12, -24, -9, 2, -60, -9, -76, -30, -33, -3, 2, 21, -6, -17, -1, 16, -8, -20, -50, -13, -2, 22, -16, 3, 12, -10, 4, 26, 5, -53, 14, 14, -59, 35, 1, -30, 5, 12, -49, -44, 27, -31, 4, 3, -44, 17, -21, 18, -33, 10, 4, -76, -5, -21, -8, -50, 3, 22, -2, 47, 9, -64, 15, 7, -34, -19, -4, -7, -39, 0, -80, -16, -28, 13, 4, -19, 10, -4, -11, 30, -16, 8, -45, -6, 7, 18, -7, 25, 22, -22, 0, 19, 0, -56, -12, 18, -25, 6, 6, 21, -12, 17, -41, -10, 21, -20, 10, -24, -40, 16, -17, 11, 45, -30, 3, -52, -31, -13, 0, 2, 8, 11, 4, 40, 18, -84, 11, -12, -43, -20, -14, 8, 1, -11, 7, -8, 8, 4, 3, -24, 10, -27, -33, 9, -23, -3, -60, -8, -4, 1, -28, -9, -10, -3, 0, 10, -1, -24, -2, -18, -19, -1, 5, 34, 32, 31, -67, -7, -29, -17, 37, 15, -18, 12, 0, 6, 11, -34, -6, -81, -8, -17, 22, 29, -3, 9, -1, 24, 18, -47, 11, -11, 3, -6, 14, 7, 6, -1, 3, -22, -9, 21, -4, 4, -16, -39, -20, 8, 0, -32, 7, -4, -11, -21, -1, -10, -9, -58, 2, 1, -22, 6, -36, 14, 12, -20, -6, 68, 12, 45, -19, 3, -11, -9, 45, -8, -27, -29, 5, -2, 9, -1, -14, 9, 40, -36, 1, -29, -37, -5, 1, 4, -7, -25, -9, 7, -1, -26, 25, 24, 1, 6, -19, 12, -22, 14, -5, 0, -8, -60, -6, -8, -23, -43, 22, 8, 4, 31, 20, 32, 2, -34, 7, -19, 0, -22, -13, -2, 10, 9, -8, -16, 0, 26, -43, 25, 13, 45, 18, -21, 20, 26, 22, 0, 17, -4, 1, 17, 9, -5, -22, 10, 9, 4, -8, 11, 0, -25, -14, -1, 24, 18, 2, -47, -119, -7, -21, 5, 9, 20, 14, -10, -5, 26, -6, 7, -17, 5, -4, -9, -8, -3, -22, 0, 8, -34, 2, -7, -14, -38, -31, 3, -17, 14, -8, 3, 13, -11, -33, 17, 12, -20, -1, -13, 9, 2, 21, -10, -5, -13, 9, 5, 37, -65, 3, 10, 4, -5, -13, 2, -7, 1, -8, -2, -1, 3, 5, -46, -75, -12, -25, -13, 26, -11, 3, -6, -13, 16, 17, -3, 23, 4, -9, 7, 7, 12, -16, 13, -5, -21, 5, 0, 9, -39, -12, 22, 0, 26, -3, -41, 5, -13, -42, 4, 19, -11, -43, -16, 7, 21, 2, 4, -13, -32, 23, -30, -39, -23, 10, -23, 22, 15, 11, 4, -27, -14, -20, -6, 1, 17, 20, 3, -52, 3, -59, 10, 64, 4, -4, -10, 11, 13, 0, 49, 9, 24, -24, -1, -7, 33, -40, 9, 8, -9, -3, 16, 18, -29, -32, 37, -30, 25, 8, -59, -25, -31, -21, -27, -7, -69, -34, 18, -5, 39, -48, 8, 3, -48, 18, 0, -39, -21, -1, -20, 7, 14, -5, -12, 13, -16, -8, 8, 32, 13, 26, 12, 16, 6, -50, -57, 11, 7, 17, -10, 35, 20, -8, 39, 12, 38, -7, -9, 5, 22, -55, 10, -7, -28, -7, 27, 1, -35, 3, -3, -27, 48, 0, -48, -16, -8, -48, 20, 11, -63, 12, 20, -24, 18, -15, 1, 13, 12, 17, -54, -21, 29, 0, -15, 14, 0, 5, 2, 5, -38, -26, -2, 22, 9, -7, 36, 21, -3, -37, -26, 1, 34, 10, 11, 23, -45, -6, 40, -1, 26, 6, -6, -4, 14, -34, -9, 14, -23, 2, -19, 6, -4, -1, -3, 0, 13, -10, -30, 57, -7, -34, 13, 10, -47, 17, -15, 0, 19, 23, -22, -9, 5, -7, -29, 25, -11, 29, -24, 41, 5, -9, 5, -43, -8, -16, -8, -8, 10, -38, 48, 20, 3, 2, -11, -9, 41, 21, 3, 14, -85, -5, 7, 12, -9, 33, 9, 4, 11, -63, 1, 20, -14, -7, -25, -5, 9, -4, 11, 16, 4, 6, -2, -13, 20, -19, 34, -2, 41, 17, -50, -9, -9, 7, -11, -33, 19, -6, -42, 53, -48, -4, 0, 22, 9, 9, 9, -32, 18, -8, 7, -6, -11, 23, 3, -5, 4, 24, 1, 20, 33, -10, -15, -3, -40, -31, 3, -30, 1, 42, -10, 6, 23, 21, 27, 30, -54, 0, 9, 21, -14, -18, -11, 16, 2, -1, -5, -12, -12, -32, 22, 0, 15, 44, -14, 1, 39, 36, 56, -10, 0, -15, 32, -16, 3, -14, -28, 23, -2, -8, 57, 2, 3, -7, 6, 47, 3, -6, -30, -15, 1, 45, 4, -29, 19, 44, -35, -9, 1, -17, 19, -40, -5, 16, -11, -15, -10, 15, -23, -23, -5, -2, -23, 36, 13, 10, -4, -43, 21, -4, 21, 10, -15, -47, 28, -14, 13, 13, -13, 5, 15, 18, -3, 0, 7, 4, 33, -12, 30, 24, 40, 7, 6, -8, -32, -48, 4, 15, 4, 31, 10, 11, 4, -33, 2, 41, -15, 24, -56, 5, -32, 21, 10, 0, 10, 12, 32, -10, 4, -9, -11, 23, 18, -30, -41, 5, -33, 14, -5, 21, 10, -5, 35, -4, -21, 68, -48, -41, -1, 9, 2, 4, 5, 43, 11, 47, -22, 28, 7, 21, 8, -44, -28, 29, 19, 40, 15, -4, -25, -3, -1, 6, 7, 76, 45, -14, -1, -16, 10, -40, -1, 1, -62, -23, -23, 27, 31, 25, 12, 0, 24, 3, 3, 5, -3, -3, -22, -60, -9, -9, -106, 15, 22, 1, 12, 23, 31, 5, -55, 44, -89, -31, -45, -3, -32, 5, -19, 30, 11, 14, -27, 0, 19, 2, -11, -6, -3, 51, 4, -78, 10, 4, -64, 22, 23, -19, -4, 4, 10, -9, 22, 0, -10, -6, 10, 16, -2, -65, -41, 3, -3, 2, -50, 23, 49, 46, 4, 1, -13, -1, -27, -49, -26, 10, -38, 22, -13, 16, -5, 17, 14, 7, -59, 9, -37, -12, -12, -22, 28, 10, -15, 55, 43, -18, 0, -2, 4, 12, -9, 5, 28, 62, -14, -14, 19, -11, -55, 2, 9, 1, 0, 57, 19, -28, 10, 35, 4, 20, 11, 15, -10, -5, -2, 13, -13, 16, 31, -3, 36, 36, 8, -4, -11, -4, -2, -5, 11, -5, -53, -12, -21, 12, 23, 23, 11, 0, -29, -4, -19, -25, 31, 2, -11, 20, -16, 24, 28, 25, -10, -14, 40, -4, -13, -21, 27, 45, 10, -7, 1, -7, 3, 12, 14, -17, 3, 73, 3, 0, -2, 26, -3, -60, 3, 7, 3, 19, -25, 7, -17, 33, 36, 4, 4, 9, 7, 0, 5, -44, 27, 30, -67, 1, -2, 31, -37, -8, 35, 38, 1, 11, -10, 51, 44, 10, 31, 8, 15, 50, 1, 3, 6, 38, 31, -14, -18, -12, 2, 49, 13, -15, -3, 23, 7, -6, -1, -14, -8, -12, 5, 53, -2, -2, -53, 5, 7, 31, 28, 7, -3, 0, -31, 4, 10, -1, 18, -77, -13, -6, 7, 0, -6, -1, 9, 5, -73, 9, -18, 8, 8, -18, -5, 21, -17, -11, 29, 13, 2, -59, 16, 6, 47, 0, -17, 13, 31, 54, 19, 22, -12, 3, 15, 29, 32, -25, -18, 13, -1, 4, 26, -14, -41, -4, -2, 24, -34, -11, 14, -73, -13, 10, 11, -14, -18, 19, 0, -3, -36, -7, 20, -25, 32, 26, 7, -3, -6, 4, 4, 6, -43, 4, -4, 3, 8, 32, 8, -13, 20, -11, -26, 42, 2, -47, -2, 0, -13, 34, 1, 24, 43, 26, -2, -8, 9, 24, -5, 28, 54, 24, -14, 36, 16, 5, -2, 20, -3, 14, -11, 8, 13, -10, 10, -14, -12, 21, 6, 5, 14, 3, 18, 7, 1, 22, 18, -18, 19, 35, -1, -9, -39, 37, -11, -44, -4, 10, -23, 2, -14, -7, -6, -23, 21, -11, -17, 33, -6, -24, -14, -6, -10, 21, -34, -2, 32, 22, 17, -14, 46, 18, 23, -37, -84, 35, 7, 12, 1, -7, 5, 25, 7, 16, 2, 38, 6, 12, 19, 0, 7, 8, 3, 16, -6, -21, -8, -9, 21, -1, 24, -23, 16, 13, -1, -2, -19, 50, 21, -19, -8, 7, -61, -26, 19, -2, 12, -24, 8, 7, -92, -8, -29, 37, -48, 19, -63, -3, -30, -46, 12, -21, -37, 2, 20, 28, 23, -19, -49, 39, 57, -9, 17, 0, 4, 21, -14, 17, 2, 28, -7, 7, 32, 27, 5, -17, -11, -43, 32, -19, -21, -25, 1, -12, -10, -5, -13, -3, 3, 1, -35, 26, 19, -40, -40, 2, -31, 9, 21, 28, -5, 7, 8, 7, -90, 9, -28, 7, -4, 12, 0, 9, -11, 4, 54, 2, -4, 13, 13, 31, 20, -3, -78, 46, 18, 14, 23, 3, -34, 27, -17, 24, 0, 53, 8, -9, -8, 37, -6, 46, -12, 7, 67, -1, -21, -20, 1, 16, -3, -9, 11, 15, 4, 1, -2, -46, -12, -6, 4, -6, -29, 41, -40, 12, 13, 14, 1, -9, 2, -6, 5, -30, -3, -11, 0, 23, 2, 27, 54, 19, -16, 3, 11, 19, -32, -18, -3, 25, 15, 20, 10, -10, -1, 7, -3, 2, -3, 48, -19, 5, 17, 31, 0, 24, 3, 34, 40, 0, -4, 7, 11, 11, 33, -12, 7, 16, -1, 14, 29, 4, 18, 27, -53, 9, 22, 22, -52, 0, 17, 7, -1, -2, -1, -2, 23, 18, 7, 12, 7, 2, -49, 44, 0, 27, 22, 30, -22, -1, 1, 31, -17, -13, 24, -11, 2, 4, 9, 17, -19, -19, 4, 0, 18, -5, -40, -34, 5, 2, -4, 40, -4, 15, -31, 27, 10, 2, 27, -38, -39, -24, -6, -9, 14, 12, 15, 5, -60, -6, -8, -3, -17, 21, 0, -42, 15, 7, 22, 39, -2, -69, 28, 13, 26, 39, -11, 18, -14, 30, 0, 28, 9, -8, 6, 17, -5, -2, 11, -15, 7, -10, 31, 41, 19, -5, -8, 42, 9, -15, 7, -66, 8, -5, -27, -27, 19, 2, 43, 0, -10, -24, -1, 3, -7, 52, -7, -5, 12, -1, 16, 17, -40, -9, 9, 15, -18, 13, 0, -3, 28, 0, -8, 1, 31, -61, 32, 24, 43, 48, -27, -24, 30, 13, -13, 23, 6, 2, -21, 20, -4, 31, 16, -33, 13, 2, 15, 38, -11, 8, 8, -4, -24, -6, -1, 9, 0, 40, 28, 13, 5, 29, 23, -3, -72, 10, 11, -33, 20, 31, 8, -12, -8, 51, 23, 4, -43, 2, 40, 29, -7, 11, -21, 1, -13, 1, -39, 32, 31, -25, 21, 23, 6, 16, -57, -6, 53, 10, 11, -5, 30, 1, 7, 20, 21, -1, 43, -33, -8, -8, 41, 33, -2, 26, -11, 49, -28, 35, 8, -17, -12, 10, 1, 0, 7, -7, 16, -4, -27, -16, 15, -39, 0, -2, -4, 0, -39, 23, 10, -16, -18, -7, 32, 11, -6, -2, 5, 13, -11, -5, -15, 33, 0, 0, -10, 17, -80, -29, -30, -88, 14, -3, -41, 24, 13, -13, 24, -3, -23, -3, 6, -3, -2, 6, 9, 9, -27, 38, 5, 39, -13, -1, 17, -38, 6, -50, 28, 3, 16, -37, -36, -19, -42, 11, 15, -31, -16, -33, -7, 9, -39, 57, 15, -7, -35, 1, 39, -18, -1, 52, 0, -12, -4, -3, -45, -9, 30, 33, 14, 8, -39, -17, -29, 3, -6, -5, -13, -4, -12, -10, 19, 6, -17, 21, 16, -17, 10, -10, -7, 25, 22, 27, -3, 33, -30, -24, 7, 31, 6, -29, -37, 21, 4, 11, -46, -43, -2, 15, 8, -53, -11, -29, -11, 9, -13, 32, 30, -8, -50, -8, 8, -1, -61, 29, -4, -5, -5, -6, -34, 5, -1, -6, -2, 19, -1, -8, -45, -19, 13, 40, -40, 16, 29, 3, 30, 7, -27, -12, 22, 0, 8, -13, 26, 20, -5, 3, 8, -19, -19, -7, -15, -9, 6, -12, 30, -16, 5, 39, -1, -17, 2, 9, -8, -42, -9, -7, 10, -2, 19, 0, 20, -12, -38, -5, 36, 9, -58, -11, 17, -14, 2, 6, -10, -13, -8, -18, -1, 27, 3, 39, -9, 26, -9, 17, -14, 15, -25, 4, 5, -16, -7, -19, 16, -24, 5, -7, 22, 15, 5, -13, 0, 3, 21, -9, -41, -43, -3, 12, 8, 34, -42, 22, 7, 16, 23, 24, 0, -26, -49, -12, -3, -14, 8, 6, 2, 8, -32, 5, 11, -11, -11, -21, 12, -20, 32, 0, -34, -5, -9, -66, -7, 35, 6, 55, 18, 28, -42, 48, 1, 26, 54, -3, -19, -28, 9, -10, -56, -65, 8, 6, -15, 50, -3, 11, -1, -6, -17, -19, 7, -84, -5, 35, 9, -12, -10, 7, -4, 7, -73, 13, -6, 12, -5, 39, -1, 8, 24, 46, 26, 21, -46, -3, 5, -12, -26, 34, -3, -17, 7, -12, 8, -4, -17, -67, 25, 22, 11, 42, 4, 1, -10, 0, -1, -10, 55, 20, -14, -10, 3, 5, -14, -62, 23, 5, -16, 44, 4, 23, -12, 18, -28, -18, -5, -75, -8, -39, -5, -3, -4, -8, 2, -4, -21, 4, -32, -17, 5, -2, 2, -12, 7, 25, 10, 22, -71, -2, 16, 6, -5, 8, 7, -18, 21, -11, -11, 21, -5, -58, 0, 20, 9, 9, -19, 17, 4, 4, 16, 8, 28, 10, -2, 20, 39, -10, -22, -30, 26, -12, 38, 19, -28, 27, 3, -22, -12, 15, -1, -68, -5, 4, -5, -12, -1, 8, 13, 3, -64, 17, -23, -23, -11, 3, 11, -3, -3, 22, 14, 26, -22, -10, 3, 12, -27, 4, 32, 4, 2, -1, -65, -1, -6, -71, -4, 15, -14, -2, -49, -35, -23, -19, -11, 10, -2, -5, 2, -13, 0, -14, -9, -25, 28, 8, 13, 44, -42, 52, 8, -19, -25, -5, 25, -71, -7, -13, 6, 15, -4, 12, -15, -1, -36, 21, -19, -52, -18, -8, -7, -3, 23, 17, -9, 20, -40, -18, 33, -10, -40, 11, 14, -31, 0, -18, -57, 12, -42, 8, 10, 4, -55, -9, -47, -42, -12, -8, -1, 20, 22, 27, -8, -13, -19, 2, -28, -20, 21, -5, 28, 11, -46, 32, -2, 3, -28, 3, -24, -60, -3, 30, -24, 16, 27, -6, 3, 0, -34, 14, 9, -43, -21, -10, 2, 0, 13, -4, 21, 14, -25, -9, 2, 3, -68, 44, 20, -10, 18, -8, -52, 26, -20, -41, -5, 34, -27, 31, -23, -6, -20, -5, -11, 0, 14, 8, -6, 16, -5, -15, -7, -9, 11, 2, -5, 25, -22, 37, 4, 10, 21, 2, -31, -29, -9, 3, 35, -3, -19, -7, -5, -2, -38, 3, -13, -27, -23, -29, 1, -12, 21, -33, 25, 4, -21, 0, 10, -13, -25, -23, 33, -40, 8, 10, -29, 38, -36, -57, -9, 23, -16, 53, 10, 37, -58, 7, 2, -30, -4, -3, -34, -32, 29, -9, 41, -73, 32, 4, 0, 30, -10, 6, 5, 0, 2, 13, -11, -48, -1, 29, 3, 1, -38, 4, 27, 17, 4, 20, -24, 13, -22, -38,
    -- layer=2 filter=0 channel=5
    0, -4, 10, 38, -19, 17, -45, 5, 1, -51, 57, -50, 24, -35, -10, 4, -42, -14, 5, 37, 6, -22, -37, -25, 3, -77, 24, -57, -37, 1, 4, 10, 22, -15, 14, -1, 18, 0, 11, -5, -8, 26, 16, 7, 8, -35, -11, 2, 21, 60, -10, -28, -25, -25, -2, -5, 8, 11, -21, -50, -20, -28, 32, 41, 2, -8, 0, -45, -17, -22, -6, 8, -35, -4, 22, -4, 8, -5, -19, 3, 24, 26, -9, 13, 5, -26, -27, 37, 36, -17, 22, -7, -5, -31, 13, 17, -31, 2, -22, 3, 27, -17, -8, 12, -10, 15, 45, -22, 1, -5, 32, -25, 41, 60, -8, -20, -37, 2, -11, -5, 18, 8, -29, -34, -11, 6, 7, 20, 8, -7, 0, 5, -4, -36, -7, -6, -18, 0, 51, 22, -14, 15, 22, -2, -20, 6, 28, 34, -7, -24, -34, -20, -20, 18, -36, 12, 22, -17, 7, 28, 4, 22, 98, 20, -2, -6, 4, 3, -5, 5, 20, -6, -4, 0, 0, 11, 38, 20, 3, 51, -3, -5, -38, 5, 24, 16, -51, 2, 17, 11, 13, 36, 3, 0, -20, 23, -14, 11, 0, -5, -13, 50, 17, -20, -4, 33, 22, 8, -32, 0, -1, 33, 37, -31, -8, -3, -2, 25, -11, 2, -7, -67, -8, 28, 26, 10, 21, -10, 5, 22, -15, -11, -9, -25, -7, 1, -11, -27, -2, 17, -12, 23, -6, -9, 14, 21, -57, 0, -15, 53, -3, -48, 26, 5, 52, 46, -5, 20, 0, 14, -35, -24, -8, -5, -12, 14, -3, 8, 7, 38, 11, 5, 1, -2, 5, 2, 24, -21, -42, 22, 7, 34, -30, -22, 0, -6, -20, 21, 20, 12, 29, -9, 24, 1, 11, -3, 0, -12, 8, -25, -3, -4, -21, -7, -28, 14, 5, 33, 41, -26, -6, -15, -10, 26, 58, 2, 9, 6, -17, -7, -2, -4, -10, 44, -32, -2, 48, 10, -14, 3, 3, 33, -6, -32, -16, 2, -25, 8, -5, 39, -2, -8, -44, 12, 10, 37, -14, 0, -3, 14, -7, 0, 42, -51, -11, -2, 38, 16, -1, 6, -20, -52, 30, -7, -1, -12, 31, 0, -33, -14, -3, -1, -34, -14, 10, -13, -5, 8, 87, -33, -29, 13, 29, -22, -10, -1, -9, 31, -10, 23, -14, 0, -10, 12, -21, -3, 0, -55, 15, 1, -54, 34, 4, 15, 11, -11, -42, -29, 27, -4, 12, 26, -2, 4, -15, 11, 50, -12, 18, 8, -3, 41, 10, 9, -4, -7, 26, 0, 4, -4, 14, -15, -54, 37, 0, -7, -31, -11, 8, -30, 0, 11, 56, -33, -25, -3, 47, -20, 5, -2, 24, 25, -28, 25, -39, 2, -6, -7, -1, -12, 15, 7, -32, -6, 34, -30, 18, 23, 17, 2, 26, -10, -2, -5, -18, -26, -19, 5, -36, -15, 2, -33, -21, -30, 46, -9, -20, 0, 4, -10, 2, -15, -2, -2, -25, -32, 4, 34, 8, -19, -28, 50, -1, 4, 9, -34, -14, -15, -4, 16, 3, -20, 5, 8, -16, 5, -16, -14, -28, -1, -42, -13, 56, 4, 2, 29, -23, -4, 3, -15, -7, 35, 30, -4, 39, -6, -7, -36, -15, -18, -26, -29, 9, 16, -14, 7, 51, -16, 8, -20, -14, 2, 6, -16, -13, -11, 4, -7, -24, -7, 32, 22, 6, -20, 4, 20, -73, 1, -15, -5, -19, -9, -8, 12, 33, 44, -3, 7, -33, 7, -16, -37, 20, -4, -5, 29, 17, -15, 16, 43, 36, 2, -11, 36, -31, 43, 12, 15, -7, -10, 9, -22, -17, -10, 33, -29, 5, 17, 4, -6, 9, -10, 10, -10, 17, 0, -19, 16, 34, -12, -1, 3, 0, 4, 51, 3, -5, 33, 28, 14, -66, -20, -6, 18, -28, 17, -1, 27, -6, 51, -3, 9, -21, 7, 23, -8, -22, -11, 13, 39, 45, -19, 27, 32, 59, -11, -7, 20, 3, 25, 26, 48, -54, -6, -2, 37, -10, 45, 37, 11, -1, 19, 0, 34, 3, 14, 46, -8, 30, -9, -41, -19, -10, -32, -1, -44, 2, 43, 20, 5, -8, 31, 48, -3, -56, -6, -8, 13, -36, 14, 1, -3, 30, 25, 2, -1, 11, 28, -15, -5, 7, 7, 5, 11, 7, -5, 6, 39, 35, -8, -28, 39, -33, 7, 25, 20, -49, -3, -7, 21, -16, 39, 16, -29, -8, 17, 0, 13, -14, 8, 21, 3, 22, 8, -6, 13, 15, -26, -7, -39, 7, 40, 0, 5, 2, 48, 26, 9, -49, 16, -3, 25, 42, 24, 0, 17, -9, 40, 0, 5, -3, 46, -13, 5, -6, -3, -35, -4, 1, -4, 3, 11, -2, -4, -20, 15, -10, 10, 40, -2, -48, -37, 20, 32, 0, 20, -3, -3, 6, 9, 26, 21, 3, 2, 34, -19, -1, -1, -19, -13, -8, -12, -8, 10, 10, 16, -42, -5, 1, 18, 7, -32, -45, -19, -28, 3, 59, -2, 4, 7, 4, -20, 5, -2, -20, 56, 8, 18, -15, -1, -9, -27, -20, 23, -1, -20, -5, 4, -65, -31, 8, 21, 20, 19, -3, -22, -3, 14, 2, -2, 15, 3, 21, -2, 17, -21, 17, -9, 8, 5, -4, 5, 0, -3, -9, 0, -3, -11, 25, -36, -57, 5, -11, -34, -30, 6, -15, -13, 6, -28, 31, -8, -31, -11, 24, -3, 4, -11, 29, 23, -40, 25, 0, 5, -12, -37, 6, 6, 14, 4, -14, -13, -7, -40, 4, 32, -4, -14, 7, -29, -14, 0, 4, -33, -31, -15, -4, 4, 10, -26, 20, -6, 31, 14, -6, 0, 3, -23, -1, 4, -5, -15, -22, 4, -12, 6, -7, -2, -16, 44, -31, 10, 30, 30, -48, 6, 12, -5, 13, -2, 5, 7, -11, 34, -1, -14, -1, -8, -20, -4, 24, 0, -5, 30, 32, 1, 31, -20, -15, 7, 41, -20, -9, -30, -16, -30, -13, -42, 1, 17, 7, -17, 2, -29, 36, -2, 3, -8, 5, -7, 0, 4, -40, -6, 0, -22, -19, -32, 29, 30, -12, 0, -8, 0, -76, -24, 2, -17, -23, 5, 2, -33, 35, 12, -7, -9, -41, 17, 19, -40, -7, 0, -11, -11, 0, 1, -7, 2, 27, -12, 38, 24, -1, 9, 12, 13, -61, -4, 7, -39, -14, 7, -5, 52, 6, -13, 4, 41, -17, 17, 4, -22, -4, -2, -20, -12, 0, -53, -3, -24, 9, -38, 38, 23, 6, -10, -8, -17, -26, -9, -14, -45, -37, 49, -5, 0, -30, 30, 2, -4, -26, -14, -1, -82, -13, 9, 20, 0, 2, 40, 9, 19, 13, -8, 55, 4, -31, 2, 0, 18, -36, -8, -10, 0, -34, -18, 8, 24, 0, -6, -6, 60, 1, 3, -12, -30, 5, 8, -28, -6, -22, -50, -9, -57, -18, -54, 49, -7, 0, -18, 11, 38, -3, -40, -55, -33, -10, 39, -38, 8, -31, 4, 0, 10, -9, 25, -4, -26, -2, -5, -6, 14, -11, 46, -15, 14, 20, 8, 16, -8, -63, -5, -12, 11, -51, 0, 17, -25, -60, -24, 18, 7, 16, 0, 2, 73, -22, 3, 26, -22, 16, -5, 5, -4, -40, -31, -6, -30, -14, 20, 15, -1, -8, -16, -2, 14, -25, -25, -31, -6, 40, 35, 3, 2, -32, -19, -4, -8, -20, 35, -1, -18, 0, -2, -18, -4, 1, 18, -10, -28, 27, -4, 4, 6, -38, 6, -24, 6, -42, -44, -22, 57, -17, -6, 7, 12, 8, 6, 28, 33, -21, 10, 10, -10, 2, 7, -6, -6, -67, -2, 0, -2, -15, 9, -13, -42, -2, -13, -7, 45, -40, -25, -9, -18, 16, 12, -19, 11, 12, -43, 2, 7, -1, 26, -17, 19, -10, -4, -32, 6, -2, 9, 4, -2, -3, -8, -57, -17, -3, 32, -6, 3, -31, -10, 1, -1, 36, 0, 11, -18, 36, 18, 40, -13, -6, 7, -4, 4, 22, 7, 16, 3, -57, 2, 0, 36, 18, -18, -25, 54, -13, -55, 5, 22, -47, -7, 10, 0, 0, 15, 2, -17, 32, -19, -12, -7, 22, 25, -44, 11, -5, -11, 7, 16, -21, -27, 8, 1, 3, -1, 19, 6, 17, 17, -16, -2, -32, -5, -26, 24, 8, -43, -18, 4, -22, -22, 0, -42, 13, -8, 25, 14, -12, 0, 21, 7, -16, 4, 6, 11, -42, 25, -16, 6, 3, -31, -15, 12, 27, -10, 21, 11, 11, -21, 13, 2, -3, -18, -5, -6, -35, 29, -7, -24, -16, 4, -45, 30, -19, 39, -19, 18, -16, 4, -14, -21, -31, 23, -17, 5, -2, 16, -48, 38, -8, -26, -22, -49, 15, 3, -3, 47, 10, 4, 13, -26, -7, 5, -4, 22, -57, 21, 2, 5, -31, 1, -6, 0, -7, -6, 6, 12, -73, -32, -1, -23, -19, 11, -19, -24, 20, -5, 8, -7, -52, 10, 13, -33, 10, 9, -39, 15, 6, 9, 5, 25, 14, 1, -6, -26, -40, -21, -38, -11, -6, -17, -43, 0, -25, -36, 7, -6, 25, -11, -11, -13, 19, 22, -2, -2, 5, 0, 15, 29, -43, -7, -9, -36, -36, -19, 16, 27, 0, 37, 28, -25, 32, -49, -47, -33, -39, 32, -7, -23, 30, -16, 1, 7, -29, 10, -1, -63, 3, 6, -21, -37, 10, 10, 16, 24, -13, -1, 59, -14, -31, 29, -44, -6, -34, -50, -7, -24, -21, -9, -6, 20, 4, -20, 16, 63, 19, -14, -1, 18, 3, 7, 7, 25, 15, -28, -8, -39, -20, -47, 36, 19, -3, -3, 15, 1, 31, 0, -81, -41, -3, 6, -50, -10, -71, 10, 1, 6, -18, 38, 14, -51, 3, 5, -24, -3, -8, -1, 0, 3, 6, 2, 6, 15, -3, 2, 9, 6, -34, 11, -1, -13, 2, 29, 18, 5, 15, -11, 28, 10, -9, -8, 4, -8, -8, -11, 0, -4, -44, 0, 8, -17, 20, -1, 1, 4, 14, -4, -1, -16, -8, -21, -65, -48, 8, 7, 17, -19, -6, -29, 2, 2, -28, 31, 6, -35, -37, 9, -15, 22, -16, 19, -6, -8, 11, -8, 43, 7, 9, 18, -27, 3, -10, -30, -33, -37, -2, -46, -13, 2, 20, 27, -5, 32, 26, 21, 10, 21, 12, 7, -14, -3, -57, 7, 1, 5, -2, -15, -4, -5, 5, 27, 17, 66, 12, -20, -10, -10, 4, 9, 0, -34, -24, -51, 5, 4, 5, 17, 6, 29, -22, 0, 9, -14, -2, 24, 1, -26, -19, 4, 4, 0, -12, 19, 31, 0, -25, -48, -5, -88, 25, -14, 0, -5, -1, 4, 25, -45, 7, 4, 16, 7, 25, 2, 25, -25, -19, 4, 6, 14, 42, 9, -21, 7, 0, -62, -16, 71, 8, 17, 8, 4, -38, -6, 17, -26, 7, -37, -4, 8, 21, 7, -18, 11, -8, 1, 2, 12, -23, -9, 12, 3, -6, -1, 5, 5, -10, 44, -6, 22, 13, -24, -56, -43, 21, -14, -5, -30, 17, -2, -2, -26, -24, -12, 19, -14, -4, 1, -11, 2, -10, -8, -6, 25, -15, 42, -17, -3, -3, -37, 2, 31, 8, 15, 28, 11, -15, -11, 2, -31, 34, 19, 8, -6, -6, 15, -2, 9, -8, -7, -24, 14, 6, -16, 19, 39, -17, 3, 5, 5, -11, 22, 19, 11, -2, 7, -31, -22, 19, -5, -8, -12, 16, 0, 6, -24, 41, 19, -9, 22, 0, 1, -9, 25, -55, 36, 7, -2, 2, 6, -3, -14, -10, 15, 15, -21, -53, -7, -5, -32, -13, -2, -6, -34, 11, -24, -12, -4, -79, 30, 7, -11, -23, 10, -6, 0, -12, 50, -5, 39, -16, 4, 2, -10, -17, 18, -3, -4, -26, 4, -20, -7, 23, -18, -11, 21, 5, 2, 21, 4, 36, 10, -35, -7, 8, -2, 12, 42, -26, 36, 0, -2, -1, -17, -1, -45, 0, 9, 17, 25, 10, 10, -3, -9, 0, 59, 21, -73, -11, -29, 3, 6, -62, -5, 11, -23, -34, 9, -19, 34, -21, 27, -15, 29, -17, 4, 27, 31, -9, -26, 2, -18, -25, 28, 1, -17, 43, 0, 5, 3, -10, -15, 8, 3, -34, 16, -28, 5, 3, -1, -1, -24, -22, 6, 7, 10, -21, -5, 7, -6, -3, -28, 25, 1, 19, -8, -40, -51, 10, 23, -16, -30, -30, -45, -1, -1, -49, 27, -6, -34, -32, -6, 12, 11, 0, 24, -16, 67, 16, 6, 7, 34, -29, 12, -25, -2, -30, 19, -24, -29, -26, 10, -12, -27, 28, 0, -9, 11, -22, 19, -8, 21, 10, -9, 15, 6, -61, 17, -6, 11, -16, -3, -4, -15, 7, 5, 36, 0, -25, -13, -36, -24, -12, 5, 21, -34, -4, -9, 4, -1, -40, 42, 10, -19, -33, 1, -11, -2, -1, 2, -8, 13, 2, 1, -5, -1, -21, 35, 20, 0, -4, -27, -30, -32, 16, -39, -11, -31, 0, -8, 18, -2, -9, 28, 6, 36, 28, 8, -6, 2, -82, 39, 0, 4, -11, 25, -31, -11, -4, 0, 17, -4, -59, -15, -20, 0, -15, -8, 3, -38, -45, -12, 4, -2, 8, 33, -7, 33, -5, 1, 19, 2, -4, -11, -9, -41, -31, -4, -53, 32, 29, 37, 37, -7, 47, -42, -1, 9, 60, -5, 5, -31, 13, -16, 34, -47, -24, -17, 12, 29, 7, 6, 6, -2, -43, 6, 9, 14, -1, -4, -30, 21, -1, -38, -19, 23, -73, -5, 3, 0, -10, -17, 15, 4, 1, -48, 6, 0, 31, 21, 9, 20, -10, -8, -6, -17, 27, -42, 3, 14, -4, -3, 20, -22, 28, 46, 4, 17, 32, 23, -11, -13, 19, -55, -32, -37, 29, -5, -9, 0, 19, -48, 28, -33, -10, 9, 10, -1, -39, -2, -8, -12, -20, 18, 12, 71, -7, -2, -20, 40, -22, 6, -17, 16, -15, -41, -14, 0, 8, 26, -13, -2, -18, 17, 2, -23, -10, -1, -35, -23, 21, 22, -14, 25, 12, 7, 28, 7, -9, 51, 1, -22, 18, -52, -18, -27, 11, -14, -2, -15, 24, 3, 18, 23, 7, -11, -6, -23, 0, -13, -5, 5, -21, -10, -10, -11, -39, 11, -5, 4, -2, 54, 5, -13, -4, 12, -20, -12, 12, 8, -21, -18, -18, -3, -6, -14, -28, -15, 10, -28, -33, 6, -2, -11, 1, 26, 8, 46, 10, -7, 55, -6, -9, 32, -15, 16, 4, -26, -29, 23, -19, -35, 8, -5, -19, 9, 5, 18, -52, 21, 1, -37, 5, -8, -4, -10, -46, 15, 0, -21, -26, 8, -20, -6, -5, 1, 10, 16, 0, 0, -4, -37, 16, -5, 15, -18, -70, -50, -10, -2, -39, -21, -5, -16, -11, -4, -7, 15, -21, 25, -27, 20, -16, -14, 8, 2, -18, 15, 20, -6, -22, 2, -4, -11, 18, -21, -42, -1, -29, 3, -15, -35, -32, 27, -7, 5, -16, 0, -22, 0, -12, 0, -11, -16, -30, -7, -10, 8, -9, -13, 27, -18, 26, -18, 5, -14, 31, -16, -4, -16, -32, -14, -7, -4, -37, 9, 7, -6, -40, 3, -32, -17, -9, 18, -31, 38, -6, -11, 53, 52, -51, -6, -32, -6, 6, -21, -52, -42, -7, 9, -16, -15, -12, 8, -4, 4, 15, 7, -60, 0, -13, 7, -15, 16, -14, -4, 4, -28, -10, 28, -2, -5, 0, 11, 4, -6, 39, -12, -2, -33, -16, -6, -36, -18, -48, 6, 7, -12, -26, 37, -7, -6, -38, -4, -27, -2, 7, 1, -12, 21, 20, 7, 38, -8, 0, 34, -12, 9, 17, -29, -48, -41, 7, -31, -6, 2, -2, 8, 23, -10, 0, 22, -41, -2, 8, -3, -23, 5, 8, -3, 1, 5, -25, 16, -19, 27, 6, -30, 31, 0, 28, -17, 5, 2, 21, 7, -29, -36, -11, 1, -4, 0, 14, 4, -22, 22, -27, 5, -15, -23, -6, -18, 3, -30, -11, 0, -5, 6, -2, 30, 2, -6, -12, -21, 3, 43, 0, -30, 13, -28, -13, 1, 40, 11, -11, 1, -25, 21, 7, 0, -7, 27, -7, 8, -7, -3, -36, 3, -17, -9, 4, -34, -44, 35, -1, -8, -22, 8, 28, -18, 9, -15, 3, -29, -2, -1, 18, 26, -15, 9, -15, -5, 41, -27, 14, -18, 3, 21, -14, 2, -31, -16, 18, 24, 6, -43, 3, -8, 17, 3, 40, -42, -7, 5, -1, -14, -10, -36, 30, -67, -21, 35, -25, -11, 28, 1, 26, 7, -3, 7, -9, 9, 6, 16, 0, -26, -25, 19, -14, 66, 43, 6, -3, -44, 17, 7, 28, 46, 6, -7, 15, 30, 2, -13, -22, 4, 1, -26, -26, -16, 7, 21, 11, 1, -22, -5, 14, 41, -5, -36, 10, -46, -50, 30, 17, -46, 14, -35, -15, -3, 6, -10, -12, -18, 18, -8, -24, -12, -1, 24, -1, 8, -1, -2, -42, -14, -18, 35, -1, 33, 1, 46, -2, 30, 4, 3, 3, -15, 30, -40, 0, 29, -12, -12, -9, 0, -17, 24, -19, -1, -1, 13, 1, 28, -4, -3, 3, 3, 40, 51, -13, 14, 31, -15, -38, 8, 10, -55, 20, -39, -10, -14, 0, 29, -20, -31, 10, 8, -8, 3, 27, 6, -33, 25, 1, 18, 8, 40, -21, -10, 15, 28, 0, -36, 3, 1, -12, 16, 21, -5, 26, -18, -3, -47, -27, -12, 5, 8, -3, 34, -7, 4, -52, -7, -21, 14, 2, 42, 18, 28, -6, -4, 33, 30, -20, 52, 39, 14, 10, 37, -11, 19, 11, 26, -8, -10, -14, -11, 25, -34, -13, 9, -12, -15, -4, 1, -12, 15, 3, -16, 3, 33, 18, 63, 16, 11, -10, -22, 23, 27, -25, 14, 17, -26, 2, -43, -30, -18, -12, 0, 8, 0, -6, 47, -16, 14, -63, -6, -2, 1, -16, 47, -5, -22, -8, -6, 16, 13, 35, 23, 65, 12, 8, -3, -13, -4, 24, -1, 7, -14, -6, -1, -8, -24, 13, -6, -8, -25, 8, -7, -40, 18, 3, 11, -9, 9, -19, 17, 14, -14, 2, -5, -3, -11, 24, 19, -29, -15, 42, -16, -23, -14, 3, 11, 4, -6, -6, 46, 14, 13, -75, 5, 8, -35, 15, -5, -19, -24, 0, 4, 5, -4, 15, 44, 54, -7, 39, -10, -3, -60, 3, -17, -7, -3, 10, 5, 35, -15, -7, 8, -34, -12, 20, 0, -7, 20, -8, 4, -3, 22, -26, -6, -19, 16, -8, -5, -16, -6, 5, 11, 11, -6, 17, 11, -16, -25, -44, 0, 1, 7, 6, 24, 9, 20, -29, 9, -27, -13, 5, 4, 8, -9, -3, 4, 32, -34, 22, 15, 38, -21, 54, -20, -19, 6, 40, -44, 14, -58, 0, 0, 32, -44, -20, 3, -43, 64, 2, 0, -1, 0, 19, 25, 7, -1, 7, -10, -10, 6, -10, 24, -21, 0, 19, 26, 34, -7, 27, -32, 25, 10, 17, -13,
    -- layer=2 filter=0 channel=6
    -1, 16, 34, -52, 9, 12, -14, -5, -18, 0, 15, -32, 23, 19, 6, -3, -64, 0, 12, -39, 11, 1, -52, -27, -6, -110, 1, -30, -47, -12, -1, 6, -70, 19, -20, 36, -24, -17, 29, 7, -4, 3, 18, -7, -5, -37, -42, 0, 56, 15, 7, 31, 24, 17, -18, -21, 7, 6, 14, -15, -45, -3, -26, 14, -2, 4, 24, -63, 37, 15, 18, -4, -18, -11, -14, 2, 27, -1, 11, -4, -8, -28, 21, -61, 24, 25, -45, 0, -3, -61, -4, 6, -54, 51, 16, -12, -77, 29, -54, 27, -57, 0, 18, -7, -6, 45, -28, 39, 6, -29, -28, 17, 44, -22, 2, 31, -11, -10, -30, -13, 13, 2, 25, -6, -39, -6, 16, 32, 0, 2, 0, -10, -24, -5, 37, 3, -34, 7, -39, 0, -3, 6, -22, 4, 22, 8, 11, -21, 20, 15, -2, 23, 16, -23, -1, -20, -63, -34, -1, 6, -40, 36, 27, -6, -40, 2, 5, -2, 1, -10, -25, 17, 2, 1, 15, 2, 19, 14, -9, 38, -19, -1, 7, -33, -10, -17, 34, 0, -30, 2, -6, 9, -10, 22, 2, -41, 1, 3, -27, 10, -12, -6, -15, -8, 8, -19, -9, -1, 10, -1, -29, -13, -1, -14, -17, -13, 16, -18, 5, 11, -19, -19, -6, 4, 34, 34, -3, 1, -106, 35, 18, 11, 23, 10, -41, 13, -11, 21, 15, -4, 14, 6, 3, 26, -8, 0, 43, -13, -6, -24, 19, 20, -10, -30, -15, 3, 2, 0, 6, -52, -8, 5, 2, -6, -19, -19, 41, -16, -14, -13, 5, -12, -24, 8, -13, 6, 12, 11, -28, 23, -3, 0, -20, 6, -7, 24, -1, -4, -31, 33, -24, 12, -68, 3, 13, -7, -4, 30, -65, 0, -8, 20, -16, 0, 44, 12, 4, 20, -30, -17, 3, -16, 20, -12, 1, -4, 8, 5, -23, 43, -4, 17, 9, -26, 23, 14, 14, 2, 15, -13, -64, 3, -12, -2, 5, -12, -35, -1, 23, -19, 6, 11, -11, -23, 17, -20, 4, 3, -29, -49, -19, 1, 4, 3, -17, 17, -49, 12, 8, 2, 5, 40, -10, -5, -9, -5, 30, -50, -12, -33, -4, 55, 12, -2, 0, -3, 23, -24, 46, 0, 0, 2, -26, -34, 9, 5, 14, 22, 11, 19, 24, 3, -38, -6, -38, -14, -1, 10, 21, -6, -59, -60, -24, -30, 46, 11, -25, -36, 7, -18, 5, -13, -34, 4, -26, 16, 7, 19, -65, 30, -26, 4, 23, 3, 7, 40, -16, 24, -8, 3, 49, -6, -5, -5, -9, 0, 3, 11, 27, -4, -14, -27, 79, -7, -17, 0, -2, -8, -10, 11, -6, -40, 0, 6, 21, -6, -1, 21, 35, -17, -13, 21, -29, -6, 19, -23, 25, 3, 23, -30, -43, 10, -4, -51, 10, -51, 4, 6, -13, 8, -25, 2, -2, 29, -17, -9, -5, 11, 8, -14, -1, -7, 7, 42, -22, 18, 76, 26, 2, -6, 22, -7, -20, -12, 0, 1, 24, 10, -31, -6, -14, 24, -9, 2, -8, -75, -12, 2, 4, -5, -9, -44, 8, 8, 22, -28, 13, -3, 3, -52, 23, -7, 30, -27, -26, 4, -12, -43, -8, -38, 15, 9, -15, 0, -33, 38, -7, 4, 3, 22, 3, 0, 20, -13, 43, 15, 2, 22, 0, 25, 35, 13, 0, 15, -43, -7, 10, 13, -14, -2, 28, -8, 12, 4, -16, 36, -5, 2, 1, -99, -2, -18, -28, -5, -16, -19, -17, -19, 0, -59, 4, -4, -21, -45, 8, -86, 7, -17, -14, 15, -1, -25, -52, 6, -30, 29, -18, -11, -72, 34, -51, -17, -53, -30, 15, -8, 22, 23, 0, 11, 2, 15, 4, -11, -13, -15, -3, -25, -50, -34, -19, 26, 0, 8, 18, -6, -26, -5, 5, 27, 3, 0, 39, -64, -9, -9, -21, 2, -17, -3, -29, -30, 21, -63, 4, -11, -52, -8, 11, -48, 9, -54, -3, 21, -15, -28, -40, -11, -35, -54, 43, 17, -31, 34, -24, -13, -117, 10, 1, 4, 3, -20, 6, 16, -2, 43, -2, 14, -6, 0, -4, 1, -24, -24, -60, 0, 24, 17, 41, 19, -4, 28, 46, 0, -1, 0, 4, -56, 1, -17, -15, 9, -35, -8, -86, -27, 5, -47, 21, 8, 6, -34, -9, -87, -36, 4, 17, -19, -18, 23, -52, -8, -27, -29, 8, 6, 1, 28, -16, 0, -120, -37, 0, 10, -37, -56, 9, 25, -3, 35, 4, -40, -59, -50, -11, -3, 5, -58, -33, -22, 50, 9, 9, 9, -21, 17, -16, 3, -4, 12, 3, -32, 5, 4, 8, 4, -2, -20, -40, -24, 11, -38, -2, -6, -34, -6, -2, -16, -44, 8, 27, -40, 4, -40, 0, -37, 20, -1, -15, -4, 14, -27, 14, 20, -59, 30, 6, -6, 2, -4, 6, -4, -13, 4, 14, -47, -22, 24, -3, -3, -24, -41, 9, 29, -3, 0, 20, 8, 14, 20, -21, -2, -10, 2, 20, -11, -21, 38, -15, 4, 17, 12, -37, -25, 0, 17, -4, 3, -28, -18, -21, -6, 26, -19, 43, -56, -22, -27, 39, -21, -15, -81, -43, 7, 25, -20, -34, -14, -7, 34, 25, 9, 25, 2, -37, 18, 0, -6, -2, 9, -14, -24, -13, -6, -16, -6, -8, 22, -17, -7, 36, 1, 27, 6, 4, 2, 9, 17, -24, -17, -22, -3, 6, 8, 16, 20, 19, -35, -12, 27, -15, -10, -28, 10, 8, -12, 7, -10, -86, 14, 0, -91, 8, -45, 16, 3, -18, -15, -30, 58, -35, 15, -14, 10, 2, 10, 58, 12, -16, -1, -1, 16, -47, 38, 33, 7, 4, -24, -14, -78, -2, -15, -12, -13, 48, 1, -33, -12, 6, -36, 6, 2, 18, -39, -10, -6, -18, 6, -27, -53, -7, -42, 7, -48, -3, -11, -71, -83, 15, 0, 13, -15, -57, 0, 24, -88, -60, -23, -1, -55, 0, 1, -25, -13, -27, -1, -59, -20, 12, -4, 7, -17, 16, 4, 8, 76, -37, 27, 30, 33, -7, 18, -38, -49, -3, 30, -42, -22, 91, 25, 24, 11, -46, 26, -8, 3, 29, -55, 21, -1, 3, -8, 13, -21, -25, -28, 8, -76, 12, 7, -69, -86, 10, -31, -15, -3, 68, 1, 0, -76, -53, -75, -37, 0, 31, 17, -20, -53, 11, 4, -72, -9, 10, -10, -11, 13, 37, 26, -13, 33, -22, 10, -20, -9, 10, -24, -20, -32, -14, 3, 18, 15, 29, 27, -9, 25, 13, 0, 8, -3, 51, -55, -3, 36, -28, -6, -44, -2, -45, -56, 28, -43, 29, 7, -116, -43, 0, -38, 22, -40, 71, -10, -11, -65, -13, -55, -13, -100, 49, 40, -18, -79, 24, -7, -165, 45, 30, 11, -22, 12, 14, 18, 0, 13, -5, 0, -49, -30, -9, -85, 10, -45, -109, -31, 37, 54, 46, 23, -48, 8, 58, -5, 1, -1, 41, -56, 0, 18, -13, 9, -56, -11, 0, -53, 46, -66, 13, -6, -49, -36, 33, -21, -20, -12, 44, 6, 6, -56, -54, -37, -71, -55, 29, 33, 38, -70, -8, 7, -75, -31, 30, 9, -15, 7, 24, 25, -11, -5, -9, -17, -8, 40, 3, 27, -4, -36, -5, -62, 23, 34, 9, 18, -18, -8, -21, -26, -2, 11, 21, -20, -15, 1, -1, -11, -30, -68, 35, -28, 27, -2, 8, -12, -66, -6, -18, 25, -25, -2, 59, -87, 0, -57, -56, -49, 8, -80, -4, -5, 29, -17, -26, -2, -39, 17, 28, -6, -12, -13, 1, 20, 5, -7, 7, -52, 23, 40, -7, -37, -34, -67, 42, 23, -30, -33, 30, 11, 31, 13, -65, 3, -8, 4, -21, -46, 27, 19, 14, 7, -1, -7, 5, -32, -5, 34, -3, -5, 20, -7, 32, 16, 37, 0, -32, -44, 21, -54, 7, -14, 21, -2, -25, -5, -3, -28, -4, 0, 23, 59, -21, 7, 31, 10, 6, 5, 0, -2, 8, -48, 36, 47, -9, 11, 17, -39, -4, 26, -22, -12, 15, 6, 13, 24, -9, -8, -1, 7, -33, -25, -11, 11, 2, 9, 22, -8, 17, -49, -11, 36, -18, 2, -8, 0, 27, -11, 23, -20, -95, -31, 3, -70, -5, -26, 21, 0, -37, -6, -12, 64, -11, -15, -28, 46, 1, -9, 36, -66, -8, -16, -5, -18, -26, 12, 44, 13, -13, 0, -5, -42, 4, -6, 4, -25, 18, 0, -4, -13, -9, -49, -8, 20, 17, 10, 17, 11, 33, -5, -2, -72, -19, -76, 14, -14, 10, -8, -18, -71, 19, 32, -28, -2, 3, -51, 10, -79, -38, -23, 22, -44, 6, 2, -10, 13, -40, 3, -74, -31, 16, -3, 21, -27, 27, 8, -12, 0, 6, 15, -9, 1, -4, -11, -20, -23, -4, 3, -76, -31, 46, 10, 42, 15, -58, -47, 4, 14, 50, -31, 23, 35, -1, 7, 13, -34, -26, -49, 25, -27, 14, -4, -22, -89, 9, 19, 14, 19, 4, -75, -14, -106, 42, -88, -2, -58, 33, 24, 2, -73, -3, 6, -80, -33, 21, -6, 14, 10, 42, 20, -10, -20, -3, 26, -48, -38, 1, -12, -9, -42, -18, 37, -51, -8, 37, -15, -12, 17, 32, -36, 8, 7, 85, -51, 27, 68, -38, -12, -36, 10, -13, -63, 63, -14, 27, 1, -47, -117, 14, -35, 9, -48, 0, -11, -26, -102, 40, -111, 13, -133, 5, 55, -69, -111, -9, 13, -119, 19, 37, -10, 2, -44, 10, 61, 0, 28, -32, 44, -33, 10, 3, -27, 0, -15, -70, 43, -38, 40, 24, 17, 4, 1, 50, -50, 0, 13, 69, -62, 2, 38, -20, 1, -34, -38, 20, -50, 37, -20, 33, 0, -54, -94, -10, -3, -35, -46, 0, -73, -30, -80, -25, -84, 0, -61, 17, 28, -9, -49, -42, 19, -26, 53, 37, 9, -4, -17, 20, 31, -11, -35, -67, 3, 1, 23, 5, -14, 12, -30, -44, -21, -19, 39, -3, 14, -4, -2, 6, -27, 0, 9, 22, -22, -2, 3, -24, -6, -21, -58, 43, -55, 40, 1, 7, -1, 0, -59, -10, 7, -29, -2, -11, -55, 26, -83, -51, -80, -6, -7, -7, -14, 13, -9, -34, -5, -29, 12, 1, -6, -33, 12, -1, 11, -7, -26, -34, -46, 26, 46, 6, 27, -14, -73, -6, -37, -60, -26, 25, 2, -20, 4, -39, -13, -3, 5, -24, -16, -29, 5, 31, -4, -9, -31, 18, -32, -13, 16, 4, 3, -36, -15, 10, 6, 1, -19, -11, -77, -4, -45, -26, -26, 27, -11, -10, -22, -12, 13, 2, 6, -31, 25, -9, -10, 36, 0, -8, 0, -11, 13, 0, -28, 14, 28, -5, -32, 9, -16, -13, 27, -20, -49, -1, -20, 41, 31, -15, 19, -6, 2, 0, -1, 15, 4, -24, -11, -7, -4, -7, 32, -29, 37, 0, 1, 21, -41, -15, 9, 37, 8, -15, -16, -9, -34, -9, -94, 22, 42, -17, -22, -8, 14, 14, 13, 23, -4, 3, 0, 34, -25, -11, 22, -8, 27, -10, 34, 0, -10, 8, 17, 4, -11, 49, 10, 0, -17, 50, 17, -4, -35, -11, -44, 7, 6, -12, -4, 2, -6, -9, -3, -28, -24, -8, -30, 12, -15, 19, 2, 11, -26, 1, 23, -13, 17, -56, -30, 11, -12, -48, -5, 10, 2, 14, -1, -15, 2, -39, 27, -62, -50, 18, 9, 1, -2, 6, 5, -4, 4, -32, 28, 10, 0, -7, 10, 28, -25, 28, -9, -9, -13, 36, 10, -5, 3, -12, -26, 2, 0, 40, 7, 19, 3, 24, -5, 42, -42, 20, -37, 11, -24, 28, -12, -9, -7, 32, 54, -21, 18, -9, -46, 46, -21, -8, 2, 9, -17, 11, 15, -13, -69, -18, -2, -93, -22, 21, -9, -13, -18, 10, -1, 8, -29, 7, -17, 6, -4, -1, 45, 17, -57, 25, 22, -59, 7, 34, 17, 0, 40, -11, -26, -9, 4, 26, -68, 8, 11, -6, -1, 12, -32, 6, -11, 34, 28, 23, -7, -47, -67, 33, -11, -12, 13, -21, -86, -9, -40, -19, -86, 59, -57, -32, 27, -71, -58, 15, 19, -47, -23, 36, -2, 24, 4, -49, 34, 0, -62, -26, -15, 14, -40, -6, 73, 26, -39, -36, 0, -41, 28, 15, 0, 76, -11, 0, -70, -6, 8, 39, -13, 2, -10, 3, -8, -3, -36, 38, -19, 29, 14, 15, -1, -5, -61, 58, -22, -22, -34, 13, -18, -2, -24, -16, -55, -4, 16, -15, 29, -28, -36, -14, 20, -31, 0, 22, -1, 27, -17, 9, 3, 6, -16, -35, -17, 69, 47, 1, -70, -17, 0, -47, 28, -41, 35, 23, -8, 42, 7, -15, 0, -7, -1, 15, -13, 15, 0, -5, -3, -11, -48, 14, -18, 35, -9, 10, 4, -14, -32, 33, 13, -4, -14, 39, -61, 18, -42, -16, -1, -10, -3, -12, 0, -3, -12, -40, 4, -56, 3, 22, -5, -18, 11, -9, 0, -4, -59, -43, -84, 40, 52, 0, 38, 13, -34, -2, 1, -36, 10, 18, 12, 0, 14, -20, 28, -9, -7, -5, -5, -2, -10, -27, -8, -10, -39, -2, 0, 15, 39, 39, 5, 3, -55, 0, -7, 2, -1, 30, -83, -15, -71, -6, -61, 29, 9, 12, -16, -1, -7, -31, 16, -32, 8, 5, -10, 3, 37, -24, 11, 8, -7, -49, -44, 44, -5, 3, -9, 14, -21, 79, -15, 3, -40, 24, 31, 11, -15, -12, -10, 1, 10, 10, 0, 12, 19, -7, -1, -21, 11, -29, 9, -6, 27, 1, -9, 32, -50, -8, 0, 33, 3, -28, -90, -48, -57, 13, -58, 10, 7, -31, -14, 13, -4, 10, 25, 12, 12, 20, -1, 0, -40, -33, -11, -11, -33, -61, -4, -12, -28, 0, 39, -4, -42, 19, -14, -25, -24, 45, 8, -15, -15, -10, -89, 3, 16, -1, 2, 10, -6, -26, 10, 4, -11, -23, -13, 7, -8, 35, 3, -37, -8, 35, 12, 38, 13, -37, -73, -33, -27, -23, -25, 24, -13, -23, -9, -30, -28, -46, 42, -56, 41, 20, -4, -28, -15, 15, -18, 0, -19, -27, 0, -13, -20, -1, -24, 22, -66, -11, 9, -2, -7, 75, 25, 27, 6, -6, -37, -10, -5, -10, -41, -12, -20, 6, -4, 1, -18, 0, -20, -12, 4, 21, -1, 1, -5, 7, 8, -8, -14, -55, -34, 20, -35, -13, -18, 7, 0, -28, 4, -20, 2, 25, 19, -63, -1, 17, -7, -13, -4, 26, -42, -10, -66, -14, -59, 30, 25, 3, -56, -16, -39, -20, 46, -2, -3, 73, 5, 21, 7, -36, 13, 1, 2, -27, -4, 10, -27, 1, 2, 3, -46, 20, 26, 10, -13, 18, 10, 1, -17, -31, 38, -6, 1, -21, -57, 18, -43, -73, -16, -30, 11, -28, 22, -17, 36, -24, 3, 4, -2, 13, 3, 0, -20, -4, -19, -11, -50, -16, -50, 37, 47, -7, -28, -23, -28, 30, 15, -30, 3, 39, 22, -7, 33, -32, -25, -6, 14, 6, 22, -3, -19, -6, 1, 10, 9, 12, 24, -3, -35, 17, -8, -12, -10, 26, 0, 16, 0, 7, -30, -3, -12, -40, -26, 19, -3, 20, -7, 15, -15, -49, 4, 11, -4, 15, -5, -24, -19, -15, -24, 1, -17, -14, -26, 56, 16, 0, 47, 13, -34, 52, -10, 20, 19, 47, -4, 28, 43, -15, 44, -8, 5, 5, -25, -1, -2, -15, -1, -9, -4, 26, -11, 17, -8, 22, -3, -20, 16, -7, 13, 16, 2, -52, -2, 12, -51, 14, -15, -27, -4, -16, 7, -13, 22, -21, 40, -20, -7, 20, 6, -10, -23, 0, 7, -3, -6, -3, -56, 35, 33, -2, -17, -12, -22, 31, 11, -3, -16, 1, 20, 4, 24, -25, 23, 0, 13, 10, -18, -2, 20, -26, 3, -44, -10, 21, -20, 8, -1, 23, -8, 18, 2, -5, -4, 43, -1, -10, -67, -38, -91, 19, -18, 8, -3, -1, 2, -8, 29, -26, 23, -34, 8, 30, -1, 6, -44, 0, -1, 4, 5, -39, -28, 62, 36, -5, -53, -4, -17, 6, 7, 21, -18, -36, 26, 8, -37, -2, 20, 4, 12, 39, -19, 31, 12, -9, 1, 18, -13, -23, 51, -21, 16, 31, -8, 45, 3, 27, -5, 27, 24, -39, -55, 2, -19, 0, -9, 33, -34, -19, 7, 6, 23, -4, 32, -31, 36, 23, -13, 28, 8, 30, -1, -5, -43, 9, -23, -9, -4, 0, 8, -19, -5, -14, -13, -7, -32, 55, 46, 0, -11, -39, -46, -6, -1, 17, -28, 9, 12, -29, -6, 33, 16, -18, -41, 4, 50, 20, 0, -36, 17, 0, 3, 0, -5, -40, -62, 1, -38, 25, -9, 42, 0, -51, 0, 29, -17, -12, 46, -46, 33, 13, -4, 12, 9, 30, -25, 0, 11, 8, -37, 11, -71, 6, 10, 23, -6, 43, -8, -7, -5, 46, 15, 6, 10, -27, -56, 1, 21, 0, -40, -10, 13, -17, -4, 10, -21, 8, -23, -5, 14, -4, 6, 1, -20, -24, -5, 10, -35, -14, -22, -8, -27, 34, -1, 24, -19, -52, 2, 5, -26, -34, 12, -24, 19, -1, -1, 16, -61, 34, -13, -4, 27, -5, -24, 16, 10, -14, -61, 0, -2, 22, 19, -7, -6, 44, 25, 12, 21, -47, 24, 8, 6, 20, -18, -26, 0, 16, -8, 3, 6, 7, -57, -14, 21, 17, -12, 44, -11, -6, 1, 27, -29, -8, -52, -24, -45, -4, -33, 30, -32, -25, 1, 3, -1, -13, 13, -92, 8, 4, 5, 11, -22, 42, -9, 3, -27, -39, -65, -1, 41, -13, -12, 14, -51, 2, 4, 24, -6, 45, 10, 20, 8, -30, -14, -11, 14, 5, -29, -32, -16, 21, 0, -7, 15, 10, -40, -15, 38, 13, -12, -19, -11, -29, 0, -9, -41, 9, -42, -2, -31, -26, -9, 33, -41, -18, 3, -28, -18, 10, 30, -77, 17, 11, -1, 32, -5, 10, -16, 0, 7, -6, -18, 32, 18, -3, -73, 37, -67, 8, 2, 33, 7, 13, -5, 36, 8, -33, 25, 0, 15, 29, -27, 10, 18, 6, 9, -15, 1, 39, -18, -6, 25, 16, 0, -35, -24, -25, 35, 25, -15, -29, -43, -27, -13, -4, 0, 45, -3, -9, 16, -42, 15, 17, 36, -34, 20, 27, -4, 38, 1, 38, -7, 3, -18, -37, -37, 42, 39, 4, -72, 11, -37, -8, 12, 11, -9, -42, 3, 32, -16, -48, 17, -8, 2, 30, -27, 12, 33, -14, 1, -32, 5, 6, -30, 0, 44, 13, 3, 33, -16, -38, -5, 21, -2, -7, -52, -6, -58, -22, -16, 38, 0, 11, 13, -33, -29, -11, 39, -84, 20, 36, 7, 44, 7, 13, 5, -3, 34, -86, -33, 37, 6, -1, -43, 34, 19, -63, -15, 15, -5, -29, 45, 31, -45, -46, 35,
    -- layer=2 filter=0 channel=7
    6, -13, -21, 23, -5, 14, -50, -7, 11, 13, 11, 17, 2, 6, -25, 0, -20, -7, 0, -4, 8, 10, 23, 16, 8, 24, -26, 36, 1, 20, -9, -29, 9, -20, 6, -36, 17, 22, -36, -13, 7, 0, 19, -28, -4, 29, -5, 15, -43, -10, 7, -34, -9, 12, 25, 19, -11, -25, -20, -9, 21, -24, -49, 20, -9, 5, -14, 2, -5, 0, 2, 6, 17, 0, -39, -17, 23, -3, -15, -15, -42, 20, -6, 0, -6, 0, 4, 1, 16, 23, 0, 36, 20, -11, -45, -8, 12, -32, -45, -30, -47, -6, -31, 7, 8, -57, 16, -42, 3, 2, 19, 24, -20, -20, 1, -29, 8, 18, 28, -7, -13, -24, 16, -16, 12, 28, 10, 19, -5, -1, 21, 17, 39, 29, -1, 5, 25, -8, -32, -27, -3, 3, -23, 2, -10, 23, -6, 5, 9, -4, 0, -25, 12, -5, -13, 24, -13, 21, -9, -37, 44, -33, -27, -8, -20, -2, -31, -4, -15, 15, -18, -42, -1, -13, -23, -13, 0, -10, -6, -7, 8, 8, 65, -12, -4, -14, 59, 13, -11, 14, -2, -28, -2, 1, 30, 1, 16, 7, -13, -5, 48, -28, -13, 19, -7, -28, 12, -2, -5, 35, 19, 7, -15, 14, -17, -20, 10, -26, -4, 28, 8, 81, -1, -23, -5, -31, -57, -22, 0, -2, -20, 5, -6, 13, 53, -31, -6, 3, -18, -10, 33, -61, -2, -66, -21, 10, 51, -6, -6, -39, 21, 18, 4, 7, -8, -14, 2, -11, 25, 13, -4, 14, -4, 7, 36, -8, 0, -8, -12, 5, -23, 1, 20, 39, 14, -1, -20, 1, 1, 18, -5, -55, 19, 37, 37, 28, -45, -4, -16, -52, -25, -37, -4, 16, -33, -2, 11, -13, 20, -28, 6, 25, -37, 12, 16, -7, 0, -65, -17, 29, 13, -2, -18, -3, -11, -15, 25, -7, -11, 11, -9, 0, 26, -36, -10, 16, -12, -3, 12, -3, 24, -63, 7, 3, -2, 2, -23, 13, 23, 0, 10, -43, 6, 37, 15, -18, 17, 36, 22, 2, -39, -13, -34, -31, 5, -42, 17, 9, -17, -3, 0, -3, 6, -33, -2, 20, -14, -24, 30, 13, 14, -24, -7, 25, 30, 6, 3, 7, -53, -54, 31, 20, 8, 18, 2, -12, -6, -85, -11, 11, -35, -5, -9, -15, -42, 1, -16, 18, -35, 0, -4, -29, 5, -10, 31, -14, 61, 21, -23, 42, -3, 37, 22, -23, 9, -12, -24, -26, 11, -47, 3, 12, -33, -11, 0, -33, -45, -42, 5, -4, -42, 4, -34, -43, -4, 35, 0, 1, 50, 4, -11, -19, 39, 14, 10, 20, 10, -22, -4, -21, 15, -27, 1, -11, -49, -4, -18, 0, 40, -29, 18, -17, 2, 7, 43, 30, 19, -14, 9, -28, 5, 25, 10, 3, -4, 17, 1, 21, 9, 4, -8, -4, 8, -5, -20, 2, 27, 11, 11, -2, 16, -27, -1, -7, -3, -10, 39, 70, -1, -15, 8, -19, 12, 20, -19, 12, -28, -7, -9, -16, -24, 33, 15, -8, 25, 9, 0, 1, -21, 4, -6, 16, 9, -43, 18, 26, 15, -2, -2, 27, -37, -12, 12, -12, 19, 17, -3, 41, 26, 43, 12, -4, -24, 12, -1, 14, -36, 11, -4, -27, 0, -5, 1, -3, -3, -11, 7, -6, 19, 0, -5, 21, 0, 35, 7, 13, 20, 9, 30, -2, -22, 18, 1, -9, 1, 7, -9, -16, 7, 52, -3, 25, -8, 3, -19, -9, -42, -17, -11, 25, 2, -2, -47, 6, 13, 31, -3, -29, 13, -33, -22, 60, 12, 13, 11, -58, -25, -5, 59, -20, -54, -4, -1, -21, 7, -8, -13, -22, -32, -11, -5, -6, -4, 12, -40, -3, 2, -28, -9, 23, 57, -9, 11, -2, 60, -20, 5, 15, -13, -44, -3, 6, 8, 47, -38, 4, -45, 7, -1, -13, 16, -12, -20, 11, -23, -6, 31, 35, -21, 31, -7, -8, -26, -58, 7, -27, -9, -18, 15, 4, -47, -14, 68, -7, 40, -3, 32, 7, -14, 11, -12, 22, 2, -23, 4, -2, -3, -38, 50, 36, 5, 14, -9, 4, -25, -12, 27, -9, 48, 13, 11, 8, -37, -19, 2, -3, -12, 19, -27, 3, -55, -5, -21, 1, 58, -1, -1, 29, -26, 7, -48, 4, -35, 33, -46, -11, -4, 3, -20, -32, 4, -18, 41, 0, 35, 0, 5, 17, -5, 2, 31, -30, -17, 12, -21, 17, -8, -12, -5, 9, -37, 2, 63, 79, -1, -3, -20, 49, -27, -30, 7, -15, -10, -26, 7, -13, -11, 24, 7, 4, -14, -22, -21, -15, -8, -5, 2, 1, 8, -35, 5, -18, -14, 2, -28, 22, -18, -7, -6, 3, 8, 45, -25, -5, 21, -4, 14, -25, -11, -5, 17, -19, 9, 4, -28, -13, -4, 6, -33, -48, 13, -23, -1, 22, -19, -17, -5, -11, -9, 9, 0, 12, 42, -5, 46, -3, 2, -6, -1, 16, 12, 14, -9, -2, 20, -9, 41, -15, 7, 9, 7, -10, -21, 4, -6, -12, 40, 9, -14, 36, -18, 23, -3, 44, -5, -1, 12, -2, -26, 68, -11, 11, -1, -9, 10, -12, 32, 11, 0, -4, 5, -9, -45, 22, 64, -33, -8, -22, 68, -55, -41, -95, -2, -36, -14, -18, 35, 5, 2, -15, 63, 36, 7, 37, -6, -19, 11, -5, 15, -36, 42, -6, -34, -2, 6, -18, 3, -23, 18, -34, 7, -2, 28, 32, 19, 10, 9, -21, 21, 13, 36, 30, -60, 85, -2, 12, -4, 17, -7, -21, 31, -17, 14, -58, -4, -2, -3, 41, 76, -36, -12, -1, 2, -30, 65, 79, -5, -63, -8, 11, 29, 26, -44, 4, -67, -7, -20, 2, -55, 72, -1, 0, -36, -12, -2, -25, -12, 0, -8, -4, 16, 5, 11, 25, -16, -2, 16, 35, -12, 18, -12, -5, 24, 29, -12, 1, 0, 53, -7, 11, -4, 13, -3, -15, 2, 4, 1, -52, 19, 3, -8, -7, 2, 19, 4, 0, -3, -5, 40, 24, -2, 16, 20, -2, 54, -3, -7, 22, -63, -4, -28, -3, 13, 18, -4, -1, -82, 21, -71, -87, -19, 5, -24, -6, -6, 38, -33, 13, 6, 6, 38, 73, -31, -1, -29, 8, -6, -33, -39, -26, 0, 13, 0, -62, -19, 0, -1, -11, 18, 61, -3, -19, -3, 9, -10, 5, -39, 38, 12, -8, -10, -9, 12, 6, -7, 30, 11, -12, -15, -30, 16, -13, 15, -21, 5, -14, -14, -42, -9, 0, -152, 25, -58, -62, -7, 1, 34, 46, 26, 12, -71, 78, -19, 6, 12, 38, 22, 24, -65, 13, -15, -42, -28, -35, -5, 43, 32, -3, -23, 0, 10, -45, 15, 47, 19, 2, -28, -6, 21, -14, -27, -19, -1, 0, 3, 26, 17, 15, 7, -26, 24, -8, -71, -4, 37, -53, 8, -2, 9, -2, -82, -50, 8, 2, -124, 25, -32, -48, -49, -10, 13, 26, 40, 7, -63, 74, -21, 5, -11, 30, -18, 23, -41, 20, -26, 4, -52, -44, -15, 25, 46, -27, -3, -28, -47, 13, -6, 42, -3, 6, -7, 5, 16, 3, -16, -21, -1, 25, -26, 23, 24, 22, -2, -68, 28, -23, -42, 25, 37, -46, -21, -30, -19, -30, 19, 27, 0, -7, -37, 26, -7, -1, -45, -4, -34, -20, 3, -7, -14, 11, 6, 2, 8, -7, -25, 25, 0, 49, 25, 6, -9, -7, -9, 13, 31, -3, 11, 1, -15, 4, 7, 25, 18, -22, 4, -2, 1, -15, 31, -19, 3, 37, -19, -2, -8, -6, -5, 17, 12, 22, 15, -19, 27, -9, 17, 13, 19, -4, -24, 9, 2, -8, 34, 32, 23, 7, -9, -6, 24, -6, -3, -2, -7, -55, 26, -9, -42, 57, -13, 3, 21, 18, 24, 0, 26, 50, -3, 70, 13, -14, 11, -17, 6, -78, -22, 5, -25, -4, 13, 3, -42, -26, 78, -39, -12, -24, 43, -25, -51, -84, 11, 7, -24, 1, 64, -22, -36, -17, 47, 3, -9, 28, 24, -32, 2, -1, 19, -11, -1, 13, -10, -4, -19, 1, 14, 2, 25, -15, 21, -8, -6, 8, 36, -54, 15, 13, 30, -1, 8, 35, -10, 45, -26, 21, -22, 28, -3, -12, -3, 0, 31, -18, 17, -2, -4, 24, 41, 8, -6, -11, 13, 13, 32, 4, 0, -25, 10, 44, 8, -26, -51, 27, -65, -2, -13, -5, 10, 55, -1, 5, -16, 33, 0, -5, -34, 1, -3, -14, 26, 12, 29, 22, 10, -4, -39, -4, -43, 20, -25, 9, 16, -8, -44, -14, -40, -13, -15, 36, -10, 16, 8, -19, -20, 14, -8, -60, 27, -1, -14, 11, -40, 23, -2, -9, -21, 5, 26, 53, -8, -65, 7, 47, 35, -6, -15, -16, -85, -22, -20, -45, -31, 55, -5, 0, -87, 48, -55, -81, -42, -7, -26, 54, -4, 47, -16, 52, -2, 7, -1, 10, -32, 7, -39, 24, -24, -53, -28, -42, -45, 18, -12, 14, -20, 13, 40, -16, 2, 18, 26, -9, -4, 2, -33, 0, -77, -18, -2, -2, -4, 23, 9, 13, 1, -31, 20, -9, -41, 0, 11, -16, -32, 31, -24, -29, -46, 19, -1, -9, -118, 17, -22, -76, 3, 7, 40, 103, -43, 20, -57, 59, -1, -14, 18, 35, 4, -32, -67, 36, -39, -29, -16, -6, -21, 0, 42, 27, -9, -24, 30, 6, 64, 2, 30, 0, -26, -6, -46, 29, -84, -21, -10, 21, -11, -1, -15, 18, 4, 5, 39, 6, -76, 2, 46, 37, 0, 35, 22, -29, 5, -33, -11, -9, -89, 0, -44, -29, -47, 2, -6, 47, -7, 33, -64, 3, -8, -7, -11, 8, -7, -14, -35, 23, -24, 0, -7, -18, -28, -20, 17, 41, 10, -21, -28, 34, -17, -11, 49, -61, -24, -8, -21, 23, -42, -33, -8, 47, -59, 17, 8, 25, 3, 4, -11, 59, -1, -35, 20, 16, -46, 1, 5, -37, 5, 6, -3, -5, -47, 35, -3, 15, -24, -2, -15, -9, -27, 54, -36, -21, 9, 4, 24, 40, -20, 24, 1, 9, -36, -39, -24, -47, 33, 27, 26, 29, 3, -21, 45, -27, -19, -6, 15, -9, 3, 8, -3, -15, 18, -19, -10, -13, -44, -3, -24, -35, -7, 2, 21, -11, -17, -16, -6, -16, 33, 10, 1, -7, 31, 15, 7, 4, 7, 40, 6, -1, -7, -6, 0, 11, -4, 2, 0, -35, 13, 0, 2, 60, 7, -5, 11, 20, -6, -30, -28, 45, 15, 28, 3, 14, -11, 1, -10, -64, -6, 1, 37, 0, 10, 0, -22, 25, 27, -5, -11, -43, 30, -11, -46, -101, -1, 2, -30, 2, 75, -14, -42, 10, 43, -8, 4, 11, 58, -20, 4, -10, 24, 3, 4, 4, -9, 8, -14, 46, 11, 12, 19, -11, 5, -13, 0, 21, 16, -41, 24, -10, 42, 72, 1, 72, -41, 33, 9, 2, 3, 45, -6, 17, -2, -11, 36, -16, 3, 10, -7, 5, -3, 30, 6, 32, -17, 19, 37, 41, 2, -41, 9, 31, 63, -2, -7, 54, -121, 9, -24, 3, -7, 54, -6, -7, 7, 30, 1, 26, -83, -10, 5, 9, 17, 22, 23, -20, -3, -3, 7, -26, 26, 17, 11, 11, -60, 9, -76, -65, -2, -71, -2, 38, 64, 21, -16, 36, 1, 4, 56, -29, 8, 0, 36, 1, -42, 18, -9, 55, -64, 4, 33, 54, -12, -47, -48, 50, 45, -14, -11, 28, -102, 2, -11, -80, 13, 37, 6, 4, 16, 26, -6, 6, -21, -2, 19, 51, 1, 55, 10, -18, -8, -10, -39, -1, -21, -21, 25, 17, 3, -23, -46, -84, -10, -2, -11, 50, 9, -1, -16, 44, 26, -19, 32, -54, 8, 3, -25, -1, 17, -3, 6, 18, -34, 11, -11, 14, 2, -59, -42, 42, -18, 23, -31, 16, -38, 11, -32, -17, 28, 19, -10, -3, 13, 43, 14, 1, 16, 3, 22, -10, -26, 44, 2, -32, -9, 8, -18, 36, -40, 5, 8, 22, 24, -12, -16, 18, -40, 40, -12, 25, 4, -26, 22, 5, 6, -39, -12, -84, -25, -7, -72, 20, 46, -42, 4, 28, -16, -15, 11, -31, -9, -26, -32, 54, -15, -32, 13, 19, -43, 33, -35, 18, 56, 63, -6, -19, -8, 29, 35, 20, -4, -3, 8, 4, -52, 55, -16, -7, -2, -5, 26, 22, -39, -24, -17, 46, -32, -17, -19, -1, -12, 33, -33, 19, 10, -4, 18, 23, 13, -49, 31, -48, -5, 5, -36, 18, -18, -10, -3, 6, -46, 3, -2, -58, -2, -40, -33, 42, 26, -2, 21, 10, -46, 14, -28, 1, 48, 21, 0, -2, 12, 53, 34, -8, -1, -3, 2, -5, -36, 21, -11, -14, 11, -3, -9, 30, -12, 14, 22, 17, -35, -47, -82, -21, 2, -4, 25, 24, 42, -17, 56, -20, 13, -15, 63, -23, 5, -3, -12, 0, -24, 6, 4, 0, -9, -28, -43, -62, 9, 36, -8, 3, 40, -1, 10, -2, 5, 23, -2, 2, 19, -51, 1, -16, -18, 8, 20, -9, -6, 4, -13, 10, -81, 25, -13, -9, 25, -10, -35, 44, 22, -12, 32, 42, -2, -11, -11, 51, 13, 31, 15, 51, 7, 7, 12, -40, 31, -13, 51, 15, 17, -11, -16, -11, -16, -18, 2, -22, 16, 7, -54, -145, 9, -45, -3, -38, 70, 9, -3, 25, 27, 29, 5, -7, 48, -30, -2, 4, -5, 7, 22, -33, -3, -6, 8, 59, -9, 25, -9, 29, 11, 3, 7, 5, 50, -36, -9, 4, 0, 76, 7, 107, -27, 36, 10, 32, -20, 39, -19, -2, -6, 28, 20, -4, 2, 2, -11, 22, 28, 40, -3, 46, -22, 48, 48, 7, -3, -65, 37, 64, 15, 12, 42, 55, -58, -4, 0, -16, 0, 28, -9, -9, -7, 16, 21, -22, -49, -3, 8, 0, -26, 21, -8, -43, 2, 4, 0, -30, -15, -56, 3, 15, -14, 24, -6, -18, -30, -17, 1, -6, 59, 14, -21, 9, -34, 1, -4, -42, 1, -7, 30, -7, -6, 28, 0, 13, -16, 21, 12, 5, -6, -73, -52, 28, -18, -17, -4, 0, -124, -4, 0, -59, -3, 17, 10, -19, 20, 33, 38, 15, -27, 9, 18, -1, -24, 31, 1, -47, -13, -5, -10, -37, 14, -61, 52, 30, -4, 31, -18, -10, 12, -21, -2, 26, 38, 18, -26, -4, 24, -8, 0, -16, 1, 0, 33, -4, -5, 21, -9, 28, -65, 18, 31, 12, -9, -31, -41, 10, 18, 18, -22, 8, -68, 23, 7, -17, 31, -18, -6, -5, 56, 26, 28, 36, -39, -7, -4, 8, -21, 5, 39, -25, 27, -14, -51, -27, -6, -9, 52, 4, 26, 2, -31, 73, 0, -12, 10, 14, 19, 21, 16, -41, 25, 1, 3, -10, 31, 4, -31, 30, 23, 28, -2, 35, -32, 64, -14, -54, -8, 6, -2, 62, -22, -7, -26, 3, -72, 21, 32, -24, 14, -10, 2, -10, 48, 17, 34, 23, -14, 1, -4, 5, -69, 13, 21, 19, 10, -7, -74, 0, -7, -40, 38, 12, 49, -10, -24, -16, 17, -16, -20, 27, 0, -11, 40, -79, 31, -19, 17, 0, 16, 5, 6, 31, 12, 12, 3, -35, -17, -12, -37, -59, 10, -66, 2, 40, -11, 2, -23, 20, -49, 8, -34, -34, -25, -57, -11, 3, 6, 41, 5, -3, -49, 8, 33, 10, -52, 81, -6, -9, 6, 0, -32, -9, 1, -1, 6, 34, 8, -17, -26, -17, -17, -30, -23, 11, 10, -28, 16, -51, -8, -11, 41, -28, 0, 7, 9, 36, -53, 10, 7, 15, -27, 16, 9, -100, 8, 13, -23, 37, -7, -6, -24, -20, -12, 43, -1, -53, -1, -43, 2, -6, -32, 11, 4, -52, -13, 0, 0, 23, -68, 39, -15, 20, 28, 0, -12, 39, 14, -21, -17, 39, 27, 20, 14, 51, -8, 12, 4, -10, 30, 29, -4, -36, 68, -3, 15, -22, -3, -10, 18, 8, -3, 19, 2, -1, 12, -1, -6, -91, -1, 1, 3, -16, -22, -1, -9, 27, -26, 32, -8, 2, 36, -7, 5, -3, -9, -3, 6, -36, -9, -6, -88, 54, -69, 24, -12, 28, 22, 0, -30, 11, -53, -62, -34, 18, 0, 17, -35, 65, -45, 9, -2, 48, -21, 27, -44, -1, -30, 39, 39, 14, 8, 0, -41, 44, 6, 13, -6, 57, -4, 53, 6, -40, 2, 10, 32, 34, 36, -46, 58, 49, -60, -5, -5, 7, 6, 26, 10, -11, -16, -21, 11, -16, -64, 1, -3, 18, -26, 24, -4, -20, -7, -12, -29, -25, -25, -40, -45, 24, -9, 62, -10, 19, -59, 9, 8, 49, -2, 12, -67, -4, -50, -2, 10, -31, -4, -5, 17, 45, -13, 8, 1, 3, -49, 50, 28, -29, -5, -34, -16, -12, 45, -39, 0, 21, -57, -33, -18, -34, -13, 49, 0, 5, 5, -1, 13, -2, -8, -2, 28, -15, -11, 33, 5, -26, -4, -7, 4, -27, -35, -35, -24, 26, -15, -28, -43, 29, -39, -29, 0, 17, -28, -15, -14, -13, 23, 0, 12, -52, -26, -7, 21, 26, -16, 16, 0, -22, -56, 2, 8, 21, -7, -16, -40, 9, -7, 0, -11, 1, -55, -35, -1, -31, -15, 37, -8, -4, 12, 56, 17, 1, -29, 4, -2, -22, -6, -23, 21, -48, 1, 9, -17, -51, -38, -7, -6, 26, 10, -34, -19, 0, -36, -39, -18, 7, 16, 25, 5, -37, 16, -13, 48, -63, -7, 0, -5, 20, -20, 4, -12, -4, -32, -4, 7, 10, 0, -24, -34, 31, 21, 3, -17, 3, -38, -8, 12, -23, -28, -12, 1, -6, 23, 17, 36, 8, -51, 7, -29, 4, -50, 26, 4, -28, 14, 4, 2, -20, -8, -34, 4, 10, 16, -8, -52, 51, -21, -31, 0, 48, 0, 9, 11, -72, 25, -16, 27, -24, -3, -3, -3, 31, -20, -5, -7, -34, 11, -9, -13, -29, -12, 24, -1, 44, 19, -11, 3, 22, -3, -19, 19, -22, -10, -43, -1, -2, 2, -7, -19, -4, -30, -3, -9, 17, -93, 13, -11, 11, 4, -13, 2, -38, -47, -41, 4, -4, -42, -30, -25, 45, -21, -21, -25, 13, -22, -11, 26, -17, 30, -9, 65, -12, 7, 2, -2, 25, -37, -8, 8, -29, 10, -10, 0, -113, -5, 36, 7, 49, 46, -15, -18, 22, -5, -14, 2, -18, -8, -23, -7, 7, 4, 16, 8, -40, -20, 0, 1, 34, -65, 33, -7, 11, 24, -13, -13, 27, 0, -25, -31, 31, 4, 26, 4, 66, -22, -6, -19, 23, 27, 42, 15, -37, -12, -6, 31, -34, 1, -2, -28, 22, -14, 0, 8, 3, 47, -1, 2, -86, 4, -42, 9, 8, -9, -56, -22, 35, 5, 10, -10, 0, 17, -20,
    -- layer=2 filter=0 channel=8
    1, -5, -28, -120, -52, 3, 52, 8, 14, 31, -57, 4, -21, 18, 29, -11, 22, 63, -8, -52, 2, -11, 21, 22, -18, 33, -2, 47, 28, 4, -13, -8, -58, -15, 4, -18, -17, 6, -39, -2, 1, -51, -3, -2, 8, 31, 5, 1, -91, 0, 4, -35, 4, -7, -41, 14, 3, 0, 13, 42, -1, 24, -16, -3, 1, -6, -19, -43, -32, -4, 29, 3, 17, 29, -30, 24, -15, 19, -7, 0, 8, 30, 2, -25, -6, 2, 40, -11, -28, 2, -1, 13, 16, -17, 8, -27, -31, 0, 38, 0, 32, 16, -23, -6, 11, -12, -50, 11, -5, 34, -14, 8, 4, -40, -13, -34, 22, 37, -42, 6, -8, -15, -15, 41, 11, 4, -29, -14, -9, 5, -23, -26, 14, 0, 0, -2, 12, 12, -48, 8, -22, 22, -14, -4, -41, 8, -7, -65, 5, 5, 12, -14, -15, -25, 9, 10, 0, -12, 23, -17, -25, -20, -50, -14, -11, 17, -40, -8, 5, -7, -44, 7, 0, 0, 2, -17, -44, -49, -10, -47, 3, -2, -19, 25, -21, -15, -38, 4, 15, -19, -9, -74, -6, -1, -18, -15, 3, -3, -15, 6, 3, -15, -59, -14, 2, 5, -10, 7, -77, -18, 0, -45, -17, 66, 2, -16, -12, -24, 3, 8, 3, 0, 8, 15, -48, -13, -6, -33, -7, 4, -15, 6, -9, 26, -34, -11, -10, 10, -26, -9, 11, -19, 4, 0, 0, -18, 0, 15, -30, 10, 2, -6, 15, -8, 12, -49, 3, 0, -3, -24, -2, 1, 27, 8, 0, 30, -12, 38, -34, 28, -21, -1, -20, 2, -11, -49, -24, 13, -6, 0, -6, -1, 0, 22, -4, 42, -16, 6, -53, 33, -41, -18, -1, 3, -28, 0, 9, 4, -56, 2, -3, 8, -31, -12, 13, -17, -1, -4, 20, 7, -9, 6, -13, 34, -36, -11, 1, -27, 22, -26, 5, -8, -17, -21, -20, -5, 31, 2, 12, 55, -36, 43, -7, 25, 21, -8, -12, 17, -2, -91, -21, 35, 16, 39, 0, -10, 19, 29, 4, 30, 8, 27, -42, 0, -41, 45, 0, 11, -6, -9, 2, 60, -50, 11, 0, 22, 0, 2, -14, 52, 0, -33, 24, 32, -54, 1, 8, 34, -57, 13, 8, 13, 10, 0, 1, 2, -22, -50, -10, -9, 32, -10, 11, 49, -1, 41, -18, 28, 38, -6, 18, 54, -23, -55, 0, -28, 20, 50, -4, -26, 4, 20, 16, 3, 3, -1, -26, -28, 15, 10, 10, 11, -12, 8, 4, -25, 0, 11, 7, 19, 18, 23, -35, 5, 7, 10, 14, 10, -86, 13, 11, 26, -42, 9, 4, 12, 2, 2, -3, -3, -6, -14, 0, 3, 5, -10, 6, 47, -51, 6, -5, 30, 4, -3, -11, 6, -8, -16, -7, 28, 41, 21, 22, -12, 13, -12, 2, -66, -33, -20, -9, 3, 16, 27, -47, 12, -6, 0, 11, -56, -33, 15, -12, 22, 49, -4, -35, 17, 2, -6, 3, 16, -23, 11, -29, -14, -17, 50, 5, 6, 3, -12, 4, -14, 38, -17, 8, 19, 0, -4, 8, 36, -54, 3, 0, 12, 19, -13, 9, -18, 1, -32, 1, 25, 18, 3, 0, -11, 9, 6, 9, -3, 19, 0, -11, -8, -59, 19, 13, 13, 5, -13, 9, 48, -13, 21, -4, 30, -5, 7, -15, 40, -1, -4, 23, 3, -7, 0, 8, 40, -30, 21, 7, -22, 18, -21, 0, -10, 9, -4, 5, 15, 9, -5, 39, 0, -52, 16, -9, -1, -10, -10, 0, 8, 6, -22, 10, 9, 22, -30, -19, -33, 36, 14, 9, 8, -27, -26, -11, 3, -18, -33, -37, 1, -24, 0, 15, 65, -21, 24, -13, -36, -22, -34, -8, 0, 1, -29, 0, 10, -15, 4, -25, 6, 3, -7, -16, -6, -2, -7, 9, 6, 0, -7, 0, -8, 9, -1, 20, -31, -67, 0, -8, -3, -41, -4, -33, -6, -1, -22, -21, 24, 3, -16, 1, 5, 1, 34, -4, 11, -21, 0, -1, -24, -50, -8, 14, -24, 19, -13, 7, -20, 19, 11, -1, -20, -18, -15, -52, 0, -2, -18, -15, 44, 28, 5, -26, -19, 22, -7, -5, 9, -26, 16, -9, -5, 2, 6, 39, 11, 19, -3, 26, -16, -70, 15, 19, -1, -9, -5, -24, 1, -6, -3, -5, 29, -5, -34, -16, -19, -2, 43, -15, 0, -34, -9, -4, 1, -5, -11, -37, 16, 15, 5, 13, 21, 26, 20, 2, -19, -2, -9, -23, -6, -4, -52, -13, 26, 2, -8, -31, -12, -4, 6, 0, -10, -37, -9, 4, 9, 9, -44, 8, -9, 19, 10, 28, -4, -34, 23, -4, 0, -9, -11, -9, 6, -8, -79, -15, 1, -9, 33, 17, -12, 17, 38, 9, 28, -1, 2, -63, 31, -25, 22, -18, -2, -8, 5, 17, 30, -21, 9, -1, 0, -18, 1, -33, -12, 0, 9, -6, 21, -6, -3, -11, -11, -8, -3, 2, 0, 17, 18, 7, 3, 11, -62, 3, 12, 38, -3, 14, 47, -28, 0, 2, 15, -18, -11, 13, 46, 14, -55, 5, -1, 28, 31, 4, 10, 13, 20, 0, 10, 21, -19, -33, 25, 3, -15, -19, 17, -43, -13, -2, -15, -14, 32, 7, 0, -27, 17, 18, 39, 11, 38, 25, 22, -5, -9, -33, 1, -15, 0, 11, -12, 44, 12, -11, -3, -7, -26, -7, -13, 18, -6, 9, 23, -53, 27, -25, 7, -27, 1, -8, 79, 25, -50, -3, -4, 27, 0, 6, -44, 34, 72, 0, -41, -48, -16, -13, 3, -27, 1, -21, 40, -7, -5, 3, -44, -38, 13, 11, 10, 10, 3, -39, 7, -2, 57, 10, -24, 7, 20, -42, -34, 5, -2, 2, 18, -16, 10, 1, -12, 16, -32, 6, 0, 8, 8, 28, 14, -90, 12, 1, -6, 20, -7, -20, 11, 13, -32, -7, 8, -9, 4, -19, -7, 27, 11, -14, -7, -59, 25, -40, 87, -17, 42, -46, 15, 15, -13, 12, 18, -6, 1, 10, -7, 8, -19, -57, -13, -4, 2, -2, -13, -2, -7, 13, -15, -10, -16, 22, -4, -34, -7, -11, -1, -32, 10, 11, -14, -5, -3, 20, 26, -33, -17, -19, -17, -6, -7, -4, -9, -1, -33, -1, 3, 18, 1, 2, -16, 24, 23, 0, 13, -28, 2, 1, 16, -23, -2, -19, 14, -11, 6, 10, 65, 43, -16, 3, -12, 20, -23, -26, 20, 10, 25, 0, 11, 14, -3, -17, -43, -6, -58, -13, -13, -53, 20, 6, 13, -15, -1, 44, -23, 13, -3, 34, -4, -65, 32, -9, -25, -21, 1, -25, -1, 5, -37, -12, 31, 14, -18, -7, 15, 19, 15, -7, -21, -21, -24, -28, -30, 13, -4, 7, 0, 1, -5, 9, 54, 50, -4, -2, -25, -13, -16, -17, -14, 10, 20, -11, 21, 76, -1, 5, -17, -31, -25, -26, -4, -36, -4, 9, 6, -10, 2, 18, 9, 13, -3, 19, 17, -17, 27, -21, -46, -26, 1, 6, 4, -11, 6, 2, 75, -11, 8, 5, -19, 30, 20, -26, 21, 31, 6, -12, -31, -34, 9, -34, -2, -28, -6, -12, 44, 37, 2, -7, -14, -3, 31, -10, 6, -6, -31, 3, 9, 24, -29, 7, -22, -10, 27, -7, 11, -49, -5, 2, -12, -14, -47, -7, 9, 6, 1, 8, 40, -57, -9, -38, -2, -22, -9, -14, 28, -8, -49, -7, 0, -11, 15, 9, 0, -7, 15, -17, 20, -32, -23, -25, -37, -27, 2, -104, 23, -8, 5, 20, 50, 13, 35, -8, 6, 0, 21, -14, -75, -5, -44, 18, 18, -9, -8, -23, -20, -32, -31, -4, 8, 0, -11, -1, -10, 6, -58, -13, 6, 5, 0, 16, 54, -12, 5, -24, 15, -15, 0, 24, 9, 6, -53, 6, 2, 27, 54, 19, 11, 18, 39, 10, -16, -27, 0, -22, 47, -9, -41, -38, 38, -33, 1, -2, 12, -35, 12, -5, 3, 6, -5, -48, -1, 8, -25, 12, -14, 7, -5, -72, 11, -75, -35, 7, -29, 12, -13, -5, 9, -28, -23, -18, -6, 4, 0, 16, -12, -6, 12, 0, 21, -23, 1, -43, 5, -1, -7, -11, 0, 31, 37, 1, -29, -8, 27, -2, 5, -25, -10, -25, 63, 13, -21, -32, -19, 0, -2, 1, 1, -18, 4, -5, 17, 20, 18, -19, -10, -10, 14, -9, 3, -17, 21, -30, -43, 16, 14, 10, 8, 6, 33, -8, 2, -9, -10, 28, -12, 13, -6, 4, 6, -27, 4, 11, -14, -11, 3, 37, 9, -17, 0, -8, 40, 1, 21, 0, -25, 2, 16, -4, 15, -21, 9, -12, 8, 71, 21, -4, 4, 0, 0, 34, 40, 19, 4, 1, -13, 24, -17, -21, -22, -8, 31, -38, -26, -7, -12, -19, -24, 33, 0, 7, 14, -20, 45, -1, -3, -46, 3, 24, -10, 17, -3, 10, -2, -43, 51, -46, -32, -29, -3, 8, -14, 3, -24, -6, 10, 11, -5, 2, -23, 41, -4, -15, -29, -1, 10, -19, -14, 14, 7, -28, -20, 15, -2, 6, 14, 62, 3, -9, -6, 27, 2, -19, -4, 3, -1, -13, 39, 70, 8, -16, -5, 3, -8, 12, 1, 9, 13, 7, 4, -63, -33, 10, -27, 18, -8, 6, -30, 0, 31, 0, -51, -28, 7, -54, -9, -9, -54, 16, 33, 1, 7, 27, 18, 13, 12, -20, 37, -40, -9, -54, -30, 37, 19, -47, -72, -16, -9, 26, 48, 44, 3, -5, -24, 22, 5, 4, -16, -1, -30, -60, 35, 0, -12, -1, -21, -43, -8, 5, 10, -62, 23, -1, -2, -22, 9, -1, -32, 8, 5, 1, -9, -34, 22, -21, -28, -14, -5, -18, 21, 2, -27, 16, 16, 3, -3, 10, 36, -8, -17, -16, -28, -16, 14, -28, -48, 0, 4, -48, -8, -12, 6, 5, 67, 58, 5, 7, -35, 14, 3, 2, -12, -6, -60, 0, 3, -32, 6, -6, 31, -34, -23, -9, 19, -63, 9, 1, 0, 28, -47, 7, -4, 27, 7, -17, -17, -25, -24, -37, 13, -27, 0, -39, 56, 24, -37, -5, 6, -25, 6, 18, 8, -16, 7, -14, 2, 1, 7, -10, 37, -30, 2, -64, -16, -5, 7, -3, 41, 14, 27, 8, -10, 7, 11, -2, -14, -9, -7, 21, 8, -20, -43, -14, 6, -25, -43, -2, 9, -27, -16, -3, -10, 7, -6, 11, 0, 4, 9, 3, 7, 8, -47, -37, 4, -41, 0, 31, 15, 32, 0, 19, -34, 6, -5, -14, 10, -4, 47, -1, -42, -7, -17, 22, 40, -26, -44, -19, 26, -36, 10, 11, 33, 22, 2, 4, 5, -23, 38, 66, 22, -1, 0, 11, -15, -4, 1, -62, 8, -38, -23, 7, -8, -19, -3, -2, -18, -97, -6, -13, 5, 31, 0, 15, -7, 31, 5, -10, -13, -36, 5, -48, -8, 0, 24, 10, -9, -8, 8, 24, -35, -6, 48, -31, 36, -18, -38, 4, -34, 46, -65, -53, -18, -15, -2, 11, -27, 14, -29, 8, -27, 36, 4, -23, -9, -9, 15, -1, -46, -14, 30, -43, -73, 53, -4, -24, 25, -35, 57, 5, -5, -1, 3, 7, 14, 13, -6, -6, -6, -11, -3, 11, -20, -41, -1, -75, 3, -19, 14, 2, 9, -7, 27, 29, 26, -19, 25, -18, -22, -36, 1, 6, -10, -8, -20, -46, -26, 27, -5, -28, 14, 33, 20, -6, -36, 46, 10, -49, -40, -4, 5, 11, 26, -17, -5, -23, 23, 0, 9, 3, -2, -8, 4, -4, -1, 6, 0, -38, -20, 17, 6, -8, -6, -7, -10, -19, 23, -5, -5, -106, -32, -30, 2, 1, 28, 15, 4, 26, 50, 25, 11, 7, -43, -28, -7, 8, 0, 34, -21, -34, -41, -5, -9, -16, 17, 19, 13, -13, -22, 39, 42, -45, -38, 8, 18, 2, -23, -6, 30, 14, 45, 7, -57, -11, 20, 35, 33, -1, 11, -37, -66, -72, -17, 9, 0, 29, -18, -57, -15, -78, -37, -10, -2, -47, -43, -2, -32, 12, 17, 29, 8, 41, 58, 52, -15, 18, 16, -56, -12, -31, 19, 32, -65, -39, 5, -14, -6, 0, 30, 35, 11, -8, -17, 26, 34, -45, -32, -9, -24, -38, -15, 30, 7, 19, 31, -6, -69, 10, 25, -13, 3, 5, 0, 11, -49, -30, 7, 12, 7, 18, -26, -12, -12, -33, -21, 12, -7, 9, -9, -19, -20, 27, -22, -26, 36, 53, 46, 49, -40, 17, -18, -11, -5, -13, -3, 17, -20, -38, -9, 16, -11, 25, 19, 40, 21, 0, -10, 22, 2, -23, -8, -9, -47, 20, 11, 32, 0, -2, 6, -3, -12, 1, 0, 2, 7, 2, 6, -19, -35, -52, 0, 6, -9, -7, 1, 55, 0, 6, -7, 33, 2, 20, 31, -3, 11, -11, 18, -2, 33, 30, 22, -9, -22, -16, -36, 6, 19, 21, 25, 11, 3, -1, -23, -13, 3, -25, -6, 48, 14, 1, -15, 40, -13, -3, -25, 2, -5, 35, 14, 22, -12, -1, 22, -16, -24, -35, 25, 1, 35, 5, 6, -51, -21, -38, 1, 2, -11, -22, -2, 17, 16, -33, -3, -43, 5, 18, 57, -3, 26, -24, -41, -10, 10, 2, -6, -18, 31, -13, -9, -1, -59, 48, 31, -33, -12, 19, -19, -45, -10, 6, 10, 8, 4, -4, 0, -3, -14, 25, 41, -3, 34, 32, 10, 41, -29, -67, -28, -25, -30, 0, 3, -22, 36, -5, -5, -78, 12, -10, 12, 6, 4, 5, -12, 37, 17, -38, -3, -43, -4, -52, 1, 11, 74, 2, -31, -3, -20, 2, 1, 9, 13, -9, -48, 5, -11, -3, -57, -19, -47, -83, -43, -50, 6, 3, -31, -16, 3, 6, -43, 46, 23, -71, 14, 5, 39, -26, -20, 9, 45, -29, -64, 42, -2, -11, -1, -31, 3, 2, -6, -15, 32, -52, 7, 22, -2, -21, -8, 32, -10, 19, 17, 3, -4, -56, -20, -34, 64, -4, 0, -11, -14, 35, 26, 0, -18, -23, -39, -14, 20, 53, -27, -10, -21, 0, -2, -19, 7, -5, -33, 0, 43, -6, -28, 29, 0, -44, -44, 0, 38, 17, 0, -5, -7, 5, 26, 35, -18, -7, 34, -14, 1, -5, 11, 5, -32, -70, 15, 39, 0, -17, 1, 54, -69, 3, 5, 14, 5, -101, -29, -42, -7, 5, -1, 20, 11, 24, 48, 12, -17, -3, -87, -34, 9, 38, 38, 70, -28, -47, 31, 0, 6, -20, -27, 9, 22, -5, 20, 25, 15, -57, -6, -3, 18, -4, -48, -38, 6, 11, 54, 4, -40, -4, 32, 66, 13, 7, -3, 34, -125, -106, 33, 4, -10, -13, -8, 7, -86, -47, 0, 18, 3, -89, -16, -26, -45, 32, -79, 25, 27, 24, 64, 38, -13, 44, -110, -34, 12, 1, 71, -12, -61, -95, 9, -19, -2, -13, -72, 5, -31, -5, 4, 43, 20, -44, 15, -13, 31, -28, -36, 33, 38, 46, 55, 0, -43, -19, 26, 22, 25, -3, 0, -21, -76, -56, 0, 1, 2, -37, -26, 18, -46, -47, -6, 5, 4, -61, -28, -9, 4, 10, -59, -16, 48, 40, 56, 6, 0, 4, -88, 45, 21, -40, 71, 14, -33, -22, -4, -3, 2, 6, -28, 21, -12, -9, 14, 45, 52, -39, 19, -3, -15, 6, -3, 31, -6, 20, 10, -19, -79, -18, 31, 22, 41, 12, -11, -1, -22, -72, -16, -2, -5, -34, 4, 44, -5, -22, -14, -13, 4, 14, -8, -11, 18, 5, -51, 35, 35, 32, 81, 34, -10, -25, -75, 54, 26, 20, 59, 4, -6, 0, 2, 8, 7, -25, 1, 26, 20, -5, 0, 38, 33, 13, -49, 2, 7, -5, -2, 0, 12, 13, -9, -53, -58, -20, 25, 24, 25, -9, 12, -71, 20, -38, 20, -13, -9, -23, -8, 66, 25, -53, -26, -32, 0, 9, 33, 11, 27, 19, -60, -4, 26, -9, 33, 56, -15, -5, 17, 0, -50, 74, 50, 37, -6, -1, -40, -51, 9, 12, 32, 6, -11, 6, 22, -26, -3, 75, 36, -7, -24, 10, 24, 75, 6, -2, -61, -35, -4, 4, -18, 16, 6, -5, 1, -135, 34, -7, 39, 23, -6, 20, -54, 53, 30, -46, -29, -46, 7, 0, -24, 45, 103, 63, -15, 67, -20, -17, -67, 5, -6, -47, -51, 56, -71, -2, 21, -68, -63, 10, -5, -48, -1, 27, 0, -14, -32, -4, 0, 49, 38, -50, 1, -6, -54, -69, -48, -27, 53, -132, -132, -8, -37, 2, -31, -65, -15, -4, -5, -33, -5, -19, 37, 15, -10, -30, -29, 27, -18, 8, -29, -14, 3, -85, 3, -10, 75, 28, 11, 30, -23, 13, 22, -6, -13, -31, -88, 21, -13, 21, 24, -4, -18, 50, -27, -13, 11, -18, -49, -29, -14, 12, 5, 37, 37, -39, -11, 2, 64, -30, -1, -68, 1, 0, 11, -2, -1, -16, 32, -6, -6, -4, 9, -11, -6, -35, 33, 14, 7, -20, -27, 38, -56, 15, 8, 33, 1, -122, -5, -32, 72, 7, -15, 36, 8, 54, 4, 15, 8, -24, -136, 8, -4, 16, 41, -24, 1, 4, -6, 5, -1, -24, -76, -3, -3, 11, -18, 71, 30, -18, -35, 6, 34, -12, -55, -52, -6, 6, 5, -26, -2, -8, 45, 22, 13, 11, 2, 38, -35, -59, 39, 35, 0, -1, -9, 77, -48, 20, -12, 7, -6, -69, -17, -14, 8, 13, -37, 25, 20, 61, 31, 40, 0, -14, -171, 50, 0, 39, 39, -45, -12, -67, -6, 1, -7, -7, -41, 16, 0, 0, 11, 28, 40, -32, -18, -1, -17, -7, -49, -23, -16, -10, 22, 21, -20, -25, 51, 27, -5, 4, 8, 10, -43, -36, 18, 30, 6, -22, -43, 65, -46, 0, 31, -40, 1, -10, -37, -20, 2, 0, -95, 28, 3, 22, 39, 40, -13, -3, -113, 23, 5, 27, 49, 19, 7, -3, 0, 2, 11, -7, -58, 2, 10, 7, 9, 33, -14, -29, -6, 4, -4, 3, -23, -49, 3, 0, 17, -10, -14, -22, 28, 42, 6, 6, 4, -20, 11, -54, 25, 24, 0, -10, -7, 89, -66, -20, -19, -17, -1, -57, -24, 0, -4, 21, -41, 17, 31, 47, 41, 50, -4, -14, -79, 13, -15, 84, 29, -2, 37, 26, 4, -19, 9, -18, -7, -11, 11, -4, 22, 44, 13, 26, -21, 8, -22, 9, 0, -56, 1, -6, -14, -3, -36, -8, 29, 55, 28, 9, 4, -156, 35, -21, 41, -16, 6, 0, -6, 80, -24, -89, -13, -112, -2, -3, 0, 75, 41, 75, -22, 26, 10, -32, 0, 74, 14, 1, -30, -64, -120, 64, 37, -44, -29, 64, -25, -69, -3, 23, -5, -40, -30, -1, 40, -34, 20, 47, -12, 8, -33, -13, -35, 13, 11, -59, -104, -14, -54, 24, -45, -6, -43,
    -- layer=2 filter=0 channel=9
    -11, -15, -16, 22, -20, 15, -50, -7, 36, 30, 14, -45, 17, 20, -6, -8, -90, 22, -5, 4, -11, 9, 20, 4, 7, 33, -3, -35, 63, -46, 0, 2, 23, -22, -2, -5, -33, 27, -10, 3, 34, 31, -55, -21, 3, 38, -9, 29, 2, 0, 7, -40, 4, 21, 27, 2, -35, -43, -39, -66, 41, 17, -30, -57, 1, -14, 17, 5, 5, 9, -64, -6, 10, 16, 77, -4, 41, 27, -19, 4, -23, -19, 1, 24, -11, -10, -7, -3, -6, 35, 20, -31, 25, -2, 27, 0, 15, -28, -17, 6, 12, 4, -12, 6, 25, 8, -11, -6, 0, 0, -27, 13, 1, 33, -7, 20, 15, 17, -11, 0, -42, 21, -23, -54, 24, -20, 0, 12, -8, -4, 7, 7, -26, -29, -21, 1, 25, -7, 43, -39, 2, 6, -22, 0, -1, 20, 4, 6, -22, 11, 14, 9, 6, 10, -12, 0, 5, 6, -20, 4, 15, 11, -13, 4, 35, -16, -12, 0, -4, -22, 38, -17, 6, -7, 28, 25, -30, -4, 0, -9, 5, -9, 0, 34, 0, 37, 32, -30, -1, 14, -30, 34, -2, -4, 9, -9, 25, -17, 14, 9, 11, -30, 41, -53, 15, 14, 7, 0, -50, -12, 19, 8, -21, -31, 2, 32, 22, 21, -36, 7, 8, 3, 9, -6, -15, 23, 22, 2, -19, -34, -14, -3, -20, -19, 51, -28, 5, 24, 39, 56, -7, -5, -12, 24, 13, -5, -40, 13, 27, 20, 37, 5, 17, 28, -11, 51, 5, -24, 8, -1, 40, -22, 14, -11, -14, -20, 34, -4, 25, 14, -13, 7, -29, -28, 11, 17, -7, -13, -4, 9, 2, 40, -5, -24, -8, -32, -10, -1, 6, -21, 18, 6, 5, -23, -18, -3, -11, 0, 20, -41, 7, 4, 18, 39, -11, -9, -13, -6, -11, -5, -23, 30, -15, 15, -4, -14, -3, 36, -37, 2, 8, -10, 4, 16, 30, -2, -41, -6, -3, -31, 30, 2, 37, 35, 8, -9, -63, 0, 15, 87, 6, -14, 19, -23, -20, 11, 0, -12, 2, -37, 6, -23, 44, -89, -16, -3, 26, -19, -35, -3, 2, -10, -10, -23, -4, 20, -7, 39, -27, -45, 3, -12, 8, 21, -20, 8, -64, -8, 19, -5, 33, -17, -26, 3, -1, -4, -1, -9, 0, 19, -8, -1, 29, -10, 15, 23, 26, 50, -16, 8, -56, -18, 0, 44, 0, 8, 4, -32, 15, 5, 8, -8, 29, -17, -12, -44, 29, -58, 28, -25, 42, 20, -20, -7, 24, 29, -61, -12, -2, 39, -2, 32, -24, -18, -3, -11, 20, 32, -37, 37, -61, 1, 28, 15, 23, -13, -19, -32, -1, -2, 19, 25, 6, 7, -25, -10, 19, -23, -5, -15, -10, 12, -5, 1, 4, -6, -19, 26, -13, -1, -13, 2, 5, -10, -31, -3, 11, -8, -9, 23, -15, 2, -55, -16, 3, 9, -19, -10, -19, -2, 6, 17, -5, -24, 6, -3, -8, -48, -4, 22, -13, 26, 26, 0, -41, -17, -14, 3, 12, 26, -20, -7, 0, -7, 28, 13, 32, 4, -7, -1, 15, -6, -6, 34, 10, -1, -48, 0, -6, 6, 19, 7, 13, 2, -10, -3, 6, -6, -24, 6, 14, 13, 16, 32, -15, 15, 2, -10, 7, 23, 5, 0, 16, -16, -29, 9, 8, 11, 27, 1, -6, -34, 0, 17, 19, 14, 9, 12, 0, 42, -48, -54, -6, -2, 0, 12, 3, -18, 19, -21, 26, -21, -6, -3, 2, -29, -2, -9, -36, 6, -43, -4, 2, -4, 26, -6, -5, 12, -12, 12, 26, 22, -12, 2, -1, 21, 6, 11, -28, -15, -7, 2, 9, -7, -12, 1, 0, -7, 32, 16, -1, -7, 38, -28, 3, -23, 0, -7, 3, 34, 35, -3, -1, 1, -34, -4, -1, -3, 22, 2, -3, -7, 0, 17, 28, -17, 9, -11, -4, -13, -4, 23, -26, 5, -31, -6, -25, -8, 7, 0, 15, -20, -23, 34, 3, 16, -42, -23, 19, 20, -12, -11, -7, -21, -1, -13, 8, 6, -15, 2, -5, -5, 36, 1, 7, 40, 39, -39, -4, -57, 3, -37, 3, 0, 29, 6, 3, 25, -30, -4, -8, 22, 0, 22, -1, -8, -11, -26, -9, 2, 19, -7, 6, -31, 17, 38, -40, -8, 0, 0, 2, 4, 16, 17, 30, -7, -2, 29, 15, 28, -16, 15, 14, 21, -27, -3, 13, -60, 29, -28, -6, -12, -21, 1, 5, -23, 70, 1, 1, -4, 44, 14, -2, -83, 0, -28, -6, 7, -31, 6, -20, 24, -8, 11, -8, 9, -23, 20, 7, -15, -2, -1, 18, -11, 6, 0, -3, -15, 7, -20, 4, 15, -16, -12, 13, -10, 15, 14, 2, 14, -1, 0, -10, 42, 6, -3, 5, 21, -24, 9, 37, -26, 4, -32, 4, -7, -6, -13, -2, -7, 19, -5, 0, -19, 11, 0, 8, -74, -7, -33, 4, 4, -11, 16, -37, 42, 16, 0, 0, -8, 1, -17, 4, -8, 7, -13, 11, 13, -32, -7, 1, 0, 0, 7, 21, -10, 18, 1, 19, 20, -4, 9, 0, -11, -7, 22, 9, -2, 18, -4, 14, -10, -22, 21, 1, -21, 13, 6, 6, -8, -12, 3, 20, 3, -2, 6, -3, 25, -1, 25, -9, -41, -13, 22, -5, 0, -33, 35, 6, 47, -22, 22, 35, -5, -6, 5, -3, -2, 19, 1, 37, -28, -2, -1, -8, -22, 7, 18, -22, -1, -6, -7, -36, -14, -17, 40, -29, 6, -10, -13, 8, -8, -80, 3, 3, -10, 35, -24, -12, 2, -8, -6, 24, -46, -8, 7, -19, 3, 20, -2, 6, -3, 1, -10, -13, -11, 3, 31, 20, 26, 38, -37, -17, -22, -13, -20, -13, 0, -19, 15, 0, -8, -2, 1, 23, 19, 24, 9, 0, 15, 4, 7, -45, -21, -30, -14, 18, 27, 3, 4, 2, 0, 25, -2, 23, -14, -38, 12, 8, 33, 6, -18, -8, 6, -45, -22, 30, 16, -16, 10, 23, 11, 6, -19, 7, 7, 17, 29, 3, -29, -6, -64, 2, 9, -37, -13, -16, 10, -52, -41, -27, 4, 0, -7, -11, -7, -11, 5, 13, 49, 17, 7, 8, 3, -8, 24, -41, 26, -20, 0, 0, -13, 18, -17, 24, 52, -1, -4, 13, -18, -21, 11, -5, 55, -7, -1, 0, 4, 12, -34, 7, 0, -37, -1, 6, -12, -11, 13, -6, -29, 16, 27, -13, -48, 9, -69, 4, -1, -44, -6, -6, 9, -35, -21, -10, -4, 14, 22, 2, -18, 21, 13, 40, 20, -1, 4, -8, 29, -21, 40, -22, -1, -26, -8, -35, -56, 2, -6, 24, 30, 0, -2, 28, 3, 11, -8, -12, 74, 0, -7, 5, -34, 30, -4, 48, -20, -21, -5, 28, 32, -12, 12, -12, 22, 22, 45, 14, -49, 1, -15, 8, 36, -20, -4, 21, 7, -24, -6, -17, -17, -30, -15, -1, -9, 15, 1, 37, 26, 17, 2, 0, 8, -20, 30, -34, -26, -27, -1, 1, 5, 39, -12, 17, 41, -19, 22, 24, 17, 30, 1, 25, 41, -21, -13, 10, -32, 59, -26, 21, 1, -31, -4, 23, 56, -7, 24, 10, 2, 22, 19, 6, -66, 3, 0, -19, 22, -30, -5, -10, 8, -15, -33, -7, -20, -2, -28, -6, -1, -17, 32, 11, 13, 3, -5, 14, 15, 12, 9, -56, -22, -22, 2, -26, 5, 14, -22, 13, 15, -2, 23, 26, 6, 52, 2, -11, 19, -40, 0, -5, 0, -6, -39, 6, -9, -41, 5, 21, -36, 4, -23, 2, -39, 32, -19, -1, -119, -3, -26, -5, 4, 63, 21, -9, 23, 2, -52, -13, 11, 31, -47, 3, -18, 9, 14, -4, 11, -17, 5, -27, -23, -9, 5, 2, -14, -32, 7, 21, 35, -15, -19, 16, 0, 27, 18, 19, 12, 0, 9, 11, 13, -32, -24, 7, -4, 35, 6, -12, -19, -9, 5, 8, 41, -16, -19, -11, -25, 1, 2, 8, -27, 1, 43, -3, 35, 54, 0, 9, -7, 0, -2, -32, -2, -83, -30, -9, -13, -20, -32, 17, -40, 0, 1, -20, -50, -10, 68, -39, -9, 0, 6, -3, -23, 34, 49, 0, -24, -10, -13, 15, -28, -103, 17, -1, 9, 26, -11, -12, -20, 11, -6, 8, -69, -23, -10, -65, -1, 12, -15, -3, -3, 20, -34, -5, -43, -8, -21, -6, -13, 38, -39, -4, -53, -23, -6, -6, 7, -1, 9, 6, -10, 3, -10, 0, 45, 34, -1, 27, -21, 6, 22, -50, -18, -46, -12, -42, 30, 57, -32, 71, 3, 9, -12, 12, -33, 23, 26, 0, 88, -28, -7, -49, -76, -32, -42, 2, 54, -45, 2, 16, -3, 8, -12, 7, -34, 8, 31, 0, -74, 10, -78, 45, -33, -44, 46, 23, 52, -72, -63, -2, -5, 11, 0, 9, -14, 52, 0, 21, 40, 34, 0, 13, -17, -2, 19, -41, -21, -34, 7, -14, -38, 33, 11, 11, 14, -16, 11, 15, -6, 55, -34, -7, 48, -13, 12, -47, 11, -8, -19, 7, 42, -42, -9, 55, 6, 3, 5, 6, -23, 2, 6, 14, -59, -4, -77, -29, 13, -19, 13, 64, 25, -54, -48, 8, -12, -7, -17, -2, -11, 23, 30, 53, 69, 8, 4, 16, -1, -29, 54, -33, -2, 6, 0, -34, -6, -7, 0, 4, 42, -22, 6, 15, 36, 95, -36, 3, 53, 0, 22, -16, -46, -8, -13, 17, 43, 8, 3, 19, 57, -26, 39, 5, -7, 0, -6, 10, -55, 5, -57, -23, 37, 56, 12, 46, 4, -51, 3, 20, -12, -19, -38, -7, -2, 55, 53, 49, 43, 28, 3, -6, -4, -19, 24, 9, 23, -22, 8, -64, -5, 0, -15, 26, 56, -57, -1, -7, 34, 107, -14, -6, 50, -26, 13, 16, -9, -11, -13, 6, 47, -13, -12, 28, 31, -14, 9, 7, -26, 1, -14, 8, -81, 1, -14, 10, 33, -20, -5, 47, 8, -17, -34, 11, 1, 44, -58, 4, -18, -13, 11, 21, 17, 21, -8, 11, 7, -19, 12, -56, 4, -26, -10, -65, -2, 1, -36, 29, 29, -12, 0, 13, 82, 35, -5, 13, 47, -42, -2, -16, -58, 8, -10, 3, 37, -34, -11, 0, 15, 16, 12, -10, -20, 34, -4, 10, -96, -6, -53, -20, 10, -8, 1, 9, -9, -25, -24, 14, -2, 18, 10, -3, 3, -26, -12, 14, -31, -16, 3, 1, -21, -10, -8, -33, -12, 6, -2, 18, 1, -34, -32, -21, 10, 12, 29, 15, 28, -44, 9, -15, 13, -10, -12, 16, 6, 34, -14, -20, -32, -18, 7, -4, 26, 0, -25, -11, -5, 21, 6, 18, -27, -3, -17, -9, 15, 45, -12, 5, -44, -14, 3, -62, 17, -74, 1, 2, -4, -25, -5, -16, -61, 6, 8, -49, -45, 13, 34, -5, -43, 6, -11, 10, 8, -24, 20, -55, -27, 15, -2, 20, 14, -123, 22, -46, -7, 23, -13, 40, -15, -3, 7, -8, -38, -25, 1, -78, 2, -7, -19, 1, -19, 22, -46, 10, -37, -6, 9, -34, -24, -38, -22, -13, -59, 3, 0, -21, 12, -39, 33, 7, 2, 26, -10, 16, 0, 40, 0, -4, -24, 17, 20, -34, 35, -14, -2, -1, 32, 29, 8, -9, -17, -36, 10, 29, -22, -10, 25, -4, 71, -52, -15, -29, -35, 0, -34, 0, 20, -40, 10, 19, -16, -4, -6, 0, -16, 20, -6, 31, -44, -8, -13, -16, -2, -119, 12, 0, -1, -29, -13, 14, 8, 19, 15, -4, -10, 38, -33, 42, 25, 29, 5, -7, -76, -7, -26, -8, -10, -23, 0, -6, -21, 37, -19, -21, 7, -20, 13, 14, -9, -51, 0, -16, 45, -6, 13, -62, 42, -1, -20, 29, 90, -27, -4, -4, 4, 7, 13, -10, -20, 2, -40, 36, -14, -6, -59, -7, -13, -66, -18, 39, -16, -45, -33, 42, 23, 28, 7, 0, -4, 27, -18, 10, 45, 12, -9, -22, -42, 20, 12, 6, 0, 1, -5, -15, -54, 12, -36, 47, 3, 16, 0, 4, 8, 22, -47, -28, 48, -34, 17, -26, -34, -13, -3, -3, 48, -9, 0, 8, 1, -33, -11, -6, 3, -9, -34, 12, -43, -1, -70, -18, 41, -77, 10, 40, -21, 17, -1, 49, 12, 39, -38, -3, -15, 13, -13, 13, 34, 28, -2, -9, -46, -21, -12, -11, -7, -21, -2, -37, 4, 36, -40, 33, 28, -16, -23, 3, 11, 38, 0, -29, 54, -81, -2, 4, -50, 18, -10, -26, 44, -26, -10, -13, 25, -13, -12, 4, -2, 17, -17, 7, -39, 2, -28, 0, 33, -85, -29, 33, -24, -25, 10, 58, 19, -39, -80, 5, -8, 25, -7, 41, -8, 31, -6, 4, -75, -10, 7, -9, -12, -22, -1, -20, 13, 26, -41, 23, 22, -27, 25, 25, -7, -22, 38, -18, 65, -56, 4, -5, -6, 34, 4, -35, 45, -45, -6, -19, 21, -17, -7, -8, 0, 32, 2, 21, -30, 2, 26, -21, -14, -78, 13, -5, -33, -17, 9, 40, 28, -73, -11, -7, -11, 4, 0, 36, -47, 19, -10, -63, -53, 20, -10, -55, 39, -9, 1, -78, -17, -57, -29, -15, 0, -27, 48, 41, -23, -39, 0, -61, 27, 30, 22, -39, -10, -31, 16, -9, -61, -23, -6, -18, 4, 57, -23, -8, -22, 35, -4, 4, -20, -7, -43, -21, -7, -28, -5, -6, -39, -36, 13, -30, 26, -15, 40, 4, -3, 0, -23, 3, -37, 17, 1, -35, -41, -7, -12, 34, -35, -29, -5, -6, 13, -23, -19, -75, -13, -13, -9, -18, -18, -101, 43, -72, -3, -17, -14, 26, -100, -29, 7, -11, -6, 9, -6, -72, 2, -3, 8, 4, -43, -10, -74, 11, -28, 4, -49, -15, -9, -5, -85, -42, -6, 10, 12, -48, 7, 40, -12, -11, -2, -37, -33, 14, -58, 35, 8, -5, -41, 24, -20, -1, -12, -36, -4, 21, 34, 5, -17, -32, -46, 12, 24, 9, -13, -70, 12, -32, 39, -28, -33, 4, 0, -7, -10, 13, -17, -9, -6, -26, -16, 5, -7, -7, -12, 54, -73, 46, -69, -5, -45, -29, -34, -14, -29, -40, -49, 8, 37, -20, 27, 25, -7, 2, -14, -37, -40, 0, -20, 7, -10, -4, -59, 6, -16, -24, -14, -17, 3, 8, 24, 21, -35, 0, -11, 0, 16, 9, -29, -26, 5, 22, 16, 18, -8, -33, -27, -38, 2, -17, 23, -38, 0, -19, -46, 15, -3, -9, 18, 25, -104, 24, -17, -7, 21, 16, -18, -96, -2, -20, -41, -12, 7, -23, 22, 41, 9, -5, -4, -22, 7, 2, -3, 23, -10, -31, -29, 7, 22, -18, 4, -10, 3, 8, 14, 8, -5, -14, 24, 25, -12, 15, -1, -10, -11, 8, 30, 11, 0, 3, -36, 15, 15, 27, 38, 3, 5, -8, -51, -18, -22, -2, -9, 13, -42, 0, 0, -12, -51, -1, -11, -125, -43, -25, -45, -12, 7, -25, 39, 60, -13, 12, -7, -19, -78, -7, 2, 34, 9, -10, -20, 13, 7, 31, 14, -21, 5, 22, 19, 17, -17, -14, 1, -13, -20, 2, 4, -40, 5, -12, 35, -26, 2, -26, -6, 9, 2, 30, 67, -19, -9, -4, -66, -4, 1, -5, -41, 5, -42, 6, -53, -12, -11, 10, -8, -93, 28, -10, -32, -2, 16, 17, 29, 84, 1, -10, 0, -22, -41, 10, -43, 59, 7, 4, -65, 5, 3, -4, -21, -16, -8, 14, 20, 60, -38, -6, -1, -36, 10, 52, -12, -37, 23, -11, 20, -13, -18, -33, -7, 3, -23, -8, 16, -22, 7, 3, -59, -35, 9, 10, -27, 55, -25, 16, -27, -2, 15, 24, -14, 38, -5, -30, -22, -23, 5, 19, 36, 57, -10, -7, -7, -26, -24, 29, -43, 35, -6, -52, -52, 26, -1, 10, -29, 10, 9, -17, 8, -3, -40, -67, 6, -54, 42, 46, -50, -67, 16, -58, 20, 28, -12, -59, -25, 9, 20, -5, -42, -2, -4, -19, -17, -18, -1, -6, 16, 31, -43, 2, -2, -4, -10, -7, 5, -17, -54, -33, -17, -6, 16, -32, 50, 11, 21, 0, 2, -10, -33, -35, -1, 37, -1, -22, 63, 10, -73, 59, 6, -41, -5, -10, 13, 0, -76, -61, -32, -25, -10, -47, -4, 19, 14, -7, -7, -22, 19, 44, -82, -32, -1, 9, -17, 30, 5, -19, -35, 20, 6, 6, -24, -31, -71, -2, -18, -1, -59, 17, -16, 1, -44, -36, 47, 19, 41, -27, -9, 107, -64, 7, 0, -4, -6, 12, -51, 62, -5, 1, 39, 0, -5, 26, 2, -18, 1, 29, 44, 25, -63, -24, -26, 5, -1, 37, -34, -8, 27, -24, 68, -13, -28, -4, -58, -20, -21, -45, 4, -22, -2, -19, -43, -21, -10, 4, -35, 55, -57, 19, 15, -11, -53, -2, -18, -63, -12, -58, -31, 27, 15, -20, 30, 72, -23, 0, -4, -37, -32, 32, -37, 50, 7, 2, 6, -57, 1, -31, 45, -27, -9, 9, 1, 35, -41, -59, -34, -4, -7, 22, -7, 11, 39, -16, 41, -6, -58, -42, -7, 68, -53, -5, -2, -48, -4, 5, -38, -19, 14, 2, 10, 29, -31, 20, -1, -12, -34, 21, 6, -18, -25, -40, -41, 13, 12, 11, 35, 56, -2, -3, 2, -36, -28, 11, 2, 33, 5, 2, 56, 12, 23, 0, 45, -33, -12, 3, 8, 23, -29, -11, -8, -39, -26, -18, 7, 45, 25, -2, 16, 8, -27, -29, -36, 13, -44, -17, 14, -42, 6, 12, -47, -15, 4, 3, -52, 26, -17, 4, 19, -4, -42, 26, 2, -43, -4, -34, -38, 28, 15, 20, 30, 91, 9, -6, -2, -32, -8, 1, -8, 68, -15, -13, 53, 27, -35, 15, 65, -27, 5, 19, 6, 23, -22, -28, 10, -26, -14, 23, 5, 71, 21, -2, 44, 1, -12, -11, -5, 6, -22, -8, 54, -37, 8, -4, -56, 8, -13, 4, -38, 48, -36, 23, 22, 6, -38, 45, -6, 0, -14, -42, -35, 8, 0, 19, 28, 80, -8, -4, -22, -53, -72, 14, -32, 61, 3, -5, 54, -27, 33, -20, -1, -18, 7, 32, 16, 27, -32, -58, -17, 1, 0, 26, -18, 28, 27, -3, 61, 21, -10, -61, 1, -50, -32, 13, 21, -47, 3, -21, -41, -14, 1, -5, -7, 39, -20, 6, 2, -8, -43, -16, -26, 2, -16, -46, -14, -10, 16, 9, 37, 64, 22, -3, -20, 3, -75, 18, -32, 41, 7, -19, 35, -14, 18, -6, -7, -2, -12, -22, 20, -37, 17, -84, -38, -5, -15, -1, -45, 12, 20, -37, 9, 60, -3, -91, -31, -16, 2, 3, -5, -17, 5, -23, -29, 34, 0, 0, -26, -1, -20, -5, 5, 0, -21, 0, 19, 8, -18, -38, -13, -67, -5, -24, 12, 68, 27,

    others => 0);
end iwght_package;
