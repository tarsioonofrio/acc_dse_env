library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 325, 0, 623, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 182, 0, 914, 0, 0, 0, 0, 207, 0, 0, 0, 0, 0, 0, 0, 0, 294, 0, 0, 110, 0, 161, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110, 0, 0, 0, 0, 647, 0, 0, 673, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 111, 41, 0, 0, 246, 38, 0, 0, 0, 0, 118, 81, 0, 0, 0, 362, 0, 0, 0, 0, 0, 125, 0, 0, 0, 446, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 371, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 71, 806, 0, 0, 0, 15, 0, 0, 321, 0, 0, 1077, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1483, 376, 0, 0, 0, 0, 0, 0, 0, 358, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 334, 0, 0, 0, 789, 0, 983, 0, 0, 0, 0, 0, 0, 607, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 161, 0, 0, 0, 451, 0, 210, 0, 0, 0, 0, 0, 0, 482, 0, 0, 159, 0, 0, 0, 0, 0, 747, 0, 13, 0, 0, 0, 0, 1471, 0, 430, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 308, 0, 0, 0, 0, 0, 384, 0, 67, 0, 0, 386, 0, 0, 0, 0, 511, 0, 0, 181, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 152, 0, 0, 0, 0, 0, 0, 4, 273, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 55, 104, 307, 0, 340, 72, 0, 0, 0, 0, 0, 0, 0, 0, 0, 335, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 814, 0, 206, 0, 0, 0, 0, 0, 576, 0, 0, 0, 611, 0, 0, 0, 0, 0, 0, 0, 0, 107, 414, 0, 0, 69, 0, 0, 0, 0, 163, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 202, 211, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 186, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 155, 0, 475, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 748, 205, 0, 0, 0, 0, 0, 0, 0, 630, 0, 0, 0, 0, 835, 409, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 352, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1197, 181, 0, 0, 0, 0, 0, 0, 0, 0, 0, 404, 0, 0, 0, 0, 0, 0, 0, 77, 0, 0, 0, 0, 17, 0, 0, 0, 0, 180, 0, 0, 0, 703, 1131, 0, 0, 128, 0, 107, 0, 0, 0, 281, 0, 0, 0, 0, 0, 0, 0, 0, 441, 0, 365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 625, 0, 0, 0, 0, 0, 0, 0, 0, 342, 0, 528, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 427, 0, 0, 0, 868, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 342, 0, 0, 29, 0, 0, 0, 0, 0, 268, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 972, 47, 0, 0, 0, 191, 0, 0, 0, 0, 0, 264, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 438, 0, 25, 613, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1440, 222, 0, 289, 0, 0, 0, 0, 419, 0, 0, 0, 0, 0, 0, 0, 0, 0, 546, 292, 0, 0, 0, 652, 539, 0, 0, 0, 223, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 449, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 435, 0, 0, 0, 0, 0, 0, 0, 0, 317, 0, 0, 0, 0, 0, 0, 0, 132, 0, 0, 436, 0, 0, 0, 0, 0, 0, 0, 254, 279, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 271, 0, 0, 0, 0, 0, 557, 0, 0, 0, 0, 0, 0, 0, 0, 284, 0, 0, 0, 0, 0, 0, 0, 0, 0, 193, 507, 0, 0, 0, 0, 0, 378, 191, 0, 0, 58, 0, 0, 0, 0, 0, 157, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 183, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 593, 0, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 440, 0, 0, 0, 427, 0, 0, 0, 0, 0, 0, 84, 0, 0, 55, 0, 25, 0, 0, 0, 0, 0, 0, 871, 0, 0, 283, 0, 0, 1011, 0, 224, 698, 0, 0, 0, 194, 0, 0, 0, 0, 0, 0, 0, 517, 0, 0, 0, 0, 0, 142, 0, 0, 0, 0, 0, 0, 128, 0, 0, 0, 0, 0, 0, 0, 0, 107, 0, 0, 0, 179, 0, 0, 593, 341, 0, 0, 0, 0, 0, 0, 0, 118, 0, 0, 0, 0, 0, 0, 0, 0, 4, 40, 0, 0, 0, 0, 325, 9, 0, 379, 434, 0, 0, 0, 226, 0, 0, 0, 177, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 252, 0, 0, 287, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 234, 102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 380, 48, 0, 0, 0, 0, 1519, 0, 0, 0, 149, 0, 108, 0, 553, 0, 0, 0, 0, 0, 34, 0, 0, 1, 0, 383, 0, 0, 0, 0, 299, 22, 142, 46, 0, 85, 0, 0, 96, 0, 0, 0, 0, 0, 254, 0, 0, 0, 74, 0, 0, 563, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 357, 0, 0, 122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 255, 0, 0, 0, 0, 0, 0, 0, 340, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 336, 0, 0, 0, 0, 0, 0, 0, 403, 0, 0, 0, 0, 269, 0, 0, 0, 280, 0, 0, 0, 0, 0, 0, 462, 0, 0, 0, 0, 0, 0, 0, 0, 338, 0, 0, 313, 0, 0, 67, 0, 0, 0, 0, 0, 0, 0, 1, 172, 0, 0, 0, 154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 496, 0, 0, 0, 0, 0, 155, 0, 0, 323, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 593, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 259, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 275, 0, 0, 120, 0, 0, 0, 596, 0, 0, 0, 0, 0, 0, 0, 0, 141, 0, 38, 0, 0, 0, 0, 398, 300, 0, 0, 60, 0, 0, 0, 0, 0, 0, 89, 0, 0, 0, 477, 0, 0, 0, 0, 365, 0, 430, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 217, 0, 0, 0, 0, 82, 0, 0, 0, 0, 206, 0, 0, 76, 0, 0, 0, 0, 345, 754, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 418, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 183, 0, 0, 0, 0, 0, 0, 0, 71, 0, 0, 0, 0, 0, 0, 0, 0, 211, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 276, 292, 0, 0, 0, 0, 0, 0, 0, 0, 0, 875, 0, 173, 0, 835, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 99, 0, 0, 0, 0, 0, 0, 0, 839, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 578, 0, 0, 0, 0, 389, 0, 0, 0, 115, 0, 0, 0, 0, 0, 525, 0, 0, 0, 0, 0, 0, 0, 16, 0, 571, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 267, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 704, 0, 0, 0, 0, 0, 233, 11, 587, 669, 0, 0, 136, 480, 0, 0, 0, 0, 0, 0, 0, 307, 0, 0, 0, 0, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 461, 0, 0, 64, 0, 0, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 255, 119, 149, 0, 0, 0, 0, 0, 0, 0, 399, 738, 0, 0, 0, 208, 0, 0, 264, 0, 0, 117, 0, 0, 0, 0, 0, 0, 643, 0, 0, 0, 0, 661, 0, 0, 0, 0, 0, 0, 656, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 732, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 442, 0, 163, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 801, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 306, 0, 0, 0, 36, 364, 0, 473, 0, 0, 0, 0, 108, 0, 0, 0, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 53, 0, 0, 0, 0, 0, 0, 341, 0, 0, 0, 0, 161, 0, 263, 0, 3083, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 206, 0, 0, 0, 0, 154, 0, 184, 0, 155, 0, 0, 0, 0, 149, 0, 0, 0, 0, 156, 0, 67, 0, 0, 410, 260, 0, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 882, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 222, 0, 0, 28, 0, 0, 0, 1033, 0, 0, 0, 0, 0, 0, 0, 162, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 204, 321, 0, 0, 0, 0, 0, 0, 199, 0, 0, 116, 1007, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 748, 0, 0, 0, 0, 0, 96, 0, 0, 0, 29, 0, 0, 0, 0, 0, 523, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 378, 0, 0, 118, 0, 0, 0, 0, 64, 0, 0, 106, 0, 0, 3, 0, 0, 0, 0, 0, 0, 207, 0, 0, 0, 0, 0, 0, 0, 334, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1189, 0, 189, 0, 0, 0, 0, 457, 0, 0, 0, 0, 0, 0, 0, 0, 0, 698, 0, 0, 335, 0, 0, 0, 0, 0, 337, 0, 0, 0, 0, 0, 0, 452, 0, 0, 0, 0, 0, 0, 1164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 32, 375, 0, 0, 0, 0, 0, 0, 0, 0, 620, 0, 0, 0, 243, 0, 0, 0, 0, 0, 0, 317, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 104, 0, 0, 62, 0, 85, 0, 0, 0, 420, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 214, 0, 0, 0, 0, 0, 0, 0, 0, 189, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 256, 0, 0, 0, 0, 447, 344, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 348, 0, 0, 72, 0, 0, 0, 0, 0, 88, 0, 0, 0, 0, 0, 0, 0, 356, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 576, 0, 889, 0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 608, 0, 0, 0, 0, 0, 92, 315, 0, 0, 0, 411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 223, 0, 0, 26, 0, 259, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 390, 206, 0, 0, 0, 0, 0, 0, 0, 0, 0, 185, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
