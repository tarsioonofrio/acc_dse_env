library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    241, 239, 243, 248, 245, 251, 252, 252, 248, 239, 237, 247, 259, 270, 273, 267, 252, 232, 216, 194, 183, 181, 185, 196, 202, 209, 213, 213, 208, 193, 
    243, 245, 247, 250, 251, 257, 258, 257, 250, 241, 240, 259, 264, 262, 260, 252, 228, 204, 169, 153, 141, 137, 138, 144, 165, 182, 202, 212, 211, 200, 
    244, 251, 255, 253, 254, 257, 261, 258, 252, 246, 249, 285, 259, 235, 223, 205, 178, 142, 120, 114, 105, 101, 100, 109, 119, 150, 175, 195, 206, 203, 
    224, 232, 246, 256, 257, 260, 262, 260, 253, 230, 246, 260, 219, 183, 162, 138, 121, 90, 87, 95, 95, 86, 82, 75, 82, 102, 127, 163, 194, 205, 
    174, 184, 194, 233, 258, 265, 265, 264, 261, 234, 252, 240, 188, 154, 125, 94, 70, 61, 85, 113, 113, 98, 86, 76, 80, 70, 85, 120, 168, 197, 
    145, 127, 143, 207, 255, 265, 263, 260, 255, 234, 215, 186, 162, 135, 85, 63, 60, 63, 90, 129, 140, 117, 88, 89, 77, 54, 44, 81, 142, 188, 
    141, 83, 90, 203, 258, 263, 257, 252, 233, 226, 183, 160, 161, 136, 83, 61, 63, 58, 87, 126, 148, 122, 95, 89, 74, 54, 35, 48, 107, 170, 
    148, 85, 99, 206, 256, 250, 245, 237, 254, 235, 186, 155, 170, 141, 96, 67, 64, 57, 69, 116, 156, 133, 107, 87, 72, 58, 44, 39, 71, 132, 
    161, 79, 144, 229, 253, 228, 213, 190, 249, 231, 184, 166, 178, 148, 98, 77, 55, 60, 51, 105, 170, 149, 118, 81, 70, 72, 55, 38, 39, 92, 
    160, 92, 165, 249, 263, 229, 171, 160, 210, 249, 204, 185, 185, 159, 113, 85, 65, 52, 42, 127, 186, 156, 126, 77, 74, 78, 71, 49, 32, 57, 
    143, 90, 168, 251, 261, 245, 177, 145, 174, 224, 193, 180, 207, 187, 140, 101, 84, 60, 44, 161, 193, 163, 118, 71, 74, 78, 70, 54, 42, 54, 
    144, 84, 162, 238, 237, 248, 211, 131, 135, 200, 182, 194, 231, 222, 159, 119, 103, 60, 65, 184, 198, 153, 102, 63, 63, 74, 71, 70, 66, 80, 
    147, 89, 168, 207, 203, 230, 226, 145, 126, 169, 166, 194, 226, 216, 164, 134, 123, 64, 80, 180, 190, 140, 103, 77, 65, 73, 78, 89, 94, 110, 
    152, 114, 182, 170, 160, 192, 227, 166, 130, 152, 182, 223, 238, 187, 157, 136, 121, 75, 95, 173, 173, 134, 91, 64, 56, 67, 90, 110, 125, 133, 
    161, 136, 186, 165, 131, 139, 211, 171, 134, 108, 174, 217, 186, 148, 129, 133, 124, 98, 114, 176, 166, 142, 113, 74, 56, 71, 100, 131, 144, 156, 
    174, 147, 178, 177, 117, 103, 162, 188, 146, 111, 163, 199, 165, 130, 107, 113, 121, 118, 140, 150, 131, 130, 101, 49, 38, 63, 101, 144, 159, 185, 
    183, 151, 171, 190, 129, 90, 121, 179, 144, 127, 137, 131, 153, 129, 110, 110, 104, 128, 175, 148, 126, 122, 84, 49, 41, 75, 113, 156, 187, 213, 
    192, 162, 167, 187, 144, 84, 92, 150, 146, 133, 120, 91, 131, 117, 130, 121, 94, 121, 154, 112, 107, 97, 51, 29, 50, 102, 148, 194, 219, 228, 
    193, 183, 173, 181, 160, 97, 87, 126, 150, 118, 73, 87, 117, 130, 174, 150, 99, 107, 109, 97, 74, 37, 15, 0, 46, 103, 169, 216, 224, 216, 
    176, 201, 181, 178, 165, 102, 83, 147, 185, 173, 104, 109, 122, 155, 197, 178, 124, 101, 96, 68, 38, 10, 0, 0, 30, 74, 132, 159, 155, 143, 
    145, 201, 184, 182, 174, 119, 102, 204, 220, 167, 120, 79, 85, 127, 144, 133, 99, 65, 46, 19, 0, 0, 0, 0, 0, 12, 52, 72, 63, 51, 
    86, 154, 168, 183, 181, 131, 145, 249, 252, 186, 91, 52, 58, 71, 72, 67, 48, 31, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 80, 115, 157, 176, 135, 198, 259, 242, 163, 62, 19, 15, 16, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 60, 121, 160, 160, 230, 253, 191, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 72, 104, 159, 239, 240, 109, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 53, 134, 237, 204, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 94, 178, 145, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 28, 103, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 34, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    41, 45, 39, 41, 45, 47, 44, 43, 44, 46, 39, 40, 48, 48, 50, 49, 44, 33, 23, 12, 10, 14, 19, 26, 32, 37, 39, 41, 41, 36, 
    43, 54, 47, 46, 49, 47, 45, 46, 46, 52, 42, 42, 48, 42, 44, 46, 32, 23, 8, 3, 0, 0, 3, 4, 12, 18, 29, 39, 41, 39, 
    43, 54, 54, 50, 51, 45, 44, 45, 49, 59, 32, 37, 40, 33, 25, 20, 9, 5, 4, 4, 0, 0, 1, 4, 3, 11, 16, 29, 36, 37, 
    28, 34, 41, 46, 50, 47, 44, 46, 50, 56, 10, 0, 2, 8, 0, 0, 3, 7, 11, 0, 0, 0, 0, 0, 0, 2, 7, 18, 29, 37, 
    0, 1, 9, 30, 48, 51, 47, 49, 53, 63, 24, 0, 0, 5, 1, 0, 8, 25, 12, 0, 0, 0, 0, 0, 0, 0, 2, 15, 20, 32, 
    0, 0, 12, 27, 44, 50, 47, 44, 42, 42, 30, 9, 4, 3, 7, 5, 4, 19, 6, 0, 0, 0, 0, 0, 0, 0, 0, 16, 19, 25, 
    0, 0, 28, 44, 43, 46, 46, 42, 28, 34, 25, 24, 13, 0, 0, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 8, 19, 17, 
    0, 0, 18, 28, 39, 40, 48, 45, 42, 42, 45, 24, 1, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 
    0, 0, 6, 0, 27, 33, 47, 24, 6, 0, 34, 12, 0, 0, 0, 0, 0, 0, 19, 20, 0, 0, 0, 1, 0, 0, 0, 0, 14, 18, 
    0, 0, 0, 0, 22, 43, 49, 25, 0, 0, 0, 2, 0, 0, 0, 0, 0, 5, 32, 17, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 
    0, 0, 0, 0, 13, 50, 53, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 37, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 40, 42, 59, 4, 0, 0, 13, 0, 0, 0, 0, 0, 16, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 3, 0, 0, 0, 26, 32, 45, 15, 0, 2, 16, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 13, 25, 41, 24, 14, 13, 0, 0, 0, 0, 0, 0, 8, 18, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 6, 
    0, 1, 0, 0, 0, 0, 11, 23, 34, 8, 0, 0, 0, 0, 0, 0, 0, 23, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 24, 
    0, 0, 0, 0, 0, 0, 0, 3, 35, 10, 0, 0, 0, 0, 0, 0, 0, 9, 18, 0, 0, 0, 0, 0, 0, 0, 0, 3, 20, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 18, 0, 0, 0, 0, 0, 0, 0, 0, 21, 9, 0, 0, 0, 0, 2, 14, 6, 21, 36, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 11, 0, 0, 0, 0, 0, 3, 9, 0, 0, 0, 10, 40, 41, 38, 41, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 32, 22, 20, 18, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 27, 10, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    72, 79, 84, 78, 76, 79, 80, 75, 71, 77, 84, 82, 76, 71, 68, 65, 66, 67, 66, 64, 60, 59, 61, 64, 68, 63, 58, 52, 47, 44, 
    67, 71, 76, 77, 79, 82, 81, 79, 79, 91, 105, 94, 76, 69, 70, 71, 65, 56, 60, 66, 64, 56, 49, 50, 56, 59, 58, 56, 52, 48, 
    68, 72, 76, 73, 76, 82, 80, 77, 84, 128, 169, 128, 84, 76, 72, 59, 43, 58, 90, 106, 103, 82, 66, 51, 50, 57, 60, 61, 58, 52, 
    72, 73, 75, 73, 74, 79, 77, 74, 81, 134, 174, 135, 83, 57, 44, 29, 43, 86, 126, 151, 155, 139, 105, 88, 63, 39, 47, 63, 67, 58, 
    61, 47, 62, 76, 75, 75, 76, 73, 72, 83, 121, 133, 89, 50, 46, 55, 58, 95, 157, 185, 175, 153, 142, 125, 80, 45, 35, 57, 73, 64, 
    57, 24, 56, 85, 78, 72, 75, 73, 69, 68, 79, 110, 118, 91, 72, 76, 76, 109, 175, 197, 168, 145, 139, 122, 94, 54, 23, 39, 69, 70, 
    96, 54, 75, 97, 82, 72, 78, 88, 83, 73, 94, 139, 153, 125, 96, 95, 93, 96, 146, 192, 171, 130, 108, 105, 91, 63, 30, 18, 52, 74, 
    153, 134, 147, 128, 91, 76, 99, 159, 180, 154, 156, 177, 176, 141, 103, 98, 92, 70, 103, 178, 188, 140, 104, 98, 96, 76, 42, 10, 25, 63, 
    210, 196, 212, 176, 105, 74, 131, 244, 300, 240, 194, 206, 195, 158, 117, 91, 72, 63, 110, 180, 207, 178, 121, 98, 104, 96, 67, 17, 0, 40, 
    232, 242, 251, 208, 127, 78, 110, 223, 318, 293, 241, 238, 217, 172, 130, 102, 72, 63, 151, 227, 227, 186, 128, 108, 113, 108, 89, 54, 14, 18, 
    214, 243, 278, 224, 139, 93, 61, 147, 275, 270, 230, 257, 255, 188, 152, 133, 89, 90, 188, 256, 233, 179, 128, 103, 115, 118, 103, 84, 55, 28, 
    214, 248, 270, 206, 136, 101, 67, 94, 188, 216, 221, 276, 295, 231, 172, 158, 120, 113, 201, 267, 232, 167, 121, 94, 95, 110, 121, 114, 93, 59, 
    231, 260, 253, 180, 128, 105, 75, 70, 135, 207, 236, 270, 289, 250, 197, 168, 136, 132, 213, 265, 224, 170, 128, 101, 99, 118, 138, 135, 111, 80, 
    248, 269, 271, 182, 116, 114, 93, 73, 125, 219, 290, 294, 261, 241, 206, 164, 132, 139, 207, 251, 224, 172, 121, 102, 111, 126, 145, 140, 106, 86, 
    269, 277, 298, 214, 132, 137, 131, 99, 111, 215, 299, 283, 223, 185, 164, 158, 139, 130, 182, 231, 211, 165, 128, 104, 112, 131, 133, 117, 99, 87, 
    293, 293, 317, 249, 160, 158, 175, 121, 114, 172, 206, 232, 192, 144, 141, 135, 134, 136, 129, 149, 188, 168, 105, 71, 79, 104, 110, 104, 98, 85, 
    318, 307, 324, 283, 185, 170, 204, 175, 129, 113, 140, 162, 154, 148, 145, 129, 146, 136, 100, 121, 147, 118, 74, 53, 62, 87, 109, 109, 97, 88, 
    332, 316, 323, 303, 214, 162, 196, 209, 168, 115, 116, 139, 145, 178, 185, 143, 137, 161, 154, 116, 81, 74, 52, 46, 73, 86, 110, 110, 96, 89, 
    325, 317, 316, 305, 238, 176, 202, 229, 200, 128, 91, 120, 170, 233, 246, 179, 128, 134, 131, 101, 66, 39, 31, 55, 83, 96, 102, 100, 87, 80, 
    315, 311, 304, 296, 239, 191, 254, 294, 239, 192, 156, 179, 243, 280, 292, 244, 155, 105, 77, 67, 69, 54, 61, 79, 95, 119, 116, 107, 95, 89, 
    311, 316, 302, 286, 232, 219, 321, 409, 358, 270, 223, 224, 249, 273, 281, 243, 179, 115, 77, 76, 87, 104, 112, 118, 122, 136, 146, 145, 130, 126, 
    287, 317, 309, 298, 266, 277, 355, 428, 417, 297, 201, 192, 202, 209, 210, 193, 167, 147, 128, 120, 123, 135, 150, 160, 164, 173, 184, 180, 175, 173, 
    232, 284, 306, 305, 288, 316, 388, 410, 332, 244, 188, 157, 157, 156, 158, 163, 154, 143, 141, 148, 157, 158, 165, 179, 190, 190, 192, 194, 191, 186, 
    183, 221, 270, 275, 288, 354, 405, 357, 263, 202, 167, 154, 151, 146, 144, 143, 144, 146, 148, 156, 167, 172, 181, 195, 205, 202, 200, 201, 203, 215, 
    185, 171, 200, 241, 292, 369, 386, 300, 218, 181, 168, 164, 158, 152, 150, 148, 148, 152, 157, 164, 178, 189, 199, 203, 200, 200, 202, 217, 239, 254, 
    201, 173, 163, 199, 279, 372, 366, 271, 193, 168, 172, 168, 160, 154, 153, 152, 156, 160, 167, 176, 186, 198, 202, 199, 192, 190, 210, 244, 251, 237, 
    206, 186, 172, 167, 226, 331, 336, 241, 179, 166, 175, 181, 170, 159, 155, 154, 159, 167, 176, 181, 183, 193, 199, 197, 190, 202, 229, 235, 214, 198, 
    209, 192, 186, 173, 169, 237, 267, 200, 161, 159, 168, 180, 184, 173, 162, 162, 171, 179, 182, 186, 186, 181, 181, 193, 212, 235, 240, 228, 196, 173, 
    207, 192, 189, 183, 164, 161, 193, 172, 134, 137, 150, 161, 169, 171, 171, 175, 182, 192, 200, 197, 185, 176, 179, 204, 243, 267, 266, 236, 185, 152, 
    213, 189, 185, 183, 176, 157, 150, 146, 127, 123, 127, 133, 140, 145, 147, 158, 180, 205, 217, 203, 185, 176, 181, 211, 257, 283, 267, 219, 185, 154, 
    
    -- channel=4
    25, 23, 27, 24, 11, 7, 11, 11, 11, 12, 14, 18, 20, 23, 24, 20, 16, 24, 44, 63, 71, 69, 59, 46, 29, 13, 13, 16, 15, 11, 
    19, 13, 18, 17, 9, 6, 10, 11, 5, 0, 0, 0, 18, 24, 19, 17, 31, 54, 60, 52, 51, 67, 80, 86, 83, 58, 28, 13, 8, 2, 
    6, 0, 8, 14, 9, 13, 17, 18, 7, 0, 0, 0, 2, 22, 41, 84, 115, 78, 12, 0, 0, 0, 0, 28, 45, 60, 52, 27, 16, 13, 
    22, 27, 28, 28, 20, 23, 26, 24, 17, 0, 27, 69, 69, 90, 131, 137, 100, 26, 0, 0, 0, 0, 0, 0, 0, 29, 64, 45, 20, 12, 
    74, 122, 104, 47, 16, 13, 18, 13, 14, 34, 112, 173, 90, 62, 70, 48, 0, 0, 0, 0, 0, 10, 0, 0, 0, 28, 46, 47, 28, 13, 
    59, 90, 70, 39, 20, 17, 14, 9, 13, 39, 61, 47, 0, 0, 0, 0, 0, 0, 0, 0, 2, 30, 21, 17, 35, 31, 15, 25, 37, 30, 
    0, 0, 0, 0, 17, 19, 9, 0, 9, 34, 7, 0, 0, 0, 0, 0, 0, 0, 24, 40, 22, 15, 35, 53, 43, 10, 10, 16, 32, 31, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 26, 15, 12, 35, 42, 23, 31, 28, 0, 0, 18, 8, 0, 0, 5, 34, 51, 
    0, 0, 0, 0, 16, 27, 0, 0, 0, 0, 0, 0, 15, 26, 0, 0, 29, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 52, 
    36, 0, 0, 14, 25, 16, 24, 42, 79, 83, 23, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 15, 38, 12, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 38, 34, 4, 24, 50, 142, 155, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 68, 70, 20, 8, 15, 0, 0, 0, 0, 
    40, 0, 2, 101, 92, 28, 26, 0, 35, 104, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 74, 58, 16, 21, 27, 0, 0, 0, 0, 
    10, 0, 0, 106, 98, 47, 40, 8, 13, 35, 0, 0, 50, 76, 0, 0, 26, 0, 0, 20, 66, 28, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 58, 20, 24, 35, 0, 0, 0, 0, 0, 68, 129, 69, 38, 34, 0, 0, 34, 54, 40, 33, 9, 0, 0, 0, 0, 10, 0, 
    0, 0, 1, 16, 0, 0, 10, 0, 0, 0, 0, 94, 102, 91, 82, 80, 51, 0, 0, 38, 48, 17, 32, 26, 8, 10, 26, 52, 25, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 39, 132, 235, 188, 74, 56, 42, 9, 0, 40, 127, 95, 48, 45, 44, 36, 45, 40, 20, 0, 0, 
    0, 0, 0, 32, 16, 0, 0, 0, 0, 30, 129, 103, 54, 0, 0, 0, 0, 0, 5, 58, 83, 130, 124, 78, 36, 14, 0, 0, 0, 0, 
    22, 0, 1, 26, 22, 0, 10, 40, 0, 0, 30, 15, 0, 0, 0, 0, 0, 11, 0, 0, 7, 121, 99, 2, 0, 0, 0, 0, 0, 15, 
    40, 4, 5, 19, 31, 0, 0, 0, 42, 58, 5, 0, 0, 0, 0, 0, 0, 59, 115, 111, 111, 85, 41, 0, 0, 0, 0, 8, 36, 38, 
    36, 12, 8, 27, 65, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 107, 139, 100, 5, 0, 0, 0, 8, 36, 74, 76, 72, 
    13, 18, 6, 26, 58, 0, 0, 0, 0, 0, 0, 0, 0, 31, 106, 111, 72, 31, 2, 0, 0, 0, 0, 0, 0, 0, 33, 55, 49, 38, 
    51, 69, 11, 4, 0, 0, 0, 0, 59, 109, 106, 140, 184, 226, 238, 212, 150, 83, 19, 0, 0, 0, 0, 0, 0, 0, 1, 6, 2, 0, 
    102, 158, 74, 41, 12, 0, 0, 27, 198, 264, 193, 100, 94, 101, 93, 82, 49, 18, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 101, 112, 100, 33, 0, 0, 148, 249, 184, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 64, 109, 9, 0, 26, 202, 200, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 6, 0, 0, 0, 
    0, 0, 11, 54, 19, 0, 90, 174, 89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 26, 0, 0, 0, 11, 
    1, 0, 0, 1, 30, 89, 177, 162, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 19, 1, 0, 0, 0, 56, 95, 
    0, 0, 0, 0, 21, 122, 250, 184, 64, 35, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 53, 49, 
    0, 0, 0, 0, 0, 39, 134, 136, 36, 32, 32, 39, 43, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    11, 0, 0, 0, 0, 0, 10, 32, 11, 0, 0, 18, 38, 56, 57, 33, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 25, 0, 
    
    -- channel=5
    117, 117, 112, 108, 111, 109, 109, 108, 108, 106, 106, 111, 118, 121, 120, 116, 110, 110, 108, 109, 110, 111, 113, 106, 103, 102, 104, 107, 103, 98, 
    116, 119, 115, 109, 109, 109, 109, 108, 104, 86, 84, 93, 108, 115, 112, 105, 107, 96, 96, 85, 86, 97, 107, 118, 115, 113, 107, 104, 100, 96, 
    106, 113, 114, 112, 110, 113, 111, 113, 108, 67, 55, 51, 88, 104, 110, 119, 110, 89, 63, 35, 27, 35, 60, 73, 98, 108, 111, 106, 103, 98, 
    101, 112, 119, 118, 117, 118, 117, 117, 120, 127, 97, 80, 101, 121, 120, 117, 95, 73, 41, 20, 9, 13, 16, 31, 57, 85, 110, 109, 102, 96, 
    112, 127, 140, 129, 118, 114, 114, 115, 119, 146, 132, 108, 90, 85, 81, 72, 61, 51, 37, 27, 28, 31, 28, 34, 32, 64, 96, 111, 105, 96, 
    70, 96, 127, 131, 121, 118, 114, 110, 109, 118, 105, 80, 51, 29, 30, 31, 44, 56, 47, 32, 34, 44, 55, 46, 45, 46, 76, 104, 111, 103, 
    12, 22, 67, 93, 113, 116, 110, 91, 95, 80, 75, 53, 30, 26, 37, 40, 44, 74, 80, 59, 35, 46, 64, 60, 50, 40, 60, 94, 110, 108, 
    0, 0, 22, 56, 95, 110, 77, 39, 0, 1, 20, 37, 27, 34, 43, 53, 57, 72, 87, 74, 34, 30, 42, 51, 42, 31, 37, 77, 109, 114, 
    0, 0, 11, 53, 87, 113, 75, 41, 0, 0, 2, 31, 29, 25, 39, 38, 59, 55, 58, 45, 14, 20, 24, 35, 41, 32, 29, 47, 92, 116, 
    4, 22, 18, 49, 82, 100, 126, 99, 66, 30, 33, 23, 22, 22, 28, 33, 44, 37, 41, 19, 8, 30, 34, 49, 40, 36, 26, 28, 52, 95, 
    17, 35, 35, 46, 84, 90, 118, 112, 110, 74, 61, 36, 10, 12, 20, 21, 20, 24, 54, 22, 30, 39, 45, 57, 53, 47, 30, 23, 29, 63, 
    6, 31, 42, 57, 104, 104, 91, 92, 95, 64, 65, 39, 7, 0, 17, 24, 12, 27, 56, 34, 37, 40, 47, 55, 62, 53, 40, 24, 27, 45, 
    0, 25, 21, 52, 105, 116, 93, 93, 84, 49, 43, 43, 36, 22, 25, 34, 23, 45, 55, 36, 23, 25, 30, 33, 43, 40, 32, 26, 40, 49, 
    3, 26, 0, 23, 65, 103, 83, 77, 66, 38, 9, 21, 30, 59, 54, 44, 35, 60, 64, 38, 34, 35, 41, 41, 38, 38, 40, 48, 56, 70, 
    1, 18, 0, 0, 20, 68, 55, 82, 57, 78, 62, 40, 52, 66, 71, 60, 53, 64, 78, 49, 35, 30, 39, 51, 54, 57, 68, 72, 74, 82, 
    0, 10, 0, 0, 18, 40, 42, 51, 72, 109, 112, 100, 88, 66, 67, 51, 44, 81, 104, 93, 73, 48, 42, 65, 74, 71, 73, 69, 79, 80, 
    0, 4, 7, 0, 12, 34, 41, 15, 57, 88, 87, 86, 52, 40, 36, 32, 44, 62, 55, 88, 95, 76, 78, 72, 81, 78, 72, 72, 85, 90, 
    6, 5, 11, 0, 0, 31, 52, 27, 24, 47, 54, 71, 33, 24, 2, 15, 54, 60, 25, 41, 61, 75, 72, 47, 49, 60, 72, 80, 90, 98, 
    26, 12, 15, 3, 0, 14, 18, 32, 32, 38, 63, 55, 35, 25, 0, 0, 48, 85, 95, 78, 68, 73, 56, 56, 46, 69, 81, 89, 93, 98, 
    40, 14, 21, 18, 12, 15, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 53, 82, 80, 56, 30, 17, 25, 32, 63, 73, 78, 80, 75, 
    37, 11, 20, 17, 6, 4, 8, 0, 0, 0, 0, 1, 27, 38, 42, 26, 20, 25, 19, 14, 7, 0, 0, 0, 8, 22, 35, 37, 32, 31, 
    44, 27, 17, 0, 0, 0, 4, 0, 0, 0, 40, 80, 91, 100, 93, 65, 48, 30, 9, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    65, 63, 42, 25, 0, 12, 3, 24, 37, 41, 52, 46, 44, 45, 43, 28, 17, 13, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 62, 66, 46, 22, 34, 23, 36, 24, 28, 6, 0, 0, 0, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 60, 44, 34, 27, 30, 15, 23, 10, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 43, 49, 44, 16, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 72, 72, 37, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 
    0, 0, 0, 0, 54, 91, 62, 33, 23, 14, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 4, 48, 38, 31, 15, 20, 24, 21, 17, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 7, 7, 3, 7, 11, 14, 24, 28, 30, 23, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    86, 89, 88, 80, 79, 76, 75, 75, 77, 79, 78, 80, 88, 94, 93, 89, 83, 88, 96, 107, 109, 108, 104, 91, 81, 72, 72, 75, 71, 64, 
    82, 87, 88, 80, 78, 75, 77, 73, 68, 48, 42, 52, 77, 89, 85, 81, 94, 96, 98, 80, 78, 89, 107, 121, 113, 100, 80, 69, 63, 58, 
    74, 77, 79, 83, 81, 83, 82, 83, 74, 9, 0, 0, 54, 82, 102, 129, 138, 97, 39, 0, 0, 0, 26, 54, 83, 87, 88, 77, 70, 63, 
    82, 90, 94, 91, 88, 90, 90, 88, 90, 85, 96, 88, 101, 133, 155, 158, 100, 44, 0, 0, 0, 0, 0, 0, 19, 66, 96, 85, 71, 61, 
    125, 137, 140, 103, 83, 84, 83, 82, 90, 156, 167, 133, 97, 91, 73, 45, 17, 7, 0, 0, 0, 8, 0, 0, 2, 46, 73, 84, 76, 62, 
    80, 94, 99, 90, 83, 86, 82, 81, 85, 116, 108, 65, 17, 0, 0, 0, 0, 13, 12, 7, 16, 25, 33, 32, 24, 22, 50, 75, 86, 75, 
    0, 0, 0, 27, 72, 87, 80, 62, 76, 70, 45, 4, 0, 0, 2, 8, 17, 53, 68, 58, 23, 25, 56, 55, 35, 5, 24, 66, 85, 78, 
    0, 0, 0, 0, 49, 79, 42, 0, 0, 0, 0, 0, 6, 21, 22, 32, 39, 69, 81, 63, 15, 6, 17, 25, 11, 0, 0, 44, 83, 96, 
    0, 0, 0, 2, 46, 92, 34, 0, 0, 0, 0, 15, 20, 5, 10, 11, 48, 29, 13, 3, 0, 0, 0, 1, 3, 0, 0, 13, 65, 98, 
    0, 0, 0, 10, 35, 77, 115, 129, 111, 44, 26, 7, 4, 0, 5, 0, 19, 0, 0, 0, 0, 16, 21, 23, 11, 2, 0, 0, 9, 64, 
    8, 20, 13, 15, 44, 56, 133, 149, 163, 104, 72, 19, 0, 0, 0, 0, 0, 0, 0, 0, 30, 45, 38, 37, 27, 21, 0, 0, 0, 17, 
    0, 1, 32, 54, 92, 74, 80, 90, 119, 84, 53, 5, 0, 0, 0, 0, 0, 0, 18, 32, 46, 39, 31, 36, 47, 35, 7, 0, 0, 0, 
    0, 0, 26, 56, 88, 89, 76, 86, 94, 28, 7, 20, 48, 26, 0, 7, 2, 6, 31, 38, 22, 7, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 1, 0, 9, 31, 72, 60, 53, 41, 0, 0, 9, 47, 74, 47, 44, 21, 20, 45, 43, 24, 14, 28, 16, 2, 0, 0, 15, 18, 14, 
    0, 3, 0, 0, 0, 37, 21, 39, 22, 58, 55, 82, 79, 77, 88, 64, 29, 20, 57, 44, 36, 18, 19, 26, 29, 39, 53, 55, 34, 27, 
    0, 0, 0, 0, 0, 10, 9, 22, 36, 129, 185, 165, 122, 69, 65, 42, 14, 37, 111, 131, 87, 36, 30, 59, 68, 68, 63, 33, 27, 36, 
    0, 0, 1, 0, 0, 0, 15, 0, 25, 101, 122, 100, 37, 2, 5, 2, 0, 34, 55, 79, 93, 106, 97, 68, 64, 35, 17, 4, 28, 51, 
    2, 0, 6, 0, 0, 5, 43, 9, 2, 29, 22, 53, 0, 0, 0, 0, 17, 33, 0, 6, 66, 88, 69, 12, 0, 0, 4, 29, 55, 70, 
    33, 4, 8, 0, 0, 0, 0, 8, 6, 34, 45, 44, 4, 0, 0, 0, 17, 77, 111, 108, 91, 72, 35, 20, 0, 16, 43, 71, 81, 87, 
    48, 8, 13, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 107, 108, 50, 0, 0, 0, 0, 42, 71, 88, 86, 83, 
    39, 4, 10, 22, 7, 0, 0, 0, 0, 0, 0, 0, 19, 64, 78, 54, 21, 20, 2, 0, 0, 0, 0, 0, 0, 7, 26, 26, 22, 18, 
    64, 39, 12, 0, 0, 0, 0, 0, 0, 35, 87, 135, 169, 186, 175, 134, 78, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    99, 98, 58, 25, 0, 0, 0, 59, 134, 132, 93, 68, 65, 64, 57, 28, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 75, 86, 78, 6, 0, 26, 115, 113, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 74, 61, 9, 0, 67, 95, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 39, 35, 50, 70, 29, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 78, 116, 104, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 30, 
    0, 0, 0, 0, 69, 141, 139, 64, 20, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 67, 63, 38, 6, 5, 12, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 21, 23, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    153, 150, 143, 142, 148, 152, 152, 153, 152, 145, 139, 143, 153, 157, 158, 158, 152, 146, 138, 131, 126, 127, 130, 132, 135, 139, 142, 146, 147, 148, 
    160, 155, 144, 140, 148, 153, 153, 154, 154, 140, 134, 139, 149, 154, 151, 145, 137, 124, 119, 114, 110, 113, 114, 116, 123, 135, 144, 150, 152, 151, 
    157, 155, 149, 143, 147, 153, 152, 153, 152, 140, 136, 128, 136, 141, 130, 118, 107, 103, 110, 102, 99, 96, 101, 102, 110, 130, 143, 147, 150, 150, 
    141, 143, 146, 150, 151, 153, 152, 154, 154, 146, 127, 107, 120, 119, 103, 93, 100, 108, 97, 87, 89, 95, 93, 97, 107, 109, 129, 142, 145, 145, 
    115, 124, 147, 161, 158, 154, 155, 157, 156, 126, 109, 122, 116, 101, 102, 117, 111, 95, 87, 84, 85, 86, 92, 99, 92, 101, 121, 135, 141, 139, 
    98, 104, 151, 173, 163, 156, 156, 151, 148, 136, 120, 120, 120, 111, 106, 108, 102, 95, 94, 86, 80, 87, 95, 90, 96, 105, 108, 120, 135, 140, 
    96, 107, 135, 158, 160, 156, 151, 140, 133, 122, 123, 117, 105, 98, 95, 99, 100, 93, 90, 90, 87, 88, 87, 90, 98, 104, 112, 110, 127, 144, 
    83, 104, 125, 133, 151, 154, 137, 123, 113, 106, 108, 93, 79, 83, 85, 93, 99, 89, 81, 95, 94, 87, 86, 95, 102, 104, 106, 108, 120, 140, 
    81, 85, 101, 130, 144, 145, 124, 109, 88, 76, 55, 64, 67, 80, 88, 87, 92, 96, 97, 91, 86, 95, 89, 89, 99, 104, 106, 102, 104, 127, 
    69, 82, 83, 125, 145, 141, 105, 65, 47, 53, 50, 59, 67, 78, 87, 87, 100, 96, 104, 91, 75, 84, 83, 93, 97, 97, 101, 105, 101, 110, 
    57, 65, 86, 119, 141, 143, 95, 41, 62, 63, 58, 65, 79, 76, 89, 96, 97, 97, 98, 76, 65, 78, 87, 91, 96, 103, 96, 99, 102, 110, 
    57, 64, 77, 99, 135, 146, 121, 67, 65, 67, 75, 79, 84, 84, 89, 94, 97, 87, 78, 68, 74, 82, 93, 91, 90, 97, 99, 100, 104, 119, 
    64, 64, 60, 82, 132, 150, 134, 89, 78, 91, 91, 66, 71, 79, 86, 83, 90, 83, 73, 72, 75, 86, 92, 91, 94, 100, 101, 99, 109, 128, 
    60, 55, 63, 83, 109, 140, 138, 108, 96, 94, 82, 56, 51, 79, 90, 80, 86, 91, 78, 72, 81, 92, 88, 89, 98, 95, 97, 105, 114, 139, 
    53, 45, 63, 83, 86, 115, 129, 132, 104, 85, 76, 58, 56, 77, 75, 88, 110, 102, 86, 83, 82, 80, 91, 92, 92, 92, 96, 110, 129, 146, 
    44, 38, 55, 76, 79, 90, 108, 115, 103, 84, 41, 70, 92, 84, 91, 90, 106, 116, 99, 79, 95, 98, 89, 86, 86, 89, 99, 119, 139, 140, 
    43, 36, 47, 71, 72, 71, 95, 106, 101, 75, 67, 90, 99, 101, 97, 89, 111, 109, 83, 97, 107, 86, 86, 94, 100, 115, 129, 136, 139, 138, 
    53, 43, 48, 70, 77, 60, 73, 91, 90, 82, 87, 103, 91, 97, 90, 81, 94, 111, 111, 98, 73, 89, 103, 95, 112, 125, 138, 137, 135, 142, 
    63, 55, 55, 65, 74, 60, 59, 76, 88, 89, 76, 84, 84, 90, 84, 76, 80, 99, 97, 85, 83, 95, 97, 95, 105, 121, 129, 131, 134, 140, 
    73, 61, 58, 62, 72, 67, 70, 68, 56, 85, 90, 79, 87, 65, 61, 76, 74, 77, 78, 82, 99, 96, 89, 82, 79, 96, 100, 105, 107, 108, 
    71, 61, 58, 57, 66, 72, 80, 81, 70, 65, 78, 68, 49, 35, 44, 56, 70, 76, 74, 88, 93, 93, 81, 66, 68, 70, 80, 91, 87, 87, 
    57, 60, 54, 57, 76, 82, 65, 43, 62, 48, 35, 42, 33, 33, 38, 43, 59, 79, 83, 79, 75, 68, 62, 58, 58, 62, 70, 69, 67, 67, 
    45, 62, 57, 63, 76, 72, 47, 32, 19, 31, 62, 54, 50, 52, 54, 63, 70, 70, 69, 68, 68, 62, 58, 58, 59, 59, 57, 59, 60, 58, 
    46, 59, 63, 57, 64, 73, 47, 27, 25, 63, 71, 66, 63, 63, 64, 65, 68, 68, 68, 67, 64, 63, 61, 60, 60, 58, 55, 54, 52, 57, 
    61, 57, 52, 65, 71, 60, 36, 27, 52, 70, 62, 60, 58, 60, 63, 67, 70, 71, 70, 65, 63, 63, 61, 58, 54, 54, 51, 52, 59, 62, 
    62, 62, 51, 58, 63, 48, 37, 49, 73, 64, 61, 59, 60, 64, 64, 65, 65, 65, 62, 60, 59, 59, 54, 50, 52, 51, 52, 60, 58, 45, 
    59, 62, 57, 47, 41, 44, 54, 65, 76, 65, 60, 65, 63, 64, 63, 60, 58, 57, 57, 54, 52, 55, 57, 57, 55, 55, 58, 48, 42, 44, 
    57, 58, 55, 49, 34, 36, 66, 71, 77, 72, 65, 64, 67, 65, 60, 58, 57, 57, 54, 54, 58, 57, 56, 60, 63, 60, 45, 37, 52, 63, 
    52, 54, 52, 52, 50, 40, 66, 88, 73, 72, 69, 67, 67, 67, 67, 64, 59, 55, 57, 58, 58, 61, 62, 66, 63, 52, 43, 52, 61, 62, 
    58, 54, 51, 53, 64, 66, 67, 79, 77, 74, 69, 65, 68, 71, 71, 65, 62, 63, 64, 59, 59, 66, 66, 63, 55, 49, 42, 45, 60, 67, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 47, 63, 53, 23, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 49, 56, 39, 44, 60, 32, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 27, 14, 22, 0, 0, 4, 55, 35, 12, 33, 72, 75, 1, 0, 0, 0, 
    99, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 42, 19, 37, 0, 0, 0, 44, 42, 8, 16, 61, 75, 49, 0, 0, 0, 
    137, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 63, 52, 26, 41, 20, 0, 0, 15, 55, 37, 20, 35, 65, 72, 13, 0, 0, 
    124, 25, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 31, 56, 59, 47, 55, 26, 0, 0, 1, 53, 69, 25, 20, 51, 73, 68, 0, 0, 
    98, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 43, 50, 51, 53, 79, 15, 0, 0, 24, 54, 79, 20, 9, 43, 68, 85, 32, 0, 
    117, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 21, 70, 31, 46, 96, 5, 0, 0, 55, 64, 79, 23, 0, 31, 57, 77, 59, 0, 
    125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 84, 38, 20, 95, 0, 0, 0, 79, 74, 70, 33, 8, 7, 34, 60, 53, 9, 
    109, 0, 52, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 34, 28, 82, 0, 0, 0, 79, 73, 73, 49, 25, 3, 12, 44, 37, 0, 
    91, 0, 75, 131, 0, 0, 0, 0, 0, 0, 0, 2, 38, 25, 13, 33, 67, 0, 0, 0, 65, 66, 70, 41, 14, 3, 0, 22, 6, 0, 
    87, 0, 55, 165, 25, 0, 0, 0, 0, 0, 0, 35, 74, 20, 0, 13, 33, 0, 0, 0, 41, 63, 74, 47, 0, 0, 0, 0, 0, 0, 
    97, 0, 29, 160, 105, 0, 0, 1, 0, 0, 0, 0, 49, 5, 5, 15, 0, 0, 0, 0, 0, 55, 81, 45, 1, 0, 0, 0, 0, 0, 
    101, 28, 24, 131, 159, 0, 0, 16, 2, 0, 0, 0, 1, 0, 22, 46, 0, 0, 0, 0, 0, 42, 70, 41, 0, 0, 0, 0, 0, 0, 
    77, 49, 29, 96, 170, 40, 0, 10, 31, 47, 0, 0, 0, 0, 35, 106, 0, 0, 0, 15, 22, 45, 61, 24, 0, 0, 0, 0, 0, 0, 
    26, 45, 24, 64, 154, 85, 0, 33, 52, 76, 10, 0, 0, 0, 33, 145, 33, 0, 0, 26, 71, 69, 48, 18, 0, 0, 0, 0, 0, 0, 
    0, 38, 11, 48, 140, 77, 0, 45, 134, 102, 51, 0, 0, 0, 35, 138, 108, 32, 41, 53, 79, 91, 77, 66, 15, 0, 0, 0, 0, 0, 
    0, 46, 14, 52, 136, 34, 0, 0, 151, 157, 90, 20, 1, 3, 48, 118, 124, 103, 106, 109, 106, 108, 121, 125, 113, 75, 57, 72, 88, 86, 
    0, 43, 25, 55, 112, 0, 0, 0, 103, 204, 139, 68, 62, 68, 83, 129, 144, 130, 146, 147, 149, 147, 157, 172, 182, 174, 165, 172, 186, 191, 
    47, 34, 13, 52, 56, 0, 0, 21, 162, 216, 184, 138, 135, 140, 140, 160, 174, 166, 170, 172, 180, 185, 188, 193, 199, 204, 197, 201, 213, 214, 
    176, 77, 10, 50, 1, 0, 0, 130, 223, 218, 186, 170, 175, 174, 172, 176, 185, 187, 189, 191, 198, 202, 200, 198, 199, 206, 207, 214, 216, 208, 
    257, 169, 62, 38, 0, 0, 27, 220, 241, 191, 182, 184, 189, 183, 178, 180, 187, 189, 192, 198, 203, 208, 205, 206, 204, 207, 209, 211, 209, 207, 
    276, 229, 155, 68, 0, 0, 114, 260, 226, 178, 180, 190, 198, 186, 178, 181, 186, 191, 194, 205, 210, 206, 212, 222, 228, 223, 208, 206, 221, 215, 
    276, 250, 215, 151, 0, 0, 138, 266, 190, 183, 176, 186, 205, 194, 186, 183, 186, 191, 198, 213, 222, 214, 217, 230, 238, 227, 220, 232, 249, 219, 
    281, 255, 235, 211, 113, 0, 126, 239, 178, 176, 169, 171, 191, 200, 196, 187, 188, 196, 205, 213, 227, 227, 219, 213, 215, 221, 245, 272, 286, 227, 
    280, 250, 237, 229, 197, 124, 131, 216, 193, 178, 169, 170, 174, 182, 184, 176, 182, 189, 203, 221, 228, 224, 208, 183, 176, 208, 260, 298, 293, 237, 
    265, 244, 227, 228, 213, 197, 172, 197, 208, 189, 182, 185, 181, 179, 165, 151, 155, 164, 187, 220, 222, 212, 188, 152, 142, 186, 262, 298, 270, 245, 
    
    -- channel=9
    141, 138, 133, 131, 134, 134, 135, 135, 138, 132, 123, 127, 138, 143, 147, 146, 139, 133, 126, 121, 117, 118, 120, 117, 117, 119, 126, 134, 136, 133, 
    146, 141, 135, 134, 136, 135, 135, 135, 133, 118, 110, 117, 133, 137, 133, 126, 123, 118, 120, 112, 108, 110, 114, 118, 117, 121, 125, 129, 131, 131, 
    138, 131, 127, 130, 134, 136, 135, 137, 134, 104, 82, 80, 113, 120, 116, 116, 118, 112, 95, 71, 62, 68, 86, 98, 113, 122, 125, 125, 127, 128, 
    120, 117, 122, 131, 139, 141, 141, 142, 143, 124, 96, 92, 114, 120, 120, 127, 122, 98, 65, 50, 45, 47, 52, 63, 81, 102, 121, 124, 124, 126, 
    118, 124, 139, 139, 139, 140, 140, 142, 147, 157, 154, 147, 127, 121, 120, 111, 88, 71, 62, 59, 61, 67, 67, 67, 71, 97, 114, 121, 120, 119, 
    102, 126, 148, 142, 136, 139, 138, 136, 137, 137, 127, 116, 92, 73, 69, 70, 74, 74, 69, 62, 70, 82, 83, 78, 84, 87, 100, 115, 121, 122, 
    61, 72, 93, 113, 134, 141, 134, 119, 118, 113, 104, 81, 62, 61, 68, 73, 78, 88, 88, 81, 71, 77, 88, 93, 93, 87, 94, 107, 121, 125, 
    35, 35, 43, 75, 120, 134, 112, 77, 50, 51, 56, 54, 52, 68, 78, 87, 89, 95, 104, 99, 72, 68, 80, 89, 85, 76, 80, 101, 120, 128, 
    24, 24, 28, 72, 113, 135, 98, 43, 0, 0, 11, 46, 56, 65, 73, 75, 92, 92, 85, 70, 54, 57, 58, 70, 77, 72, 72, 82, 107, 128, 
    43, 40, 35, 77, 113, 132, 123, 84, 50, 37, 43, 45, 51, 56, 68, 73, 85, 77, 63, 40, 34, 58, 68, 77, 74, 75, 73, 71, 81, 109, 
    48, 55, 52, 71, 105, 120, 132, 122, 112, 81, 68, 54, 44, 49, 65, 67, 70, 63, 55, 37, 52, 73, 83, 86, 83, 81, 69, 63, 63, 88, 
    47, 53, 55, 76, 114, 121, 120, 102, 99, 93, 86, 59, 41, 39, 53, 60, 58, 52, 57, 56, 70, 79, 83, 83, 88, 90, 79, 64, 64, 81, 
    37, 39, 47, 82, 117, 125, 122, 104, 96, 82, 60, 43, 50, 49, 53, 63, 68, 63, 60, 61, 63, 71, 73, 75, 83, 81, 71, 63, 73, 89, 
    31, 36, 41, 63, 86, 115, 114, 103, 95, 69, 37, 38, 62, 85, 73, 70, 76, 80, 76, 71, 70, 66, 68, 70, 69, 66, 68, 78, 95, 113, 
    24, 28, 34, 44, 53, 85, 86, 95, 80, 76, 44, 44, 69, 89, 98, 95, 87, 85, 97, 88, 78, 76, 89, 89, 83, 80, 86, 102, 116, 121, 
    17, 21, 26, 31, 42, 62, 74, 88, 93, 103, 110, 129, 119, 98, 101, 87, 83, 92, 103, 105, 97, 75, 71, 86, 92, 94, 102, 107, 109, 109, 
    17, 19, 30, 35, 47, 55, 63, 59, 76, 94, 114, 121, 101, 87, 79, 70, 71, 82, 102, 127, 115, 103, 111, 108, 109, 107, 110, 107, 112, 121, 
    35, 28, 37, 39, 43, 48, 64, 56, 55, 74, 86, 89, 63, 55, 45, 54, 73, 83, 65, 62, 83, 114, 111, 85, 84, 89, 103, 108, 120, 131, 
    55, 40, 45, 45, 43, 43, 52, 61, 54, 61, 71, 78, 66, 47, 27, 38, 70, 98, 101, 90, 95, 100, 88, 74, 59, 74, 91, 104, 113, 118, 
    60, 39, 46, 50, 50, 43, 24, 7, 24, 50, 55, 36, 25, 8, 14, 21, 35, 82, 116, 121, 105, 79, 63, 57, 56, 73, 71, 79, 83, 81, 
    48, 30, 39, 48, 55, 49, 26, 0, 0, 0, 0, 0, 6, 19, 38, 36, 31, 47, 60, 62, 50, 34, 20, 18, 29, 48, 61, 66, 64, 63, 
    44, 35, 31, 34, 32, 18, 8, 6, 17, 13, 42, 77, 90, 99, 103, 91, 79, 67, 46, 26, 25, 30, 33, 31, 35, 40, 45, 45, 44, 42, 
    70, 65, 45, 37, 24, 20, 12, 33, 63, 89, 99, 88, 86, 87, 88, 77, 63, 56, 52, 46, 44, 41, 41, 38, 35, 35, 38, 39, 35, 30, 
    62, 82, 73, 63, 50, 42, 28, 54, 76, 80, 53, 39, 35, 36, 43, 45, 48, 52, 51, 47, 44, 40, 34, 29, 24, 25, 24, 24, 22, 19, 
    27, 51, 71, 68, 45, 25, 36, 65, 83, 61, 40, 38, 39, 43, 48, 50, 49, 47, 42, 37, 31, 27, 24, 24, 27, 34, 29, 23, 14, 6, 
    27, 35, 52, 61, 45, 32, 45, 61, 64, 43, 39, 40, 43, 45, 44, 42, 40, 36, 34, 33, 29, 27, 26, 32, 42, 44, 36, 22, 14, 22, 
    29, 29, 29, 42, 58, 63, 68, 58, 54, 40, 39, 38, 35, 39, 42, 42, 39, 36, 34, 34, 37, 43, 44, 41, 39, 30, 20, 16, 39, 59, 
    26, 28, 26, 30, 60, 92, 102, 82, 69, 55, 47, 40, 35, 31, 34, 38, 38, 35, 34, 36, 38, 41, 45, 43, 30, 13, 9, 27, 52, 57, 
    25, 30, 29, 28, 43, 77, 98, 91, 69, 69, 66, 61, 56, 47, 40, 32, 27, 24, 26, 30, 35, 43, 43, 33, 14, 3, 6, 20, 26, 41, 
    32, 31, 32, 34, 37, 47, 58, 63, 56, 57, 60, 65, 72, 70, 66, 59, 49, 37, 27, 26, 34, 41, 36, 28, 17, 13, 17, 29, 38, 43, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 4, 7, 13, 11, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 23, 12, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 38, 37, 32, 6, 0, 0, 0, 0, 0, 0, 3, 13, 0, 0, 0, 
    0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 19, 1, 4, 25, 30, 17, 15, 3, 0, 0, 17, 13, 7, 9, 20, 21, 13, 0, 0, 
    6, 16, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 15, 15, 0, 0, 15, 27, 23, 32, 38, 27, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 24, 24, 37, 28, 0, 0, 25, 38, 40, 32, 33, 26, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 32, 39, 42, 40, 32, 0, 0, 0, 23, 28, 21, 17, 23, 29, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 37, 38, 27, 0, 0, 0, 0, 9, 15, 14, 19, 19, 25, 29, 
    0, 15, 0, 0, 0, 0, 0, 38, 6, 0, 0, 0, 0, 0, 2, 5, 25, 26, 8, 0, 0, 0, 3, 25, 22, 12, 16, 19, 15, 13, 
    6, 30, 0, 0, 0, 0, 0, 37, 59, 6, 0, 0, 0, 0, 0, 1, 0, 4, 2, 0, 0, 5, 22, 31, 29, 29, 21, 19, 7, 0, 
    2, 18, 0, 0, 0, 0, 0, 6, 31, 6, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 10, 27, 32, 36, 39, 29, 12, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 24, 2, 0, 0, 0, 0, 0, 0, 7, 20, 8, 0, 0, 1, 4, 16, 22, 17, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 21, 10, 9, 11, 17, 16, 3, 0, 6, 23, 29, 27, 9, 3, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 1, 26, 32, 29, 15, 1, 3, 7, 6, 0, 13, 31, 40, 29, 15, 12, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 38, 42, 66, 57, 30, 35, 23, 4, 0, 8, 51, 51, 11, 18, 46, 56, 49, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 9, 0, 0, 12, 52, 44, 10, 1, 0, 3, 6, 0, 0, 11, 40, 51, 59, 64, 50, 29, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 28, 3, 0, 0, 9, 28, 0, 0, 0, 0, 9, 10, 0, 0, 2, 55, 70, 45, 9, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 1, 12, 0, 0, 17, 12, 25, 5, 0, 0, 0, 0, 29, 51, 57, 60, 65, 66, 57, 15, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 1, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 85, 83, 56, 34, 38, 28, 17, 3, 4, 7, 15, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 35, 39, 30, 30, 32, 41, 41, 39, 35, 34, 49, 52, 47, 46, 48, 52, 
    60, 19, 0, 0, 0, 0, 0, 0, 0, 9, 50, 94, 113, 120, 127, 121, 96, 77, 66, 51, 49, 57, 69, 75, 77, 76, 76, 73, 75, 75, 
    104, 98, 46, 3, 0, 0, 0, 0, 30, 89, 111, 97, 97, 98, 98, 100, 91, 81, 84, 85, 82, 83, 86, 85, 79, 74, 77, 80, 82, 84, 
    90, 103, 92, 49, 4, 0, 0, 2, 70, 108, 82, 68, 67, 67, 71, 77, 84, 85, 87, 90, 88, 85, 81, 75, 68, 69, 73, 76, 73, 66, 
    78, 85, 93, 83, 28, 0, 0, 27, 90, 97, 75, 72, 77, 80, 78, 79, 82, 81, 81, 83, 81, 75, 70, 75, 81, 90, 95, 88, 66, 54, 
    91, 87, 86, 83, 63, 11, 0, 30, 78, 73, 78, 76, 76, 83, 82, 78, 77, 77, 78, 82, 86, 90, 88, 87, 97, 106, 101, 84, 72, 83, 
    97, 93, 85, 80, 81, 83, 57, 51, 80, 74, 74, 72, 66, 67, 76, 84, 87, 85, 83, 88, 92, 97, 103, 102, 99, 92, 85, 86, 104, 120, 
    86, 98, 93, 84, 88, 109, 131, 101, 99, 101, 95, 83, 74, 65, 65, 72, 73, 75, 79, 85, 91, 95, 100, 99, 84, 69, 69, 82, 99, 107, 
    83, 95, 99, 87, 84, 90, 111, 116, 95, 105, 107, 106, 107, 96, 83, 73, 68, 64, 61, 65, 77, 89, 89, 80, 62, 50, 52, 77, 88, 91, 
    87, 87, 96, 93, 85, 81, 83, 94, 90, 95, 98, 100, 108, 110, 112, 106, 94, 80, 68, 64, 72, 80, 79, 74, 61, 60, 68, 87, 99, 98, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=12
    75, 76, 71, 65, 69, 69, 68, 65, 64, 67, 72, 75, 73, 68, 65, 61, 61, 71, 76, 78, 80, 81, 81, 73, 68, 62, 57, 53, 48, 45, 
    69, 71, 67, 62, 69, 69, 69, 65, 64, 61, 67, 68, 68, 65, 63, 61, 68, 68, 77, 76, 77, 82, 85, 88, 86, 78, 65, 57, 50, 46, 
    62, 68, 66, 63, 68, 73, 69, 69, 72, 77, 82, 58, 61, 71, 76, 80, 72, 67, 76, 70, 65, 60, 66, 68, 82, 87, 81, 70, 60, 52, 
    70, 82, 79, 70, 71, 73, 69, 69, 80, 138, 139, 83, 76, 90, 85, 73, 61, 84, 96, 98, 89, 77, 62, 57, 68, 75, 90, 86, 69, 54, 
    85, 99, 106, 87, 73, 67, 65, 65, 76, 137, 136, 105, 75, 62, 57, 52, 61, 98, 122, 126, 120, 108, 90, 88, 60, 60, 83, 98, 81, 59, 
    58, 68, 111, 110, 80, 67, 64, 62, 68, 86, 87, 84, 65, 36, 42, 54, 73, 117, 149, 136, 114, 106, 116, 99, 69, 50, 64, 95, 96, 71, 
    25, 31, 91, 103, 82, 69, 68, 63, 68, 60, 76, 96, 86, 63, 74, 82, 84, 125, 167, 153, 104, 96, 108, 94, 73, 48, 51, 80, 99, 84, 
    36, 60, 108, 94, 77, 73, 70, 74, 52, 42, 85, 124, 105, 82, 81, 92, 89, 101, 145, 160, 112, 83, 78, 82, 70, 51, 35, 56, 94, 99, 
    80, 127, 144, 112, 79, 79, 103, 158, 118, 89, 106, 138, 112, 82, 77, 75, 76, 68, 120, 146, 116, 91, 68, 74, 80, 66, 39, 29, 69, 102, 
    132, 187, 175, 124, 82, 67, 146, 235, 234, 162, 146, 141, 112, 88, 77, 67, 57, 58, 138, 156, 131, 113, 79, 92, 93, 80, 53, 26, 39, 78, 
    150, 208, 202, 133, 92, 57, 104, 192, 250, 185, 165, 165, 125, 92, 79, 76, 40, 71, 190, 181, 152, 116, 86, 100, 106, 96, 69, 45, 36, 53, 
    136, 207, 207, 141, 114, 75, 45, 123, 192, 155, 164, 195, 155, 101, 93, 96, 49, 99, 213, 190, 150, 105, 87, 93, 107, 102, 90, 69, 58, 44, 
    136, 212, 177, 123, 125, 101, 43, 94, 145, 139, 170, 211, 195, 139, 119, 115, 70, 131, 211, 187, 133, 97, 81, 78, 89, 98, 103, 88, 81, 56, 
    153, 216, 152, 101, 108, 117, 56, 74, 116, 160, 187, 200, 178, 171, 150, 120, 77, 142, 206, 175, 135, 110, 90, 83, 92, 107, 117, 105, 83, 69, 
    167, 209, 161, 98, 94, 127, 76, 89, 109, 203, 247, 198, 154, 156, 147, 120, 93, 133, 183, 163, 135, 104, 85, 93, 110, 124, 129, 103, 78, 75, 
    176, 208, 192, 113, 108, 136, 112, 86, 114, 217, 239, 196, 158, 126, 124, 111, 98, 137, 164, 160, 151, 112, 76, 85, 110, 119, 110, 84, 82, 75, 
    187, 213, 216, 135, 113, 144, 154, 85, 110, 146, 148, 146, 108, 103, 101, 97, 116, 126, 84, 121, 156, 115, 78, 73, 92, 102, 90, 76, 79, 68, 
    206, 214, 223, 160, 110, 141, 174, 131, 106, 85, 98, 126, 96, 117, 96, 86, 136, 131, 71, 90, 97, 78, 61, 50, 67, 84, 90, 86, 79, 74, 
    219, 213, 220, 181, 117, 127, 157, 158, 133, 81, 99, 118, 122, 163, 121, 78, 120, 147, 140, 112, 73, 62, 51, 77, 86, 104, 104, 92, 83, 81, 
    232, 207, 214, 193, 131, 133, 165, 141, 101, 65, 92, 98, 150, 189, 155, 97, 88, 105, 111, 92, 70, 50, 51, 88, 107, 137, 133, 118, 111, 107, 
    245, 208, 211, 188, 126, 142, 233, 199, 118, 84, 114, 160, 213, 232, 217, 163, 120, 88, 55, 57, 68, 70, 83, 94, 120, 141, 146, 135, 125, 124, 
    266, 234, 218, 181, 120, 170, 275, 281, 241, 183, 182, 222, 241, 244, 231, 186, 154, 119, 93, 89, 104, 119, 131, 133, 142, 150, 160, 149, 140, 140, 
    268, 268, 250, 212, 165, 237, 288, 297, 251, 182, 172, 167, 164, 163, 160, 144, 135, 127, 128, 132, 138, 140, 145, 147, 149, 152, 158, 155, 153, 150, 
    206, 249, 269, 228, 208, 285, 302, 262, 174, 144, 130, 123, 120, 118, 123, 125, 129, 128, 132, 139, 143, 144, 145, 154, 156, 155, 154, 154, 151, 151, 
    155, 194, 238, 215, 240, 300, 288, 189, 141, 138, 134, 135, 131, 129, 129, 127, 127, 127, 132, 138, 142, 147, 155, 167, 169, 171, 168, 166, 170, 181, 
    155, 159, 184, 205, 277, 326, 250, 138, 130, 135, 141, 138, 131, 130, 129, 126, 127, 131, 137, 146, 156, 166, 172, 170, 170, 168, 174, 189, 205, 208, 
    159, 152, 151, 183, 283, 338, 238, 138, 137, 138, 143, 138, 127, 127, 131, 133, 136, 139, 146, 152, 159, 173, 176, 166, 156, 155, 185, 205, 204, 192, 
    158, 154, 152, 157, 233, 300, 232, 156, 151, 150, 157, 151, 140, 131, 126, 128, 135, 141, 148, 150, 153, 160, 161, 158, 153, 169, 186, 183, 161, 160, 
    155, 154, 157, 149, 164, 211, 179, 151, 134, 145, 159, 163, 163, 149, 140, 137, 140, 141, 143, 146, 145, 146, 147, 158, 172, 188, 178, 165, 129, 143, 
    157, 151, 153, 152, 144, 147, 138, 128, 117, 126, 135, 141, 152, 154, 158, 160, 161, 164, 163, 149, 139, 139, 148, 175, 204, 209, 187, 159, 137, 138, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 53, 3, 0, 0, 0, 0, 0, 4, 42, 49, 46, 17, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 67, 74, 53, 32, 25, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 75, 73, 40, 28, 25, 9, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 33, 9, 0, 0, 11, 30, 59, 66, 41, 18, 7, 0, 0, 0, 0, 0, 0, 
    59, 13, 4, 20, 0, 0, 0, 0, 10, 29, 21, 53, 78, 52, 16, 0, 1, 0, 0, 30, 60, 43, 13, 0, 0, 0, 0, 0, 0, 0, 
    100, 74, 82, 70, 0, 0, 0, 58, 157, 162, 113, 96, 101, 55, 27, 2, 0, 0, 0, 30, 76, 68, 38, 0, 0, 0, 0, 0, 0, 0, 
    129, 105, 126, 92, 6, 0, 6, 85, 193, 202, 145, 110, 113, 77, 30, 11, 0, 0, 0, 78, 126, 94, 53, 11, 2, 7, 0, 0, 0, 0, 
    134, 104, 142, 112, 22, 0, 0, 26, 118, 173, 123, 107, 123, 98, 40, 15, 0, 0, 24, 127, 149, 89, 40, 7, 7, 13, 5, 0, 0, 0, 
    123, 97, 158, 123, 21, 0, 0, 0, 52, 98, 81, 105, 144, 127, 68, 43, 25, 11, 51, 141, 137, 76, 29, 5, 3, 0, 4, 5, 0, 0, 
    128, 112, 158, 112, 11, 0, 0, 0, 8, 56, 83, 150, 174, 145, 88, 68, 43, 27, 67, 143, 121, 61, 28, 1, 0, 0, 11, 24, 11, 0, 
    146, 132, 156, 110, 21, 0, 0, 0, 0, 48, 104, 186, 169, 126, 101, 71, 35, 26, 67, 122, 120, 79, 44, 15, 2, 18, 32, 33, 0, 0, 
    169, 151, 162, 126, 55, 15, 6, 0, 0, 71, 173, 198, 155, 89, 67, 47, 22, 8, 43, 93, 89, 61, 26, 6, 5, 25, 34, 6, 0, 0, 
    193, 176, 184, 152, 99, 40, 47, 23, 9, 48, 124, 118, 79, 39, 29, 26, 5, 20, 42, 46, 50, 71, 38, 0, 0, 1, 1, 0, 0, 0, 
    209, 196, 198, 168, 117, 65, 67, 60, 41, 33, 35, 28, 23, 11, 24, 34, 18, 22, 2, 0, 26, 38, 3, 0, 0, 0, 0, 0, 0, 0, 
    206, 199, 197, 176, 132, 83, 82, 94, 62, 38, 11, 13, 34, 32, 58, 67, 36, 32, 32, 26, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    180, 190, 183, 175, 140, 88, 67, 115, 114, 54, 25, 5, 34, 74, 111, 92, 53, 36, 49, 36, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    158, 187, 173, 173, 150, 94, 78, 122, 135, 64, 22, 31, 84, 143, 169, 134, 74, 33, 3, 0, 0, 0, 0, 0, 10, 32, 32, 25, 16, 6, 
    157, 199, 178, 167, 132, 78, 120, 217, 223, 183, 138, 139, 178, 208, 207, 176, 123, 55, 4, 0, 0, 7, 29, 47, 57, 65, 69, 67, 59, 52, 
    168, 204, 190, 172, 134, 114, 175, 278, 308, 254, 176, 138, 143, 150, 142, 118, 92, 62, 43, 39, 48, 59, 72, 82, 85, 89, 96, 95, 89, 86, 
    154, 174, 183, 196, 162, 158, 226, 306, 274, 179, 97, 67, 67, 67, 66, 64, 65, 63, 58, 63, 73, 75, 79, 85, 90, 95, 95, 97, 97, 91, 
    113, 127, 150, 166, 151, 170, 262, 294, 206, 110, 74, 67, 71, 69, 64, 60, 59, 56, 56, 62, 71, 78, 80, 93, 103, 109, 107, 109, 105, 104, 
    110, 101, 117, 122, 140, 200, 282, 240, 137, 75, 79, 82, 79, 70, 63, 58, 54, 55, 60, 68, 78, 88, 101, 114, 120, 119, 114, 112, 125, 145, 
    117, 96, 91, 107, 139, 220, 271, 194, 94, 74, 80, 81, 78, 68, 65, 63, 64, 69, 74, 85, 98, 108, 115, 118, 112, 101, 101, 127, 161, 165, 
    118, 102, 94, 101, 144, 197, 237, 169, 84, 74, 80, 81, 78, 73, 70, 71, 73, 79, 88, 92, 97, 103, 108, 107, 97, 94, 123, 156, 158, 122, 
    124, 105, 102, 100, 117, 153, 157, 124, 72, 70, 78, 85, 88, 84, 75, 68, 74, 84, 92, 94, 96, 96, 91, 86, 91, 117, 143, 147, 118, 86, 
    129, 105, 101, 102, 91, 94, 83, 69, 49, 46, 60, 76, 83, 83, 80, 81, 87, 92, 98, 102, 96, 84, 77, 83, 109, 146, 168, 155, 109, 83, 
    124, 105, 96, 98, 90, 77, 64, 52, 44, 36, 41, 47, 53, 62, 64, 69, 82, 98, 114, 115, 97, 82, 79, 96, 137, 172, 182, 148, 101, 73, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    322, 332, 335, 337, 339, 343, 343, 341, 338, 329, 326, 335, 352, 366, 369, 362, 342, 309, 277, 249, 236, 238, 253, 270, 283, 294, 304, 307, 298, 279, 
    330, 344, 347, 346, 344, 348, 347, 348, 343, 339, 337, 341, 348, 358, 361, 346, 302, 249, 205, 178, 166, 166, 177, 195, 220, 251, 285, 304, 302, 287, 
    337, 354, 361, 356, 352, 350, 351, 349, 345, 353, 353, 351, 333, 322, 302, 263, 208, 180, 159, 146, 131, 131, 137, 140, 162, 197, 240, 276, 291, 287, 
    305, 313, 335, 347, 352, 350, 352, 351, 343, 324, 290, 284, 263, 229, 188, 155, 148, 135, 128, 110, 100, 102, 109, 124, 124, 143, 177, 230, 270, 285, 
    215, 206, 250, 319, 353, 360, 359, 360, 348, 284, 240, 206, 197, 166, 137, 124, 124, 114, 108, 95, 80, 70, 88, 91, 92, 91, 125, 184, 246, 281, 
    143, 130, 186, 282, 347, 364, 365, 359, 341, 290, 247, 215, 197, 172, 137, 115, 98, 92, 97, 105, 96, 85, 77, 76, 71, 64, 90, 145, 211, 264, 
    139, 122, 188, 278, 335, 356, 354, 345, 308, 265, 234, 213, 185, 145, 100, 80, 72, 68, 77, 96, 116, 107, 81, 75, 63, 67, 72, 111, 177, 242, 
    129, 130, 182, 275, 326, 337, 336, 338, 316, 285, 236, 188, 156, 117, 88, 66, 58, 52, 73, 97, 123, 121, 106, 89, 82, 80, 83, 92, 136, 197, 
    102, 98, 163, 241, 307, 304, 296, 272, 286, 250, 215, 162, 140, 122, 101, 79, 55, 71, 101, 130, 147, 134, 120, 101, 91, 88, 87, 87, 105, 151, 
    67, 48, 128, 221, 302, 298, 230, 141, 130, 157, 168, 164, 152, 143, 109, 98, 69, 89, 125, 151, 151, 114, 100, 86, 83, 85, 84, 88, 97, 129, 
    37, 28, 93, 206, 299, 325, 217, 123, 69, 114, 140, 166, 170, 158, 134, 108, 96, 106, 114, 130, 112, 90, 79, 68, 75, 73, 80, 83, 100, 125, 
    44, 40, 74, 162, 256, 325, 275, 174, 106, 119, 152, 168, 174, 169, 148, 121, 103, 105, 91, 105, 88, 85, 73, 64, 59, 63, 72, 84, 102, 141, 
    69, 58, 65, 119, 205, 294, 291, 195, 131, 151, 168, 158, 125, 125, 132, 115, 94, 75, 82, 90, 93, 93, 86, 75, 70, 80, 83, 93, 108, 157, 
    80, 68, 76, 94, 166, 242, 270, 207, 159, 161, 174, 141, 98, 79, 99, 96, 94, 81, 82, 90, 97, 89, 74, 71, 75, 86, 94, 102, 131, 188, 
    78, 74, 87, 83, 126, 174, 231, 205, 167, 133, 122, 92, 87, 71, 72, 83, 101, 117, 119, 114, 96, 93, 75, 60, 57, 64, 84, 118, 178, 231, 
    74, 70, 78, 75, 82, 112, 173, 178, 163, 77, 39, 40, 48, 82, 74, 79, 112, 145, 123, 92, 86, 95, 83, 55, 43, 55, 96, 169, 229, 266, 
    66, 54, 54, 67, 52, 73, 102, 168, 150, 96, 63, 77, 112, 126, 103, 85, 115, 146, 159, 121, 79, 56, 50, 44, 54, 98, 166, 241, 280, 296, 
    59, 46, 42, 62, 57, 54, 58, 105, 126, 123, 116, 105, 142, 148, 130, 92, 86, 128, 178, 142, 90, 57, 45, 69, 103, 169, 230, 271, 290, 293, 
    60, 57, 51, 61, 60, 52, 54, 69, 91, 92, 99, 95, 121, 140, 137, 101, 84, 86, 82, 61, 46, 38, 40, 44, 100, 178, 247, 271, 275, 268, 
    59, 75, 70, 61, 52, 49, 87, 111, 124, 122, 100, 133, 130, 128, 123, 107, 94, 82, 34, 7, 5, 18, 31, 7, 34, 72, 123, 139, 139, 128, 
    31, 71, 77, 61, 52, 70, 102, 155, 163, 157, 110, 75, 40, 26, 15, 13, 27, 36, 38, 13, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 11, 55, 68, 89, 119, 115, 114, 70, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 35, 82, 106, 115, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 50, 82, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 77, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=16
    264, 261, 262, 262, 262, 262, 262, 262, 261, 262, 262, 262, 263, 263, 265, 264, 263, 262, 259, 258, 255, 260, 262, 264, 263, 262, 262, 262, 262, 263, 
    266, 264, 264, 264, 264, 264, 264, 264, 263, 263, 264, 264, 264, 264, 267, 266, 263, 260, 251, 247, 232, 248, 252, 262, 265, 263, 263, 263, 264, 265, 
    265, 263, 263, 263, 263, 263, 263, 263, 263, 263, 263, 263, 263, 264, 266, 265, 261, 253, 242, 226, 214, 235, 248, 260, 264, 263, 263, 263, 264, 265, 
    267, 264, 264, 264, 264, 264, 264, 264, 263, 264, 264, 263, 263, 261, 259, 252, 238, 224, 219, 190, 190, 214, 237, 258, 265, 264, 264, 264, 265, 265, 
    261, 259, 262, 262, 264, 266, 266, 264, 264, 265, 263, 262, 257, 256, 252, 237, 214, 194, 183, 156, 155, 183, 213, 247, 266, 266, 264, 264, 265, 266, 
    253, 257, 260, 261, 265, 267, 267, 265, 266, 267, 262, 260, 242, 252, 252, 224, 196, 180, 171, 157, 156, 170, 199, 237, 265, 266, 265, 265, 267, 267, 
    244, 250, 255, 258, 264, 268, 267, 267, 266, 267, 267, 257, 233, 254, 253, 226, 195, 187, 187, 175, 174, 177, 201, 239, 261, 263, 262, 264, 266, 268, 
    167, 177, 190, 212, 239, 265, 267, 266, 266, 266, 273, 250, 235, 258, 257, 238, 221, 219, 213, 201, 197, 191, 191, 208, 217, 219, 228, 244, 262, 268, 
    140, 141, 152, 175, 215, 260, 263, 262, 264, 264, 271, 250, 244, 258, 262, 250, 238, 241, 230, 216, 200, 190, 181, 176, 173, 174, 186, 217, 258, 268, 
    142, 140, 149, 167, 219, 254, 250, 248, 251, 253, 253, 240, 238, 246, 252, 251, 248, 248, 241, 230, 209, 195, 185, 169, 161, 153, 153, 211, 256, 267, 
    146, 147, 155, 172, 222, 239, 229, 220, 221, 221, 196, 160, 161, 169, 176, 186, 202, 217, 240, 233, 209, 195, 186, 178, 175, 159, 158, 216, 250, 260, 
    134, 135, 142, 163, 194, 217, 217, 211, 220, 210, 152, 92, 90, 98, 110, 133, 165, 206, 244, 236, 221, 217, 210, 206, 203, 180, 185, 209, 219, 236, 
    83, 90, 101, 120, 160, 183, 178, 190, 216, 202, 113, 49, 53, 72, 102, 133, 158, 200, 227, 220, 206, 194, 183, 173, 171, 164, 170, 170, 172, 195, 
    20, 41, 58, 87, 119, 126, 145, 183, 209, 200, 129, 89, 89, 99, 117, 126, 141, 171, 182, 174, 159, 147, 138, 132, 139, 149, 154, 148, 152, 176, 
    0, 13, 69, 132, 122, 114, 146, 190, 210, 212, 183, 165, 160, 173, 191, 180, 173, 170, 165, 155, 142, 128, 121, 120, 123, 132, 143, 145, 143, 162, 
    0, 33, 158, 194, 159, 152, 181, 203, 216, 227, 227, 225, 220, 243, 235, 200, 176, 156, 152, 144, 135, 127, 125, 126, 121, 123, 129, 131, 131, 142, 
    0, 79, 191, 189, 161, 165, 182, 189, 201, 216, 226, 220, 209, 213, 181, 150, 128, 123, 117, 108, 110, 115, 111, 103, 97, 104, 114, 121, 124, 122, 
    7, 112, 158, 148, 140, 145, 152, 154, 155, 159, 165, 154, 152, 150, 131, 120, 110, 117, 107, 90, 95, 101, 94, 81, 78, 84, 84, 83, 86, 92, 
    21, 70, 78, 73, 74, 78, 80, 83, 85, 89, 95, 93, 98, 92, 81, 73, 77, 80, 57, 39, 44, 46, 37, 23, 21, 29, 37, 49, 67, 89, 
    5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 9, 8, 10, 14, 21, 22, 9, 0, 0, 0, 0, 0, 0, 15, 34, 51, 71, 90, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 27, 48, 63, 79, 102, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 31, 52, 68, 77, 96, 120, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 1, 15, 28, 42, 54, 71, 88, 99, 115, 134, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 68, 59, 50, 46, 46, 46, 47, 50, 57, 73, 89, 98, 102, 109, 126, 150, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 125, 124, 112, 106, 98, 90, 85, 87, 94, 97, 96, 99, 111, 122, 140, 165, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 69, 147, 162, 145, 132, 116, 103, 93, 87, 85, 92, 103, 113, 121, 130, 150, 173, 
    46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 112, 130, 106, 87, 79, 80, 80, 83, 93, 111, 122, 124, 126, 136, 158, 176, 
    62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 72, 95, 81, 69, 65, 76, 92, 108, 117, 123, 126, 128, 135, 145, 164, 181, 
    70, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 51, 66, 62, 67, 82, 102, 121, 128, 125, 123, 128, 134, 141, 152, 168, 185, 
    75, 36, 17, 7, 1, 0, 0, 0, 0, 0, 0, 0, 5, 24, 49, 63, 76, 100, 121, 130, 135, 129, 123, 126, 133, 142, 148, 157, 171, 187, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 17, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 17, 0, 0, 0, 24, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 4, 0, 5, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 2, 5, 0, 0, 0, 0, 0, 4, 6, 12, 28, 15, 18, 28, 22, 14, 10, 14, 20, 25, 25, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 9, 0, 0, 0, 0, 0, 0, 5, 11, 33, 23, 0, 24, 40, 45, 46, 42, 33, 25, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 8, 9, 11, 0, 0, 0, 0, 1, 7, 10, 34, 54, 16, 19, 38, 40, 37, 25, 9, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 9, 7, 10, 9, 5, 6, 5, 6, 9, 9, 21, 58, 69, 76, 82, 62, 38, 20, 11, 5, 9, 15, 12, 4, 0, 0, 0, 0, 0, 
    0, 0, 8, 9, 9, 6, 5, 7, 8, 8, 8, 10, 34, 62, 70, 69, 49, 31, 22, 23, 25, 25, 18, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 10, 9, 6, 6, 8, 9, 9, 8, 4, 13, 30, 26, 27, 29, 33, 33, 29, 21, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 16, 13, 10, 10, 12, 14, 15, 15, 10, 12, 23, 21, 23, 34, 40, 37, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 18, 18, 16, 16, 19, 21, 22, 24, 23, 23, 30, 34, 34, 34, 25, 17, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    429, 428, 428, 428, 428, 428, 428, 428, 428, 429, 429, 429, 430, 430, 429, 427, 426, 428, 428, 429, 430, 429, 428, 428, 428, 428, 428, 429, 430, 430, 
    431, 429, 429, 429, 429, 429, 429, 429, 428, 429, 429, 429, 430, 430, 428, 425, 423, 424, 414, 406, 411, 416, 424, 428, 429, 429, 429, 429, 430, 430, 
    431, 430, 430, 430, 430, 430, 429, 428, 428, 429, 429, 428, 429, 430, 428, 426, 423, 415, 385, 368, 387, 407, 424, 429, 429, 429, 429, 430, 431, 431, 
    432, 430, 430, 430, 430, 430, 430, 429, 430, 431, 430, 429, 429, 429, 423, 413, 401, 387, 362, 346, 369, 398, 416, 429, 430, 430, 431, 432, 433, 433, 
    426, 426, 427, 429, 431, 431, 431, 431, 431, 432, 430, 425, 426, 426, 406, 379, 365, 356, 343, 323, 328, 365, 403, 428, 432, 430, 431, 432, 434, 435, 
    422, 424, 425, 428, 432, 432, 433, 433, 433, 434, 423, 408, 418, 422, 398, 368, 355, 350, 336, 315, 309, 338, 392, 429, 434, 431, 433, 434, 436, 436, 
    428, 431, 430, 431, 433, 434, 433, 434, 433, 435, 413, 392, 408, 419, 408, 389, 380, 378, 370, 361, 353, 361, 395, 430, 437, 435, 436, 437, 438, 438, 
    354, 364, 376, 401, 426, 432, 431, 431, 432, 434, 416, 392, 402, 423, 420, 406, 411, 416, 414, 414, 409, 395, 385, 390, 394, 395, 411, 432, 440, 440, 
    268, 276, 303, 365, 418, 425, 423, 426, 430, 431, 427, 412, 410, 425, 431, 425, 425, 431, 427, 407, 383, 359, 339, 324, 314, 321, 369, 422, 440, 440, 
    284, 287, 303, 354, 401, 406, 404, 410, 416, 419, 419, 414, 413, 421, 428, 432, 433, 434, 414, 380, 360, 346, 331, 316, 288, 284, 343, 412, 438, 440, 
    352, 358, 364, 371, 384, 378, 359, 372, 387, 362, 327, 321, 330, 341, 353, 367, 389, 418, 421, 404, 394, 383, 373, 363, 333, 327, 361, 403, 432, 440, 
    324, 329, 343, 355, 369, 357, 345, 371, 370, 287, 208, 195, 205, 216, 239, 281, 352, 417, 440, 433, 421, 412, 401, 398, 391, 377, 373, 383, 406, 426, 
    220, 219, 244, 295, 331, 347, 366, 383, 370, 286, 188, 154, 168, 200, 248, 303, 358, 395, 407, 393, 375, 356, 336, 333, 341, 332, 319, 322, 350, 390, 
    148, 166, 212, 241, 242, 282, 335, 366, 375, 339, 274, 246, 273, 309, 321, 316, 318, 325, 320, 296, 272, 258, 246, 242, 253, 272, 282, 287, 319, 366, 
    115, 209, 251, 223, 209, 236, 285, 339, 380, 390, 372, 363, 374, 368, 334, 309, 298, 294, 286, 272, 254, 248, 248, 247, 258, 285, 308, 315, 323, 337, 
    123, 281, 327, 298, 277, 282, 317, 360, 397, 414, 411, 409, 419, 409, 374, 340, 325, 328, 331, 330, 322, 315, 310, 309, 311, 315, 318, 314, 300, 300, 
    182, 310, 372, 371, 349, 350, 364, 379, 394, 406, 399, 395, 400, 395, 373, 341, 334, 330, 319, 328, 338, 327, 307, 292, 282, 271, 269, 275, 276, 276, 
    237, 303, 348, 350, 347, 348, 352, 354, 357, 358, 352, 341, 327, 312, 302, 304, 302, 280, 265, 274, 282, 271, 249, 230, 229, 231, 232, 237, 243, 244, 
    210, 252, 265, 265, 273, 282, 284, 286, 289, 294, 299, 298, 290, 274, 261, 261, 263, 253, 231, 216, 216, 212, 200, 189, 188, 192, 193, 202, 219, 238, 
    118, 137, 142, 149, 155, 159, 166, 175, 186, 196, 208, 224, 233, 227, 218, 214, 215, 210, 191, 174, 168, 165, 159, 158, 163, 172, 181, 199, 217, 234, 
    18, 27, 52, 60, 54, 49, 48, 51, 58, 68, 84, 108, 125, 130, 133, 139, 141, 133, 123, 118, 117, 118, 124, 138, 161, 185, 192, 194, 207, 229, 
    0, 0, 27, 49, 35, 12, 0, 0, 0, 0, 0, 26, 62, 67, 63, 68, 71, 70, 72, 77, 90, 110, 140, 172, 191, 194, 183, 185, 208, 242, 
    0, 0, 10, 59, 53, 19, 0, 0, 0, 0, 0, 19, 107, 131, 114, 102, 103, 107, 112, 123, 142, 165, 183, 183, 170, 166, 180, 199, 224, 264, 
    0, 0, 0, 5, 23, 5, 0, 0, 0, 0, 0, 6, 147, 218, 202, 185, 179, 175, 170, 167, 162, 152, 137, 132, 149, 175, 192, 209, 246, 288, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 181, 189, 170, 160, 148, 131, 112, 93, 90, 109, 136, 156, 171, 195, 232, 271, 307, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 87, 70, 59, 48, 40, 41, 57, 86, 120, 145, 160, 181, 213, 250, 287, 321, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 0, 0, 0, 14, 52, 87, 117, 140, 161, 180, 198, 222, 256, 297, 330, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 70, 106, 133, 151, 165, 181, 197, 212, 233, 265, 303, 336, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 47, 77, 108, 140, 158, 167, 178, 191, 207, 225, 248, 279, 312, 340, 
    52, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 24, 57, 79, 97, 114, 136, 155, 163, 172, 184, 197, 213, 235, 258, 285, 316, 341, 
    
    -- channel=20
    6, 4, 5, 5, 5, 5, 5, 5, 5, 6, 7, 7, 6, 6, 6, 6, 5, 3, 5, 8, 8, 7, 7, 5, 6, 6, 5, 4, 4, 6, 
    11, 8, 8, 8, 8, 8, 9, 10, 11, 11, 12, 12, 12, 11, 12, 14, 15, 20, 45, 64, 63, 47, 29, 14, 11, 12, 10, 10, 10, 11, 
    10, 7, 7, 7, 7, 7, 7, 8, 8, 7, 7, 8, 8, 8, 7, 5, 11, 31, 76, 90, 67, 36, 14, 8, 6, 7, 6, 5, 6, 7, 
    10, 8, 8, 8, 8, 8, 9, 9, 6, 5, 5, 7, 8, 10, 23, 46, 67, 81, 91, 58, 12, 6, 0, 5, 7, 5, 5, 4, 4, 5, 
    23, 19, 17, 13, 8, 6, 6, 6, 4, 4, 9, 18, 17, 17, 42, 85, 113, 111, 94, 66, 51, 72, 44, 17, 9, 8, 8, 7, 7, 7, 
    27, 16, 15, 13, 9, 6, 4, 3, 3, 5, 26, 46, 33, 23, 42, 42, 19, 6, 6, 7, 20, 39, 32, 15, 8, 7, 7, 6, 6, 7, 
    0, 0, 0, 0, 7, 10, 8, 7, 8, 7, 35, 45, 21, 10, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 5, 5, 5, 6, 
    179, 185, 158, 93, 35, 14, 14, 14, 14, 13, 26, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 121, 115, 77, 32, 9, 7, 
    207, 210, 190, 120, 50, 26, 24, 17, 14, 14, 13, 0, 0, 0, 2, 0, 0, 0, 4, 37, 91, 131, 158, 173, 190, 182, 122, 48, 11, 8, 
    0, 0, 0, 0, 0, 43, 53, 46, 37, 36, 39, 27, 12, 22, 21, 12, 2, 8, 35, 64, 76, 55, 22, 1, 10, 10, 0, 0, 5, 9, 
    0, 0, 0, 0, 0, 63, 93, 89, 82, 136, 216, 245, 234, 220, 200, 173, 128, 64, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 
    162, 158, 155, 129, 95, 65, 21, 0, 25, 146, 249, 281, 283, 281, 262, 205, 109, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 67, 48, 
    234, 238, 223, 176, 141, 90, 0, 0, 0, 66, 40, 0, 0, 0, 0, 0, 0, 0, 40, 96, 130, 164, 182, 182, 172, 151, 155, 172, 133, 89, 
    97, 36, 0, 9, 90, 117, 82, 60, 67, 18, 0, 0, 0, 0, 0, 0, 0, 100, 196, 230, 243, 239, 214, 182, 169, 156, 118, 65, 18, 21, 
    34, 0, 0, 0, 24, 22, 23, 46, 23, 0, 0, 0, 0, 0, 0, 87, 129, 130, 101, 60, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 53, 82, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 63, 76, 93, 118, 98, 25, 0, 1, 43, 54, 45, 48, 80, 113, 130, 143, 157, 154, 126, 88, 
    0, 0, 122, 132, 109, 121, 140, 158, 169, 177, 174, 159, 166, 203, 206, 176, 148, 154, 178, 173, 180, 194, 197, 180, 156, 133, 96, 61, 38, 19, 
    27, 169, 204, 188, 188, 195, 190, 177, 162, 149, 136, 116, 102, 89, 56, 47, 60, 76, 55, 39, 70, 95, 79, 44, 19, 20, 22, 17, 11, 1, 
    262, 288, 253, 239, 233, 229, 224, 216, 201, 184, 167, 152, 134, 108, 76, 66, 77, 96, 90, 81, 85, 81, 65, 50, 38, 32, 22, 6, 0, 0, 
    119, 120, 101, 104, 135, 164, 181, 195, 209, 223, 226, 222, 221, 221, 214, 198, 183, 174, 162, 141, 118, 92, 67, 38, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 31, 58, 81, 86, 57, 31, 48, 83, 102, 111, 103, 79, 49, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 8, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 14, 0, 0, 0, 
    33, 33, 36, 79, 112, 87, 56, 33, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 65, 69, 30, 0, 0, 0, 0, 
    0, 1, 12, 38, 83, 88, 68, 44, 18, 2, 0, 0, 47, 138, 122, 68, 47, 47, 67, 102, 135, 144, 108, 37, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 19, 33, 31, 18, 5, 0, 0, 0, 16, 95, 165, 168, 176, 196, 205, 177, 112, 26, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 9, 11, 4, 0, 0, 0, 0, 0, 24, 100, 142, 161, 142, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 122, 136, 82, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 4, 3, 0, 2, 0, 1, 1, 2, 3, 2, 2, 2, 2, 2, 1, 
    2, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 5, 6, 7, 6, 19, 19, 28, 15, 13, 6, 3, 4, 3, 4, 3, 3, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 2, 2, 4, 9, 21, 30, 32, 18, 10, 4, 1, 2, 2, 2, 2, 1, 
    2, 3, 2, 2, 2, 2, 2, 2, 2, 1, 1, 2, 2, 4, 9, 17, 21, 24, 13, 23, 19, 13, 6, 3, 2, 2, 1, 1, 1, 1, 
    8, 8, 6, 5, 3, 2, 1, 1, 1, 1, 3, 4, 5, 7, 13, 25, 35, 33, 20, 31, 43, 43, 28, 12, 3, 3, 2, 2, 2, 1, 
    10, 5, 5, 5, 4, 2, 0, 0, 1, 1, 12, 10, 17, 10, 0, 0, 0, 0, 0, 3, 21, 36, 31, 15, 2, 2, 2, 2, 1, 1, 
    0, 0, 0, 0, 3, 4, 3, 2, 2, 2, 8, 10, 21, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 
    79, 76, 62, 37, 21, 7, 7, 5, 5, 5, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 32, 48, 45, 28, 14, 3, 1, 
    90, 94, 88, 63, 38, 13, 11, 8, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 28, 45, 58, 68, 79, 79, 59, 31, 6, 1, 
    0, 0, 0, 0, 14, 21, 27, 22, 16, 15, 8, 9, 8, 8, 4, 1, 0, 0, 2, 6, 10, 8, 0, 0, 5, 13, 29, 15, 4, 2, 
    0, 0, 0, 0, 0, 30, 44, 43, 44, 62, 83, 105, 101, 94, 85, 73, 47, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 
    68, 69, 66, 51, 34, 17, 9, 12, 16, 42, 87, 127, 131, 130, 120, 93, 59, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 26, 19, 
    103, 111, 102, 89, 64, 28, 4, 0, 0, 0, 0, 9, 3, 0, 0, 0, 0, 2, 18, 36, 50, 62, 74, 79, 72, 68, 65, 71, 61, 46, 
    54, 34, 35, 48, 60, 75, 64, 35, 4, 0, 0, 0, 0, 0, 0, 0, 23, 56, 78, 89, 96, 95, 90, 88, 83, 70, 47, 35, 29, 29, 
    39, 0, 0, 0, 30, 57, 53, 31, 2, 0, 0, 0, 0, 0, 0, 38, 52, 47, 31, 14, 3, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 29, 36, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 10, 16, 25, 37, 23, 13, 0, 0, 6, 15, 19, 16, 16, 29, 43, 55, 62, 65, 59, 47, 38, 
    0, 9, 35, 38, 36, 41, 47, 52, 53, 53, 46, 51, 55, 62, 67, 57, 52, 47, 58, 69, 67, 65, 63, 64, 60, 50, 41, 34, 28, 21, 
    55, 70, 74, 70, 67, 65, 63, 57, 52, 44, 35, 27, 14, 11, 12, 20, 18, 9, 11, 21, 27, 30, 24, 19, 17, 20, 24, 26, 26, 20, 
    133, 130, 118, 109, 105, 102, 101, 97, 91, 83, 72, 57, 41, 31, 27, 31, 33, 33, 34, 36, 36, 35, 35, 31, 28, 29, 28, 27, 25, 21, 
    89, 91, 82, 78, 86, 97, 107, 116, 122, 126, 120, 110, 101, 96, 92, 83, 78, 71, 69, 64, 57, 50, 43, 30, 15, 6, 8, 16, 24, 21, 
    44, 53, 33, 17, 11, 27, 45, 65, 79, 88, 85, 61, 48, 43, 56, 63, 61, 55, 49, 39, 28, 14, 0, 0, 0, 0, 13, 24, 26, 15, 
    66, 74, 72, 55, 32, 25, 32, 46, 56, 63, 66, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 30, 36, 33, 27, 16, 10, 
    66, 76, 98, 104, 95, 78, 68, 64, 65, 65, 72, 84, 39, 0, 0, 0, 0, 0, 0, 0, 4, 30, 52, 64, 63, 48, 30, 18, 13, 11, 
    41, 60, 82, 96, 99, 91, 80, 72, 70, 67, 68, 109, 132, 123, 86, 64, 63, 67, 76, 88, 101, 100, 80, 54, 36, 28, 22, 18, 15, 12, 
    30, 50, 70, 77, 82, 79, 73, 70, 69, 68, 68, 87, 127, 155, 144, 132, 137, 137, 133, 117, 91, 63, 41, 29, 28, 31, 29, 23, 15, 11, 
    30, 48, 66, 70, 73, 72, 69, 68, 68, 68, 67, 75, 112, 146, 149, 144, 141, 120, 89, 58, 33, 24, 28, 32, 34, 32, 31, 28, 20, 13, 
    36, 52, 59, 63, 65, 65, 65, 65, 66, 66, 64, 71, 110, 151, 154, 129, 102, 70, 42, 24, 22, 29, 37, 37, 30, 25, 21, 21, 16, 12, 
    41, 48, 47, 50, 51, 52, 53, 54, 53, 52, 50, 50, 77, 103, 92, 60, 37, 31, 33, 35, 37, 40, 40, 38, 32, 25, 21, 16, 12, 9, 
    36, 38, 36, 35, 34, 32, 31, 30, 28, 26, 24, 22, 28, 36, 32, 23, 21, 33, 46, 51, 45, 40, 37, 34, 33, 28, 26, 23, 19, 14, 
    
    -- channel=22
    3, 4, 4, 4, 4, 4, 4, 4, 5, 5, 6, 6, 5, 5, 5, 6, 6, 3, 5, 4, 6, 3, 5, 5, 5, 4, 4, 4, 4, 4, 
    6, 7, 7, 7, 7, 7, 7, 8, 9, 9, 10, 10, 9, 9, 10, 12, 15, 17, 40, 43, 56, 34, 25, 12, 8, 9, 8, 8, 8, 8, 
    6, 6, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 7, 6, 4, 4, 11, 25, 59, 60, 57, 27, 12, 7, 5, 5, 5, 5, 5, 4, 
    5, 6, 6, 6, 6, 6, 6, 6, 5, 4, 4, 6, 6, 9, 18, 36, 52, 61, 47, 33, 17, 12, 7, 7, 5, 4, 4, 4, 4, 3, 
    18, 17, 14, 11, 7, 5, 4, 4, 4, 4, 8, 12, 12, 16, 35, 64, 78, 71, 40, 43, 63, 70, 48, 21, 5, 7, 7, 6, 6, 4, 
    21, 14, 11, 10, 8, 5, 3, 3, 4, 5, 26, 27, 28, 20, 16, 10, 0, 0, 0, 0, 25, 43, 33, 20, 4, 5, 5, 4, 4, 5, 
    0, 0, 0, 0, 3, 6, 7, 7, 8, 8, 28, 20, 25, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 2, 2, 4, 
    153, 150, 123, 75, 35, 11, 12, 14, 12, 12, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 65, 94, 89, 58, 27, 4, 3, 
    160, 164, 144, 89, 50, 20, 21, 18, 12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 69, 100, 122, 136, 149, 141, 93, 45, 7, 3, 
    0, 0, 0, 0, 0, 34, 46, 42, 34, 30, 17, 17, 17, 21, 12, 4, 0, 2, 23, 36, 34, 14, 0, 0, 0, 1, 10, 3, 4, 4, 
    0, 0, 0, 0, 0, 53, 78, 79, 78, 116, 166, 203, 195, 181, 164, 144, 99, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 
    129, 132, 131, 112, 76, 43, 14, 1, 29, 111, 177, 226, 229, 228, 212, 164, 86, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 55, 38, 
    190, 200, 184, 148, 99, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 77, 106, 132, 147, 148, 130, 133, 139, 137, 110, 81, 
    73, 29, 1, 37, 89, 104, 88, 67, 24, 0, 0, 0, 0, 0, 0, 0, 41, 123, 167, 186, 192, 182, 164, 152, 142, 120, 77, 45, 26, 33, 
    21, 0, 0, 0, 24, 51, 67, 48, 0, 0, 0, 0, 0, 0, 7, 82, 106, 93, 58, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 58, 72, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 34, 49, 55, 75, 56, 28, 0, 0, 2, 30, 37, 31, 35, 62, 85, 108, 124, 127, 112, 81, 54, 
    0, 30, 87, 83, 84, 99, 113, 124, 129, 129, 117, 116, 132, 142, 142, 116, 112, 118, 125, 129, 134, 136, 133, 124, 108, 81, 54, 34, 22, 16, 
    105, 153, 154, 148, 145, 142, 137, 128, 117, 103, 84, 73, 53, 35, 22, 29, 36, 26, 17, 31, 49, 52, 33, 16, 9, 10, 18, 22, 20, 5, 
    228, 226, 206, 194, 189, 186, 182, 173, 161, 148, 133, 117, 88, 65, 51, 57, 59, 56, 58, 63, 62, 53, 43, 37, 32, 27, 19, 10, 3, 1, 
    105, 110, 102, 100, 120, 143, 159, 173, 187, 197, 197, 191, 181, 177, 170, 154, 141, 130, 121, 106, 86, 68, 52, 28, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 14, 47, 74, 93, 95, 66, 48, 41, 67, 82, 85, 74, 56, 34, 9, 0, 0, 0, 0, 0, 0, 6, 1, 0, 
    37, 47, 37, 17, 0, 0, 0, 3, 17, 27, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 47, 28, 0, 0, 0, 
    34, 56, 86, 106, 105, 78, 55, 40, 31, 26, 38, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 75, 101, 81, 32, 0, 0, 0, 0, 
    0, 21, 57, 86, 102, 93, 70, 48, 34, 28, 32, 97, 149, 159, 126, 102, 95, 103, 121, 149, 174, 166, 112, 39, 0, 0, 0, 0, 0, 0, 
    0, 2, 30, 43, 55, 58, 49, 37, 30, 29, 27, 64, 133, 198, 229, 233, 243, 249, 238, 192, 119, 43, 0, 0, 0, 4, 1, 0, 0, 0, 
    0, 1, 22, 29, 36, 38, 34, 29, 27, 27, 27, 38, 83, 151, 210, 233, 234, 189, 109, 22, 0, 0, 0, 3, 11, 4, 1, 3, 1, 0, 
    1, 5, 7, 15, 18, 20, 20, 21, 21, 22, 21, 28, 73, 152, 204, 189, 120, 35, 0, 0, 0, 0, 10, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 64, 70, 17, 0, 0, 0, 0, 13, 19, 15, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 32, 32, 20, 5, 0, 3, 1, 1, 2, 4, 4, 
    
    -- channel=23
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 42, 42, 42, 43, 42, 42, 42, 43, 43, 40, 40, 42, 44, 44, 43, 43, 43, 43, 43, 43, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 43, 44, 43, 41, 41, 37, 41, 40, 43, 43, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 43, 42, 42, 43, 44, 44, 42, 38, 36, 35, 48, 46, 47, 43, 41, 42, 42, 42, 43, 42, 
    42, 42, 42, 42, 42, 42, 43, 42, 43, 43, 42, 41, 42, 43, 44, 43, 40, 36, 40, 48, 55, 51, 42, 41, 42, 43, 43, 42, 42, 42, 
    41, 41, 40, 41, 42, 43, 43, 42, 41, 41, 41, 40, 42, 43, 39, 35, 41, 45, 54, 55, 48, 47, 43, 44, 45, 44, 43, 42, 43, 42, 
    43, 41, 41, 43, 45, 45, 44, 41, 39, 39, 40, 39, 45, 46, 43, 44, 52, 56, 55, 51, 47, 50, 54, 52, 46, 45, 45, 45, 44, 43, 
    47, 42, 43, 46, 48, 47, 43, 40, 38, 38, 40, 41, 53, 49, 51, 57, 58, 57, 55, 57, 57, 55, 52, 53, 49, 47, 47, 47, 47, 45, 
    40, 41, 44, 48, 52, 49, 43, 38, 39, 40, 47, 50, 52, 52, 53, 49, 51, 51, 49, 52, 55, 53, 43, 42, 46, 46, 48, 51, 50, 46, 
    50, 51, 57, 65, 66, 50, 43, 39, 40, 43, 52, 55, 47, 47, 49, 47, 41, 41, 42, 39, 38, 40, 43, 44, 45, 49, 57, 62, 53, 48, 
    71, 69, 64, 63, 59, 48, 44, 41, 41, 46, 52, 51, 43, 43, 44, 45, 41, 40, 38, 35, 49, 60, 63, 62, 56, 54, 62, 62, 54, 49, 
    63, 61, 52, 35, 33, 46, 43, 41, 46, 46, 40, 42, 42, 43, 43, 42, 42, 46, 52, 60, 72, 73, 67, 61, 54, 56, 55, 44, 48, 49, 
    37, 34, 30, 25, 36, 47, 45, 53, 51, 35, 31, 50, 52, 51, 49, 50, 55, 63, 61, 61, 57, 53, 48, 47, 53, 50, 37, 33, 41, 47, 
    35, 32, 31, 42, 57, 63, 63, 52, 47, 54, 61, 71, 71, 71, 73, 74, 64, 47, 39, 38, 36, 37, 36, 41, 49, 41, 30, 37, 43, 49, 
    55, 56, 68, 69, 52, 57, 57, 43, 52, 75, 83, 79, 85, 89, 75, 50, 27, 18, 24, 28, 33, 41, 46, 49, 51, 53, 55, 56, 54, 58, 
    66, 83, 82, 58, 63, 65, 50, 48, 65, 80, 83, 73, 66, 49, 32, 31, 35, 39, 45, 52, 59, 65, 71, 70, 68, 70, 72, 68, 58, 52, 
    72, 89, 66, 63, 84, 69, 54, 53, 57, 57, 59, 53, 48, 44, 51, 63, 65, 67, 66, 66, 66, 65, 63, 63, 63, 60, 55, 51, 42, 42, 
    76, 50, 42, 67, 65, 50, 39, 31, 26, 30, 38, 42, 47, 53, 64, 57, 52, 51, 42, 42, 45, 41, 39, 40, 40, 37, 40, 48, 53, 58, 
    44, 3, 20, 32, 26, 18, 12, 9, 9, 15, 25, 27, 24, 27, 34, 35, 31, 21, 25, 32, 32, 31, 34, 36, 43, 55, 62, 63, 61, 56, 
    9, 7, 18, 14, 11, 11, 10, 8, 9, 11, 18, 17, 18, 26, 31, 31, 30, 34, 38, 33, 32, 41, 47, 48, 51, 58, 58, 55, 54, 58, 
    35, 39, 33, 29, 23, 18, 19, 22, 24, 23, 20, 14, 15, 18, 22, 23, 25, 31, 29, 25, 31, 40, 43, 41, 43, 51, 55, 58, 62, 63, 
    72, 68, 62, 55, 47, 42, 45, 47, 47, 44, 36, 26, 16, 12, 16, 23, 27, 25, 26, 31, 39, 44, 45, 46, 52, 62, 66, 62, 61, 66, 
    98, 97, 96, 89, 78, 74, 77, 79, 78, 76, 67, 53, 44, 40, 42, 44, 44, 42, 45, 50, 55, 57, 58, 62, 61, 56, 53, 57, 68, 76, 
    108, 102, 105, 108, 93, 85, 89, 95, 97, 98, 92, 81, 77, 66, 66, 65, 64, 64, 63, 65, 66, 64, 61, 52, 38, 36, 53, 71, 77, 79, 
    110, 107, 100, 96, 89, 86, 92, 98, 104, 106, 100, 88, 89, 74, 50, 49, 52, 50, 44, 42, 40, 32, 25, 28, 46, 69, 78, 75, 79, 79, 
    110, 111, 104, 91, 86, 85, 93, 104, 109, 109, 106, 82, 57, 44, 2, 0, 0, 0, 0, 0, 1, 14, 42, 72, 85, 82, 79, 81, 81, 75, 
    115, 109, 111, 104, 94, 91, 96, 105, 110, 109, 110, 96, 55, 8, 0, 0, 0, 0, 0, 5, 40, 67, 83, 87, 82, 82, 87, 87, 80, 74, 
    121, 111, 112, 109, 104, 101, 103, 109, 111, 110, 110, 107, 75, 13, 0, 0, 0, 0, 20, 59, 84, 90, 85, 83, 88, 93, 90, 84, 80, 76, 
    123, 121, 117, 116, 114, 114, 114, 114, 113, 113, 112, 110, 86, 32, 0, 0, 12, 58, 85, 90, 90, 90, 89, 94, 98, 96, 90, 84, 80, 76, 
    132, 138, 129, 126, 126, 126, 124, 122, 119, 118, 118, 119, 107, 73, 52, 61, 86, 98, 95, 87, 87, 95, 102, 103, 100, 95, 91, 86, 80, 74, 
    146, 149, 142, 136, 136, 136, 135, 131, 128, 128, 130, 135, 134, 121, 108, 99, 97, 98, 94, 90, 91, 102, 109, 105, 98, 95, 92, 85, 79, 74, 
    
    -- channel=24
    5, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 5, 3, 0, 0, 0, 2, 1, 0, 0, 2, 
    5, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 14, 0, 0, 0, 0, 1, 1, 1, 0, 0, 1, 
    4, 0, 1, 1, 1, 1, 2, 2, 0, 1, 1, 1, 0, 0, 0, 0, 8, 21, 60, 30, 0, 0, 0, 0, 2, 1, 1, 0, 0, 1, 
    4, 0, 0, 0, 0, 1, 2, 2, 0, 0, 2, 3, 1, 1, 9, 14, 24, 43, 78, 48, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 6, 10, 0, 6, 39, 53, 49, 60, 80, 62, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 20, 18, 0, 9, 61, 83, 75, 79, 95, 87, 49, 0, 0, 0, 3, 2, 1, 0, 0, 0, 
    10, 16, 17, 5, 0, 0, 0, 0, 0, 0, 38, 27, 0, 3, 56, 73, 63, 74, 93, 93, 78, 39, 0, 0, 10, 8, 7, 4, 1, 1, 
    10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 39, 31, 0, 0, 35, 46, 31, 47, 65, 65, 68, 57, 32, 12, 14, 1, 0, 0, 0, 2, 
    52, 36, 0, 0, 0, 0, 0, 0, 0, 2, 24, 26, 0, 0, 14, 26, 18, 27, 52, 61, 67, 64, 58, 49, 40, 7, 0, 0, 0, 2, 
    99, 82, 48, 0, 0, 3, 0, 0, 0, 5, 14, 15, 0, 4, 8, 14, 18, 29, 69, 90, 84, 85, 81, 87, 97, 41, 0, 0, 0, 3, 
    77, 58, 49, 15, 6, 30, 5, 0, 0, 47, 40, 5, 0, 0, 0, 0, 0, 1, 58, 89, 75, 77, 73, 83, 114, 56, 0, 0, 0, 2, 
    48, 22, 13, 8, 12, 44, 30, 0, 41, 154, 133, 52, 41, 29, 7, 0, 0, 0, 26, 54, 45, 51, 51, 44, 68, 48, 13, 13, 0, 0, 
    73, 53, 15, 0, 4, 10, 8, 6, 81, 218, 211, 113, 89, 64, 43, 12, 0, 0, 18, 36, 33, 38, 38, 13, 11, 26, 34, 29, 0, 0, 
    89, 75, 33, 37, 29, 0, 0, 0, 67, 166, 180, 115, 78, 57, 55, 33, 8, 11, 37, 55, 55, 50, 50, 33, 18, 27, 50, 49, 0, 0, 
    30, 0, 49, 105, 61, 0, 0, 0, 21, 71, 89, 65, 40, 57, 83, 64, 49, 58, 72, 93, 101, 87, 81, 76, 61, 48, 58, 68, 43, 29, 
    0, 0, 49, 130, 73, 0, 0, 0, 2, 21, 36, 27, 14, 67, 114, 107, 83, 81, 91, 99, 109, 102, 97, 91, 78, 65, 60, 66, 68, 54, 
    0, 0, 33, 91, 49, 19, 9, 15, 16, 23, 40, 30, 24, 62, 87, 88, 73, 83, 87, 66, 76, 94, 100, 90, 76, 76, 71, 67, 73, 68, 
    0, 1, 64, 71, 58, 58, 55, 60, 61, 60, 70, 71, 79, 99, 88, 76, 83, 116, 119, 84, 92, 116, 127, 118, 97, 96, 90, 77, 71, 67, 
    22, 77, 94, 94, 98, 106, 105, 107, 108, 104, 108, 119, 136, 150, 133, 116, 114, 148, 152, 128, 129, 141, 141, 136, 118, 107, 93, 73, 61, 56, 
    68, 88, 92, 101, 111, 117, 113, 106, 104, 104, 108, 120, 136, 143, 134, 131, 131, 146, 150, 142, 142, 139, 133, 130, 120, 108, 90, 65, 50, 42, 
    109, 78, 86, 113, 125, 121, 110, 99, 89, 87, 90, 106, 128, 134, 125, 123, 135, 146, 147, 144, 139, 131, 123, 114, 101, 92, 85, 61, 34, 21, 
    115, 64, 49, 93, 133, 133, 119, 106, 93, 87, 82, 86, 133, 172, 158, 142, 148, 155, 149, 141, 130, 119, 104, 88, 79, 75, 68, 40, 14, 0, 
    89, 57, 4, 24, 88, 111, 110, 103, 89, 80, 69, 15, 54, 170, 194, 171, 161, 157, 142, 121, 100, 87, 77, 63, 49, 40, 35, 17, 0, 0, 
    80, 64, 16, 0, 31, 65, 83, 88, 78, 68, 63, 0, 0, 26, 108, 101, 90, 84, 75, 58, 40, 32, 33, 29, 14, 7, 13, 0, 0, 0, 
    104, 73, 46, 15, 18, 42, 63, 72, 67, 59, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    135, 92, 56, 44, 34, 43, 57, 61, 59, 55, 56, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    151, 111, 58, 53, 49, 52, 58, 58, 57, 55, 55, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 
    142, 110, 60, 56, 57, 59, 60, 58, 57, 56, 57, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 1, 
    118, 86, 56, 53, 57, 60, 58, 56, 55, 56, 58, 56, 13, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 6, 
    90, 52, 42, 43, 47, 50, 50, 49, 47, 49, 50, 45, 25, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=25
    22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 23, 23, 22, 22, 22, 23, 24, 24, 23, 20, 20, 21, 23, 23, 22, 22, 22, 22, 22, 22, 
    24, 25, 25, 25, 25, 25, 25, 25, 25, 26, 26, 26, 26, 25, 26, 27, 27, 26, 32, 31, 37, 31, 31, 27, 26, 25, 25, 25, 25, 25, 
    23, 24, 23, 23, 23, 23, 24, 24, 24, 24, 24, 24, 24, 24, 25, 26, 26, 28, 41, 51, 55, 41, 32, 25, 23, 24, 24, 24, 24, 23, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 23, 23, 23, 23, 24, 27, 30, 33, 36, 42, 47, 41, 29, 21, 22, 23, 24, 24, 23, 23, 23, 
    26, 26, 25, 25, 25, 24, 24, 24, 23, 22, 23, 24, 25, 27, 34, 48, 58, 58, 50, 46, 46, 45, 36, 28, 24, 25, 25, 23, 23, 22, 
    30, 26, 24, 25, 25, 25, 23, 21, 21, 21, 29, 31, 37, 33, 35, 42, 46, 44, 39, 45, 57, 63, 51, 35, 24, 24, 24, 24, 24, 23, 
    19, 16, 18, 21, 24, 25, 24, 21, 21, 21, 32, 38, 44, 33, 31, 22, 12, 8, 3, 2, 2, 10, 19, 23, 24, 23, 23, 23, 23, 23, 
    59, 60, 55, 45, 36, 28, 26, 25, 24, 25, 27, 30, 32, 26, 20, 12, 8, 1, 0, 0, 0, 0, 11, 34, 49, 49, 42, 34, 26, 24, 
    128, 129, 118, 89, 57, 32, 29, 27, 27, 28, 24, 19, 17, 22, 19, 12, 9, 11, 15, 20, 38, 58, 76, 88, 98, 97, 80, 53, 30, 25, 
    23, 27, 31, 36, 36, 38, 40, 36, 33, 35, 30, 25, 22, 25, 25, 22, 19, 20, 31, 47, 65, 70, 62, 56, 57, 61, 61, 42, 30, 26, 
    0, 0, 0, 0, 10, 45, 54, 54, 55, 63, 74, 85, 81, 76, 70, 63, 50, 40, 30, 24, 13, 0, 0, 0, 0, 0, 7, 14, 27, 26, 
    54, 50, 45, 40, 42, 46, 47, 46, 47, 76, 120, 151, 150, 147, 138, 121, 92, 58, 25, 8, 0, 0, 3, 2, 0, 0, 6, 28, 40, 35, 
    117, 120, 115, 105, 82, 53, 27, 8, 15, 38, 60, 75, 75, 69, 55, 36, 23, 18, 28, 38, 46, 58, 67, 73, 66, 60, 66, 78, 73, 59, 
    90, 83, 76, 71, 76, 85, 70, 48, 43, 24, 0, 0, 0, 0, 0, 0, 2, 42, 74, 93, 107, 114, 115, 115, 114, 106, 91, 79, 66, 58, 
    73, 40, 19, 31, 73, 85, 81, 72, 54, 18, 0, 0, 0, 0, 14, 59, 81, 85, 80, 74, 67, 60, 49, 41, 37, 29, 16, 8, 14, 31, 
    67, 23, 0, 0, 10, 4, 7, 9, 4, 0, 0, 0, 8, 16, 29, 35, 24, 13, 0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 36, 56, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 11, 28, 38, 45, 35, 22, 3, 0, 5, 9, 13, 10, 10, 22, 37, 50, 65, 82, 88, 83, 74, 
    0, 2, 40, 40, 31, 30, 36, 41, 45, 51, 54, 55, 63, 77, 84, 74, 67, 71, 88, 94, 90, 89, 96, 101, 101, 95, 84, 69, 56, 49, 
    29, 64, 77, 77, 76, 75, 71, 68, 66, 64, 60, 53, 48, 51, 51, 49, 47, 45, 43, 47, 58, 65, 60, 53, 46, 45, 46, 47, 51, 51, 
    137, 137, 122, 111, 103, 98, 97, 93, 87, 79, 70, 56, 39, 29, 27, 32, 38, 41, 40, 43, 52, 55, 52, 50, 50, 56, 59, 57, 54, 52, 
    135, 135, 126, 118, 120, 126, 133, 139, 142, 142, 135, 121, 105, 95, 93, 91, 87, 82, 82, 81, 77, 72, 66, 61, 56, 50, 45, 44, 50, 54, 
    85, 89, 75, 61, 60, 75, 91, 106, 117, 125, 123, 107, 95, 89, 95, 95, 90, 83, 78, 74, 69, 60, 45, 30, 22, 24, 35, 49, 57, 52, 
    102, 103, 95, 76, 56, 56, 68, 81, 90, 97, 94, 61, 26, 2, 12, 29, 37, 36, 32, 28, 23, 16, 11, 13, 27, 48, 62, 60, 51, 43, 
    113, 118, 122, 120, 112, 102, 99, 98, 100, 101, 102, 85, 35, 0, 0, 0, 0, 0, 0, 0, 0, 16, 41, 71, 88, 80, 61, 48, 44, 40, 
    88, 104, 112, 117, 119, 116, 113, 110, 106, 103, 103, 111, 100, 81, 49, 30, 26, 28, 39, 56, 77, 96, 102, 89, 67, 54, 53, 52, 47, 43, 
    78, 92, 104, 104, 102, 102, 103, 104, 104, 102, 103, 105, 92, 81, 69, 62, 70, 79, 91, 101, 102, 87, 65, 51, 51, 60, 63, 56, 48, 45, 
    81, 90, 102, 103, 101, 100, 102, 103, 103, 102, 103, 98, 70, 42, 26, 27, 51, 70, 78, 70, 56, 44, 46, 60, 71, 71, 66, 61, 54, 48, 
    91, 98, 101, 104, 104, 103, 103, 103, 103, 103, 103, 99, 80, 61, 55, 64, 78, 75, 59, 49, 48, 55, 65, 72, 71, 65, 60, 59, 54, 48, 
    103, 103, 98, 101, 102, 102, 101, 100, 99, 98, 98, 96, 90, 85, 81, 73, 61, 53, 50, 58, 69, 78, 81, 76, 70, 63, 58, 53, 48, 44, 
    102, 99, 92, 91, 93, 92, 89, 85, 83, 82, 82, 80, 80, 73, 62, 48, 49, 61, 69, 74, 79, 84, 82, 76, 72, 68, 63, 58, 53, 48, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 29, 23, 20, 20, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    66, 66, 52, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 21, 7, 0, 0, 0, 
    93, 95, 85, 57, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 36, 52, 59, 67, 68, 52, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 0, 0, 5, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 5, 15, 61, 97, 91, 83, 73, 59, 40, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    69, 69, 67, 51, 22, 0, 0, 0, 0, 14, 84, 142, 142, 139, 130, 104, 56, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    120, 119, 120, 94, 56, 28, 0, 0, 0, 0, 14, 36, 34, 13, 0, 0, 0, 0, 0, 6, 26, 43, 55, 63, 63, 55, 52, 62, 55, 30, 
    97, 65, 37, 31, 43, 62, 50, 22, 7, 0, 0, 0, 0, 0, 0, 0, 0, 25, 59, 77, 89, 96, 91, 81, 77, 70, 51, 33, 17, 10, 
    99, 34, 0, 0, 12, 27, 23, 15, 0, 0, 0, 0, 0, 0, 0, 17, 43, 45, 35, 22, 9, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 28, 38, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 21, 24, 9, 0, 9, 29, 44, 37, 31, 44, 61, 74, 77, 81, 78, 65, 50, 
    0, 0, 44, 54, 49, 48, 52, 59, 64, 67, 62, 61, 66, 79, 91, 87, 80, 74, 89, 102, 102, 100, 102, 102, 97, 84, 69, 54, 43, 34, 
    68, 99, 112, 110, 110, 110, 106, 100, 94, 87, 80, 72, 62, 56, 51, 52, 56, 56, 55, 61, 72, 79, 76, 70, 61, 55, 53, 48, 40, 28, 
    165, 181, 168, 161, 162, 161, 158, 152, 146, 138, 133, 125, 112, 96, 84, 81, 81, 85, 87, 89, 94, 91, 87, 85, 78, 68, 55, 43, 31, 21, 
    109, 129, 122, 110, 122, 140, 149, 154, 161, 167, 174, 177, 172, 166, 161, 153, 143, 136, 134, 128, 120, 109, 97, 83, 62, 36, 17, 15, 18, 14, 
    55, 69, 68, 40, 25, 43, 64, 83, 99, 112, 122, 124, 107, 98, 117, 129, 130, 124, 116, 103, 87, 69, 42, 12, 0, 0, 10, 18, 12, 0, 
    78, 79, 83, 72, 41, 34, 41, 55, 67, 76, 83, 78, 34, 0, 0, 0, 3, 8, 4, 0, 0, 0, 0, 0, 18, 32, 26, 13, 0, 0, 
    69, 84, 90, 99, 97, 84, 78, 75, 74, 74, 77, 80, 63, 0, 0, 0, 0, 0, 0, 0, 0, 3, 33, 48, 47, 32, 11, 0, 0, 0, 
    31, 66, 79, 83, 91, 89, 85, 82, 77, 73, 74, 79, 75, 65, 22, 0, 0, 2, 17, 38, 56, 66, 58, 31, 4, 0, 0, 0, 0, 0, 
    15, 49, 72, 71, 73, 75, 75, 75, 74, 72, 72, 67, 41, 25, 5, 0, 20, 41, 59, 62, 50, 23, 0, 0, 0, 0, 5, 0, 0, 0, 
    19, 45, 68, 70, 71, 72, 72, 72, 71, 71, 72, 63, 29, 0, 0, 0, 26, 41, 29, 2, 0, 0, 0, 0, 3, 5, 3, 2, 0, 0, 
    31, 48, 57, 64, 66, 67, 68, 68, 68, 69, 71, 65, 43, 26, 25, 22, 22, 6, 0, 0, 0, 0, 0, 5, 3, 0, 0, 0, 0, 0, 
    31, 40, 36, 43, 48, 51, 52, 53, 52, 52, 54, 50, 37, 25, 20, 3, 0, 0, 0, 0, 0, 6, 10, 6, 2, 0, 0, 0, 0, 0, 
    17, 17, 15, 18, 23, 24, 22, 19, 18, 16, 14, 10, 2, 0, 0, 0, 0, 0, 0, 0, 6, 12, 9, 3, 1, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 6, 7, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 2, 4, 3, 4, 7, 9, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 6, 7, 8, 8, 9, 10, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 7, 8, 10, 10, 10, 10, 9, 10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 4, 6, 7, 7, 6, 6, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    280, 280, 280, 280, 280, 280, 280, 280, 281, 282, 282, 282, 282, 282, 280, 279, 279, 279, 282, 282, 283, 282, 282, 281, 281, 280, 280, 281, 282, 281, 
    282, 282, 282, 282, 282, 282, 282, 282, 283, 283, 283, 283, 284, 284, 282, 281, 282, 283, 288, 289, 297, 289, 289, 285, 282, 283, 283, 283, 284, 283, 
    282, 282, 282, 282, 282, 282, 282, 281, 281, 281, 281, 281, 282, 282, 281, 279, 280, 281, 271, 275, 288, 285, 288, 283, 281, 281, 281, 282, 283, 282, 
    282, 283, 282, 282, 283, 283, 282, 281, 282, 282, 281, 281, 283, 284, 286, 288, 286, 279, 244, 253, 271, 282, 285, 284, 281, 282, 282, 283, 283, 283, 
    284, 284, 283, 283, 283, 283, 281, 281, 282, 282, 283, 282, 285, 286, 280, 277, 277, 269, 239, 252, 276, 295, 299, 292, 284, 283, 284, 285, 285, 284, 
    286, 283, 283, 286, 286, 284, 282, 282, 282, 283, 284, 277, 290, 285, 257, 237, 236, 233, 220, 222, 241, 273, 301, 300, 287, 285, 286, 287, 287, 286, 
    287, 284, 284, 287, 288, 286, 285, 284, 284, 285, 270, 263, 290, 276, 246, 227, 225, 220, 205, 197, 198, 229, 277, 297, 293, 289, 290, 290, 290, 288, 
    322, 322, 317, 309, 301, 289, 285, 285, 285, 288, 253, 252, 279, 273, 254, 242, 252, 248, 239, 238, 242, 258, 289, 306, 312, 310, 306, 302, 295, 290, 
    273, 280, 293, 313, 315, 291, 284, 284, 285, 288, 258, 260, 274, 281, 271, 267, 275, 275, 283, 289, 294, 293, 291, 287, 288, 295, 311, 315, 299, 292, 
    147, 156, 188, 262, 294, 285, 285, 287, 288, 291, 280, 283, 287, 291, 288, 288, 289, 288, 283, 266, 253, 238, 218, 205, 197, 213, 277, 305, 300, 293, 
    186, 186, 201, 251, 266, 272, 276, 285, 293, 296, 302, 319, 322, 322, 321, 319, 312, 303, 265, 231, 218, 206, 196, 185, 158, 180, 254, 286, 297, 297, 
    290, 293, 299, 297, 277, 248, 235, 260, 262, 226, 223, 258, 269, 275, 281, 284, 297, 305, 274, 258, 258, 255, 257, 248, 218, 237, 270, 288, 304, 306, 
    252, 260, 269, 282, 278, 248, 244, 259, 229, 136, 102, 120, 127, 133, 150, 185, 248, 284, 293, 298, 301, 296, 293, 295, 290, 290, 279, 284, 301, 312, 
    153, 148, 179, 217, 229, 258, 288, 288, 242, 141, 91, 82, 100, 133, 167, 212, 261, 282, 286, 277, 269, 254, 242, 245, 250, 245, 224, 225, 256, 287, 
    118, 135, 163, 149, 162, 214, 248, 257, 242, 197, 172, 168, 199, 229, 236, 248, 249, 234, 210, 184, 165, 156, 152, 151, 160, 171, 176, 186, 228, 260, 
    121, 205, 176, 118, 125, 156, 185, 215, 240, 250, 255, 263, 282, 254, 211, 194, 184, 180, 170, 157, 148, 150, 158, 165, 185, 209, 228, 235, 247, 249, 
    161, 255, 225, 199, 195, 213, 230, 257, 279, 294, 290, 298, 313, 283, 253, 227, 230, 242, 248, 255, 255, 250, 248, 251, 258, 259, 255, 244, 230, 222, 
    212, 259, 275, 280, 285, 291, 296, 301, 304, 305, 289, 293, 291, 282, 277, 267, 268, 249, 248, 268, 271, 256, 235, 226, 219, 207, 198, 194, 192, 191, 
    236, 249, 255, 259, 263, 265, 265, 259, 256, 254, 247, 241, 219, 205, 200, 210, 208, 180, 170, 184, 187, 177, 160, 153, 154, 159, 164, 171, 179, 181, 
    206, 209, 205, 204, 207, 209, 213, 214, 215, 217, 218, 215, 201, 190, 186, 190, 187, 174, 165, 161, 156, 150, 145, 145, 149, 153, 154, 160, 169, 178, 
    86, 98, 104, 105, 110, 117, 127, 138, 150, 160, 170, 181, 186, 186, 184, 181, 176, 162, 152, 144, 137, 132, 128, 126, 127, 129, 133, 145, 161, 173, 
    9, 30, 42, 32, 14, 14, 20, 31, 39, 50, 62, 74, 85, 88, 100, 112, 111, 100, 94, 91, 89, 90, 90, 97, 113, 125, 131, 142, 158, 173, 
    17, 35, 68, 70, 34, 7, 0, 0, 0, 0, 10, 32, 35, 8, 7, 22, 27, 30, 33, 38, 49, 67, 94, 121, 135, 133, 131, 143, 160, 187, 
    7, 18, 64, 87, 69, 38, 15, 0, 0, 0, 4, 80, 120, 85, 35, 22, 24, 31, 40, 57, 83, 109, 126, 130, 128, 129, 134, 149, 177, 210, 
    0, 0, 19, 37, 36, 21, 6, 0, 0, 0, 0, 75, 158, 170, 115, 84, 84, 87, 93, 102, 109, 108, 100, 96, 106, 126, 144, 170, 200, 227, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 82, 106, 63, 39, 50, 58, 62, 60, 55, 56, 74, 98, 120, 141, 163, 191, 215, 235, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 45, 4, 0, 0, 0, 4, 18, 38, 68, 103, 126, 138, 153, 175, 204, 226, 242, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 48, 11, 0, 0, 0, 26, 56, 87, 114, 131, 139, 146, 158, 176, 204, 227, 245, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 30, 1, 0, 3, 42, 77, 105, 124, 134, 142, 151, 160, 170, 186, 208, 230, 245, 
    30, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 21, 31, 56, 87, 111, 127, 129, 135, 146, 157, 169, 181, 198, 220, 239, 249, 
    
    -- channel=29
    282, 280, 280, 280, 280, 280, 280, 280, 280, 281, 282, 282, 281, 282, 282, 280, 277, 277, 281, 283, 284, 283, 280, 280, 280, 281, 280, 280, 281, 282, 
    282, 280, 280, 280, 280, 280, 280, 280, 280, 280, 280, 280, 280, 280, 280, 278, 276, 280, 288, 279, 275, 277, 274, 278, 280, 280, 279, 280, 280, 281, 
    283, 280, 281, 281, 281, 281, 281, 280, 279, 279, 280, 279, 279, 280, 278, 276, 278, 281, 271, 247, 232, 253, 265, 278, 281, 279, 279, 280, 280, 281, 
    282, 281, 281, 281, 281, 281, 281, 280, 279, 280, 281, 281, 280, 281, 285, 285, 279, 271, 243, 220, 217, 247, 268, 279, 282, 280, 281, 281, 282, 283, 
    281, 280, 280, 280, 280, 280, 281, 280, 281, 282, 285, 283, 279, 281, 281, 266, 245, 232, 220, 212, 217, 234, 254, 275, 282, 280, 281, 282, 283, 284, 
    271, 276, 278, 278, 279, 281, 281, 283, 284, 285, 289, 276, 265, 275, 265, 234, 211, 205, 199, 189, 182, 195, 224, 263, 283, 280, 280, 282, 283, 285, 
    276, 283, 283, 282, 281, 282, 283, 285, 287, 287, 279, 258, 244, 261, 258, 236, 223, 224, 219, 205, 197, 204, 235, 269, 286, 284, 283, 285, 285, 286, 
    273, 273, 267, 259, 270, 281, 282, 283, 285, 286, 271, 250, 242, 262, 263, 254, 253, 260, 263, 263, 271, 274, 280, 284, 281, 273, 267, 275, 284, 286, 
    147, 151, 163, 188, 240, 278, 276, 277, 281, 281, 270, 261, 259, 274, 277, 275, 277, 284, 293, 294, 283, 260, 235, 218, 206, 199, 206, 244, 280, 286, 
    117, 115, 134, 181, 239, 270, 266, 267, 273, 276, 276, 274, 276, 279, 281, 283, 286, 289, 282, 254, 213, 187, 169, 163, 158, 142, 168, 231, 277, 285, 
    227, 226, 236, 254, 264, 262, 244, 234, 255, 277, 261, 243, 248, 253, 258, 263, 260, 265, 262, 241, 221, 217, 218, 215, 200, 183, 206, 257, 279, 284, 
    245, 249, 258, 257, 249, 227, 204, 205, 234, 224, 155, 104, 114, 122, 130, 140, 174, 227, 266, 273, 271, 274, 273, 262, 250, 252, 262, 271, 268, 276, 
    140, 142, 136, 162, 198, 203, 212, 241, 251, 192, 96, 33, 27, 30, 59, 112, 185, 251, 286, 288, 280, 267, 252, 239, 237, 240, 234, 220, 218, 241, 
    50, 46, 72, 126, 153, 158, 194, 237, 237, 186, 124, 89, 100, 145, 201, 234, 251, 257, 243, 218, 191, 163, 141, 132, 133, 137, 140, 143, 164, 206, 
    0, 28, 110, 131, 100, 94, 134, 177, 198, 204, 201, 206, 226, 254, 251, 216, 185, 168, 149, 130, 113, 99, 97, 101, 109, 124, 148, 170, 198, 217, 
    0, 72, 173, 162, 115, 120, 153, 195, 228, 255, 266, 266, 271, 263, 227, 187, 166, 169, 180, 182, 181, 181, 186, 188, 195, 211, 224, 225, 215, 198, 
    16, 170, 251, 239, 227, 241, 258, 276, 287, 292, 283, 274, 278, 281, 263, 238, 236, 246, 249, 242, 250, 253, 244, 228, 212, 198, 180, 164, 154, 152, 
    131, 232, 257, 255, 262, 271, 275, 277, 276, 272, 260, 251, 241, 229, 208, 201, 202, 198, 177, 170, 182, 183, 159, 136, 120, 113, 112, 118, 128, 132, 
    174, 202, 197, 195, 201, 207, 210, 209, 206, 205, 203, 204, 193, 176, 157, 160, 165, 158, 142, 133, 133, 126, 110, 100, 100, 104, 106, 108, 112, 121, 
    71, 76, 88, 100, 110, 119, 123, 129, 134, 144, 154, 169, 177, 176, 166, 160, 159, 153, 140, 124, 110, 99, 92, 88, 89, 86, 84, 89, 101, 115, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 28, 53, 82, 95, 94, 91, 93, 88, 75, 64, 57, 52, 51, 49, 53, 66, 82, 90, 95, 103, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 12, 13, 8, 4, 6, 10, 23, 46, 77, 99, 98, 85, 84, 99, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 2, 14, 39, 79, 111, 112, 90, 76, 74, 85, 115, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 89, 108, 84, 74, 73, 76, 87, 100, 104, 95, 70, 48, 48, 65, 82, 105, 141, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 129, 127, 121, 116, 107, 91, 67, 35, 10, 9, 29, 53, 72, 93, 124, 161, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 57, 66, 63, 52, 26, 0, 0, 0, 0, 31, 56, 66, 79, 105, 139, 172, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 46, 11, 0, 0, 0, 0, 7, 36, 51, 60, 67, 84, 112, 145, 177, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 46, 55, 55, 61, 75, 92, 117, 148, 180, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 45, 50, 50, 58, 71, 86, 106, 129, 158, 188, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 24, 38, 47, 44, 47, 60, 75, 93, 113, 138, 165, 190, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    85, 85, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 85, 87, 90, 88, 84, 78, 76, 76, 81, 84, 86, 85, 84, 84, 84, 84, 84, 
    83, 82, 82, 82, 82, 82, 82, 82, 81, 81, 81, 81, 81, 82, 85, 87, 84, 76, 57, 46, 42, 58, 71, 80, 82, 81, 81, 81, 81, 82, 
    83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 82, 83, 86, 87, 79, 61, 30, 22, 23, 54, 71, 81, 84, 83, 83, 83, 83, 84, 
    84, 84, 84, 84, 83, 83, 83, 83, 84, 85, 84, 82, 81, 80, 73, 58, 39, 21, 15, 17, 35, 54, 74, 81, 84, 85, 84, 84, 84, 84, 
    78, 80, 81, 82, 84, 85, 85, 85, 86, 87, 82, 75, 73, 70, 51, 19, 0, 0, 0, 0, 0, 10, 42, 70, 83, 84, 83, 82, 82, 84, 
    67, 74, 76, 78, 82, 85, 87, 88, 88, 88, 73, 64, 61, 64, 51, 29, 14, 6, 3, 0, 0, 1, 26, 56, 78, 81, 80, 79, 81, 84, 
    59, 65, 67, 72, 78, 84, 87, 88, 87, 87, 71, 68, 61, 71, 70, 61, 55, 52, 52, 54, 63, 61, 58, 58, 65, 70, 71, 73, 77, 81, 
    0, 0, 0, 14, 54, 81, 86, 85, 83, 81, 83, 84, 81, 87, 85, 81, 72, 67, 68, 66, 64, 49, 23, 8, 0, 7, 25, 50, 70, 79, 
    0, 0, 0, 0, 31, 74, 83, 83, 80, 74, 87, 89, 90, 84, 84, 81, 72, 63, 41, 13, 0, 0, 0, 0, 0, 0, 0, 27, 63, 76, 
    54, 53, 54, 54, 56, 66, 71, 70, 65, 59, 61, 59, 61, 57, 61, 61, 57, 49, 22, 0, 0, 0, 2, 11, 9, 9, 19, 42, 61, 72, 
    88, 97, 100, 80, 69, 51, 43, 39, 32, 0, 0, 0, 0, 0, 0, 0, 0, 16, 36, 49, 63, 76, 90, 92, 91, 93, 70, 62, 55, 64, 
    0, 0, 0, 0, 10, 35, 55, 57, 32, 0, 0, 0, 0, 0, 0, 0, 0, 19, 56, 66, 68, 65, 58, 61, 75, 74, 48, 24, 21, 36, 
    0, 0, 0, 0, 0, 20, 57, 65, 47, 20, 0, 0, 0, 2, 36, 66, 67, 56, 37, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 6, 17, 53, 77, 99, 116, 128, 120, 87, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 55, 39, 23, 28, 25, 23, 41, 83, 111, 130, 120, 82, 34, 0, 0, 0, 0, 0, 3, 17, 29, 37, 43, 51, 62, 60, 37, 8, 
    16, 65, 89, 109, 121, 140, 130, 109, 96, 92, 83, 73, 56, 46, 45, 44, 50, 55, 66, 73, 82, 83, 75, 67, 56, 40, 19, 0, 0, 0, 
    66, 58, 63, 73, 102, 112, 99, 69, 44, 27, 14, 5, 0, 0, 0, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 24, 31, 36, 
    24, 17, 16, 29, 34, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 40, 43, 40, 43, 51, 64, 
    23, 13, 12, 30, 59, 62, 52, 41, 33, 25, 14, 26, 41, 60, 46, 21, 12, 12, 21, 37, 56, 70, 72, 65, 51, 43, 52, 64, 74, 82, 
    35, 13, 0, 4, 20, 34, 35, 35, 37, 38, 27, 29, 63, 119, 162, 164, 160, 157, 152, 145, 129, 97, 59, 42, 49, 68, 77, 81, 82, 77, 
    72, 43, 22, 27, 35, 40, 37, 37, 40, 45, 39, 11, 47, 116, 182, 206, 205, 193, 164, 125, 91, 73, 77, 95, 106, 99, 84, 76, 70, 63, 
    83, 60, 43, 49, 58, 58, 52, 47, 46, 48, 48, 43, 109, 221, 294, 302, 264, 214, 163, 133, 127, 138, 145, 134, 109, 86, 73, 64, 58, 53, 
    77, 66, 51, 51, 52, 53, 50, 49, 49, 50, 48, 63, 152, 292, 372, 355, 282, 221, 192, 185, 180, 164, 135, 104, 83, 74, 66, 56, 48, 44, 
    67, 66, 64, 57, 52, 50, 50, 51, 52, 51, 47, 56, 118, 219, 270, 257, 220, 199, 190, 179, 153, 122, 98, 87, 82, 78, 71, 58, 51, 44, 
    70, 80, 87, 78, 67, 62, 63, 66, 68, 67, 63, 65, 93, 149, 191, 200, 194, 185, 175, 149, 113, 86, 76, 78, 78, 73, 69, 62, 54, 47, 
    86, 105, 112, 105, 96, 92, 94, 99, 102, 102, 101, 105, 120, 153, 182, 185, 174, 162, 152, 129, 100, 79, 74, 75, 72, 67, 59, 52, 44, 40, 
    
    -- channel=32
    143, 134, 110, 119, 163, 182, 189, 194, 206, 218, 217, 224, 240, 248, 254, 248, 239, 249, 256, 261, 260, 254, 264, 267, 262, 253, 264, 267, 257, 258, 
    159, 150, 124, 134, 179, 200, 206, 209, 223, 234, 227, 230, 242, 252, 256, 255, 245, 250, 252, 254, 233, 234, 266, 274, 267, 258, 269, 271, 259, 262, 
    172, 162, 136, 145, 193, 213, 218, 218, 233, 246, 234, 233, 241, 248, 250, 255, 246, 247, 252, 239, 200, 217, 262, 274, 270, 260, 271, 275, 258, 266, 
    184, 171, 146, 153, 202, 223, 232, 230, 245, 255, 240, 235, 241, 240, 236, 240, 239, 237, 243, 198, 144, 197, 257, 273, 272, 261, 269, 271, 255, 266, 
    194, 177, 150, 154, 208, 230, 242, 239, 254, 259, 241, 238, 245, 235, 219, 220, 220, 227, 230, 171, 122, 175, 225, 248, 264, 261, 266, 265, 254, 267, 
    205, 188, 153, 160, 216, 239, 247, 249, 265, 262, 243, 241, 253, 239, 209, 205, 179, 174, 158, 87, 66, 108, 138, 167, 205, 239, 261, 264, 255, 264, 
    191, 179, 139, 149, 197, 219, 223, 239, 257, 251, 237, 236, 247, 226, 195, 181, 147, 130, 115, 79, 66, 87, 99, 108, 149, 188, 223, 236, 230, 239, 
    150, 142, 110, 120, 155, 164, 172, 192, 209, 206, 200, 201, 203, 187, 183, 157, 108, 71, 49, 38, 28, 40, 46, 51, 122, 160, 194, 196, 171, 187, 
    91, 93, 79, 86, 110, 111, 117, 136, 145, 151, 147, 149, 142, 136, 141, 113, 67, 46, 41, 33, 31, 47, 54, 67, 100, 134, 170, 177, 122, 134, 
    41, 53, 56, 57, 74, 70, 70, 74, 90, 105, 99, 97, 92, 94, 99, 81, 63, 57, 57, 50, 51, 66, 99, 143, 141, 145, 158, 160, 101, 78, 
    16, 36, 37, 38, 59, 56, 45, 51, 79, 85, 73, 61, 56, 60, 56, 47, 45, 49, 54, 59, 55, 84, 143, 177, 170, 152, 174, 167, 114, 50, 
    13, 37, 34, 40, 54, 36, 20, 32, 62, 69, 61, 56, 57, 59, 52, 50, 51, 56, 64, 77, 80, 125, 184, 206, 205, 155, 168, 165, 115, 39, 
    21, 41, 34, 35, 38, 23, 20, 46, 74, 86, 83, 74, 75, 75, 71, 68, 76, 81, 91, 100, 112, 157, 193, 206, 215, 167, 144, 140, 83, 29, 
    36, 46, 47, 47, 42, 44, 48, 63, 78, 92, 97, 91, 92, 92, 90, 88, 96, 103, 108, 109, 116, 155, 178, 190, 195, 177, 137, 118, 72, 39, 
    38, 47, 55, 55, 52, 52, 59, 74, 89, 101, 108, 112, 114, 115, 108, 107, 111, 120, 126, 121, 118, 146, 168, 179, 177, 175, 147, 110, 102, 99, 
    39, 52, 62, 53, 56, 65, 85, 96, 104, 112, 114, 114, 114, 116, 113, 109, 115, 129, 143, 125, 116, 137, 156, 164, 163, 163, 143, 110, 125, 133, 
    34, 37, 47, 50, 52, 71, 86, 93, 96, 96, 98, 101, 109, 117, 123, 118, 119, 127, 138, 122, 117, 141, 152, 156, 153, 153, 141, 132, 152, 152, 
    27, 28, 37, 50, 54, 71, 83, 88, 89, 90, 97, 104, 110, 115, 121, 122, 121, 129, 142, 135, 135, 149, 152, 151, 140, 134, 122, 114, 110, 105, 
    39, 23, 23, 38, 58, 70, 82, 88, 86, 93, 97, 102, 107, 110, 109, 108, 102, 105, 134, 141, 139, 143, 143, 134, 118, 107, 96, 83, 63, 54, 
    27, 24, 43, 63, 75, 82, 81, 76, 71, 84, 96, 108, 111, 106, 85, 69, 63, 76, 118, 135, 126, 120, 118, 107, 94, 80, 63, 47, 31, 28, 
    27, 49, 60, 63, 63, 68, 63, 51, 53, 68, 80, 102, 113, 101, 69, 49, 39, 58, 99, 107, 100, 95, 88, 74, 54, 42, 31, 17, 18, 15, 
    19, 49, 56, 57, 59, 58, 41, 30, 33, 42, 57, 90, 111, 92, 52, 34, 23, 43, 76, 83, 76, 65, 49, 34, 24, 21, 7, 4, 8, 0, 
    14, 49, 59, 61, 68, 58, 32, 22, 28, 26, 45, 73, 79, 59, 35, 33, 37, 48, 58, 52, 41, 30, 26, 17, 14, 3, 0, 0, 0, 0, 
    16, 45, 55, 55, 61, 42, 15, 11, 13, 10, 24, 46, 52, 48, 41, 37, 32, 29, 29, 27, 23, 16, 10, 0, 1, 0, 0, 0, 0, 0, 
    2, 20, 29, 27, 29, 16, 2, 8, 18, 25, 32, 33, 25, 18, 16, 15, 11, 11, 16, 19, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 4, 6, 3, 0, 4, 11, 11, 8, 5, 1, 2, 7, 11, 8, 4, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 2, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 15, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    375, 338, 332, 378, 417, 423, 423, 433, 439, 430, 425, 433, 440, 445, 441, 428, 431, 446, 453, 441, 430, 438, 448, 447, 439, 446, 452, 441, 440, 451, 
    376, 340, 333, 375, 415, 421, 418, 428, 435, 426, 417, 423, 432, 439, 441, 429, 430, 439, 428, 394, 391, 422, 445, 447, 439, 446, 454, 440, 436, 450, 
    373, 337, 327, 367, 406, 417, 409, 415, 427, 418, 404, 411, 418, 423, 433, 425, 424, 429, 394, 347, 360, 410, 440, 444, 435, 440, 448, 435, 433, 446, 
    371, 330, 318, 359, 397, 407, 399, 407, 420, 409, 396, 401, 402, 396, 405, 404, 409, 416, 367, 307, 326, 393, 435, 441, 428, 427, 434, 428, 429, 438, 
    365, 320, 304, 345, 384, 398, 394, 399, 407, 399, 389, 394, 389, 360, 356, 366, 382, 390, 331, 275, 304, 360, 399, 420, 412, 408, 415, 411, 419, 428, 
    356, 308, 291, 335, 372, 384, 384, 388, 392, 386, 381, 386, 377, 349, 335, 325, 309, 299, 261, 203, 200, 238, 275, 328, 367, 384, 394, 388, 391, 405, 
    326, 287, 271, 308, 331, 337, 349, 358, 361, 358, 360, 362, 360, 352, 321, 274, 230, 208, 204, 175, 156, 157, 160, 220, 297, 334, 343, 328, 328, 350, 
    262, 241, 218, 234, 249, 258, 278, 287, 293, 295, 302, 304, 304, 309, 295, 255, 221, 204, 185, 173, 169, 149, 131, 158, 219, 273, 275, 244, 241, 259, 
    184, 175, 158, 168, 186, 186, 193, 207, 216, 217, 224, 233, 244, 256, 255, 230, 208, 198, 185, 174, 170, 175, 190, 186, 192, 236, 239, 195, 177, 184, 
    138, 141, 150, 172, 169, 150, 146, 168, 184, 179, 186, 208, 226, 231, 227, 212, 199, 192, 187, 173, 185, 225, 237, 230, 215, 244, 261, 199, 155, 153, 
    148, 155, 161, 181, 175, 149, 156, 196, 215, 207, 206, 223, 233, 227, 217, 200, 188, 190, 194, 188, 214, 274, 304, 293, 231, 220, 271, 224, 152, 147, 
    170, 164, 156, 170, 168, 160, 173, 203, 234, 239, 225, 231, 243, 236, 219, 207, 203, 208, 216, 222, 247, 291, 328, 335, 282, 216, 238, 222, 139, 127, 
    173, 173, 157, 149, 153, 158, 174, 212, 250, 268, 266, 265, 272, 268, 258, 257, 255, 257, 259, 263, 275, 294, 309, 316, 303, 230, 189, 177, 111, 94, 
    195, 196, 185, 186, 195, 208, 236, 263, 281, 299, 311, 313, 314, 312, 308, 309, 308, 301, 278, 258, 258, 274, 287, 288, 287, 240, 155, 133, 119, 94, 
    225, 231, 234, 247, 264, 274, 288, 307, 323, 332, 338, 344, 347, 339, 321, 313, 314, 298, 256, 220, 226, 251, 271, 278, 279, 255, 192, 174, 184, 153, 
    247, 258, 254, 244, 266, 302, 324, 336, 344, 347, 344, 339, 331, 320, 300, 285, 291, 289, 256, 222, 228, 246, 260, 273, 273, 267, 252, 243, 237, 208, 
    240, 223, 215, 223, 257, 301, 327, 333, 329, 321, 313, 307, 302, 299, 295, 286, 286, 293, 280, 255, 252, 263, 269, 272, 273, 270, 253, 230, 235, 245, 
    195, 199, 227, 255, 268, 284, 303, 302, 296, 297, 301, 305, 306, 304, 301, 288, 278, 292, 297, 283, 279, 286, 284, 274, 264, 242, 211, 184, 176, 200, 
    216, 230, 251, 266, 277, 280, 277, 281, 293, 303, 306, 306, 303, 291, 273, 254, 251, 275, 293, 291, 286, 288, 274, 245, 217, 192, 165, 138, 127, 145, 
    246, 244, 258, 275, 289, 291, 277, 276, 284, 290, 295, 297, 282, 242, 202, 180, 199, 252, 283, 281, 268, 249, 223, 195, 175, 154, 126, 113, 104, 78, 
    261, 273, 276, 279, 276, 266, 249, 234, 235, 250, 275, 289, 260, 202, 163, 150, 167, 218, 244, 233, 216, 197, 181, 161, 135, 110, 98, 93, 71, 41, 
    249, 267, 269, 268, 248, 213, 192, 183, 182, 208, 254, 278, 262, 215, 172, 154, 149, 165, 186, 186, 176, 162, 136, 111, 98, 86, 75, 59, 43, 28, 
    216, 247, 255, 257, 233, 189, 169, 170, 178, 196, 226, 239, 225, 192, 160, 147, 146, 154, 160, 150, 131, 113, 103, 98, 84, 67, 51, 39, 28, 13, 
    201, 233, 241, 242, 228, 194, 170, 167, 167, 164, 163, 166, 162, 156, 151, 147, 142, 136, 124, 107, 96, 95, 96, 87, 64, 47, 39, 30, 20, 12, 
    171, 190, 190, 184, 177, 160, 139, 133, 128, 127, 131, 134, 132, 129, 123, 114, 105, 99, 98, 94, 85, 71, 67, 68, 54, 37, 30, 27, 22, 21, 
    104, 112, 114, 110, 107, 103, 103, 106, 107, 102, 98, 95, 95, 95, 91, 85, 88, 98, 92, 75, 61, 54, 49, 46, 40, 30, 25, 25, 27, 22, 
    50, 51, 54, 57, 59, 61, 67, 71, 73, 71, 69, 70, 74, 78, 74, 73, 92, 100, 77, 57, 50, 46, 36, 31, 28, 25, 26, 29, 27, 11, 
    24, 19, 20, 27, 34, 36, 40, 47, 53, 57, 61, 66, 68, 67, 60, 56, 82, 99, 73, 47, 40, 32, 25, 24, 23, 24, 27, 30, 16, 0, 
    15, 13, 15, 22, 28, 33, 37, 44, 52, 56, 56, 57, 58, 55, 44, 37, 63, 87, 66, 38, 27, 24, 21, 19, 20, 22, 28, 25, 0, 0, 
    19, 20, 24, 29, 34, 37, 41, 45, 47, 49, 48, 44, 37, 26, 10, 2, 33, 67, 53, 26, 20, 19, 16, 14, 15, 20, 26, 7, 0, 0, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 6, 30, 39, 21, 3, 4, 4, 0, 0, 10, 0, 0, 
    9, 19, 0, 0, 0, 0, 0, 0, 0, 12, 14, 8, 19, 16, 17, 13, 0, 8, 50, 117, 106, 41, 7, 12, 11, 0, 5, 19, 6, 4, 
    5, 20, 0, 0, 0, 6, 8, 0, 2, 17, 16, 10, 25, 27, 26, 21, 6, 17, 71, 117, 74, 16, 10, 16, 18, 5, 18, 29, 6, 3, 
    5, 22, 0, 0, 0, 7, 12, 0, 5, 21, 18, 8, 28, 50, 62, 66, 32, 34, 100, 118, 17, 0, 9, 23, 30, 20, 32, 36, 10, 10, 
    21, 42, 13, 0, 2, 11, 10, 0, 6, 30, 19, 3, 29, 67, 82, 95, 64, 67, 111, 93, 31, 47, 78, 63, 51, 34, 41, 41, 20, 27, 
    24, 47, 9, 0, 0, 15, 20, 2, 18, 36, 18, 8, 28, 31, 15, 63, 131, 211, 253, 170, 127, 233, 291, 236, 140, 51, 38, 56, 46, 48, 
    74, 75, 27, 4, 62, 83, 79, 56, 67, 64, 38, 39, 54, 36, 13, 68, 140, 172, 174, 114, 62, 118, 179, 195, 185, 129, 110, 132, 114, 106, 
    172, 150, 107, 117, 190, 191, 175, 168, 172, 156, 131, 135, 133, 112, 107, 120, 80, 21, 0, 0, 0, 0, 0, 0, 0, 94, 151, 198, 180, 181, 
    172, 156, 127, 113, 144, 147, 151, 175, 180, 176, 172, 174, 155, 133, 141, 126, 55, 12, 10, 23, 18, 0, 0, 0, 0, 0, 22, 74, 99, 130, 
    64, 50, 14, 0, 0, 27, 55, 50, 40, 54, 59, 45, 31, 40, 66, 55, 19, 5, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 37, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 4, 29, 21, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 49, 20, 23, 
    0, 0, 0, 26, 68, 36, 0, 0, 0, 0, 0, 0, 4, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 7, 102, 64, 41, 
    0, 15, 12, 12, 39, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 51, 57, 41, 58, 162, 124, 35, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 44, 48, 39, 41, 55, 73, 100, 74, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 37, 44, 76, 97, 81, 58, 42, 32, 27, 30, 0, 0, 0, 0, 
    0, 0, 0, 15, 22, 7, 0, 0, 0, 3, 16, 32, 51, 64, 67, 55, 41, 28, 24, 0, 0, 0, 0, 18, 28, 23, 0, 0, 0, 0, 
    30, 64, 90, 70, 28, 13, 8, 9, 31, 56, 68, 66, 56, 39, 15, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 18, 17, 27, 80, 80, 
    64, 58, 0, 0, 0, 0, 22, 59, 67, 54, 28, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 2, 7, 30, 58, 92, 122, 141, 103, 
    0, 0, 0, 0, 0, 0, 24, 36, 5, 0, 0, 0, 0, 11, 53, 95, 88, 40, 19, 10, 4, 19, 46, 77, 105, 122, 131, 123, 97, 84, 
    0, 0, 0, 0, 19, 18, 7, 0, 0, 0, 0, 13, 54, 123, 173, 181, 129, 53, 21, 28, 49, 83, 119, 130, 116, 108, 90, 56, 35, 64, 
    3, 0, 0, 0, 4, 32, 61, 68, 88, 100, 66, 32, 46, 79, 78, 43, 0, 0, 66, 104, 119, 124, 120, 105, 81, 71, 59, 40, 50, 79, 
    22, 13, 13, 14, 46, 101, 131, 119, 102, 78, 33, 9, 13, 2, 0, 0, 0, 8, 93, 115, 96, 87, 85, 79, 71, 60, 47, 50, 70, 67, 
    0, 21, 21, 14, 32, 49, 30, 0, 0, 0, 0, 59, 106, 94, 44, 19, 19, 26, 47, 56, 66, 71, 59, 37, 27, 30, 30, 33, 36, 18, 
    0, 0, 7, 14, 24, 3, 0, 0, 0, 22, 69, 127, 137, 106, 63, 34, 24, 28, 47, 62, 61, 51, 26, 4, 8, 28, 26, 16, 5, 0, 
    33, 72, 96, 112, 124, 109, 72, 69, 78, 81, 84, 72, 44, 19, 13, 32, 57, 67, 63, 50, 31, 17, 14, 30, 47, 33, 12, 6, 0, 0, 
    105, 143, 157, 144, 133, 114, 85, 58, 39, 21, 13, 19, 32, 45, 56, 60, 36, 5, 4, 14, 20, 26, 25, 33, 40, 18, 0, 0, 0, 0, 
    63, 74, 72, 56, 42, 30, 21, 21, 30, 40, 45, 44, 38, 34, 33, 18, 0, 0, 0, 27, 27, 19, 16, 18, 15, 0, 0, 0, 0, 11, 
    7, 6, 4, 7, 12, 13, 16, 24, 29, 23, 15, 5, 0, 0, 3, 0, 0, 1, 42, 32, 14, 13, 14, 10, 1, 0, 0, 0, 12, 43, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 32, 30, 8, 25, 47, 19, 8, 14, 11, 3, 0, 0, 0, 5, 40, 56, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 29, 44, 57, 70, 61, 28, 32, 42, 16, 9, 10, 1, 1, 2, 0, 0, 27, 55, 39, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 5, 6, 1, 0, 0, 1, 4, 23, 34, 38, 28, 5, 0, 0, 1, 0, 0, 3, 5, 
    0, 0, 3, 10, 0, 0, 0, 2, 2, 0, 6, 9, 13, 9, 6, 2, 3, 8, 16, 27, 44, 30, 8, 1, 1, 7, 5, 0, 7, 5, 
    0, 0, 8, 18, 5, 3, 3, 9, 8, 2, 9, 12, 16, 24, 27, 25, 15, 18, 17, 23, 42, 26, 9, 6, 8, 16, 15, 5, 10, 9, 
    0, 4, 17, 30, 15, 11, 7, 14, 13, 8, 12, 15, 17, 31, 43, 45, 39, 26, 11, 29, 61, 55, 41, 26, 20, 24, 25, 18, 18, 17, 
    3, 5, 19, 28, 20, 16, 16, 22, 20, 16, 16, 20, 11, 8, 25, 38, 77, 88, 67, 78, 107, 136, 144, 107, 65, 36, 30, 34, 35, 35, 
    26, 19, 37, 45, 50, 46, 48, 46, 39, 36, 31, 34, 23, 16, 18, 28, 56, 69, 59, 48, 51, 78, 112, 131, 107, 80, 64, 69, 72, 74, 
    74, 61, 80, 94, 101, 103, 102, 96, 88, 85, 77, 72, 62, 59, 41, 28, 17, 8, 1, 0, 0, 0, 3, 46, 58, 82, 88, 93, 112, 112, 
    89, 79, 81, 83, 85, 94, 101, 100, 101, 100, 98, 86, 75, 69, 51, 35, 24, 18, 17, 23, 22, 12, 12, 21, 32, 36, 43, 41, 83, 87, 
    53, 43, 30, 24, 22, 42, 54, 52, 48, 47, 48, 36, 27, 24, 20, 22, 20, 18, 13, 15, 2, 0, 0, 0, 35, 34, 21, 3, 27, 46, 
    13, 11, 14, 17, 10, 12, 13, 7, 0, 0, 0, 1, 2, 2, 9, 14, 15, 11, 3, 0, 0, 0, 0, 0, 0, 40, 35, 25, 14, 38, 
    6, 7, 29, 44, 32, 24, 24, 20, 4, 0, 0, 1, 1, 0, 0, 0, 4, 2, 0, 0, 5, 18, 18, 6, 0, 37, 40, 41, 31, 46, 
    13, 13, 24, 28, 26, 21, 15, 13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 21, 35, 39, 13, 37, 68, 64, 58, 52, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 44, 47, 46, 40, 26, 22, 51, 52, 49, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 17, 32, 50, 64, 58, 46, 34, 28, 3, 0, 0, 0, 0, 
    0, 0, 3, 17, 12, 1, 0, 0, 0, 0, 0, 1, 11, 16, 19, 22, 19, 11, 0, 8, 18, 25, 26, 28, 27, 7, 0, 0, 0, 0, 
    16, 29, 33, 29, 25, 9, 0, 0, 0, 8, 13, 14, 13, 10, 1, 2, 3, 0, 0, 0, 0, 4, 15, 18, 22, 18, 27, 51, 57, 34, 
    22, 16, 0, 0, 0, 0, 9, 15, 13, 10, 1, 0, 0, 0, 0, 0, 5, 11, 2, 2, 8, 9, 13, 15, 29, 40, 56, 74, 82, 71, 
    0, 0, 0, 0, 0, 0, 6, 2, 0, 0, 0, 0, 0, 9, 29, 42, 41, 35, 17, 12, 15, 20, 30, 43, 56, 64, 70, 67, 73, 90, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 28, 50, 71, 80, 71, 51, 27, 22, 34, 49, 55, 59, 62, 61, 55, 49, 57, 78, 
    3, 0, 0, 0, 2, 11, 20, 35, 46, 41, 29, 14, 12, 21, 32, 32, 41, 51, 49, 54, 60, 60, 58, 55, 55, 53, 51, 58, 60, 64, 
    23, 4, 0, 3, 20, 37, 52, 55, 51, 44, 31, 10, 0, 0, 0, 2, 28, 50, 60, 59, 54, 53, 53, 54, 56, 51, 55, 63, 64, 59, 
    22, 13, 7, 3, 2, 8, 17, 13, 1, 12, 27, 39, 39, 34, 31, 30, 36, 40, 42, 47, 50, 51, 45, 45, 42, 43, 49, 53, 53, 51, 
    14, 10, 7, 9, 0, 0, 0, 10, 22, 42, 60, 68, 63, 51, 43, 36, 35, 41, 47, 50, 50, 48, 40, 39, 37, 45, 48, 46, 44, 43, 
    44, 48, 51, 58, 53, 48, 48, 50, 56, 59, 58, 52, 40, 34, 38, 46, 53, 55, 53, 45, 42, 41, 49, 53, 48, 48, 48, 45, 42, 42, 
    80, 84, 84, 81, 75, 68, 58, 50, 43, 40, 41, 45, 49, 52, 55, 52, 41, 37, 33, 39, 45, 47, 54, 52, 49, 47, 44, 42, 41, 47, 
    65, 66, 66, 60, 55, 52, 51, 50, 51, 54, 56, 54, 51, 47, 47, 40, 28, 23, 27, 43, 48, 48, 48, 47, 46, 44, 43, 40, 47, 53, 
    48, 49, 51, 50, 50, 52, 55, 54, 51, 48, 44, 40, 37, 37, 41, 45, 45, 38, 35, 45, 50, 47, 48, 46, 44, 43, 42, 45, 56, 62, 
    51, 48, 46, 43, 41, 40, 39, 38, 35, 33, 34, 37, 41, 46, 54, 60, 58, 45, 37, 47, 48, 48, 48, 45, 46, 46, 44, 55, 60, 69, 
    43, 40, 39, 37, 37, 36, 37, 39, 42, 45, 51, 55, 61, 67, 75, 78, 71, 51, 42, 48, 49, 48, 47, 45, 47, 46, 52, 59, 63, 69, 
    
    -- channel=38
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 21, 18, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 17, 8, 6, 0, 3, 11, 50, 80, 74, 47, 11, 4, 0, 3, 3, 4, 6, 14, 
    0, 0, 0, 2, 0, 0, 0, 1, 4, 1, 11, 15, 26, 19, 18, 7, 7, 21, 55, 65, 56, 37, 16, 11, 7, 13, 17, 9, 11, 14, 
    0, 0, 0, 11, 1, 4, 3, 4, 10, 5, 13, 15, 32, 42, 52, 49, 28, 36, 51, 43, 44, 28, 16, 17, 16, 25, 30, 16, 16, 20, 
    0, 7, 8, 26, 13, 11, 1, 7, 16, 13, 15, 13, 29, 56, 76, 78, 58, 57, 52, 35, 62, 80, 74, 55, 37, 35, 39, 28, 28, 31, 
    3, 10, 7, 20, 16, 18, 17, 21, 27, 22, 18, 19, 20, 13, 27, 56, 129, 170, 144, 127, 167, 233, 249, 195, 118, 54, 43, 48, 50, 53, 
    50, 35, 33, 53, 82, 83, 81, 72, 68, 56, 45, 52, 36, 12, 25, 61, 120, 135, 93, 65, 71, 116, 163, 181, 157, 123, 108, 120, 113, 117, 
    133, 102, 113, 149, 180, 174, 168, 165, 154, 142, 129, 130, 111, 99, 83, 62, 23, 0, 0, 0, 0, 0, 0, 18, 54, 112, 139, 160, 175, 183, 
    141, 119, 118, 126, 125, 133, 152, 161, 162, 160, 162, 151, 129, 117, 92, 55, 17, 0, 3, 12, 10, 0, 0, 0, 15, 30, 48, 47, 113, 131, 
    57, 38, 6, 0, 0, 33, 57, 54, 50, 52, 57, 39, 27, 33, 29, 15, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 4, 0, 18, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 23, 1, 28, 
    0, 0, 10, 40, 36, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 20, 35, 66, 27, 39, 
    0, 0, 7, 22, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 41, 51, 9, 43, 84, 105, 78, 47, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 59, 57, 51, 27, 30, 72, 60, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 17, 26, 54, 72, 81, 64, 49, 39, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 20, 4, 0, 0, 0, 0, 0, 7, 23, 28, 34, 33, 23, 8, 0, 0, 0, 0, 13, 28, 27, 0, 0, 0, 0, 0, 
    13, 51, 66, 50, 25, 4, 0, 0, 10, 28, 36, 33, 23, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 17, 6, 12, 60, 81, 34, 
    43, 28, 0, 0, 0, 0, 13, 35, 36, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 6, 26, 50, 83, 112, 121, 89, 
    0, 0, 0, 0, 0, 0, 14, 4, 0, 0, 0, 0, 0, 5, 43, 69, 62, 43, 12, 3, 8, 18, 38, 62, 88, 100, 100, 90, 86, 101, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 43, 87, 127, 135, 95, 56, 23, 19, 43, 74, 94, 97, 83, 72, 60, 37, 41, 95, 
    0, 0, 0, 0, 0, 10, 30, 55, 77, 71, 44, 14, 20, 34, 33, 17, 12, 36, 64, 85, 97, 96, 81, 60, 55, 52, 39, 39, 56, 73, 
    15, 0, 0, 0, 31, 65, 87, 88, 81, 53, 25, 0, 0, 0, 0, 0, 0, 57, 87, 83, 66, 53, 56, 57, 56, 40, 38, 55, 59, 42, 
    11, 10, 1, 0, 4, 4, 0, 0, 0, 0, 9, 51, 59, 43, 28, 22, 28, 33, 33, 38, 47, 54, 40, 23, 17, 21, 32, 33, 27, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 89, 113, 99, 66, 36, 18, 15, 26, 42, 52, 47, 30, 6, 7, 15, 26, 25, 17, 11, 7, 
    44, 64, 77, 90, 79, 64, 59, 65, 70, 72, 64, 45, 23, 10, 15, 33, 53, 59, 51, 28, 15, 16, 26, 37, 34, 26, 17, 11, 7, 3, 
    108, 125, 125, 116, 101, 83, 63, 42, 23, 14, 14, 24, 37, 46, 52, 49, 25, 4, 0, 10, 25, 27, 34, 36, 28, 16, 10, 6, 1, 9, 
    64, 66, 60, 48, 36, 28, 25, 27, 34, 42, 46, 45, 38, 29, 24, 6, 0, 0, 0, 23, 26, 21, 23, 23, 16, 9, 6, 1, 9, 23, 
    18, 18, 21, 21, 21, 24, 31, 34, 32, 24, 14, 5, 0, 1, 8, 10, 12, 20, 18, 20, 20, 21, 23, 17, 10, 7, 5, 6, 28, 42, 
    19, 13, 11, 7, 4, 1, 0, 0, 0, 0, 0, 0, 10, 20, 32, 39, 40, 33, 13, 16, 22, 23, 19, 14, 12, 11, 8, 24, 41, 48, 
    2, 0, 0, 0, 0, 0, 0, 0, 5, 14, 24, 34, 44, 54, 65, 68, 59, 40, 17, 21, 21, 18, 15, 14, 15, 11, 17, 37, 43, 36, 
    
    -- channel=39
    42, 44, 41, 40, 36, 34, 32, 33, 32, 31, 33, 38, 38, 37, 42, 40, 39, 38, 38, 37, 39, 46, 44, 42, 40, 40, 39, 38, 38, 37, 
    45, 49, 45, 44, 40, 39, 37, 39, 38, 38, 38, 36, 37, 37, 43, 41, 41, 39, 38, 36, 41, 48, 42, 42, 39, 39, 40, 38, 35, 36, 
    49, 54, 49, 47, 43, 46, 44, 42, 45, 45, 42, 40, 40, 36, 44, 42, 40, 39, 36, 40, 53, 52, 39, 41, 40, 39, 40, 39, 37, 36, 
    52, 55, 51, 53, 48, 50, 48, 50, 54, 50, 47, 43, 43, 37, 44, 44, 42, 45, 49, 54, 55, 46, 39, 44, 44, 43, 44, 42, 39, 37, 
    54, 57, 51, 57, 52, 55, 55, 55, 57, 54, 51, 48, 51, 42, 43, 50, 49, 50, 49, 56, 64, 51, 42, 47, 49, 49, 53, 47, 41, 41, 
    53, 57, 51, 56, 51, 51, 51, 52, 55, 55, 53, 53, 55, 51, 53, 56, 49, 47, 60, 59, 48, 48, 50, 53, 55, 53, 57, 55, 49, 50, 
    48, 54, 50, 48, 40, 37, 42, 45, 50, 52, 50, 49, 57, 67, 59, 42, 38, 40, 64, 68, 54, 61, 61, 68, 73, 60, 54, 50, 49, 58, 
    47, 56, 48, 37, 36, 38, 43, 41, 46, 50, 46, 44, 48, 55, 54, 52, 62, 72, 73, 70, 76, 81, 72, 65, 57, 60, 56, 53, 53, 59, 
    56, 62, 57, 51, 59, 59, 53, 50, 52, 52, 49, 47, 47, 51, 58, 65, 68, 67, 64, 65, 66, 76, 90, 82, 58, 62, 65, 61, 61, 59, 
    69, 73, 78, 82, 76, 70, 67, 65, 64, 61, 62, 61, 55, 50, 56, 67, 69, 69, 73, 76, 78, 89, 77, 69, 78, 81, 89, 69, 65, 68, 
    78, 84, 84, 81, 70, 67, 72, 78, 70, 66, 70, 66, 53, 48, 57, 66, 69, 76, 82, 86, 87, 89, 75, 72, 72, 64, 88, 77, 62, 75, 
    75, 72, 69, 71, 68, 73, 75, 63, 59, 62, 55, 51, 49, 50, 57, 65, 74, 77, 79, 83, 80, 67, 61, 70, 74, 60, 65, 79, 65, 80, 
    60, 68, 71, 64, 66, 69, 56, 49, 54, 58, 55, 50, 52, 57, 61, 68, 72, 72, 76, 77, 71, 59, 53, 56, 70, 65, 51, 76, 72, 77, 
    58, 68, 69, 65, 62, 57, 58, 54, 49, 49, 53, 52, 49, 52, 55, 59, 59, 62, 66, 64, 61, 59, 60, 56, 58, 66, 51, 72, 98, 86, 
    55, 61, 63, 61, 55, 44, 36, 34, 36, 37, 39, 44, 47, 49, 45, 44, 48, 51, 55, 58, 66, 69, 66, 60, 58, 68, 72, 87, 104, 89, 
    45, 51, 52, 39, 31, 31, 27, 26, 27, 31, 37, 42, 48, 53, 54, 51, 53, 59, 66, 73, 79, 73, 61, 59, 57, 67, 87, 95, 83, 70, 
    44, 35, 35, 39, 41, 41, 35, 29, 28, 31, 37, 45, 55, 64, 72, 73, 68, 70, 74, 75, 68, 61, 55, 55, 57, 64, 69, 59, 60, 78, 
    32, 38, 55, 61, 49, 35, 35, 33, 34, 43, 53, 61, 68, 72, 73, 70, 61, 63, 68, 63, 56, 54, 55, 56, 61, 60, 58, 60, 65, 70, 
    53, 64, 61, 45, 36, 33, 34, 42, 55, 65, 65, 63, 61, 58, 55, 58, 60, 63, 63, 59, 53, 51, 53, 56, 59, 61, 69, 74, 76, 75, 
    57, 44, 35, 35, 41, 47, 48, 53, 58, 55, 55, 55, 55, 51, 50, 59, 68, 74, 67, 60, 55, 50, 51, 60, 74, 83, 85, 89, 90, 69, 
    51, 46, 44, 47, 48, 48, 50, 44, 43, 47, 57, 62, 60, 57, 67, 81, 80, 77, 67, 59, 58, 60, 72, 86, 90, 89, 94, 98, 87, 79, 
    61, 52, 49, 49, 49, 45, 51, 52, 50, 57, 67, 65, 67, 75, 82, 86, 77, 62, 63, 71, 78, 87, 89, 87, 89, 95, 99, 93, 90, 98, 
    58, 55, 54, 54, 55, 58, 68, 72, 71, 68, 62, 57, 61, 69, 70, 72, 74, 75, 83, 89, 90, 90, 91, 96, 95, 94, 93, 94, 100, 101, 
    59, 60, 58, 59, 65, 72, 74, 75, 76, 67, 52, 50, 58, 69, 81, 87, 87, 85, 85, 85, 90, 102, 106, 99, 87, 88, 94, 97, 98, 98, 
    62, 60, 55, 55, 63, 70, 65, 65, 70, 74, 79, 84, 85, 85, 88, 89, 83, 80, 87, 97, 103, 100, 93, 91, 89, 92, 95, 98, 97, 97, 
    62, 61, 64, 67, 72, 77, 79, 84, 92, 97, 96, 93, 86, 85, 89, 91, 91, 97, 100, 98, 93, 92, 91, 90, 95, 98, 97, 98, 100, 97, 
    81, 82, 88, 92, 96, 97, 96, 95, 94, 95, 94, 92, 91, 94, 101, 104, 104, 98, 89, 91, 94, 94, 91, 92, 98, 98, 98, 99, 100, 97, 
    96, 96, 97, 100, 103, 103, 99, 97, 98, 99, 102, 104, 103, 101, 103, 100, 93, 92, 91, 95, 97, 91, 89, 94, 98, 98, 97, 99, 99, 98, 
    100, 100, 101, 102, 104, 105, 104, 104, 105, 106, 103, 101, 99, 100, 102, 96, 89, 94, 97, 98, 91, 88, 91, 94, 97, 97, 97, 98, 98, 104, 
    103, 103, 103, 103, 104, 102, 101, 101, 101, 101, 100, 100, 100, 101, 101, 95, 90, 96, 99, 93, 90, 90, 90, 93, 96, 98, 100, 97, 100, 114, 
    
    -- channel=40
    143, 160, 87, 34, 71, 88, 76, 57, 58, 68, 43, 15, 21, 16, 36, 38, 5, 7, 10, 27, 13, 0, 0, 22, 24, 0, 14, 31, 0, 0, 
    126, 144, 72, 13, 47, 71, 62, 32, 38, 54, 33, 3, 12, 6, 22, 35, 3, 6, 29, 43, 0, 0, 0, 15, 20, 0, 7, 32, 0, 0, 
    113, 129, 56, 0, 24, 48, 48, 9, 16, 43, 24, 0, 10, 1, 3, 29, 1, 12, 74, 76, 0, 0, 0, 8, 17, 0, 0, 25, 0, 0, 
    100, 122, 44, 0, 7, 26, 34, 0, 0, 31, 18, 0, 12, 11, 0, 15, 0, 16, 116, 93, 0, 0, 0, 3, 17, 0, 0, 12, 0, 0, 
    83, 117, 35, 0, 0, 3, 16, 0, 0, 20, 9, 0, 19, 38, 0, 0, 0, 11, 142, 102, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    68, 111, 25, 0, 0, 0, 0, 0, 0, 5, 0, 0, 16, 47, 15, 26, 16, 21, 110, 101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    50, 88, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 43, 84, 92, 83, 102, 117, 71, 66, 25, 0, 0, 0, 0, 0, 0, 0, 
    32, 61, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 125, 127, 121, 122, 124, 108, 115, 74, 0, 0, 0, 0, 6, 0, 0, 
    39, 59, 43, 10, 26, 14, 0, 0, 0, 0, 0, 1, 11, 19, 77, 127, 117, 111, 122, 125, 101, 88, 50, 26, 0, 0, 27, 67, 0, 0, 
    63, 79, 60, 50, 84, 78, 41, 20, 39, 52, 36, 44, 65, 83, 115, 126, 110, 104, 118, 128, 76, 37, 41, 53, 48, 0, 3, 119, 72, 48, 
    77, 102, 70, 52, 109, 116, 62, 38, 79, 111, 90, 82, 110, 135, 138, 126, 105, 93, 105, 113, 37, 0, 9, 56, 99, 0, 0, 127, 114, 69, 
    87, 117, 88, 62, 110, 108, 66, 44, 71, 117, 124, 110, 128, 155, 151, 130, 114, 97, 99, 88, 12, 0, 0, 10, 86, 35, 0, 95, 142, 63, 
    101, 121, 111, 94, 113, 102, 77, 69, 81, 107, 135, 133, 136, 153, 146, 132, 130, 116, 106, 78, 9, 0, 0, 0, 36, 82, 0, 52, 132, 59, 
    122, 125, 123, 111, 127, 119, 103, 103, 106, 111, 125, 132, 134, 143, 132, 113, 116, 114, 106, 67, 1, 0, 0, 0, 12, 91, 106, 43, 85, 75, 
    131, 115, 120, 107, 110, 122, 117, 111, 112, 116, 119, 121, 123, 132, 129, 101, 90, 97, 112, 68, 0, 0, 0, 0, 16, 81, 135, 44, 49, 107, 
    128, 111, 121, 111, 82, 93, 115, 121, 120, 123, 126, 124, 120, 117, 120, 99, 70, 82, 119, 82, 2, 0, 0, 10, 28, 57, 80, 10, 12, 88, 
    139, 127, 121, 112, 83, 79, 106, 128, 133, 129, 127, 123, 116, 107, 101, 95, 63, 59, 95, 78, 17, 18, 30, 35, 40, 46, 49, 9, 0, 27, 
    159, 128, 114, 112, 112, 104, 110, 131, 136, 125, 118, 111, 104, 97, 87, 90, 68, 43, 67, 66, 33, 32, 51, 54, 54, 57, 56, 42, 22, 0, 
    171, 127, 109, 112, 119, 130, 128, 125, 121, 115, 107, 98, 92, 93, 90, 87, 57, 25, 50, 61, 48, 45, 63, 72, 65, 69, 75, 70, 47, 2, 
    157, 134, 123, 128, 124, 133, 139, 114, 98, 99, 96, 95, 110, 123, 110, 93, 33, 0, 40, 66, 64, 66, 76, 84, 78, 85, 89, 70, 67, 67, 
    119, 140, 143, 137, 133, 131, 134, 113, 92, 82, 72, 91, 140, 166, 130, 104, 44, 0, 46, 74, 76, 83, 88, 92, 90, 93, 86, 68, 79, 99, 
    87, 129, 138, 133, 151, 155, 130, 117, 109, 73, 44, 79, 137, 171, 135, 103, 71, 35, 61, 82, 87, 96, 102, 94, 89, 97, 90, 81, 87, 98, 
    72, 114, 127, 129, 171, 185, 138, 120, 120, 87, 54, 79, 114, 131, 111, 93, 84, 71, 83, 94, 99, 100, 99, 96, 100, 103, 96, 92, 92, 89, 
    73, 105, 121, 121, 156, 175, 134, 114, 111, 94, 77, 88, 102, 106, 98, 93, 91, 87, 92, 99, 100, 99, 89, 90, 108, 107, 94, 96, 92, 86, 
    77, 95, 112, 109, 121, 133, 116, 104, 104, 96, 92, 93, 96, 98, 94, 95, 96, 89, 92, 98, 99, 98, 82, 84, 110, 106, 92, 93, 94, 87, 
    89, 95, 105, 103, 108, 108, 102, 96, 95, 93, 89, 88, 88, 90, 92, 97, 94, 92, 105, 101, 94, 92, 87, 89, 103, 99, 90, 91, 92, 92, 
    100, 97, 95, 93, 98, 96, 87, 84, 86, 85, 85, 87, 92, 93, 95, 89, 69, 91, 123, 107, 90, 92, 93, 94, 97, 92, 88, 86, 88, 97, 
    93, 90, 83, 82, 85, 86, 81, 81, 87, 90, 90, 90, 94, 93, 92, 76, 45, 85, 139, 106, 85, 92, 92, 93, 91, 88, 87, 80, 92, 100, 
    82, 82, 77, 80, 84, 85, 84, 85, 88, 91, 91, 90, 94, 92, 89, 69, 35, 83, 139, 102, 86, 90, 92, 92, 90, 87, 82, 83, 100, 94, 
    80, 81, 79, 82, 85, 84, 82, 83, 84, 85, 87, 89, 94, 90, 84, 61, 24, 72, 129, 100, 85, 89, 89, 92, 92, 83, 79, 97, 99, 77, 
    
    -- channel=41
    9, 16, 20, 18, 9, 9, 11, 11, 10, 11, 15, 18, 17, 16, 18, 18, 21, 19, 17, 21, 27, 31, 24, 20, 18, 18, 17, 17, 17, 16, 
    21, 26, 27, 25, 18, 18, 20, 21, 20, 21, 25, 26, 28, 24, 25, 22, 24, 24, 33, 45, 51, 44, 26, 22, 20, 21, 19, 20, 21, 22, 
    24, 31, 31, 32, 26, 25, 24, 26, 27, 26, 29, 30, 32, 28, 30, 25, 25, 29, 43, 60, 64, 43, 24, 22, 23, 24, 25, 23, 24, 23, 
    26, 34, 36, 39, 31, 32, 32, 35, 36, 32, 33, 31, 35, 38, 42, 40, 34, 40, 47, 52, 50, 34, 26, 28, 29, 32, 35, 30, 26, 23, 
    34, 41, 42, 48, 39, 38, 36, 38, 41, 38, 37, 35, 40, 49, 61, 64, 54, 50, 57, 67, 66, 51, 44, 42, 39, 42, 46, 40, 34, 33, 
    39, 44, 44, 49, 42, 40, 39, 42, 47, 45, 42, 42, 44, 47, 57, 62, 75, 83, 81, 79, 89, 113, 119, 97, 71, 51, 49, 49, 48, 52, 
    46, 47, 44, 44, 45, 46, 49, 49, 53, 52, 47, 49, 50, 42, 37, 52, 86, 110, 114, 100, 99, 127, 148, 145, 113, 77, 65, 71, 72, 75, 
    82, 75, 72, 77, 88, 89, 85, 80, 82, 79, 71, 70, 71, 68, 62, 64, 61, 50, 38, 31, 30, 35, 44, 71, 82, 96, 97, 104, 107, 102, 
    104, 97, 96, 102, 107, 106, 107, 107, 107, 103, 100, 96, 90, 84, 76, 68, 55, 47, 49, 53, 54, 54, 43, 35, 43, 61, 77, 84, 103, 104, 
    84, 81, 75, 66, 60, 71, 81, 81, 76, 75, 79, 70, 59, 55, 59, 63, 60, 61, 66, 67, 56, 40, 26, 38, 65, 56, 52, 41, 60, 75, 
    53, 51, 46, 43, 42, 51, 55, 44, 28, 32, 37, 31, 25, 30, 42, 47, 48, 50, 47, 40, 29, 12, 0, 0, 29, 56, 67, 59, 54, 74, 
    36, 42, 59, 69, 66, 59, 45, 32, 24, 23, 25, 32, 37, 39, 45, 50, 52, 48, 44, 36, 31, 31, 35, 31, 26, 47, 61, 76, 67, 82, 
    42, 52, 60, 65, 67, 58, 49, 50, 48, 38, 26, 21, 19, 17, 12, 11, 11, 15, 20, 22, 28, 39, 54, 60, 48, 54, 68, 89, 88, 91, 
    34, 39, 36, 28, 20, 11, 6, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 15, 32, 49, 58, 61, 58, 52, 55, 75, 97, 98, 78, 
    12, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 8, 17, 27, 35, 42, 60, 78, 88, 81, 67, 55, 48, 45, 42, 39, 36, 29, 
    19, 19, 20, 24, 24, 20, 10, 8, 11, 15, 21, 29, 38, 45, 52, 56, 58, 56, 56, 58, 55, 50, 47, 48, 46, 41, 25, 6, 0, 5, 
    33, 42, 58, 63, 55, 38, 23, 17, 20, 30, 42, 52, 60, 63, 56, 49, 40, 32, 22, 15, 16, 26, 37, 42, 47, 47, 46, 57, 72, 62, 
    51, 62, 54, 27, 13, 17, 30, 39, 46, 52, 51, 45, 37, 32, 27, 28, 33, 39, 34, 28, 29, 33, 38, 41, 50, 56, 69, 87, 98, 86, 
    35, 22, 3, 0, 4, 21, 37, 47, 46, 34, 24, 20, 22, 30, 45, 59, 63, 59, 47, 40, 38, 40, 47, 58, 72, 86, 96, 100, 103, 100, 
    0, 0, 13, 30, 37, 35, 32, 31, 28, 26, 32, 39, 52, 70, 92, 108, 100, 78, 54, 46, 49, 58, 73, 89, 98, 98, 93, 88, 86, 96, 
    35, 24, 25, 27, 31, 35, 42, 49, 60, 64, 63, 54, 56, 72, 89, 91, 82, 73, 67, 71, 81, 90, 96, 95, 91, 91, 91, 87, 86, 98, 
    56, 38, 35, 36, 47, 63, 80, 85, 85, 80, 66, 48, 40, 40, 39, 40, 50, 68, 90, 99, 97, 93, 89, 91, 97, 97, 95, 95, 101, 102, 
    56, 52, 49, 46, 52, 63, 72, 66, 54, 49, 49, 55, 59, 56, 55, 61, 72, 81, 86, 86, 87, 92, 93, 93, 88, 86, 90, 93, 96, 91, 
    49, 47, 43, 43, 42, 39, 36, 39, 44, 54, 71, 92, 101, 99, 90, 81, 74, 72, 77, 88, 99, 102, 87, 75, 73, 83, 87, 86, 84, 81, 
    63, 65, 68, 75, 77, 73, 70, 79, 93, 104, 107, 99, 84, 73, 73, 78, 84, 90, 97, 96, 90, 85, 85, 87, 87, 88, 87, 86, 82, 79, 
    102, 111, 116, 118, 116, 111, 104, 98, 92, 85, 80, 79, 79, 84, 94, 100, 96, 89, 81, 80, 83, 87, 91, 92, 92, 88, 84, 84, 82, 81, 
    109, 112, 112, 107, 101, 95, 90, 86, 87, 89, 93, 96, 97, 96, 97, 93, 75, 62, 67, 84, 89, 86, 85, 88, 88, 85, 83, 82, 84, 87, 
    88, 89, 92, 94, 94, 95, 96, 98, 99, 99, 96, 91, 84, 79, 82, 85, 80, 76, 80, 88, 86, 82, 85, 87, 85, 83, 81, 81, 89, 99, 
    90, 88, 89, 90, 90, 89, 88, 87, 83, 79, 76, 79, 83, 85, 91, 96, 94, 89, 85, 86, 83, 84, 86, 85, 85, 85, 82, 85, 96, 111, 
    86, 83, 82, 79, 78, 77, 77, 79, 82, 86, 90, 95, 101, 103, 107, 109, 103, 93, 84, 84, 84, 83, 83, 85, 87, 86, 87, 91, 104, 112, 
    
    -- channel=42
    1, 3, 12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 5, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 0, 1, 0, 16, 35, 18, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 70, 92, 83, 86, 110, 124, 104, 41, 0, 0, 0, 0, 0, 
    6, 7, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 51, 73, 83, 74, 60, 68, 86, 105, 89, 39, 8, 3, 8, 3, 
    63, 53, 49, 55, 65, 61, 55, 40, 34, 32, 28, 27, 27, 30, 28, 37, 46, 38, 28, 27, 27, 21, 11, 7, 13, 34, 32, 47, 56, 53, 
    90, 78, 75, 71, 68, 67, 69, 69, 65, 62, 66, 67, 64, 60, 58, 61, 56, 48, 47, 55, 57, 39, 11, 0, 0, 6, 0, 2, 43, 54, 
    71, 56, 45, 32, 20, 32, 51, 53, 37, 32, 44, 43, 38, 38, 44, 46, 43, 44, 43, 43, 33, 3, 0, 0, 0, 1, 0, 0, 12, 39, 
    41, 27, 27, 35, 26, 33, 33, 21, 0, 0, 9, 25, 31, 36, 46, 49, 44, 42, 33, 21, 3, 0, 0, 0, 0, 0, 7, 0, 11, 53, 
    36, 32, 40, 58, 65, 59, 47, 39, 35, 28, 20, 34, 46, 44, 43, 41, 36, 32, 25, 8, 0, 0, 0, 0, 0, 0, 0, 22, 20, 67, 
    46, 47, 47, 52, 60, 61, 50, 39, 36, 31, 18, 10, 10, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 60, 60, 65, 
    31, 27, 18, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 19, 13, 4, 0, 0, 0, 6, 42, 55, 31, 
    22, 15, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 6, 8, 13, 25, 35, 28, 30, 42, 47, 24, 8, 0, 0, 0, 0, 0, 0, 0, 
    37, 27, 30, 45, 56, 50, 26, 20, 20, 22, 26, 34, 40, 44, 45, 41, 38, 23, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 70, 79, 76, 61, 51, 40, 32, 38, 48, 54, 54, 48, 37, 24, 11, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 24, 30, 
    76, 81, 56, 23, 10, 16, 41, 55, 59, 55, 42, 27, 13, 2, 0, 0, 2, 9, 4, 0, 0, 0, 0, 0, 9, 20, 38, 52, 64, 63, 
    35, 29, 22, 18, 25, 32, 39, 49, 39, 20, 10, 8, 10, 20, 35, 53, 59, 44, 17, 6, 3, 5, 13, 27, 49, 59, 65, 69, 68, 69, 
    25, 17, 27, 42, 45, 41, 32, 32, 35, 28, 28, 28, 34, 58, 91, 104, 96, 69, 27, 15, 24, 38, 55, 63, 64, 67, 65, 59, 55, 65, 
    66, 40, 36, 38, 39, 47, 59, 67, 78, 83, 68, 41, 31, 41, 60, 60, 49, 49, 51, 56, 66, 70, 69, 68, 68, 68, 68, 64, 65, 75, 
    81, 57, 51, 49, 54, 73, 97, 101, 93, 84, 67, 37, 20, 16, 15, 20, 32, 51, 70, 75, 70, 68, 71, 75, 78, 74, 73, 73, 78, 80, 
    67, 60, 55, 50, 47, 51, 62, 58, 45, 36, 40, 55, 68, 70, 61, 54, 54, 54, 57, 61, 70, 78, 74, 66, 62, 67, 72, 70, 71, 68, 
    56, 51, 46, 49, 48, 41, 37, 42, 52, 67, 80, 93, 96, 86, 72, 61, 57, 59, 65, 73, 77, 76, 68, 61, 56, 68, 75, 71, 65, 62, 
    80, 86, 88, 96, 100, 98, 89, 86, 87, 88, 86, 79, 70, 62, 59, 66, 78, 84, 80, 72, 69, 67, 69, 74, 74, 74, 72, 70, 67, 62, 
    112, 123, 126, 120, 114, 109, 99, 86, 73, 66, 63, 66, 74, 79, 80, 82, 78, 64, 54, 61, 68, 70, 74, 75, 77, 74, 69, 67, 65, 63, 
    94, 97, 100, 94, 87, 82, 80, 79, 77, 79, 82, 81, 80, 75, 71, 68, 62, 46, 42, 66, 74, 69, 70, 72, 73, 69, 67, 64, 62, 65, 
    70, 71, 75, 76, 76, 76, 78, 80, 80, 75, 71, 67, 65, 61, 59, 64, 68, 62, 59, 71, 71, 68, 71, 72, 70, 69, 65, 61, 63, 72, 
    69, 66, 67, 66, 65, 64, 63, 62, 61, 59, 58, 61, 66, 68, 69, 76, 81, 72, 64, 69, 70, 70, 72, 70, 71, 71, 68, 62, 68, 79, 
    62, 59, 58, 58, 59, 59, 59, 59, 62, 66, 71, 76, 83, 87, 89, 94, 97, 82, 68, 70, 71, 71, 69, 70, 72, 71, 68, 67, 74, 80, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    
    -- channel=44
    238, 214, 240, 277, 281, 282, 284, 290, 290, 278, 283, 293, 293, 294, 280, 279, 291, 298, 302, 295, 291, 298, 296, 285, 284, 296, 291, 281, 289, 297, 
    245, 217, 242, 281, 286, 280, 280, 291, 291, 276, 282, 291, 294, 296, 286, 280, 290, 300, 305, 289, 293, 305, 298, 287, 286, 300, 294, 281, 292, 302, 
    242, 216, 241, 278, 284, 278, 275, 288, 287, 271, 273, 282, 286, 291, 288, 279, 288, 296, 272, 245, 281, 304, 299, 287, 285, 300, 295, 277, 292, 298, 
    238, 212, 236, 275, 280, 274, 268, 284, 284, 265, 265, 277, 274, 284, 291, 284, 287, 290, 239, 215, 271, 298, 299, 289, 283, 297, 292, 276, 291, 295, 
    238, 205, 230, 271, 275, 269, 260, 278, 276, 259, 260, 273, 260, 261, 274, 277, 290, 280, 206, 200, 279, 306, 309, 296, 281, 289, 285, 276, 289, 289, 
    230, 191, 216, 256, 263, 258, 254, 271, 264, 252, 254, 268, 244, 223, 236, 247, 283, 278, 207, 204, 264, 301, 324, 318, 292, 282, 275, 270, 282, 280, 
    227, 183, 213, 250, 259, 253, 258, 266, 254, 248, 251, 260, 240, 227, 222, 206, 211, 202, 170, 158, 169, 184, 219, 274, 292, 289, 273, 260, 271, 276, 
    226, 190, 217, 245, 247, 249, 261, 262, 251, 252, 254, 254, 245, 252, 224, 180, 150, 135, 123, 113, 117, 98, 97, 165, 214, 253, 245, 224, 249, 258, 
    192, 173, 179, 188, 188, 201, 216, 218, 218, 223, 229, 223, 224, 235, 208, 172, 157, 154, 145, 143, 144, 120, 127, 146, 164, 189, 171, 141, 185, 193, 
    139, 128, 126, 135, 129, 138, 148, 157, 159, 159, 168, 169, 181, 188, 173, 160, 156, 153, 140, 132, 131, 131, 145, 132, 160, 187, 157, 101, 120, 136, 
    116, 114, 129, 146, 126, 111, 119, 142, 134, 128, 143, 162, 173, 169, 161, 156, 151, 148, 138, 124, 149, 181, 173, 137, 128, 186, 184, 125, 99, 127, 
    134, 125, 146, 164, 140, 123, 146, 175, 171, 159, 161, 179, 182, 168, 159, 152, 152, 155, 152, 144, 188, 227, 231, 204, 137, 170, 184, 135, 95, 125, 
    147, 132, 136, 135, 125, 132, 154, 177, 191, 181, 168, 171, 169, 158, 145, 143, 143, 152, 156, 164, 204, 224, 231, 227, 172, 159, 176, 132, 93, 107, 
    137, 128, 119, 105, 102, 113, 138, 159, 176, 182, 183, 186, 184, 180, 181, 186, 183, 187, 188, 197, 221, 221, 218, 210, 188, 143, 131, 100, 84, 79, 
    148, 143, 136, 140, 145, 154, 176, 196, 209, 217, 224, 229, 231, 225, 227, 233, 234, 224, 200, 193, 207, 209, 209, 198, 193, 137, 79, 67, 67, 55, 
    177, 185, 187, 200, 213, 224, 225, 231, 239, 244, 249, 254, 257, 247, 232, 225, 223, 204, 156, 145, 165, 182, 192, 194, 196, 156, 120, 140, 127, 87, 
    197, 201, 193, 192, 215, 233, 239, 241, 245, 247, 246, 242, 235, 224, 205, 199, 202, 193, 153, 148, 169, 179, 188, 191, 193, 179, 180, 203, 193, 162, 
    175, 165, 160, 163, 190, 215, 237, 240, 233, 228, 219, 211, 204, 202, 199, 198, 205, 212, 195, 189, 197, 195, 195, 190, 194, 189, 185, 181, 180, 188, 
    134, 148, 171, 191, 202, 210, 213, 208, 206, 207, 208, 212, 215, 219, 224, 217, 218, 225, 213, 205, 206, 207, 203, 197, 192, 176, 158, 137, 139, 178, 
    154, 175, 197, 212, 215, 206, 194, 196, 211, 218, 225, 227, 226, 216, 207, 196, 208, 228, 218, 209, 210, 211, 195, 177, 162, 144, 121, 104, 110, 129, 
    202, 199, 199, 202, 209, 207, 200, 209, 222, 228, 230, 221, 191, 152, 134, 126, 165, 213, 218, 209, 200, 184, 163, 146, 133, 116, 102, 105, 95, 71, 
    216, 208, 204, 206, 204, 194, 189, 187, 183, 197, 217, 210, 164, 117, 104, 107, 147, 183, 187, 177, 164, 150, 135, 123, 112, 97, 95, 95, 72, 47, 
    198, 200, 198, 197, 170, 140, 136, 136, 130, 163, 201, 210, 184, 152, 138, 132, 140, 147, 145, 141, 136, 127, 107, 99, 87, 78, 76, 64, 50, 37, 
    178, 185, 186, 188, 153, 122, 122, 134, 145, 171, 186, 182, 164, 147, 139, 130, 129, 132, 130, 120, 110, 104, 95, 90, 71, 65, 61, 52, 42, 35, 
    178, 188, 189, 191, 170, 153, 148, 148, 148, 149, 143, 131, 119, 116, 121, 123, 124, 122, 113, 97, 90, 85, 93, 91, 67, 57, 55, 50, 42, 40, 
    158, 162, 158, 152, 141, 131, 124, 117, 109, 105, 104, 108, 112, 116, 116, 107, 96, 96, 88, 84, 80, 73, 79, 73, 59, 52, 51, 48, 47, 47, 
    92, 91, 93, 90, 86, 86, 92, 96, 98, 100, 100, 99, 98, 95, 90, 82, 87, 91, 77, 74, 70, 64, 61, 55, 52, 50, 49, 48, 51, 44, 
    49, 48, 55, 62, 67, 71, 79, 83, 83, 81, 79, 79, 79, 78, 73, 78, 105, 101, 71, 63, 63, 56, 51, 48, 49, 50, 49, 52, 50, 30, 
    44, 42, 45, 50, 54, 56, 59, 63, 65, 67, 70, 75, 79, 78, 71, 76, 105, 94, 62, 58, 55, 47, 47, 45, 49, 51, 52, 55, 34, 12, 
    41, 41, 44, 48, 52, 54, 57, 63, 69, 72, 75, 76, 76, 71, 60, 64, 93, 84, 58, 52, 47, 44, 42, 43, 47, 49, 56, 44, 13, 0, 
    
    -- channel=45
    251, 228, 206, 225, 269, 285, 285, 285, 295, 294, 285, 284, 293, 294, 293, 286, 280, 293, 304, 306, 289, 280, 289, 294, 291, 289, 298, 299, 288, 296, 
    248, 223, 202, 222, 264, 277, 275, 274, 285, 285, 276, 274, 285, 288, 287, 286, 278, 290, 306, 289, 253, 256, 285, 293, 292, 289, 300, 298, 288, 294, 
    241, 218, 196, 214, 254, 269, 269, 263, 274, 275, 264, 263, 275, 280, 278, 284, 275, 284, 279, 237, 205, 238, 284, 294, 291, 286, 297, 292, 283, 291, 
    240, 215, 189, 204, 245, 256, 255, 250, 262, 266, 254, 254, 264, 270, 263, 270, 261, 272, 269, 207, 178, 232, 282, 290, 287, 278, 283, 283, 279, 290, 
    234, 209, 181, 191, 233, 245, 246, 242, 254, 255, 243, 246, 253, 248, 226, 229, 240, 247, 227, 172, 164, 226, 264, 270, 273, 261, 261, 266, 267, 280, 
    225, 196, 165, 175, 224, 235, 238, 235, 243, 240, 232, 239, 234, 212, 198, 207, 222, 223, 184, 143, 138, 174, 196, 198, 222, 236, 243, 250, 243, 253, 
    215, 183, 164, 180, 224, 224, 222, 227, 229, 223, 219, 228, 222, 211, 208, 195, 152, 114, 82, 61, 50, 51, 58, 85, 144, 203, 225, 224, 205, 211, 
    170, 150, 144, 156, 172, 173, 180, 193, 194, 191, 195, 203, 196, 193, 190, 164, 117, 94, 87, 80, 77, 63, 31, 43, 93, 141, 172, 158, 144, 155, 
    94, 90, 77, 75, 88, 94, 103, 115, 122, 126, 132, 137, 140, 151, 155, 133, 109, 103, 100, 92, 76, 63, 70, 85, 103, 97, 121, 103, 81, 89, 
    39, 41, 35, 46, 69, 70, 55, 58, 78, 85, 80, 90, 113, 131, 126, 107, 91, 82, 75, 64, 49, 56, 90, 103, 111, 99, 115, 121, 71, 63, 
    34, 54, 61, 72, 90, 65, 43, 63, 91, 104, 101, 114, 138, 145, 131, 109, 93, 82, 80, 71, 76, 115, 160, 160, 137, 116, 108, 135, 77, 46, 
    66, 76, 73, 75, 80, 65, 74, 107, 132, 137, 135, 133, 139, 136, 116, 96, 89, 88, 93, 94, 110, 154, 195, 198, 165, 139, 112, 116, 79, 27, 
    83, 80, 68, 57, 59, 55, 68, 96, 124, 138, 140, 142, 145, 143, 128, 119, 119, 122, 125, 130, 145, 168, 184, 187, 170, 149, 129, 85, 47, 3, 
    89, 84, 77, 63, 68, 81, 105, 134, 158, 172, 182, 188, 191, 191, 190, 187, 190, 188, 182, 166, 157, 158, 162, 166, 163, 140, 102, 31, 0, 0, 
    124, 118, 124, 134, 150, 173, 190, 204, 215, 220, 222, 224, 227, 223, 219, 209, 203, 194, 171, 128, 102, 118, 138, 153, 159, 137, 83, 24, 23, 39, 
    145, 157, 169, 172, 173, 190, 212, 224, 231, 234, 233, 230, 223, 210, 191, 173, 159, 155, 132, 97, 86, 116, 140, 154, 161, 145, 124, 121, 128, 109, 
    161, 158, 139, 121, 137, 172, 207, 228, 234, 226, 211, 194, 176, 163, 149, 148, 153, 156, 152, 137, 134, 148, 158, 157, 157, 151, 147, 142, 136, 117, 
    126, 95, 91, 114, 149, 183, 201, 205, 193, 177, 166, 162, 161, 164, 168, 168, 165, 165, 170, 168, 165, 169, 168, 164, 161, 152, 133, 110, 91, 84, 
    102, 105, 137, 173, 186, 189, 180, 161, 155, 163, 173, 182, 189, 191, 186, 170, 147, 146, 165, 170, 171, 177, 175, 164, 135, 109, 82, 51, 35, 57, 
    143, 152, 165, 173, 175, 173, 170, 162, 167, 180, 182, 183, 187, 172, 133, 99, 84, 105, 154, 171, 172, 167, 143, 109, 78, 57, 35, 14, 14, 21, 
    146, 164, 170, 170, 175, 177, 166, 158, 155, 150, 150, 161, 156, 115, 58, 29, 44, 91, 141, 148, 130, 106, 83, 62, 44, 25, 7, 6, 2, 0, 
    122, 158, 165, 165, 167, 148, 114, 96, 90, 92, 114, 148, 147, 111, 71, 56, 65, 80, 91, 82, 70, 62, 49, 28, 9, 0, 0, 0, 0, 0, 
    98, 132, 141, 143, 133, 99, 58, 51, 59, 82, 120, 151, 147, 116, 83, 62, 52, 49, 52, 53, 43, 26, 6, 0, 0, 0, 0, 0, 0, 0, 
    87, 119, 134, 138, 126, 100, 77, 78, 88, 96, 100, 91, 70, 51, 41, 40, 44, 46, 43, 25, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    86, 110, 119, 113, 102, 85, 69, 56, 43, 30, 24, 24, 26, 30, 33, 34, 29, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 40, 36, 27, 19, 10, 5, 3, 3, 2, 5, 10, 14, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 12, 22, 31, 40, 50, 56, 59, 58, 55, 58, 60, 57, 59, 66, 73, 72, 71, 70, 70, 73, 76, 78, 
    0, 0, 0, 0, 0, 1, 11, 20, 28, 38, 40, 47, 49, 55, 58, 62, 60, 56, 41, 26, 36, 59, 79, 77, 74, 72, 75, 76, 78, 76, 
    0, 0, 0, 0, 13, 23, 31, 39, 48, 56, 56, 61, 57, 59, 60, 65, 64, 52, 26, 20, 33, 60, 79, 80, 78, 76, 76, 80, 81, 82, 
    5, 6, 10, 15, 33, 42, 52, 59, 64, 71, 70, 71, 62, 54, 47, 50, 59, 44, 25, 17, 31, 61, 75, 79, 80, 78, 78, 84, 82, 84, 
    18, 16, 20, 26, 48, 62, 76, 82, 83, 82, 78, 79, 71, 53, 39, 33, 43, 31, 16, 10, 4, 19, 37, 57, 72, 80, 84, 86, 83, 86, 
    39, 34, 40, 52, 75, 87, 98, 103, 103, 98, 92, 87, 85, 80, 65, 37, 0, 0, 0, 0, 0, 0, 0, 0, 26, 75, 94, 93, 92, 101, 
    37, 43, 51, 64, 69, 81, 90, 103, 106, 104, 98, 88, 89, 89, 65, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 65, 70, 80, 93, 
    0, 10, 9, 10, 6, 22, 34, 48, 60, 62, 60, 50, 45, 30, 14, 0, 0, 0, 0, 0, 0, 15, 37, 35, 37, 27, 35, 33, 38, 46, 
    0, 0, 0, 0, 0, 0, 0, 3, 13, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 60, 70, 75, 81, 72, 29, 19, 
    0, 0, 2, 14, 16, 5, 0, 9, 17, 14, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 81, 94, 74, 98, 110, 110, 50, 21, 
    0, 1, 9, 6, 5, 0, 13, 24, 31, 25, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 81, 116, 137, 114, 108, 104, 85, 52, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 40, 64, 82, 101, 120, 105, 106, 64, 44, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 14, 35, 53, 69, 74, 80, 104, 84, 74, 41, 20, 0, 
    0, 0, 0, 9, 10, 11, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 11, 15, 26, 54, 75, 83, 92, 76, 46, 49, 38, 35, 
    0, 0, 7, 21, 18, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 49, 72, 81, 79, 80, 87, 128, 138, 117, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 40, 65, 79, 79, 69, 60, 70, 100, 132, 142, 128, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 53, 72, 82, 79, 67, 53, 48, 55, 56, 46, 52, 65, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 8, 13, 28, 40, 48, 53, 48, 44, 34, 26, 13, 6, 5, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 21, 29, 32, 22, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 3, 0, 0, 0, 0, 0, 0, 6, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 10, 
    8, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 6, 11, 18, 
    13, 16, 14, 9, 7, 7, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 3, 0, 0, 0, 0, 4, 19, 31, 
    
    -- channel=48
    129, 141, 156, 168, 164, 161, 159, 155, 151, 164, 176, 182, 183, 180, 176, 177, 179, 179, 180, 181, 183, 183, 181, 181, 181, 185, 197, 204, 203, 221, 
    124, 133, 148, 164, 166, 171, 169, 151, 141, 154, 165, 167, 172, 163, 159, 167, 173, 169, 171, 171, 175, 178, 167, 160, 172, 183, 196, 202, 203, 222, 
    125, 132, 144, 160, 173, 199, 195, 171, 171, 169, 165, 172, 179, 175, 167, 177, 181, 177, 178, 177, 178, 187, 170, 155, 180, 195, 200, 200, 203, 223, 
    122, 132, 142, 152, 166, 201, 190, 172, 194, 191, 183, 193, 195, 183, 181, 192, 198, 199, 199, 199, 195, 204, 188, 177, 191, 199, 202, 203, 202, 223, 
    122, 132, 142, 152, 169, 195, 168, 154, 175, 169, 164, 177, 174, 166, 166, 172, 176, 175, 183, 180, 173, 182, 170, 172, 174, 181, 196, 201, 199, 220, 
    122, 130, 141, 154, 177, 206, 174, 169, 168, 163, 168, 177, 177, 171, 166, 170, 171, 173, 181, 180, 172, 173, 176, 187, 167, 172, 194, 197, 194, 215, 
    124, 129, 139, 152, 177, 196, 179, 182, 173, 168, 170, 178, 180, 176, 174, 178, 178, 186, 193, 189, 186, 182, 192, 189, 171, 178, 188, 188, 188, 208, 
    131, 132, 135, 149, 166, 167, 165, 165, 150, 151, 142, 150, 153, 150, 153, 155, 157, 160, 166, 157, 158, 159, 172, 169, 167, 179, 186, 184, 183, 203, 
    143, 142, 140, 150, 154, 156, 161, 153, 139, 142, 140, 141, 141, 143, 146, 148, 148, 150, 152, 152, 152, 152, 157, 167, 178, 179, 182, 181, 180, 200, 
    158, 155, 152, 155, 155, 157, 163, 154, 148, 148, 148, 147, 146, 150, 155, 157, 158, 159, 157, 157, 159, 154, 152, 170, 182, 181, 182, 182, 180, 201, 
    170, 162, 157, 149, 138, 135, 148, 158, 158, 158, 154, 154, 157, 161, 166, 166, 162, 159, 161, 162, 164, 165, 165, 173, 181, 185, 189, 189, 186, 206, 
    178, 170, 164, 153, 125, 103, 105, 124, 145, 162, 169, 170, 170, 174, 178, 181, 181, 179, 179, 178, 177, 180, 183, 182, 183, 184, 186, 187, 185, 206, 
    183, 187, 181, 176, 159, 131, 112, 100, 104, 125, 150, 170, 178, 183, 186, 188, 188, 187, 185, 181, 179, 179, 180, 179, 180, 181, 183, 184, 184, 205, 
    184, 188, 178, 172, 176, 166, 137, 110, 87, 91, 116, 146, 173, 188, 192, 193, 193, 194, 192, 189, 186, 186, 186, 185, 183, 184, 183, 180, 177, 198, 
    187, 194, 193, 198, 205, 205, 179, 139, 91, 57, 71, 105, 135, 165, 187, 195, 196, 195, 192, 188, 186, 186, 184, 180, 180, 181, 181, 178, 174, 192, 
    191, 203, 202, 205, 210, 215, 220, 189, 128, 67, 51, 76, 97, 119, 141, 160, 177, 186, 189, 187, 183, 184, 185, 182, 182, 182, 181, 179, 174, 190, 
    194, 209, 210, 213, 215, 215, 224, 217, 162, 81, 50, 62, 68, 85, 103, 117, 126, 137, 147, 157, 163, 175, 186, 186, 185, 183, 182, 180, 175, 190, 
    200, 215, 217, 219, 219, 220, 218, 220, 174, 72, 33, 47, 48, 56, 70, 88, 99, 101, 99, 90, 91, 118, 150, 168, 179, 184, 188, 186, 179, 193, 
    201, 216, 216, 216, 215, 217, 211, 219, 160, 61, 27, 25, 36, 50, 54, 61, 68, 73, 75, 63, 58, 77, 102, 115, 122, 139, 153, 165, 172, 190, 
    194, 210, 213, 211, 211, 212, 216, 216, 155, 84, 51, 28, 15, 34, 53, 83, 103, 91, 70, 38, 42, 63, 79, 91, 109, 146, 163, 162, 168, 184, 
    189, 204, 207, 209, 211, 212, 227, 208, 169, 146, 120, 87, 72, 77, 89, 120, 148, 148, 121, 91, 96, 105, 103, 88, 102, 139, 158, 169, 178, 188, 
    179, 191, 195, 199, 198, 197, 197, 175, 156, 163, 157, 111, 92, 86, 93, 130, 156, 153, 115, 104, 121, 122, 107, 90, 106, 133, 137, 140, 149, 165, 
    130, 129, 135, 137, 135, 133, 129, 127, 124, 124, 120, 92, 78, 77, 84, 105, 118, 114, 97, 91, 98, 103, 98, 93, 98, 104, 105, 108, 111, 128, 
    118, 115, 116, 118, 117, 114, 114, 113, 109, 110, 106, 99, 94, 88, 88, 88, 84, 78, 78, 80, 77, 75, 74, 77, 75, 69, 65, 66, 64, 87, 
    78, 64, 64, 63, 60, 57, 57, 55, 53, 52, 46, 39, 34, 29, 34, 44, 48, 41, 36, 36, 36, 35, 34, 35, 36, 37, 41, 39, 33, 52, 
    66, 45, 48, 47, 45, 48, 51, 53, 58, 53, 47, 45, 44, 45, 44, 49, 55, 53, 48, 46, 45, 43, 43, 45, 45, 46, 48, 46, 42, 56, 
    68, 48, 54, 54, 52, 51, 49, 54, 58, 51, 44, 40, 39, 41, 42, 44, 47, 47, 41, 37, 35, 33, 33, 32, 31, 31, 36, 42, 45, 67, 
    50, 26, 32, 31, 34, 34, 32, 38, 40, 33, 27, 25, 31, 36, 38, 39, 43, 41, 37, 33, 34, 37, 38, 33, 30, 30, 38, 50, 62, 82, 
    53, 30, 32, 30, 33, 34, 35, 39, 40, 38, 35, 41, 44, 46, 48, 51, 55, 51, 48, 44, 42, 40, 40, 37, 37, 41, 52, 69, 79, 85, 
    54, 32, 32, 27, 27, 29, 33, 36, 36, 34, 33, 42, 46, 46, 47, 50, 50, 48, 47, 47, 46, 41, 44, 48, 50, 56, 69, 75, 69, 59, 
    
    -- channel=49
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 20, 22, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 19, 16, 11, 10, 12, 15, 17, 13, 6, 15, 8, 5, 5, 0, 19, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 24, 0, 0, 5, 0, 0, 18, 20, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 39, 5, 0, 0, 0, 0, 1, 8, 5, 2, 0, 0, 9, 8, 1, 0, 0, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 9, 0, 0, 4, 9, 13, 4, 6, 7, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 38, 33, 35, 37, 19, 7, 1, 15, 20, 21, 25, 30, 37, 28, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 16, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 5, 4, 4, 6, 6, 4, 3, 6, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    317, 354, 369, 357, 332, 316, 305, 303, 316, 334, 337, 336, 332, 326, 328, 330, 328, 328, 331, 337, 338, 333, 333, 335, 347, 364, 375, 378, 381, 370, 
    324, 361, 381, 385, 368, 334, 284, 274, 302, 324, 338, 333, 326, 320, 322, 334, 335, 332, 337, 338, 338, 337, 331, 348, 369, 376, 384, 388, 390, 379, 
    324, 355, 375, 384, 378, 332, 252, 242, 260, 260, 273, 271, 265, 268, 272, 278, 281, 280, 287, 289, 286, 283, 291, 333, 373, 383, 386, 388, 389, 378, 
    323, 355, 371, 381, 379, 336, 271, 239, 234, 228, 235, 245, 233, 232, 239, 250, 256, 259, 264, 266, 265, 262, 282, 327, 373, 391, 389, 391, 394, 383, 
    319, 351, 365, 376, 376, 327, 269, 255, 263, 258, 252, 253, 235, 233, 251, 272, 279, 289, 288, 283, 286, 287, 297, 308, 346, 384, 390, 390, 394, 382, 
    316, 348, 364, 373, 352, 279, 226, 232, 263, 264, 254, 257, 245, 236, 250, 262, 277, 283, 276, 272, 271, 282, 287, 279, 311, 364, 387, 389, 392, 381, 
    318, 345, 363, 366, 332, 279, 235, 221, 255, 259, 262, 264, 257, 249, 255, 256, 263, 268, 262, 250, 256, 278, 280, 274, 296, 345, 379, 382, 386, 377, 
    327, 346, 360, 362, 353, 329, 292, 265, 275, 281, 282, 279, 282, 282, 286, 289, 292, 291, 281, 269, 273, 288, 312, 328, 322, 348, 380, 385, 385, 375, 
    340, 352, 360, 367, 370, 358, 332, 309, 301, 301, 300, 300, 306, 310, 314, 317, 316, 313, 308, 303, 303, 313, 345, 370, 367, 373, 384, 385, 385, 374, 
    356, 363, 369, 370, 367, 366, 357, 338, 330, 326, 326, 330, 333, 338, 340, 338, 337, 339, 336, 332, 334, 338, 353, 375, 383, 380, 379, 381, 386, 376, 
    365, 372, 362, 341, 328, 347, 371, 369, 361, 361, 358, 359, 364, 368, 371, 370, 364, 360, 360, 358, 361, 364, 363, 374, 384, 383, 383, 386, 390, 380, 
    368, 365, 330, 293, 263, 271, 307, 339, 363, 377, 380, 380, 382, 387, 390, 389, 387, 384, 382, 380, 381, 382, 383, 383, 385, 387, 387, 387, 388, 377, 
    372, 375, 347, 312, 255, 202, 205, 247, 295, 337, 364, 378, 387, 392, 395, 395, 394, 390, 384, 379, 380, 382, 382, 380, 380, 381, 381, 381, 384, 372, 
    379, 400, 391, 365, 324, 254, 186, 161, 190, 254, 317, 360, 385, 394, 395, 392, 390, 387, 382, 377, 376, 378, 380, 380, 381, 379, 378, 377, 381, 369, 
    384, 403, 402, 400, 396, 366, 288, 188, 133, 152, 216, 282, 334, 370, 387, 390, 387, 383, 379, 375, 376, 378, 378, 380, 381, 380, 379, 379, 381, 370, 
    387, 407, 408, 407, 403, 401, 376, 277, 156, 109, 123, 166, 227, 285, 327, 354, 371, 377, 378, 375, 376, 379, 380, 381, 382, 382, 382, 381, 383, 373, 
    387, 406, 407, 407, 404, 398, 395, 338, 198, 106, 95, 98, 117, 161, 212, 256, 289, 317, 334, 345, 364, 381, 384, 383, 382, 380, 380, 380, 383, 372, 
    385, 401, 402, 404, 404, 401, 396, 341, 204, 94, 73, 78, 85, 94, 109, 135, 165, 195, 216, 235, 275, 318, 346, 362, 373, 379, 381, 381, 382, 371, 
    383, 399, 395, 398, 402, 402, 381, 301, 176, 73, 45, 58, 74, 87, 93, 91, 92, 95, 100, 110, 143, 196, 234, 262, 295, 324, 346, 364, 377, 369, 
    377, 398, 390, 395, 400, 397, 354, 278, 203, 119, 63, 48, 51, 70, 112, 150, 155, 124, 87, 80, 89, 97, 109, 151, 224, 283, 317, 345, 363, 360, 
    375, 397, 392, 394, 397, 394, 368, 328, 296, 251, 170, 122, 121, 146, 208, 261, 258, 211, 180, 192, 188, 165, 152, 182, 245, 286, 308, 333, 352, 354, 
    363, 385, 382, 379, 377, 377, 377, 358, 337, 331, 299, 252, 236, 239, 263, 305, 325, 306, 271, 267, 285, 281, 262, 256, 278, 310, 323, 326, 332, 334, 
    283, 302, 294, 288, 282, 278, 274, 270, 268, 271, 267, 247, 234, 239, 251, 270, 285, 291, 280, 267, 275, 286, 288, 279, 277, 285, 292, 296, 299, 296, 
    208, 226, 220, 216, 211, 208, 204, 199, 199, 197, 193, 192, 194, 205, 221, 231, 228, 225, 228, 231, 229, 229, 237, 245, 247, 244, 240, 232, 229, 230, 
    171, 184, 186, 181, 177, 170, 163, 160, 154, 150, 148, 145, 144, 145, 154, 166, 163, 157, 155, 154, 151, 151, 153, 157, 161, 163, 158, 147, 139, 145, 
    126, 138, 138, 136, 133, 125, 121, 119, 112, 107, 104, 101, 102, 104, 104, 106, 104, 95, 87, 86, 85, 84, 84, 84, 85, 85, 83, 76, 85, 120, 
    78, 85, 85, 86, 85, 78, 74, 72, 66, 60, 58, 61, 60, 61, 62, 65, 66, 57, 49, 46, 47, 49, 49, 46, 45, 46, 50, 70, 115, 139, 
    52, 52, 52, 52, 51, 50, 50, 50, 46, 41, 42, 44, 45, 45, 47, 51, 50, 48, 44, 42, 44, 45, 46, 45, 46, 56, 91, 133, 141, 120, 
    52, 52, 52, 52, 52, 51, 50, 50, 49, 52, 62, 67, 63, 60, 65, 67, 67, 65, 63, 58, 52, 48, 45, 47, 65, 108, 145, 137, 109, 96, 
    49, 47, 49, 49, 52, 52, 49, 48, 48, 57, 68, 70, 69, 66, 68, 73, 74, 73, 70, 62, 51, 48, 49, 71, 117, 144, 128, 104, 90, 69, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 29, 38, 13, 2, 9, 13, 15, 16, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 6, 3, 17, 
    0, 0, 0, 9, 5, 27, 56, 53, 65, 99, 118, 121, 118, 116, 101, 102, 113, 109, 107, 113, 109, 110, 85, 35, 2, 4, 13, 12, 7, 17, 
    0, 0, 0, 8, 16, 34, 16, 0, 0, 24, 17, 28, 36, 20, 10, 7, 13, 8, 8, 13, 13, 10, 0, 0, 0, 2, 0, 0, 0, 13, 
    0, 0, 0, 4, 28, 75, 69, 6, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 14, 1, 5, 6, 18, 
    0, 0, 0, 7, 43, 93, 91, 59, 63, 55, 41, 49, 46, 42, 50, 64, 75, 77, 88, 93, 80, 62, 68, 88, 82, 42, 20, 21, 19, 33, 
    0, 0, 0, 5, 18, 16, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 2, 6, 27, 22, 11, 2, 0, 0, 0, 0, 17, 17, 13, 29, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 5, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 3, 18, 
    0, 0, 0, 0, 0, 0, 9, 26, 18, 20, 27, 25, 18, 5, 7, 18, 28, 30, 29, 20, 13, 14, 0, 0, 0, 0, 0, 4, 3, 17, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 10, 8, 12, 7, 14, 
    0, 0, 13, 64, 83, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 2, 
    0, 20, 58, 116, 143, 154, 150, 100, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 16, 135, 208, 179, 109, 43, 6, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 9, 10, 11, 15, 19, 23, 21, 34, 
    0, 0, 0, 0, 0, 0, 0, 6, 122, 161, 126, 55, 3, 0, 0, 6, 10, 13, 15, 13, 9, 10, 13, 11, 9, 9, 12, 14, 11, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 136, 156, 121, 63, 23, 10, 12, 18, 18, 9, 2, 2, 2, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 66, 133, 194, 202, 156, 92, 42, 12, 5, 8, 8, 6, 6, 6, 7, 9, 5, 3, 0, 12, 
    0, 4, 0, 3, 2, 6, 8, 25, 22, 0, 7, 34, 78, 147, 210, 228, 202, 154, 109, 74, 36, 6, 0, 0, 2, 8, 9, 9, 6, 17, 
    0, 8, 7, 12, 10, 6, 7, 61, 118, 77, 44, 42, 23, 24, 60, 124, 190, 243, 275, 268, 219, 155, 97, 49, 17, 0, 0, 0, 0, 13, 
    0, 11, 10, 14, 10, 9, 41, 128, 166, 94, 58, 59, 33, 21, 7, 2, 22, 67, 130, 189, 220, 248, 262, 242, 195, 140, 85, 39, 11, 12, 
    0, 20, 14, 16, 14, 20, 67, 111, 46, 0, 0, 0, 31, 27, 0, 0, 0, 0, 0, 0, 0, 21, 130, 155, 110, 75, 70, 62, 40, 35, 
    0, 16, 9, 7, 7, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    7, 31, 33, 39, 45, 52, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 18, 26, 45, 
    164, 199, 206, 218, 227, 231, 235, 240, 242, 244, 232, 181, 132, 122, 115, 142, 176, 168, 130, 96, 112, 120, 101, 79, 88, 118, 133, 138, 134, 131, 
    120, 151, 153, 149, 144, 137, 133, 131, 127, 128, 128, 121, 116, 114, 113, 111, 108, 108, 115, 118, 118, 122, 128, 129, 119, 101, 98, 112, 129, 141, 
    3, 7, 8, 1, 2, 6, 8, 6, 5, 9, 12, 10, 12, 20, 38, 66, 85, 89, 95, 102, 107, 111, 115, 122, 127, 130, 135, 139, 138, 121, 
    98, 106, 108, 109, 109, 111, 111, 107, 107, 113, 115, 111, 107, 104, 102, 102, 106, 102, 103, 110, 107, 98, 93, 99, 105, 109, 111, 100, 56, 3, 
    75, 77, 86, 86, 84, 77, 63, 57, 59, 57, 51, 48, 43, 38, 36, 31, 31, 28, 22, 18, 15, 13, 14, 14, 12, 10, 0, 0, 0, 0, 
    16, 5, 15, 15, 13, 12, 6, 7, 13, 10, 2, 0, 0, 0, 0, 0, 3, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    14, 0, 4, 3, 4, 2, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 97, 
    13, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 82, 96, 45, 
    
    -- channel=53
    3, 0, 0, 0, 0, 0, 8, 8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 4, 30, 36, 33, 15, 11, 18, 14, 15, 13, 10, 7, 4, 3, 4, 6, 12, 1, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 8, 34, 52, 59, 62, 66, 70, 66, 65, 67, 62, 66, 66, 61, 63, 62, 62, 54, 25, 1, 1, 0, 1, 0, 0, 
    1, 0, 0, 0, 0, 3, 15, 19, 25, 36, 37, 38, 37, 41, 36, 25, 25, 21, 21, 23, 22, 14, 26, 13, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 7, 39, 50, 38, 21, 28, 25, 26, 37, 42, 35, 26, 18, 17, 16, 18, 20, 9, 30, 28, 14, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 47, 78, 57, 44, 45, 41, 41, 50, 50, 50, 50, 52, 52, 57, 59, 54, 44, 51, 55, 49, 21, 4, 4, 3, 3, 
    0, 0, 0, 0, 0, 10, 23, 17, 19, 17, 16, 15, 18, 18, 20, 17, 17, 19, 26, 27, 25, 26, 7, 13, 21, 5, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 2, 8, 19, 16, 21, 18, 18, 20, 20, 14, 9, 16, 17, 23, 24, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 12, 15, 17, 12, 10, 9, 13, 12, 12, 13, 14, 16, 15, 12, 8, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 20, 28, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 37, 70, 86, 72, 38, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 47, 97, 112, 84, 44, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 
    0, 0, 0, 0, 0, 0, 0, 52, 94, 94, 61, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 32, 88, 107, 93, 61, 27, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 93, 115, 125, 108, 74, 39, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 26, 59, 71, 96, 120, 131, 125, 103, 72, 47, 24, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 2, 0, 0, 0, 0, 0, 11, 50, 70, 65, 63, 68, 84, 108, 130, 141, 140, 129, 107, 76, 44, 20, 3, 0, 0, 0, 0, 0, 
    3, 1, 4, 0, 0, 0, 20, 19, 29, 62, 71, 75, 68, 58, 53, 52, 61, 81, 100, 125, 143, 150, 142, 122, 97, 64, 35, 13, 0, 0, 
    5, 1, 5, 1, 0, 4, 15, 2, 0, 0, 12, 47, 71, 61, 32, 0, 0, 2, 8, 20, 39, 70, 103, 104, 86, 61, 44, 32, 18, 6, 
    7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 
    14, 9, 12, 13, 17, 17, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 12, 12, 
    86, 90, 92, 96, 101, 104, 108, 110, 112, 107, 88, 79, 70, 67, 68, 68, 65, 55, 47, 44, 48, 43, 34, 32, 36, 42, 46, 48, 47, 44, 
    72, 73, 70, 68, 66, 67, 66, 65, 67, 66, 64, 64, 63, 65, 61, 55, 51, 52, 55, 55, 56, 58, 60, 55, 49, 44, 47, 54, 62, 65, 
    29, 29, 25, 20, 23, 28, 30, 33, 36, 34, 35, 37, 39, 45, 53, 59, 62, 67, 71, 73, 74, 78, 82, 83, 85, 85, 84, 89, 88, 78, 
    77, 86, 84, 79, 79, 81, 84, 87, 88, 90, 90, 88, 89, 87, 88, 85, 83, 85, 88, 90, 88, 85, 85, 87, 89, 90, 89, 86, 65, 50, 
    72, 82, 82, 81, 78, 74, 74, 73, 72, 72, 71, 70, 69, 69, 69, 67, 64, 62, 62, 63, 63, 62, 59, 59, 59, 57, 50, 32, 17, 20, 
    50, 58, 57, 58, 58, 57, 59, 58, 59, 57, 54, 52, 54, 55, 56, 57, 56, 56, 55, 54, 54, 57, 56, 56, 51, 36, 17, 14, 27, 46, 
    52, 56, 54, 54, 52, 53, 56, 57, 55, 47, 42, 36, 38, 40, 41, 39, 35, 36, 37, 42, 46, 52, 56, 50, 32, 15, 16, 33, 58, 75, 
    54, 58, 57, 55, 51, 52, 54, 55, 56, 53, 50, 45, 46, 49, 52, 50, 47, 44, 43, 46, 50, 55, 50, 36, 27, 31, 44, 63, 69, 66, 
    
    -- channel=54
    1, 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 25, 48, 39, 16, 11, 16, 14, 16, 8, 4, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 3, 1, 0, 
    0, 0, 0, 0, 0, 23, 54, 89, 103, 111, 131, 132, 128, 121, 116, 121, 122, 119, 120, 119, 114, 122, 85, 57, 22, 3, 8, 6, 4, 1, 
    2, 0, 0, 0, 0, 2, 0, 28, 44, 61, 69, 62, 60, 66, 65, 59, 53, 49, 48, 46, 45, 38, 32, 24, 4, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 10, 30, 52, 57, 20, 11, 8, 23, 27, 37, 24, 15, 0, 0, 0, 0, 5, 0, 21, 39, 34, 21, 2, 2, 2, 2, 
    0, 0, 0, 0, 28, 70, 111, 102, 71, 76, 65, 71, 69, 81, 87, 91, 88, 96, 101, 97, 104, 74, 103, 103, 87, 52, 14, 12, 13, 12, 
    0, 0, 0, 0, 5, 7, 39, 33, 35, 39, 26, 19, 19, 26, 36, 37, 45, 45, 54, 57, 49, 37, 28, 23, 30, 23, 10, 8, 9, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 6, 18, 15, 14, 9, 7, 2, 0, 0, 5, 15, 12, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 14, 14, 21, 18, 7, 3, 9, 16, 20, 21, 17, 14, 16, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 2, 4, 0, 0, 
    0, 0, 6, 41, 54, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 41, 77, 111, 131, 127, 82, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 48, 139, 179, 149, 91, 38, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 8, 11, 14, 14, 12, 
    0, 0, 0, 0, 0, 0, 0, 49, 135, 149, 107, 49, 6, 0, 0, 0, 4, 6, 5, 4, 5, 5, 3, 0, 0, 0, 2, 4, 3, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 115, 154, 148, 112, 61, 20, 5, 5, 7, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 119, 166, 192, 178, 134, 79, 34, 9, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 3, 0, 0, 0, 0, 44, 76, 127, 173, 201, 202, 175, 134, 97, 61, 29, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 1, 7, 5, 2, 0, 0, 8, 20, 45, 64, 56, 53, 70, 108, 153, 195, 224, 238, 227, 192, 141, 86, 43, 14, 0, 0, 0, 0, 0, 
    9, 4, 9, 7, 5, 0, 37, 58, 57, 61, 67, 70, 54, 39, 34, 39, 62, 102, 141, 184, 215, 232, 230, 207, 170, 119, 72, 35, 10, 0, 
    17, 10, 11, 11, 8, 14, 49, 24, 0, 0, 0, 11, 61, 48, 0, 0, 0, 0, 0, 0, 2, 71, 145, 152, 120, 79, 59, 52, 35, 18, 
    16, 4, 5, 6, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 9, 
    30, 21, 26, 33, 37, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 28, 32, 33, 
    161, 170, 176, 186, 191, 195, 200, 205, 208, 197, 158, 132, 118, 119, 132, 142, 138, 107, 90, 91, 97, 85, 70, 74, 87, 99, 105, 105, 102, 94, 
    120, 123, 124, 121, 114, 110, 108, 104, 104, 102, 99, 96, 94, 95, 92, 89, 85, 90, 95, 92, 96, 102, 106, 98, 86, 77, 82, 95, 112, 112, 
    20, 16, 12, 8, 7, 12, 15, 14, 19, 21, 22, 23, 28, 45, 62, 75, 81, 86, 93, 99, 103, 108, 113, 118, 121, 122, 125, 130, 131, 112, 
    100, 108, 110, 108, 108, 109, 107, 108, 107, 110, 112, 111, 108, 104, 106, 105, 102, 101, 105, 108, 104, 99, 99, 102, 106, 109, 106, 97, 61, 17, 
    79, 87, 91, 89, 82, 74, 69, 66, 64, 65, 61, 57, 55, 54, 51, 47, 42, 39, 37, 36, 34, 32, 32, 32, 32, 30, 13, 0, 0, 0, 
    27, 32, 35, 37, 34, 29, 29, 30, 30, 28, 23, 20, 19, 21, 21, 23, 24, 23, 17, 14, 13, 17, 17, 17, 12, 0, 0, 0, 0, 24, 
    25, 25, 25, 24, 22, 22, 24, 25, 22, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 17, 11, 0, 0, 0, 0, 61, 68, 
    25, 25, 23, 21, 18, 19, 20, 21, 19, 11, 11, 10, 11, 13, 16, 16, 11, 6, 6, 13, 18, 20, 9, 0, 0, 0, 26, 69, 58, 34, 
    
    -- channel=55
    37, 29, 25, 26, 33, 45, 45, 31, 23, 27, 35, 37, 38, 37, 40, 40, 38, 37, 37, 38, 38, 35, 37, 38, 39, 38, 33, 32, 32, 49, 
    32, 26, 23, 34, 42, 46, 35, 14, 18, 16, 18, 24, 23, 24, 21, 24, 28, 23, 25, 25, 22, 28, 26, 13, 20, 22, 19, 25, 27, 48, 
    34, 33, 28, 28, 34, 29, 5, 0, 7, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 8, 22, 24, 27, 24, 44, 
    33, 35, 31, 29, 35, 30, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 5, 14, 26, 28, 25, 20, 40, 
    37, 37, 32, 32, 40, 40, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 8, 1, 0, 0, 13, 27, 31, 27, 39, 
    34, 36, 33, 36, 34, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 24, 24, 22, 36, 
    32, 33, 30, 27, 21, 6, 0, 0, 0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 12, 30, 31, 24, 38, 
    29, 31, 29, 28, 36, 28, 0, 0, 7, 13, 10, 14, 24, 22, 12, 4, 4, 10, 9, 5, 10, 10, 16, 20, 0, 7, 27, 27, 23, 41, 
    31, 31, 30, 31, 39, 31, 19, 22, 29, 32, 31, 29, 36, 35, 27, 21, 23, 27, 31, 33, 32, 33, 34, 26, 11, 20, 30, 27, 22, 43, 
    36, 35, 35, 32, 32, 30, 31, 35, 38, 38, 37, 38, 36, 33, 27, 21, 25, 34, 40, 41, 41, 36, 28, 23, 23, 27, 30, 29, 27, 44, 
    38, 38, 34, 34, 34, 34, 37, 34, 33, 37, 35, 30, 27, 24, 23, 23, 25, 30, 35, 37, 35, 31, 23, 23, 28, 29, 31, 31, 29, 44, 
    39, 34, 26, 35, 48, 46, 37, 26, 24, 25, 25, 22, 19, 17, 17, 18, 20, 23, 26, 29, 28, 25, 24, 29, 32, 32, 32, 30, 26, 40, 
    40, 33, 32, 51, 64, 49, 43, 42, 33, 25, 21, 20, 20, 20, 20, 21, 24, 26, 25, 24, 25, 25, 25, 26, 26, 26, 25, 24, 21, 38, 
    40, 40, 45, 53, 67, 66, 57, 49, 40, 36, 32, 26, 23, 20, 19, 20, 23, 24, 25, 25, 25, 24, 25, 26, 27, 26, 26, 25, 23, 39, 
    39, 34, 29, 36, 58, 74, 73, 61, 49, 42, 40, 36, 28, 22, 21, 20, 20, 22, 25, 27, 28, 28, 28, 27, 27, 26, 27, 27, 24, 38, 
    38, 36, 32, 30, 37, 47, 62, 67, 58, 58, 53, 44, 45, 42, 34, 27, 23, 22, 23, 24, 23, 23, 23, 24, 25, 26, 29, 28, 24, 38, 
    39, 38, 34, 31, 34, 34, 42, 64, 65, 69, 80, 69, 56, 51, 50, 46, 39, 30, 23, 17, 17, 19, 20, 21, 23, 26, 29, 29, 25, 35, 
    39, 38, 34, 31, 34, 34, 37, 53, 64, 73, 85, 86, 82, 69, 56, 52, 53, 50, 42, 31, 26, 25, 25, 25, 26, 27, 29, 28, 23, 32, 
    38, 36, 33, 28, 31, 33, 35, 42, 62, 78, 81, 86, 86, 84, 80, 75, 69, 64, 58, 53, 47, 50, 51, 45, 41, 35, 29, 24, 18, 27, 
    34, 31, 29, 27, 28, 29, 29, 43, 80, 86, 79, 84, 81, 75, 78, 84, 90, 93, 85, 81, 74, 66, 61, 59, 58, 52, 43, 33, 24, 30, 
    34, 28, 26, 26, 29, 29, 35, 58, 79, 80, 66, 66, 79, 79, 85, 82, 69, 67, 78, 97, 86, 76, 80, 82, 75, 51, 33, 28, 26, 34, 
    33, 26, 25, 26, 29, 32, 45, 53, 42, 47, 64, 70, 71, 61, 40, 31, 38, 54, 56, 50, 55, 62, 61, 48, 29, 26, 23, 15, 15, 28, 
    33, 27, 22, 24, 29, 31, 31, 29, 28, 34, 47, 51, 40, 29, 14, 5, 11, 25, 27, 14, 14, 22, 22, 11, 0, 0, 0, 1, 6, 22, 
    39, 36, 29, 30, 35, 38, 40, 41, 44, 46, 47, 46, 42, 37, 32, 27, 23, 21, 21, 24, 22, 19, 17, 18, 18, 16, 13, 9, 10, 27, 
    60, 54, 50, 48, 52, 57, 61, 67, 69, 68, 68, 65, 60, 51, 44, 46, 49, 50, 51, 50, 49, 48, 49, 47, 46, 45, 43, 41, 39, 56, 
    67, 66, 58, 53, 54, 57, 66, 73, 76, 77, 75, 72, 72, 72, 70, 71, 76, 79, 79, 80, 81, 80, 78, 79, 79, 78, 80, 81, 84, 112, 
    79, 80, 76, 77, 82, 85, 90, 96, 99, 97, 93, 93, 95, 96, 98, 101, 105, 107, 106, 108, 108, 108, 106, 104, 102, 102, 106, 118, 135, 149, 
    95, 95, 94, 94, 96, 101, 104, 105, 108, 108, 103, 101, 104, 108, 110, 112, 111, 113, 115, 114, 114, 114, 113, 109, 105, 106, 122, 148, 145, 130, 
    96, 98, 97, 96, 97, 100, 102, 104, 106, 104, 102, 101, 101, 105, 108, 108, 107, 110, 110, 111, 110, 112, 114, 112, 116, 133, 145, 131, 115, 131, 
    98, 104, 106, 101, 97, 98, 100, 104, 107, 107, 103, 98, 101, 105, 107, 108, 106, 105, 103, 102, 103, 110, 116, 126, 143, 145, 125, 116, 129, 134, 
    
    -- channel=56
    29, 56, 66, 109, 105, 62, 48, 43, 39, 41, 50, 49, 53, 56, 41, 46, 50, 46, 45, 41, 46, 50, 45, 40, 26, 19, 27, 35, 35, 45, 
    47, 75, 75, 101, 104, 61, 33, 0, 0, 21, 22, 29, 32, 31, 18, 18, 29, 27, 27, 25, 32, 35, 29, 31, 38, 39, 38, 40, 40, 52, 
    50, 76, 74, 85, 80, 61, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 48, 39, 35, 37, 48, 
    50, 76, 82, 91, 75, 59, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 52, 43, 41, 41, 49, 
    46, 72, 84, 94, 71, 48, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 34, 43, 42, 40, 49, 
    52, 72, 83, 87, 66, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 45, 48, 43, 53, 
    61, 77, 81, 87, 76, 26, 0, 0, 0, 4, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 45, 56, 55, 60, 
    73, 85, 80, 92, 85, 57, 33, 26, 25, 33, 25, 25, 34, 20, 15, 18, 27, 24, 27, 9, 0, 7, 0, 24, 21, 29, 52, 59, 62, 68, 
    78, 93, 82, 93, 85, 83, 96, 86, 63, 65, 64, 63, 63, 57, 54, 55, 63, 68, 65, 52, 42, 42, 20, 34, 54, 58, 61, 64, 65, 71, 
    70, 94, 79, 97, 88, 85, 108, 104, 82, 88, 81, 79, 75, 71, 76, 78, 83, 84, 84, 72, 64, 63, 48, 48, 63, 63, 61, 62, 62, 68, 
    53, 91, 83, 101, 78, 42, 61, 90, 83, 83, 78, 71, 67, 66, 71, 76, 78, 76, 75, 70, 62, 64, 64, 60, 63, 62, 59, 60, 58, 64, 
    41, 101, 109, 113, 85, 16, 0, 26, 50, 69, 75, 71, 67, 65, 70, 73, 74, 73, 73, 70, 64, 64, 66, 64, 62, 60, 56, 56, 55, 60, 
    33, 101, 124, 125, 125, 84, 14, 0, 0, 12, 42, 57, 59, 61, 64, 65, 64, 65, 69, 64, 57, 59, 64, 62, 61, 60, 57, 56, 55, 63, 
    25, 80, 92, 95, 110, 136, 113, 55, 0, 0, 0, 11, 37, 53, 59, 58, 55, 55, 61, 59, 53, 56, 63, 64, 63, 65, 63, 63, 62, 71, 
    19, 67, 64, 63, 63, 89, 136, 154, 89, 0, 0, 0, 0, 11, 39, 53, 56, 56, 59, 57, 52, 55, 61, 61, 62, 68, 67, 68, 69, 77, 
    14, 56, 52, 56, 48, 43, 81, 178, 174, 58, 0, 0, 0, 0, 0, 10, 33, 47, 57, 58, 54, 56, 62, 61, 63, 68, 66, 68, 70, 78, 
    8, 43, 35, 45, 42, 40, 44, 145, 215, 93, 16, 17, 0, 0, 0, 0, 0, 0, 22, 38, 35, 47, 63, 64, 64, 67, 63, 63, 67, 75, 
    2, 37, 26, 36, 37, 39, 39, 129, 221, 108, 12, 19, 11, 8, 1, 0, 0, 0, 0, 1, 0, 0, 17, 31, 43, 55, 59, 62, 66, 75, 
    0, 37, 25, 32, 36, 37, 58, 141, 201, 119, 28, 11, 6, 9, 15, 23, 24, 29, 40, 32, 0, 0, 0, 0, 0, 3, 18, 35, 54, 70, 
    0, 40, 31, 34, 37, 41, 91, 142, 145, 133, 102, 49, 20, 1, 0, 11, 59, 92, 83, 55, 43, 25, 10, 0, 0, 0, 7, 14, 34, 59, 
    0, 45, 36, 38, 39, 46, 87, 115, 82, 114, 171, 118, 68, 31, 0, 0, 71, 132, 101, 44, 71, 96, 84, 11, 0, 13, 32, 29, 37, 59, 
    2, 44, 36, 36, 36, 37, 49, 61, 39, 58, 126, 117, 72, 51, 0, 1, 53, 104, 99, 43, 53, 87, 91, 54, 19, 36, 52, 48, 48, 64, 
    0, 29, 27, 26, 26, 24, 24, 26, 21, 28, 54, 59, 41, 32, 23, 39, 62, 71, 79, 65, 60, 64, 74, 77, 77, 80, 80, 73, 68, 74, 
    33, 53, 58, 61, 64, 61, 63, 64, 59, 64, 71, 70, 68, 61, 56, 75, 95, 89, 84, 88, 90, 84, 81, 88, 97, 101, 103, 95, 82, 74, 
    55, 58, 67, 72, 75, 70, 66, 62, 58, 59, 63, 66, 65, 64, 57, 61, 78, 75, 66, 67, 70, 68, 64, 63, 64, 66, 72, 71, 66, 45, 
    42, 33, 40, 47, 55, 54, 44, 37, 38, 39, 39, 41, 41, 42, 42, 36, 45, 50, 43, 40, 41, 41, 41, 42, 40, 40, 43, 46, 36, 18, 
    51, 29, 34, 36, 42, 42, 28, 24, 29, 33, 35, 36, 34, 31, 29, 25, 31, 39, 36, 31, 29, 28, 31, 33, 33, 35, 34, 26, 18, 27, 
    52, 28, 32, 30, 34, 33, 23, 23, 29, 31, 31, 30, 30, 25, 18, 20, 29, 33, 32, 29, 27, 28, 28, 29, 34, 35, 24, 20, 41, 47, 
    52, 32, 39, 34, 36, 35, 29, 30, 32, 29, 29, 36, 39, 32, 21, 25, 35, 37, 35, 37, 35, 27, 28, 28, 22, 20, 32, 52, 60, 42, 
    48, 25, 32, 30, 32, 34, 30, 27, 24, 12, 12, 24, 27, 22, 10, 12, 21, 23, 25, 36, 35, 21, 25, 19, 10, 26, 56, 68, 56, 23, 
    
    -- channel=57
    23, 8, 5, 5, 14, 26, 34, 34, 28, 21, 22, 24, 27, 29, 28, 25, 25, 27, 28, 28, 26, 26, 28, 26, 20, 13, 8, 11, 15, 22, 
    21, 12, 11, 3, 0, 6, 27, 42, 39, 28, 22, 22, 20, 21, 21, 17, 14, 14, 12, 10, 15, 16, 16, 10, 0, 0, 7, 15, 18, 24, 
    24, 18, 18, 12, 4, 5, 23, 41, 41, 44, 52, 57, 59, 55, 54, 51, 51, 54, 51, 46, 53, 56, 49, 34, 13, 13, 13, 14, 15, 22, 
    26, 22, 19, 14, 8, 0, 0, 0, 0, 19, 20, 22, 26, 20, 16, 10, 11, 14, 15, 11, 17, 17, 20, 16, 11, 16, 15, 14, 14, 19, 
    28, 23, 20, 19, 15, 14, 26, 13, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 20, 10, 10, 11, 17, 
    26, 22, 19, 19, 16, 23, 54, 47, 33, 26, 27, 30, 26, 24, 29, 33, 39, 36, 38, 47, 45, 37, 42, 45, 54, 38, 24, 21, 17, 20, 
    20, 19, 17, 12, 0, 0, 0, 0, 3, 0, 5, 5, 0, 0, 0, 0, 5, 4, 7, 13, 14, 11, 3, 11, 22, 17, 17, 20, 18, 21, 
    15, 16, 16, 12, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 12, 13, 14, 21, 
    13, 14, 16, 14, 12, 6, 10, 21, 31, 33, 35, 37, 37, 31, 27, 26, 27, 30, 33, 32, 35, 37, 22, 4, 0, 9, 14, 15, 14, 21, 
    13, 11, 12, 13, 15, 13, 10, 9, 8, 9, 9, 6, 1, 0, 0, 0, 7, 11, 10, 8, 8, 7, 8, 11, 12, 15, 16, 18, 17, 21, 
    18, 16, 17, 29, 39, 34, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 16, 16, 16, 16, 14, 19, 
    22, 22, 36, 64, 85, 83, 65, 40, 22, 12, 7, 6, 6, 6, 5, 5, 7, 9, 10, 12, 11, 10, 11, 13, 13, 13, 11, 10, 10, 17, 
    21, 11, 13, 27, 50, 81, 111, 112, 81, 46, 25, 14, 10, 8, 7, 7, 8, 7, 8, 10, 12, 12, 11, 12, 14, 16, 17, 18, 18, 23, 
    21, 2, 0, 0, 0, 0, 36, 84, 107, 96, 64, 32, 13, 6, 6, 10, 12, 14, 16, 18, 19, 19, 19, 19, 18, 18, 18, 18, 16, 21, 
    22, 11, 9, 10, 2, 0, 0, 6, 54, 92, 100, 83, 56, 33, 19, 14, 15, 15, 15, 14, 14, 13, 12, 12, 11, 10, 11, 12, 11, 17, 
    21, 14, 10, 12, 14, 10, 0, 2, 29, 72, 105, 120, 120, 97, 66, 40, 24, 18, 16, 15, 14, 14, 13, 12, 13, 14, 14, 14, 12, 15, 
    23, 19, 16, 15, 16, 18, 15, 16, 26, 55, 84, 96, 115, 131, 131, 114, 87, 62, 44, 30, 21, 13, 8, 10, 14, 17, 18, 18, 15, 16, 
    25, 23, 22, 21, 20, 18, 18, 28, 46, 71, 87, 86, 85, 91, 108, 130, 142, 138, 125, 104, 80, 57, 40, 30, 23, 19, 16, 14, 12, 15, 
    25, 20, 18, 18, 17, 14, 26, 45, 75, 96, 101, 99, 88, 77, 73, 78, 94, 115, 136, 150, 152, 146, 129, 106, 82, 57, 37, 24, 14, 11, 
    24, 18, 18, 19, 17, 18, 35, 53, 57, 48, 57, 76, 86, 80, 67, 49, 39, 47, 55, 70, 83, 109, 138, 142, 125, 96, 68, 47, 30, 21, 
    25, 15, 16, 18, 18, 20, 18, 10, 0, 0, 0, 5, 34, 32, 12, 0, 0, 0, 5, 3, 0, 0, 21, 27, 13, 1, 5, 16, 25, 26, 
    27, 17, 21, 24, 27, 26, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 21, 
    71, 67, 70, 77, 81, 86, 88, 90, 93, 92, 80, 61, 46, 41, 45, 55, 61, 52, 37, 31, 38, 36, 25, 19, 27, 40, 43, 42, 45, 47, 
    106, 104, 105, 106, 107, 108, 109, 110, 113, 113, 114, 114, 109, 101, 88, 78, 72, 75, 78, 78, 76, 75, 75, 71, 64, 57, 54, 58, 71, 79, 
    50, 43, 40, 36, 37, 40, 44, 47, 50, 52, 51, 47, 45, 48, 55, 64, 70, 74, 78, 79, 82, 85, 88, 89, 90, 90, 90, 93, 101, 104, 
    90, 89, 87, 85, 88, 94, 101, 106, 109, 111, 110, 110, 111, 111, 112, 114, 118, 119, 122, 125, 124, 122, 121, 122, 124, 125, 123, 121, 115, 108, 
    111, 114, 115, 114, 113, 113, 114, 114, 115, 114, 109, 107, 105, 105, 105, 105, 103, 101, 101, 102, 101, 98, 96, 96, 97, 96, 94, 91, 82, 74, 
    84, 86, 86, 86, 87, 89, 90, 90, 93, 92, 87, 86, 89, 92, 94, 95, 95, 97, 96, 94, 94, 96, 96, 95, 92, 87, 78, 72, 74, 93, 
    89, 91, 90, 89, 90, 90, 91, 94, 95, 90, 84, 79, 81, 84, 86, 86, 85, 86, 85, 86, 88, 94, 96, 91, 84, 77, 71, 79, 110, 134, 
    87, 91, 91, 86, 84, 85, 87, 91, 92, 85, 76, 71, 75, 80, 81, 79, 76, 73, 73, 78, 85, 94, 98, 95, 86, 78, 89, 118, 131, 117, 
    
    -- channel=58
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 9, 4, 0, 0, 0, 0, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 11, 10, 2, 0, 0, 0, 0, 0, 12, 22, 20, 15, 14, 15, 10, 9, 17, 14, 12, 18, 7, 19, 28, 0, 0, 0, 0, 0, 0, 
    18, 12, 13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 11, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    15, 11, 13, 1, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 4, 4, 2, 0, 0, 34, 21, 0, 0, 0, 0, 
    10, 8, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 4, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 2, 0, 0, 0, 0, 6, 5, 11, 10, 8, 2, 0, 2, 7, 7, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 20, 37, 37, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 35, 58, 82, 90, 61, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 63, 111, 104, 66, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 76, 100, 78, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 92, 91, 66, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 63, 83, 106, 104, 75, 38, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 35, 41, 61, 85, 106, 110, 97, 72, 47, 27, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 56, 49, 43, 41, 50, 71, 95, 117, 131, 133, 118, 83, 42, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 29, 48, 63, 67, 51, 39, 32, 28, 34, 51, 76, 106, 128, 134, 127, 117, 97, 67, 38, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 56, 51, 29, 0, 0, 0, 0, 16, 10, 36, 76, 95, 77, 39, 27, 24, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 6, 5, 
    82, 83, 81, 87, 91, 95, 98, 100, 104, 106, 99, 89, 76, 73, 70, 72, 78, 76, 67, 56, 60, 62, 56, 48, 49, 60, 64, 65, 64, 53, 
    67, 74, 70, 69, 67, 66, 65, 65, 65, 66, 68, 69, 69, 70, 71, 69, 66, 69, 73, 73, 74, 77, 81, 79, 75, 70, 66, 71, 82, 75, 
    30, 31, 29, 27, 26, 29, 31, 32, 33, 36, 39, 41, 44, 50, 55, 63, 68, 73, 79, 82, 84, 86, 89, 93, 94, 94, 92, 92, 102, 91, 
    71, 79, 77, 79, 79, 77, 78, 76, 74, 79, 83, 82, 81, 80, 80, 78, 76, 75, 78, 82, 82, 80, 77, 78, 81, 82, 81, 80, 77, 51, 
    58, 67, 66, 68, 67, 64, 60, 56, 53, 56, 58, 57, 55, 53, 53, 51, 49, 46, 45, 47, 47, 47, 46, 45, 46, 47, 44, 32, 12, 0, 
    38, 44, 43, 45, 43, 42, 42, 40, 40, 42, 43, 40, 36, 37, 37, 37, 38, 40, 40, 37, 35, 35, 36, 38, 40, 40, 22, 0, 5, 30, 
    37, 42, 40, 42, 40, 38, 38, 38, 38, 34, 27, 19, 19, 20, 20, 18, 17, 19, 18, 22, 27, 32, 35, 39, 35, 18, 2, 15, 49, 64, 
    33, 40, 40, 41, 39, 37, 36, 37, 36, 35, 33, 26, 26, 26, 27, 29, 27, 24, 23, 24, 29, 36, 37, 29, 16, 12, 34, 61, 69, 51, 
    
    -- channel=59
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=60
    223, 244, 243, 216, 200, 201, 202, 204, 213, 218, 218, 214, 210, 207, 210, 207, 206, 208, 211, 215, 215, 212, 213, 214, 222, 235, 241, 244, 249, 230, 
    235, 257, 260, 237, 215, 199, 185, 183, 200, 208, 207, 213, 202, 198, 206, 205, 204, 204, 203, 208, 213, 207, 208, 212, 231, 250, 250, 254, 259, 241, 
    234, 254, 262, 255, 242, 199, 157, 160, 186, 195, 201, 204, 191, 188, 200, 197, 199, 206, 204, 206, 210, 199, 213, 233, 246, 258, 253, 255, 257, 238, 
    235, 252, 262, 263, 250, 187, 133, 127, 129, 135, 141, 141, 135, 137, 148, 143, 151, 153, 157, 159, 161, 148, 182, 221, 242, 252, 254, 255, 257, 239, 
    233, 249, 258, 261, 247, 198, 165, 145, 132, 130, 135, 123, 120, 124, 136, 140, 143, 146, 147, 148, 148, 144, 178, 210, 237, 252, 260, 259, 262, 242, 
    229, 248, 254, 252, 230, 169, 153, 153, 158, 163, 168, 154, 149, 143, 161, 174, 186, 191, 184, 185, 184, 189, 198, 207, 237, 254, 261, 261, 266, 246, 
    224, 243, 251, 249, 209, 139, 119, 125, 153, 154, 156, 152, 146, 138, 147, 149, 160, 164, 154, 153, 157, 176, 156, 157, 203, 239, 256, 260, 264, 245, 
    221, 239, 251, 246, 213, 178, 152, 149, 171, 171, 180, 176, 179, 178, 176, 169, 169, 173, 160, 160, 167, 188, 174, 177, 197, 227, 251, 255, 258, 242, 
    222, 235, 248, 245, 241, 234, 209, 201, 205, 207, 211, 204, 208, 211, 213, 214, 217, 217, 207, 207, 207, 219, 236, 241, 232, 243, 256, 256, 258, 241, 
    229, 235, 244, 245, 251, 244, 216, 204, 201, 199, 196, 196, 199, 203, 203, 202, 203, 204, 202, 202, 201, 211, 243, 256, 252, 255, 257, 255, 259, 240, 
    237, 245, 255, 253, 253, 251, 233, 219, 216, 214, 215, 217, 221, 224, 222, 219, 216, 218, 220, 223, 223, 229, 242, 250, 253, 252, 250, 250, 256, 238, 
    245, 246, 240, 229, 237, 265, 276, 264, 252, 247, 247, 248, 251, 252, 252, 249, 246, 244, 244, 246, 248, 248, 247, 251, 254, 255, 254, 255, 261, 242, 
    247, 225, 193, 162, 151, 179, 226, 263, 274, 269, 258, 251, 252, 254, 254, 252, 251, 250, 247, 248, 252, 253, 253, 254, 256, 258, 259, 260, 263, 243, 
    254, 239, 218, 184, 135, 97, 106, 156, 217, 258, 269, 263, 258, 255, 255, 256, 258, 255, 250, 248, 251, 252, 252, 252, 253, 253, 252, 253, 257, 238, 
    261, 264, 260, 249, 220, 161, 99, 78, 116, 189, 246, 275, 279, 269, 259, 253, 253, 253, 249, 247, 248, 249, 248, 249, 250, 248, 248, 249, 254, 235, 
    264, 267, 264, 261, 260, 245, 184, 105, 72, 113, 170, 218, 264, 284, 281, 266, 254, 246, 243, 245, 248, 250, 250, 253, 254, 253, 252, 252, 254, 236, 
    265, 270, 270, 266, 264, 264, 237, 154, 75, 75, 102, 122, 165, 216, 255, 276, 278, 269, 258, 250, 251, 250, 246, 248, 250, 251, 253, 253, 256, 238, 
    264, 268, 269, 266, 265, 260, 256, 188, 93, 81, 92, 88, 96, 114, 144, 184, 221, 249, 260, 267, 280, 280, 267, 255, 249, 246, 247, 248, 251, 234, 
    260, 265, 267, 263, 265, 263, 264, 184, 86, 70, 76, 86, 89, 86, 86, 91, 105, 128, 146, 178, 226, 264, 278, 279, 279, 271, 261, 253, 252, 231, 
    259, 264, 264, 263, 265, 266, 238, 144, 64, 28, 30, 60, 82, 84, 83, 71, 60, 58, 46, 57, 91, 132, 166, 196, 226, 237, 246, 255, 259, 235, 
    258, 262, 260, 260, 263, 258, 196, 128, 91, 45, 6, 11, 33, 57, 98, 112, 89, 53, 43, 61, 52, 38, 43, 95, 152, 174, 194, 222, 243, 231, 
    258, 264, 264, 262, 266, 262, 230, 208, 202, 170, 105, 80, 77, 106, 168, 204, 193, 138, 128, 146, 145, 119, 103, 144, 192, 215, 224, 231, 242, 231, 
    270, 282, 278, 276, 278, 277, 277, 276, 278, 267, 237, 225, 217, 223, 241, 249, 248, 233, 228, 228, 233, 229, 223, 225, 230, 237, 242, 245, 249, 235, 
    201, 212, 203, 197, 194, 192, 189, 185, 187, 185, 180, 179, 181, 190, 198, 196, 192, 196, 199, 199, 201, 205, 211, 208, 201, 197, 197, 198, 208, 203, 
    129, 137, 131, 124, 124, 125, 122, 121, 122, 116, 115, 117, 120, 131, 146, 154, 151, 151, 155, 156, 156, 159, 165, 168, 171, 172, 165, 159, 163, 160, 
    136, 153, 149, 143, 142, 139, 139, 140, 135, 131, 130, 128, 129, 128, 131, 130, 123, 120, 119, 120, 116, 114, 116, 118, 121, 121, 116, 110, 107, 120, 
    96, 114, 110, 107, 104, 96, 95, 93, 87, 83, 82, 82, 83, 83, 84, 84, 79, 72, 67, 67, 68, 68, 65, 63, 64, 65, 64, 65, 87, 117, 
    55, 68, 64, 66, 65, 63, 66, 65, 60, 56, 55, 57, 58, 60, 62, 66, 64, 60, 57, 56, 58, 61, 58, 56, 57, 61, 71, 101, 137, 139, 
    54, 63, 60, 61, 59, 60, 64, 62, 58, 53, 55, 54, 53, 54, 59, 59, 53, 53, 53, 55, 57, 60, 62, 63, 65, 83, 119, 143, 138, 118, 
    51, 61, 60, 58, 56, 58, 58, 57, 57, 63, 70, 67, 64, 66, 72, 72, 68, 66, 64, 60, 57, 61, 63, 71, 98, 134, 146, 129, 102, 84, 
    
    -- channel=61
    188, 237, 250, 243, 223, 196, 186, 187, 197, 210, 212, 209, 203, 202, 196, 198, 200, 198, 199, 202, 206, 207, 205, 205, 213, 232, 250, 256, 254, 244, 
    191, 240, 254, 257, 244, 234, 205, 176, 189, 218, 233, 234, 229, 222, 216, 227, 228, 225, 230, 233, 230, 234, 218, 226, 249, 258, 264, 260, 257, 245, 
    195, 236, 247, 259, 259, 243, 187, 144, 163, 181, 185, 187, 182, 177, 179, 193, 198, 193, 200, 209, 196, 199, 191, 203, 252, 266, 263, 262, 261, 248, 
    191, 231, 239, 257, 263, 249, 206, 165, 177, 155, 144, 155, 144, 149, 148, 160, 161, 156, 162, 169, 157, 158, 166, 189, 243, 261, 260, 262, 265, 254, 
    188, 227, 235, 250, 265, 254, 207, 190, 209, 196, 192, 208, 189, 182, 191, 216, 222, 226, 233, 225, 223, 224, 230, 236, 245, 258, 267, 265, 265, 258, 
    187, 227, 231, 247, 257, 215, 157, 139, 181, 187, 178, 183, 171, 163, 172, 187, 196, 201, 206, 189, 188, 192, 200, 201, 190, 225, 261, 268, 268, 258, 
    193, 228, 231, 247, 245, 202, 159, 150, 166, 176, 173, 174, 174, 174, 177, 175, 174, 177, 175, 159, 159, 171, 178, 182, 177, 214, 249, 255, 258, 253, 
    203, 232, 232, 249, 249, 243, 241, 226, 214, 216, 216, 216, 209, 214, 222, 224, 229, 236, 227, 216, 213, 212, 224, 232, 231, 245, 258, 261, 260, 251, 
    212, 236, 230, 244, 247, 249, 243, 218, 197, 200, 195, 191, 190, 196, 207, 213, 216, 210, 203, 196, 191, 197, 221, 249, 260, 257, 259, 260, 260, 248, 
    219, 242, 232, 248, 247, 240, 230, 214, 200, 197, 195, 196, 201, 209, 215, 215, 211, 206, 203, 202, 201, 207, 228, 250, 260, 257, 255, 253, 254, 246, 
    224, 256, 248, 252, 234, 221, 234, 245, 244, 242, 241, 244, 250, 255, 259, 258, 254, 247, 243, 241, 243, 247, 250, 254, 257, 255, 253, 253, 256, 248, 
    225, 255, 232, 203, 177, 177, 200, 226, 239, 252, 259, 260, 263, 266, 269, 268, 263, 258, 255, 253, 254, 256, 256, 255, 255, 257, 260, 262, 263, 254, 
    227, 244, 208, 171, 130, 112, 115, 142, 183, 218, 242, 253, 260, 265, 269, 269, 267, 265, 264, 260, 259, 261, 262, 261, 260, 260, 261, 261, 261, 250, 
    232, 267, 253, 239, 193, 136, 95, 76, 94, 140, 189, 229, 254, 269, 273, 271, 268, 264, 259, 254, 251, 252, 253, 253, 253, 254, 254, 254, 256, 247, 
    234, 271, 264, 267, 252, 220, 174, 124, 76, 72, 121, 175, 216, 244, 260, 265, 265, 262, 257, 252, 251, 253, 254, 255, 257, 257, 255, 255, 257, 247, 
    236, 273, 265, 273, 266, 261, 236, 184, 109, 38, 38, 78, 126, 176, 214, 237, 248, 254, 256, 257, 255, 257, 258, 258, 259, 259, 257, 258, 258, 249, 
    237, 273, 265, 274, 270, 265, 257, 222, 145, 42, 3, 11, 27, 65, 113, 158, 192, 216, 233, 239, 242, 254, 262, 261, 259, 257, 254, 254, 256, 250, 
    234, 269, 260, 269, 267, 264, 265, 242, 161, 46, 0, 0, 0, 5, 19, 41, 72, 109, 143, 170, 192, 219, 238, 244, 245, 249, 251, 253, 256, 250, 
    233, 269, 260, 266, 268, 269, 276, 229, 118, 15, 0, 0, 0, 0, 3, 4, 3, 5, 11, 25, 53, 100, 147, 173, 196, 219, 234, 245, 255, 252, 
    232, 270, 262, 266, 268, 273, 256, 182, 72, 8, 0, 0, 0, 0, 0, 3, 26, 29, 0, 0, 0, 4, 15, 21, 60, 128, 178, 211, 236, 246, 
    229, 268, 264, 264, 265, 263, 230, 180, 136, 109, 71, 17, 0, 1, 41, 99, 128, 100, 56, 34, 46, 41, 20, 31, 86, 149, 186, 205, 223, 233, 
    225, 266, 266, 263, 261, 261, 255, 247, 244, 232, 195, 153, 129, 142, 177, 218, 234, 205, 179, 173, 185, 178, 165, 172, 201, 228, 242, 243, 240, 237, 
    199, 233, 233, 225, 219, 214, 211, 209, 206, 203, 197, 188, 184, 187, 196, 209, 215, 214, 212, 211, 212, 215, 218, 220, 219, 218, 222, 224, 222, 216, 
    93, 115, 115, 107, 100, 94, 89, 83, 80, 77, 74, 72, 77, 93, 112, 130, 139, 138, 138, 140, 143, 146, 152, 158, 163, 163, 169, 167, 160, 151, 
    77, 95, 101, 100, 100, 95, 87, 82, 77, 74, 72, 74, 76, 82, 90, 96, 96, 90, 86, 86, 84, 83, 83, 87, 90, 93, 92, 84, 68, 52, 
    51, 63, 70, 69, 65, 57, 43, 35, 28, 24, 19, 18, 18, 17, 18, 15, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 35, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 31, 6, 0, 0, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=63
    18, 6, 12, 16, 27, 42, 50, 49, 41, 42, 47, 55, 54, 55, 56, 58, 60, 58, 57, 57, 56, 56, 56, 58, 65, 68, 69, 66, 57, 71, 
    0, 0, 0, 0, 28, 79, 102, 97, 77, 69, 74, 76, 81, 79, 81, 84, 89, 89, 87, 85, 82, 83, 79, 69, 58, 47, 45, 43, 36, 51, 
    0, 0, 0, 0, 12, 82, 140, 143, 116, 98, 94, 94, 100, 107, 108, 105, 110, 101, 95, 99, 92, 92, 91, 54, 38, 36, 42, 48, 44, 59, 
    0, 0, 0, 0, 2, 104, 186, 199, 195, 181, 170, 169, 174, 184, 177, 172, 169, 162, 153, 157, 149, 153, 144, 88, 42, 34, 43, 47, 42, 59, 
    0, 0, 0, 0, 4, 107, 157, 165, 180, 193, 190, 200, 216, 213, 202, 193, 192, 191, 190, 188, 179, 185, 162, 116, 58, 33, 36, 39, 36, 57, 
    0, 0, 0, 0, 32, 143, 169, 147, 136, 137, 130, 145, 173, 173, 151, 129, 117, 115, 127, 123, 114, 118, 100, 91, 54, 24, 25, 28, 26, 45, 
    0, 0, 0, 0, 53, 176, 211, 189, 143, 137, 138, 142, 160, 173, 169, 156, 136, 142, 154, 156, 150, 137, 138, 148, 106, 45, 19, 16, 14, 35, 
    0, 0, 0, 0, 40, 121, 156, 142, 104, 101, 97, 93, 88, 103, 119, 123, 118, 123, 135, 141, 134, 105, 124, 138, 109, 53, 25, 23, 14, 30, 
    6, 0, 0, 0, 0, 19, 30, 29, 21, 21, 16, 16, 16, 24, 34, 30, 18, 17, 29, 38, 38, 25, 35, 50, 48, 25, 17, 17, 9, 26, 
    13, 0, 0, 0, 0, 0, 6, 20, 27, 27, 32, 35, 39, 44, 44, 40, 32, 30, 33, 43, 48, 41, 26, 17, 17, 14, 14, 13, 8, 30, 
    19, 0, 0, 0, 0, 0, 13, 33, 39, 40, 42, 46, 47, 48, 49, 50, 48, 41, 38, 40, 47, 43, 26, 15, 14, 19, 24, 26, 21, 41, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 14, 14, 16, 17, 20, 21, 20, 19, 19, 21, 23, 22, 18, 17, 20, 25, 26, 21, 40, 
    30, 18, 28, 43, 43, 12, 0, 0, 0, 0, 0, 14, 21, 23, 24, 26, 28, 29, 27, 24, 22, 20, 18, 16, 14, 12, 14, 15, 11, 31, 
    30, 31, 50, 77, 113, 124, 94, 28, 0, 0, 0, 0, 25, 32, 31, 29, 28, 28, 28, 28, 26, 22, 17, 15, 16, 15, 16, 14, 8, 27, 
    28, 19, 24, 33, 71, 121, 145, 119, 48, 0, 0, 0, 0, 11, 28, 32, 30, 28, 28, 30, 31, 29, 25, 23, 22, 20, 20, 17, 8, 25, 
    32, 26, 33, 32, 41, 65, 100, 109, 86, 37, 0, 0, 0, 0, 0, 8, 27, 36, 35, 30, 26, 24, 23, 19, 16, 15, 16, 14, 7, 24, 
    37, 34, 41, 39, 43, 46, 67, 83, 82, 72, 53, 37, 4, 0, 0, 0, 0, 0, 0, 6, 15, 25, 31, 28, 22, 16, 15, 15, 8, 24, 
    45, 42, 48, 44, 45, 50, 56, 59, 52, 46, 48, 58, 58, 46, 22, 0, 0, 0, 0, 0, 0, 0, 0, 19, 27, 27, 28, 25, 16, 30, 
    49, 45, 51, 45, 43, 48, 38, 33, 34, 33, 35, 41, 57, 73, 78, 70, 47, 14, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 19, 35, 
    46, 41, 48, 44, 40, 40, 27, 51, 86, 105, 93, 57, 44, 60, 89, 122, 131, 107, 84, 66, 48, 11, 0, 0, 0, 1, 9, 13, 13, 29, 
    42, 37, 46, 44, 42, 42, 68, 115, 166, 185, 166, 142, 120, 130, 151, 164, 166, 148, 147, 146, 150, 148, 133, 123, 110, 95, 78, 57, 33, 32, 
    34, 26, 33, 32, 26, 29, 57, 81, 98, 111, 126, 144, 158, 146, 118, 84, 71, 91, 104, 107, 105, 116, 130, 109, 74, 42, 26, 23, 11, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 30, 36, 38, 37, 36, 40, 44, 44, 41, 37, 32, 26, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 2, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 12, 
    26, 10, 14, 15, 16, 22, 30, 37, 41, 38, 35, 33, 35, 39, 40, 45, 49, 52, 54, 54, 55, 57, 58, 58, 57, 55, 58, 66, 65, 55, 
    76, 62, 64, 62, 61, 65, 67, 71, 74, 72, 70, 69, 71, 73, 75, 72, 68, 67, 69, 71, 72, 70, 73, 74, 68, 60, 65, 65, 31, 13, 
    77, 61, 63, 63, 62, 64, 65, 66, 68, 74, 79, 82, 82, 84, 87, 87, 87, 84, 85, 81, 76, 73, 73, 69, 65, 62, 47, 14, 0, 10, 
    84, 68, 68, 70, 70, 71, 73, 75, 79, 85, 84, 86, 86, 87, 88, 89, 91, 91, 90, 85, 81, 77, 72, 69, 64, 38, 0, 0, 15, 56, 
    
    -- channel=64
    72, 69, 47, 22, 38, 54, 43, 45, 41, 3, 0, 34, 57, 57, 48, 60, 97, 108, 101, 105, 105, 82, 63, 115, 162, 97, 36, 65, 63, 54, 
    88, 80, 62, 42, 71, 66, 50, 54, 43, 0, 0, 37, 57, 54, 42, 67, 107, 106, 92, 100, 107, 78, 62, 127, 180, 108, 37, 65, 76, 74, 
    100, 95, 86, 65, 84, 64, 55, 61, 41, 0, 0, 22, 44, 45, 40, 69, 99, 91, 79, 94, 105, 78, 62, 138, 195, 125, 58, 82, 104, 105, 
    89, 99, 86, 80, 77, 57, 57, 59, 37, 0, 3, 24, 45, 52, 55, 76, 97, 89, 76, 84, 91, 82, 75, 139, 201, 153, 95, 113, 129, 120, 
    81, 94, 72, 78, 71, 60, 56, 52, 31, 0, 18, 53, 73, 77, 77, 70, 67, 71, 80, 62, 77, 95, 91, 140, 214, 185, 125, 129, 131, 121, 
    75, 71, 59, 81, 75, 67, 52, 46, 24, 8, 50, 102, 113, 104, 83, 45, 37, 64, 79, 42, 74, 122, 104, 151, 214, 196, 139, 132, 135, 126, 
    76, 50, 60, 99, 102, 87, 57, 54, 32, 29, 96, 139, 134, 119, 73, 31, 36, 90, 83, 46, 108, 152, 140, 167, 209, 190, 148, 137, 142, 109, 
    73, 44, 71, 129, 124, 102, 71, 61, 46, 69, 138, 150, 135, 101, 42, 32, 78, 115, 105, 96, 143, 163, 168, 168, 204, 185, 153, 143, 140, 78, 
    74, 46, 83, 151, 154, 112, 80, 66, 54, 100, 145, 146, 138, 89, 41, 73, 132, 136, 128, 150, 164, 169, 163, 160, 201, 175, 149, 148, 135, 58, 
    84, 43, 82, 149, 171, 141, 98, 72, 81, 132, 141, 138, 133, 89, 90, 141, 167, 161, 154, 164, 171, 168, 145, 169, 206, 168, 148, 154, 131, 48, 
    80, 32, 70, 137, 159, 170, 137, 98, 122, 156, 145, 141, 127, 98, 116, 155, 169, 168, 165, 161, 176, 153, 131, 174, 205, 167, 144, 148, 137, 57, 
    87, 40, 72, 123, 146, 169, 165, 138, 155, 162, 158, 159, 142, 133, 150, 157, 158, 161, 161, 159, 164, 152, 154, 186, 201, 169, 147, 154, 150, 69, 
    93, 50, 78, 112, 133, 150, 177, 176, 170, 161, 162, 172, 166, 151, 162, 168, 158, 154, 148, 151, 151, 157, 172, 186, 197, 159, 145, 160, 146, 69, 
    98, 66, 81, 113, 121, 141, 176, 195, 181, 178, 158, 144, 165, 175, 174, 175, 176, 168, 162, 155, 152, 155, 173, 194, 191, 166, 147, 157, 129, 65, 
    100, 82, 93, 120, 123, 145, 165, 180, 179, 178, 157, 127, 161, 187, 188, 189, 190, 186, 189, 187, 174, 163, 172, 190, 195, 179, 150, 149, 123, 59, 
    101, 92, 108, 115, 127, 131, 156, 154, 183, 195, 159, 137, 157, 176, 191, 201, 199, 194, 186, 190, 182, 172, 177, 180, 199, 165, 160, 148, 106, 42, 
    108, 110, 125, 131, 129, 119, 142, 137, 152, 189, 165, 164, 163, 167, 191, 189, 197, 208, 209, 211, 212, 193, 173, 178, 183, 156, 131, 126, 97, 60, 
    115, 124, 134, 130, 110, 108, 114, 139, 133, 150, 168, 183, 180, 178, 191, 199, 203, 198, 202, 202, 192, 193, 190, 183, 157, 148, 105, 103, 104, 76, 
    120, 130, 127, 121, 102, 91, 91, 126, 130, 111, 149, 164, 166, 184, 188, 203, 212, 205, 208, 211, 190, 188, 194, 183, 163, 126, 90, 91, 94, 107, 
    130, 128, 101, 116, 108, 77, 97, 116, 131, 114, 123, 145, 163, 190, 210, 211, 201, 210, 209, 197, 180, 182, 185, 178, 162, 118, 96, 87, 94, 139, 
    136, 103, 94, 125, 114, 81, 97, 117, 115, 139, 118, 123, 162, 203, 218, 218, 207, 205, 206, 193, 180, 189, 195, 185, 169, 141, 112, 97, 130, 151, 
    139, 109, 145, 188, 154, 110, 95, 116, 120, 129, 133, 121, 162, 213, 222, 216, 210, 200, 195, 186, 185, 190, 190, 195, 186, 158, 115, 124, 162, 156, 
    145, 148, 201, 235, 219, 164, 122, 125, 142, 122, 126, 150, 172, 210, 223, 221, 205, 201, 194, 180, 183, 203, 196, 199, 191, 157, 127, 136, 156, 151, 
    134, 162, 227, 264, 266, 231, 178, 155, 150, 126, 115, 160, 196, 200, 212, 203, 183, 186, 193, 185, 193, 203, 197, 190, 177, 157, 133, 127, 143, 146, 
    136, 163, 199, 241, 274, 268, 242, 212, 171, 137, 129, 146, 175, 183, 184, 163, 145, 164, 192, 185, 205, 204, 196, 178, 167, 141, 105, 104, 139, 146, 
    118, 123, 131, 179, 236, 266, 263, 257, 226, 178, 162, 171, 172, 178, 169, 137, 124, 146, 191, 202, 200, 207, 189, 163, 158, 127, 67, 94, 144, 136, 
    109, 90, 67, 113, 173, 234, 261, 268, 264, 237, 198, 186, 187, 183, 161, 134, 119, 145, 183, 199, 194, 201, 192, 165, 136, 90, 52, 112, 131, 145, 
    118, 97, 46, 56, 114, 179, 236, 268, 278, 273, 247, 218, 210, 198, 172, 151, 124, 142, 176, 182, 191, 199, 179, 156, 124, 57, 67, 114, 120, 172, 
    116, 97, 48, 40, 61, 132, 190, 239, 266, 274, 266, 253, 240, 224, 213, 198, 164, 138, 139, 149, 149, 161, 159, 150, 129, 94, 115, 122, 162, 219, 
    103, 70, 66, 70, 43, 75, 141, 198, 243, 256, 257, 263, 263, 245, 238, 239, 214, 164, 137, 135, 130, 144, 153, 161, 159, 140, 137, 140, 190, 233, 
    
    -- channel=65
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=66
    0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 15, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 1, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 1, 14, 3, 0, 0, 0, 0, 0, 12, 0, 0, 16, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 15, 25, 0, 0, 0, 0, 0, 15, 17, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 11, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 7, 34, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 1, 0, 0, 0, 0, 0, 17, 0, 7, 14, 15, 16, 0, 0, 0, 0, 0, 4, 11, 10, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 1, 0, 0, 0, 0, 0, 0, 0, 4, 8, 13, 23, 23, 9, 2, 0, 0, 0, 0, 14, 20, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 5, 10, 11, 17, 23, 21, 14, 3, 0, 0, 0, 12, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 7, 7, 13, 3, 1, 5, 13, 26, 25, 22, 13, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 41, 15, 8, 12, 5, 0, 0, 0, 1, 5, 21, 12, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 20, 0, 0, 0, 11, 14, 3, 0, 0, 0, 10, 2, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 0, 1, 0, 2, 2, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 3, 1, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 10, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 3, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 5, 3, 5, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 9, 0, 24, 0, 
    0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 6, 0, 
    
    -- channel=67
    93, 63, 32, 44, 63, 70, 79, 71, 28, 0, 13, 56, 69, 53, 58, 87, 101, 98, 105, 123, 107, 77, 108, 167, 123, 36, 32, 65, 78, 74, 
    110, 87, 58, 69, 84, 86, 91, 74, 23, 0, 8, 49, 61, 39, 50, 92, 103, 90, 101, 122, 104, 76, 111, 177, 139, 53, 58, 98, 102, 76, 
    126, 117, 87, 87, 95, 97, 98, 73, 18, 0, 0, 25, 42, 42, 58, 97, 115, 99, 97, 112, 103, 79, 118, 192, 178, 107, 99, 128, 127, 101, 
    133, 118, 95, 91, 99, 98, 93, 67, 10, 0, 0, 26, 55, 74, 76, 94, 116, 109, 85, 90, 99, 91, 132, 213, 216, 148, 128, 154, 163, 150, 
    101, 86, 86, 90, 103, 92, 78, 54, 6, 0, 28, 69, 92, 99, 89, 79, 96, 99, 56, 63, 107, 105, 143, 233, 242, 181, 160, 178, 185, 141, 
    67, 52, 82, 104, 103, 90, 65, 32, 6, 29, 79, 111, 121, 99, 51, 35, 81, 96, 56, 58, 109, 123, 158, 242, 258, 208, 188, 195, 173, 96, 
    65, 68, 108, 132, 114, 96, 70, 29, 24, 68, 113, 135, 121, 65, 19, 30, 75, 103, 91, 85, 126, 157, 173, 235, 260, 223, 203, 202, 160, 66, 
    76, 93, 154, 182, 139, 98, 79, 55, 59, 101, 144, 144, 92, 35, 29, 72, 93, 109, 130, 138, 156, 168, 175, 217, 244, 226, 210, 203, 140, 41, 
    82, 99, 175, 225, 191, 110, 66, 71, 92, 130, 161, 139, 88, 53, 67, 108, 137, 147, 150, 172, 172, 144, 158, 211, 229, 221, 218, 198, 120, 23, 
    81, 91, 173, 230, 232, 164, 70, 72, 117, 149, 163, 148, 121, 113, 128, 151, 173, 172, 166, 176, 161, 132, 159, 215, 220, 220, 224, 199, 116, 7, 
    64, 76, 153, 213, 241, 216, 147, 119, 137, 156, 158, 145, 136, 151, 172, 183, 177, 168, 165, 157, 154, 152, 165, 209, 216, 210, 217, 202, 115, 6, 
    72, 73, 133, 190, 225, 245, 226, 175, 158, 160, 151, 136, 122, 140, 174, 177, 167, 165, 167, 156, 156, 154, 162, 207, 212, 194, 213, 206, 125, 47, 
    95, 87, 131, 165, 195, 238, 241, 200, 165, 146, 142, 150, 148, 142, 148, 154, 155, 157, 159, 160, 166, 170, 172, 189, 197, 195, 205, 201, 142, 81, 
    108, 104, 137, 155, 176, 219, 235, 220, 180, 136, 124, 141, 159, 166, 171, 173, 159, 147, 151, 155, 165, 195, 210, 196, 188, 189, 202, 191, 119, 63, 
    112, 111, 145, 174, 185, 208, 229, 240, 219, 142, 101, 135, 163, 180, 196, 192, 184, 180, 181, 176, 171, 194, 222, 239, 209, 178, 195, 165, 80, 64, 
    127, 128, 156, 187, 187, 197, 203, 209, 239, 210, 143, 146, 179, 191, 189, 194, 205, 205, 201, 200, 183, 174, 209, 246, 221, 182, 176, 157, 89, 68, 
    152, 161, 173, 172, 167, 176, 183, 180, 199, 244, 221, 167, 174, 196, 205, 208, 199, 204, 211, 209, 209, 202, 192, 194, 204, 167, 136, 145, 106, 80, 
    172, 185, 170, 146, 135, 141, 165, 178, 170, 198, 239, 207, 184, 202, 223, 228, 224, 226, 223, 201, 189, 203, 201, 187, 151, 116, 111, 115, 123, 143, 
    180, 161, 145, 140, 115, 117, 146, 160, 157, 143, 183, 219, 212, 225, 236, 229, 239, 246, 233, 214, 200, 201, 200, 186, 148, 118, 104, 96, 140, 188, 
    160, 134, 142, 135, 111, 115, 133, 131, 157, 149, 128, 187, 235, 249, 259, 252, 239, 238, 236, 216, 199, 196, 191, 176, 163, 136, 118, 145, 169, 187, 
    136, 122, 141, 137, 121, 113, 143, 149, 148, 175, 154, 159, 231, 266, 264, 269, 252, 228, 220, 206, 195, 196, 195, 180, 164, 137, 148, 192, 195, 190, 
    150, 153, 181, 184, 146, 118, 150, 188, 161, 155, 181, 187, 216, 259, 269, 255, 255, 239, 205, 202, 205, 197, 195, 184, 159, 146, 163, 187, 199, 202, 
    209, 241, 252, 235, 192, 152, 156, 186, 182, 149, 173, 214, 222, 240, 256, 243, 245, 242, 217, 210, 215, 208, 195, 172, 152, 148, 153, 175, 199, 201, 
    217, 248, 291, 292, 253, 211, 183, 173, 174, 178, 186, 216, 235, 229, 223, 214, 224, 235, 220, 224, 236, 211, 181, 164, 149, 115, 122, 169, 194, 190, 
    167, 193, 255, 300, 290, 255, 223, 198, 174, 177, 200, 207, 214, 198, 163, 149, 180, 223, 233, 224, 228, 217, 186, 173, 140, 81, 85, 154, 178, 152, 
    120, 101, 147, 226, 275, 280, 257, 239, 208, 172, 175, 195, 195, 171, 136, 116, 145, 207, 235, 222, 224, 221, 193, 160, 113, 68, 81, 137, 148, 135, 
    105, 41, 35, 117, 207, 268, 293, 271, 238, 210, 182, 179, 184, 181, 174, 144, 149, 195, 213, 223, 227, 206, 181, 137, 75, 67, 93, 114, 162, 171, 
    112, 51, 0, 28, 123, 213, 278, 301, 281, 248, 222, 204, 193, 194, 195, 175, 159, 178, 199, 210, 221, 202, 151, 106, 75, 71, 69, 121, 204, 202, 
    108, 66, 26, 0, 42, 138, 220, 284, 309, 290, 266, 247, 224, 206, 199, 183, 156, 151, 168, 167, 157, 153, 149, 138, 117, 97, 112, 159, 201, 222, 
    65, 53, 66, 33, 1, 48, 142, 223, 273, 297, 301, 287, 262, 251, 252, 221, 158, 131, 127, 110, 123, 156, 191, 209, 188, 172, 189, 193, 213, 231, 
    
    -- channel=68
    0, 0, 0, 0, 0, 0, 0, 0, 29, 7, 0, 0, 0, 0, 0, 0, 7, 53, 44, 17, 23, 17, 0, 0, 30, 55, 11, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 40, 42, 1, 0, 0, 4, 0, 0, 14, 8, 0, 0, 31, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 35, 9, 0, 32, 40, 5, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 11, 0, 0, 33, 39, 3, 0, 0, 0, 0, 0, 0, 16, 27, 34, 42, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    64, 87, 72, 5, 0, 0, 20, 53, 39, 0, 0, 0, 0, 0, 0, 38, 31, 18, 54, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    62, 52, 11, 0, 0, 0, 13, 46, 26, 0, 0, 0, 0, 2, 88, 99, 33, 1, 5, 0, 0, 0, 0, 0, 6, 2, 0, 0, 4, 113, 
    17, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 12, 93, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 28, 0, 0, 55, 132, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 66, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 33, 0, 9, 92, 121, 
    0, 0, 0, 0, 0, 0, 9, 17, 0, 0, 0, 4, 27, 0, 0, 0, 0, 0, 0, 0, 0, 49, 48, 0, 0, 8, 0, 20, 89, 93, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 19, 0, 0, 0, 0, 0, 0, 0, 0, 34, 41, 0, 0, 2, 12, 0, 14, 65, 61, 
    48, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 6, 5, 0, 0, 0, 0, 0, 6, 20, 30, 0, 0, 0, 17, 28, 11, 14, 54, 37, 
    17, 0, 0, 24, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 75, 52, 18, 0, 0, 0, 0, 0, 0, 37, 6, 0, 14, 43, 0, 
    0, 0, 0, 1, 14, 8, 0, 8, 28, 28, 8, 0, 0, 0, 0, 17, 31, 26, 18, 10, 0, 0, 0, 0, 45, 2, 0, 7, 44, 0, 
    10, 0, 0, 0, 0, 0, 12, 0, 0, 18, 73, 44, 3, 0, 0, 0, 0, 0, 6, 30, 30, 0, 0, 0, 0, 0, 0, 38, 105, 50, 
    19, 0, 0, 0, 0, 0, 14, 0, 0, 0, 14, 29, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 7, 57, 104, 20, 
    0, 0, 0, 0, 0, 0, 29, 44, 42, 14, 0, 0, 0, 0, 0, 12, 28, 12, 0, 0, 0, 0, 7, 50, 47, 11, 7, 47, 30, 0, 
    0, 0, 0, 0, 47, 60, 44, 36, 43, 53, 0, 0, 0, 23, 14, 0, 0, 0, 21, 30, 33, 7, 0, 30, 104, 126, 86, 62, 0, 0, 
    0, 0, 6, 38, 59, 44, 26, 0, 12, 53, 74, 1, 0, 0, 0, 0, 0, 0, 0, 4, 17, 18, 18, 18, 60, 100, 108, 67, 18, 0, 
    0, 37, 72, 55, 40, 5, 13, 20, 32, 32, 99, 113, 0, 0, 0, 0, 12, 4, 0, 21, 15, 0, 16, 27, 35, 7, 0, 0, 0, 0, 
    41, 72, 31, 0, 0, 0, 0, 28, 32, 9, 0, 60, 36, 0, 0, 0, 0, 20, 56, 38, 11, 14, 30, 32, 28, 2, 0, 0, 0, 0, 
    68, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 11, 51, 60, 25, 14, 21, 10, 3, 6, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 6, 28, 17, 28, 35, 18, 13, 5, 0, 0, 1, 5, 0, 0, 0, 5, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 3, 34, 38, 28, 31, 23, 0, 0, 0, 19, 38, 45, 31, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 1, 23, 52, 90, 61, 27, 7, 0, 0, 10, 36, 48, 38, 56, 62, 40, 1, 2, 
    88, 139, 140, 76, 0, 0, 0, 0, 0, 0, 0, 4, 26, 78, 133, 170, 118, 53, 8, 0, 18, 51, 19, 12, 35, 74, 48, 7, 16, 52, 
    71, 126, 159, 146, 94, 21, 0, 0, 0, 0, 0, 49, 58, 68, 91, 82, 44, 18, 18, 13, 10, 37, 30, 23, 81, 106, 0, 0, 35, 44, 
    25, 69, 111, 150, 131, 63, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 39, 16, 6, 47, 96, 128, 59, 0, 0, 0, 0, 
    2, 19, 2, 46, 96, 75, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 34, 28, 59, 68, 83, 77, 0, 0, 0, 0, 0, 
    39, 26, 0, 0, 28, 99, 79, 53, 21, 0, 0, 0, 0, 0, 0, 0, 45, 58, 77, 104, 127, 138, 79, 0, 0, 0, 0, 0, 0, 0, 
    110, 58, 0, 0, 0, 70, 116, 95, 84, 65, 0, 0, 0, 0, 0, 0, 0, 0, 74, 113, 100, 43, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=69
    31, 33, 35, 45, 35, 32, 40, 43, 46, 56, 63, 52, 49, 54, 61, 67, 68, 73, 74, 61, 51, 47, 60, 54, 36, 53, 75, 57, 45, 45, 
    32, 33, 32, 47, 33, 37, 39, 41, 45, 62, 72, 70, 70, 66, 68, 60, 49, 51, 59, 56, 46, 46, 63, 55, 23, 24, 38, 26, 29, 40, 
    27, 30, 31, 47, 36, 42, 39, 41, 49, 73, 78, 82, 67, 53, 57, 53, 41, 39, 49, 53, 50, 46, 58, 46, 6, 5, 23, 26, 27, 19, 
    54, 39, 50, 49, 44, 50, 46, 48, 52, 69, 66, 59, 42, 33, 42, 53, 55, 59, 72, 70, 60, 47, 51, 44, 9, 9, 33, 36, 21, 14, 
    85, 74, 78, 53, 44, 47, 54, 56, 53, 51, 41, 27, 23, 33, 52, 66, 59, 62, 65, 75, 63, 43, 47, 47, 15, 10, 28, 26, 33, 48, 
    70, 71, 69, 48, 41, 39, 52, 56, 52, 47, 35, 25, 42, 61, 77, 92, 79, 47, 32, 56, 53, 39, 58, 48, 21, 9, 20, 25, 45, 64, 
    39, 43, 26, 20, 35, 37, 44, 36, 41, 51, 37, 42, 66, 71, 72, 66, 69, 38, 23, 40, 27, 34, 56, 59, 38, 23, 29, 35, 42, 51, 
    30, 39, 25, 0, 16, 39, 48, 28, 27, 33, 30, 54, 66, 64, 54, 36, 26, 25, 32, 32, 23, 45, 54, 72, 44, 33, 34, 43, 42, 50, 
    38, 54, 48, 18, 0, 24, 56, 56, 52, 34, 32, 42, 33, 33, 39, 37, 27, 32, 39, 36, 53, 63, 75, 83, 40, 30, 33, 37, 37, 51, 
    43, 65, 58, 36, 4, 2, 25, 55, 71, 53, 56, 43, 2, 0, 0, 13, 33, 43, 47, 60, 63, 47, 63, 64, 38, 32, 31, 29, 28, 49, 
    51, 75, 71, 51, 30, 0, 0, 11, 31, 43, 63, 57, 42, 37, 24, 20, 31, 43, 49, 62, 49, 42, 48, 49, 47, 45, 38, 34, 23, 35, 
    38, 60, 64, 63, 48, 16, 0, 8, 15, 42, 58, 51, 55, 70, 74, 69, 55, 50, 48, 38, 28, 40, 54, 59, 48, 41, 41, 37, 13, 15, 
    21, 40, 43, 58, 52, 44, 29, 41, 57, 68, 68, 57, 40, 39, 47, 59, 64, 64, 66, 51, 39, 30, 38, 57, 42, 40, 36, 33, 23, 32, 
    41, 51, 47, 44, 54, 49, 37, 26, 46, 65, 79, 81, 66, 49, 34, 29, 34, 51, 63, 71, 66, 45, 28, 23, 38, 38, 39, 45, 58, 67, 
    47, 53, 47, 28, 38, 38, 48, 40, 22, 29, 55, 81, 66, 55, 58, 49, 35, 28, 21, 24, 47, 64, 48, 19, 22, 30, 39, 47, 53, 63, 
    29, 37, 34, 41, 35, 51, 52, 82, 57, 8, 9, 39, 50, 48, 49, 56, 64, 54, 51, 38, 35, 50, 63, 65, 30, 45, 36, 29, 33, 55, 
    24, 21, 29, 51, 57, 70, 57, 75, 89, 35, 14, 20, 52, 66, 45, 42, 43, 49, 58, 63, 56, 49, 56, 67, 78, 76, 69, 47, 28, 36, 
    27, 36, 46, 53, 69, 61, 64, 46, 78, 84, 58, 37, 38, 44, 48, 47, 35, 33, 36, 44, 57, 58, 57, 49, 74, 64, 83, 74, 35, 26, 
    42, 54, 67, 59, 61, 54, 71, 61, 54, 99, 98, 71, 44, 23, 30, 38, 46, 46, 40, 38, 50, 52, 53, 53, 40, 29, 36, 35, 39, 38, 
    55, 54, 63, 41, 38, 54, 50, 70, 54, 55, 76, 84, 63, 39, 31, 25, 44, 55, 54, 48, 54, 56, 58, 57, 40, 35, 15, 8, 22, 31, 
    47, 59, 54, 33, 35, 48, 33, 27, 47, 26, 35, 53, 62, 48, 39, 35, 34, 46, 60, 59, 58, 57, 52, 50, 47, 39, 24, 32, 25, 33, 
    18, 17, 12, 9, 25, 39, 44, 23, 30, 46, 43, 47, 53, 53, 53, 48, 40, 43, 44, 51, 52, 47, 49, 54, 50, 32, 34, 40, 36, 44, 
    0, 0, 0, 0, 0, 16, 36, 48, 34, 40, 52, 55, 56, 56, 61, 52, 44, 41, 41, 38, 41, 42, 58, 64, 63, 66, 57, 45, 38, 38, 
    50, 54, 30, 7, 0, 3, 21, 39, 45, 30, 27, 40, 52, 67, 72, 72, 62, 47, 38, 43, 40, 46, 59, 58, 63, 83, 76, 60, 45, 49, 
    106, 125, 109, 67, 21, 12, 21, 22, 36, 52, 51, 58, 70, 90, 101, 108, 100, 72, 40, 54, 51, 52, 44, 51, 58, 71, 72, 67, 61, 60, 
    85, 119, 147, 128, 84, 36, 18, 17, 23, 43, 66, 76, 85, 77, 69, 81, 87, 79, 56, 43, 53, 55, 48, 63, 72, 59, 68, 60, 53, 63, 
    51, 80, 136, 148, 132, 78, 33, 15, 16, 26, 40, 51, 64, 50, 21, 13, 43, 66, 67, 54, 50, 50, 67, 82, 74, 57, 77, 40, 28, 24, 
    37, 41, 78, 120, 132, 115, 72, 29, 4, 8, 18, 28, 41, 50, 50, 35, 51, 69, 67, 61, 61, 60, 67, 70, 54, 64, 60, 53, 52, 4, 
    53, 44, 49, 69, 117, 135, 121, 81, 35, 4, 0, 10, 20, 32, 42, 59, 79, 89, 94, 96, 103, 92, 63, 27, 7, 17, 1, 36, 52, 42, 
    72, 76, 55, 44, 83, 128, 141, 130, 97, 59, 25, 9, 6, 6, 0, 0, 33, 71, 94, 98, 91, 63, 28, 0, 0, 0, 0, 8, 25, 36, 
    
    -- channel=70
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 19, 33, 49, 46, 23, 13, 1, 0, 0, 7, 22, 46, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 20, 32, 44, 35, 20, 12, 6, 6, 8, 5, 5, 0, 1, 3, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 45, 59, 40, 4, 0, 0, 0, 0, 0, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 2, 8, 5, 6, 4, 16, 6, 25, 17, 3, 0, 0, 0, 3, 14, 18, 42, 42, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    77, 60, 62, 15, 0, 7, 19, 30, 5, 0, 0, 0, 0, 0, 4, 39, 28, 31, 44, 40, 10, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    60, 37, 27, 0, 0, 0, 17, 28, 0, 0, 0, 0, 0, 18, 69, 84, 41, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 76, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 21, 62, 51, 2, 0, 0, 0, 0, 0, 0, 0, 14, 19, 0, 0, 0, 43, 50, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 46, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 19, 2, 0, 19, 42, 31, 
    0, 0, 0, 0, 0, 0, 12, 2, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 1, 42, 43, 42, 7, 0, 0, 14, 26, 17, 
    0, 17, 20, 0, 0, 0, 0, 0, 9, 12, 21, 9, 0, 0, 0, 0, 0, 0, 0, 10, 34, 17, 0, 2, 4, 2, 0, 0, 0, 9, 
    23, 36, 44, 23, 0, 0, 0, 0, 0, 0, 12, 23, 0, 0, 0, 0, 0, 0, 12, 37, 16, 0, 0, 0, 17, 16, 7, 0, 0, 0, 
    0, 5, 33, 35, 16, 0, 0, 0, 0, 0, 8, 27, 37, 50, 68, 66, 49, 30, 13, 12, 0, 0, 11, 29, 26, 6, 0, 0, 0, 0, 
    0, 0, 0, 29, 21, 8, 0, 10, 33, 50, 50, 27, 0, 0, 22, 41, 46, 42, 50, 36, 15, 3, 9, 35, 23, 0, 0, 0, 0, 0, 
    0, 0, 3, 13, 16, 17, 10, 0, 8, 46, 77, 74, 38, 15, 0, 0, 0, 22, 46, 61, 52, 24, 0, 0, 8, 0, 7, 20, 38, 37, 
    4, 1, 0, 0, 0, 0, 13, 0, 0, 10, 31, 64, 49, 29, 27, 25, 7, 0, 0, 0, 6, 37, 39, 0, 0, 0, 19, 39, 39, 12, 
    0, 0, 0, 0, 0, 24, 29, 67, 35, 0, 0, 0, 14, 23, 36, 45, 42, 30, 28, 8, 10, 37, 47, 59, 34, 36, 16, 8, 0, 0, 
    0, 0, 0, 21, 35, 64, 29, 58, 79, 8, 0, 0, 30, 64, 34, 20, 25, 35, 51, 53, 36, 29, 43, 79, 88, 101, 86, 17, 0, 0, 
    0, 0, 12, 43, 51, 41, 31, 0, 62, 71, 59, 27, 11, 30, 25, 20, 13, 4, 7, 33, 48, 44, 46, 40, 86, 83, 92, 46, 0, 0, 
    1, 42, 55, 36, 32, 12, 41, 24, 35, 101, 102, 80, 22, 0, 5, 24, 31, 29, 34, 31, 32, 33, 41, 40, 34, 0, 0, 0, 0, 0, 
    43, 37, 26, 0, 0, 0, 15, 48, 6, 30, 54, 64, 51, 14, 8, 12, 33, 50, 59, 42, 41, 48, 54, 49, 16, 0, 0, 0, 0, 0, 
    37, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 33, 27, 17, 27, 48, 64, 57, 55, 45, 37, 28, 18, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 38, 47, 46, 39, 38, 37, 34, 30, 27, 29, 27, 26, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 1, 8, 36, 46, 60, 57, 47, 35, 22, 12, 19, 20, 48, 56, 54, 35, 30, 24, 0, 0, 
    0, 18, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 61, 85, 95, 74, 42, 23, 16, 22, 39, 58, 52, 52, 76, 71, 39, 0, 0, 
    116, 149, 127, 52, 0, 0, 0, 0, 0, 0, 6, 41, 57, 103, 145, 159, 127, 71, 24, 40, 48, 56, 33, 30, 48, 79, 55, 28, 17, 35, 
    81, 131, 170, 146, 76, 0, 0, 0, 0, 0, 22, 46, 70, 80, 83, 81, 69, 64, 45, 43, 47, 39, 34, 61, 85, 62, 26, 10, 21, 21, 
    19, 71, 152, 167, 139, 54, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 31, 70, 48, 39, 41, 61, 98, 98, 25, 26, 0, 0, 0, 
    0, 0, 48, 101, 128, 104, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 49, 67, 62, 55, 62, 78, 81, 30, 6, 34, 0, 0, 0, 
    18, 0, 0, 19, 99, 131, 112, 59, 0, 0, 0, 0, 0, 0, 0, 6, 49, 86, 109, 119, 145, 127, 60, 0, 0, 0, 0, 0, 0, 3, 
    67, 29, 0, 0, 50, 125, 141, 126, 84, 36, 0, 0, 0, 0, 0, 0, 0, 25, 101, 118, 102, 37, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=71
    140, 142, 146, 158, 155, 155, 164, 161, 155, 148, 157, 167, 159, 149, 154, 167, 167, 166, 167, 170, 166, 154, 157, 167, 161, 142, 145, 153, 154, 144, 
    143, 149, 152, 161, 158, 162, 164, 160, 154, 149, 152, 154, 152, 146, 154, 165, 163, 160, 167, 172, 167, 152, 153, 163, 161, 145, 150, 155, 149, 138, 
    141, 154, 156, 163, 158, 161, 157, 155, 151, 145, 142, 145, 146, 151, 158, 163, 167, 164, 162, 164, 168, 157, 150, 158, 165, 158, 152, 150, 149, 148, 
    147, 151, 153, 158, 155, 154, 147, 152, 149, 141, 142, 154, 161, 168, 161, 155, 163, 165, 158, 156, 171, 165, 150, 153, 161, 154, 151, 157, 165, 172, 
    142, 143, 157, 156, 154, 143, 136, 148, 148, 147, 163, 181, 185, 179, 168, 158, 157, 158, 144, 150, 178, 169, 146, 148, 150, 153, 162, 163, 169, 154, 
    145, 147, 165, 163, 149, 136, 131, 141, 146, 162, 187, 200, 205, 191, 163, 151, 158, 154, 139, 150, 168, 174, 165, 151, 146, 151, 163, 154, 143, 120, 
    161, 169, 167, 156, 145, 142, 137, 137, 150, 176, 193, 210, 212, 182, 163, 166, 163, 156, 154, 147, 157, 194, 192, 160, 152, 146, 151, 137, 130, 121, 
    165, 168, 166, 160, 144, 140, 144, 144, 152, 169, 189, 209, 192, 171, 176, 183, 167, 158, 177, 168, 172, 204, 197, 175, 155, 148, 142, 132, 132, 125, 
    158, 150, 153, 162, 158, 139, 137, 151, 159, 165, 178, 174, 159, 169, 177, 175, 182, 196, 193, 182, 188, 190, 190, 191, 159, 145, 140, 134, 137, 130, 
    147, 140, 147, 155, 162, 158, 137, 150, 175, 173, 165, 143, 136, 153, 156, 164, 194, 210, 193, 182, 181, 178, 190, 193, 163, 146, 140, 142, 147, 130, 
    135, 137, 143, 150, 160, 166, 164, 171, 181, 173, 148, 116, 114, 129, 133, 149, 167, 171, 163, 153, 160, 182, 177, 170, 165, 151, 147, 152, 150, 129, 
    141, 139, 139, 149, 155, 168, 180, 166, 154, 157, 131, 99, 92, 104, 116, 124, 129, 134, 125, 112, 117, 141, 142, 157, 163, 152, 159, 162, 150, 142, 
    150, 142, 141, 145, 145, 160, 159, 143, 126, 120, 105, 106, 109, 104, 100, 104, 107, 107, 97, 86, 87, 94, 104, 128, 144, 157, 162, 162, 158, 148, 
    151, 148, 143, 142, 142, 153, 145, 131, 110, 95, 97, 106, 109, 107, 100, 98, 93, 88, 88, 87, 84, 85, 86, 91, 116, 143, 150, 161, 153, 134, 
    153, 152, 151, 152, 147, 145, 150, 140, 113, 79, 79, 102, 97, 94, 101, 94, 89, 92, 92, 91, 86, 86, 78, 81, 96, 112, 137, 147, 140, 143, 
    155, 157, 157, 159, 144, 141, 145, 128, 111, 99, 86, 94, 92, 84, 75, 78, 94, 97, 92, 92, 87, 75, 77, 86, 80, 92, 120, 149, 156, 151, 
    151, 156, 153, 149, 139, 146, 151, 140, 106, 107, 100, 72, 73, 77, 76, 81, 75, 75, 82, 83, 95, 98, 79, 66, 81, 95, 104, 156, 164, 137, 
    144, 151, 146, 141, 144, 146, 156, 155, 124, 96, 98, 76, 68, 71, 76, 83, 79, 78, 80, 76, 80, 94, 90, 80, 79, 81, 118, 152, 168, 161, 
    141, 135, 137, 155, 155, 147, 158, 153, 143, 104, 95, 101, 80, 73, 71, 63, 74, 79, 68, 69, 83, 89, 89, 85, 89, 101, 129, 135, 162, 175, 
    135, 134, 156, 163, 157, 151, 150, 144, 159, 148, 103, 107, 98, 74, 73, 67, 65, 66, 74, 76, 76, 79, 85, 84, 99, 114, 123, 144, 156, 155, 
    137, 152, 164, 158, 164, 152, 150, 159, 157, 169, 146, 105, 101, 87, 70, 71, 67, 57, 71, 79, 76, 80, 89, 91, 103, 113, 127, 152, 156, 166, 
    149, 155, 158, 173, 177, 163, 159, 170, 157, 146, 160, 127, 93, 86, 81, 64, 64, 73, 71, 78, 85, 80, 84, 96, 111, 126, 133, 141, 166, 195, 
    163, 161, 151, 170, 193, 190, 175, 167, 160, 141, 139, 137, 101, 79, 79, 66, 63, 75, 81, 78, 76, 73, 81, 95, 116, 133, 130, 149, 190, 205, 
    151, 133, 139, 169, 199, 212, 198, 177, 166, 161, 139, 120, 110, 83, 71, 68, 71, 75, 73, 72, 76, 66, 71, 92, 113, 117, 127, 173, 202, 204, 
    135, 134, 150, 172, 189, 204, 211, 205, 191, 172, 157, 128, 109, 91, 71, 73, 81, 85, 77, 67, 64, 71, 75, 91, 101, 104, 132, 188, 204, 192, 
    146, 142, 155, 168, 181, 194, 202, 217, 220, 188, 167, 165, 147, 117, 101, 107, 110, 98, 79, 64, 67, 86, 83, 79, 86, 111, 152, 190, 192, 196, 
    154, 143, 145, 163, 184, 190, 197, 200, 211, 222, 211, 201, 195, 175, 162, 144, 123, 102, 74, 72, 83, 77, 80, 87, 93, 130, 173, 172, 193, 207, 
    158, 161, 153, 155, 180, 190, 186, 186, 192, 215, 230, 226, 222, 215, 202, 178, 137, 95, 76, 70, 79, 85, 82, 97, 128, 155, 154, 174, 220, 195, 
    166, 173, 176, 154, 157, 187, 191, 184, 184, 192, 205, 219, 223, 217, 204, 185, 157, 115, 92, 83, 75, 83, 105, 132, 149, 150, 159, 193, 191, 185, 
    159, 174, 195, 178, 151, 162, 192, 196, 190, 189, 188, 193, 205, 212, 211, 191, 159, 136, 118, 101, 104, 122, 141, 155, 152, 155, 173, 174, 163, 182, 
    
    -- channel=72
    31, 92, 61, 0, 17, 49, 45, 74, 116, 71, 0, 0, 30, 51, 0, 0, 0, 0, 0, 0, 55, 54, 0, 0, 101, 98, 0, 0, 21, 32, 
    32, 80, 43, 0, 27, 54, 44, 85, 117, 48, 0, 0, 31, 52, 0, 0, 16, 27, 0, 0, 59, 53, 0, 0, 105, 114, 0, 0, 33, 68, 
    27, 59, 39, 0, 40, 47, 43, 96, 115, 38, 0, 0, 24, 36, 0, 0, 18, 39, 0, 0, 51, 45, 0, 0, 83, 109, 0, 0, 45, 81, 
    15, 30, 33, 9, 45, 44, 43, 95, 114, 38, 0, 6, 14, 18, 4, 0, 15, 36, 22, 0, 18, 33, 0, 0, 50, 99, 0, 0, 30, 57, 
    30, 9, 3, 11, 40, 57, 51, 84, 103, 21, 0, 0, 6, 15, 33, 19, 0, 40, 71, 0, 0, 31, 0, 0, 33, 90, 13, 0, 17, 61, 
    63, 19, 0, 9, 31, 61, 68, 82, 72, 0, 0, 0, 0, 35, 67, 19, 0, 31, 102, 0, 0, 19, 0, 0, 16, 78, 13, 0, 48, 110, 
    72, 13, 0, 24, 48, 51, 62, 88, 36, 0, 0, 0, 11, 73, 66, 0, 0, 16, 66, 0, 0, 0, 0, 0, 0, 55, 5, 6, 95, 160, 
    68, 0, 0, 31, 88, 64, 29, 54, 0, 0, 0, 2, 57, 86, 15, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 34, 6, 28, 133, 168, 
    74, 0, 0, 5, 94, 114, 39, 0, 0, 0, 0, 23, 88, 72, 0, 0, 0, 8, 0, 0, 0, 3, 0, 0, 0, 22, 16, 55, 155, 158, 
    86, 0, 0, 0, 51, 134, 104, 0, 0, 0, 0, 2, 57, 21, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 17, 21, 64, 161, 158, 
    92, 0, 0, 0, 5, 89, 112, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 8, 24, 4, 48, 157, 152, 
    93, 0, 0, 0, 0, 22, 54, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 33, 0, 36, 145, 117, 
    82, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 34, 123, 74, 
    62, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 115, 30, 
    53, 0, 0, 3, 0, 0, 0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 89, 126, 0, 
    35, 4, 0, 0, 9, 0, 2, 0, 0, 29, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 91, 129, 0, 
    7, 0, 0, 18, 14, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 5, 34, 99, 0, 
    0, 0, 20, 32, 31, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 32, 13, 1, 21, 0, 
    17, 24, 21, 24, 51, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 58, 34, 21, 0, 0, 
    60, 31, 0, 23, 59, 0, 0, 17, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 54, 32, 11, 0, 0, 
    83, 12, 0, 14, 54, 9, 0, 37, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 10, 0, 9, 24, 
    51, 0, 0, 19, 54, 26, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 27, 
    0, 0, 0, 13, 42, 39, 0, 0, 30, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 14, 
    0, 0, 0, 0, 4, 26, 2, 4, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 
    0, 0, 0, 0, 0, 0, 0, 5, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 10, 21, 
    18, 0, 0, 0, 0, 0, 0, 0, 11, 2, 0, 0, 0, 0, 19, 4, 0, 0, 0, 0, 0, 0, 0, 0, 25, 53, 0, 0, 29, 13, 
    51, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 37, 0, 0, 0, 0, 0, 0, 0, 3, 58, 17, 0, 0, 0, 11, 
    57, 89, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 26, 56, 1, 0, 0, 0, 0, 
    61, 57, 38, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 50, 15, 2, 0, 0, 0, 
    68, 2, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 27, 0, 0, 0, 0, 0, 0, 0, 43, 17, 0, 0, 0, 0, 
    
    -- channel=73
    91, 96, 101, 105, 104, 105, 116, 115, 113, 118, 120, 113, 109, 110, 119, 128, 132, 139, 142, 132, 122, 117, 113, 113, 114, 121, 135, 126, 111, 101, 
    93, 100, 98, 109, 109, 113, 115, 112, 112, 119, 125, 127, 126, 125, 132, 132, 128, 130, 135, 128, 118, 116, 114, 114, 111, 103, 105, 93, 90, 96, 
    96, 103, 99, 114, 113, 113, 110, 111, 112, 122, 129, 137, 130, 122, 119, 114, 107, 104, 111, 121, 123, 114, 108, 107, 97, 80, 77, 85, 96, 99, 
    102, 99, 112, 122, 117, 111, 110, 115, 115, 124, 128, 129, 118, 106, 104, 117, 126, 124, 126, 133, 134, 115, 100, 98, 91, 79, 93, 107, 106, 92, 
    128, 129, 139, 126, 115, 109, 116, 122, 115, 114, 112, 107, 102, 107, 119, 128, 130, 129, 129, 141, 136, 111, 97, 97, 93, 92, 106, 105, 100, 96, 
    135, 140, 139, 118, 102, 101, 114, 120, 115, 110, 109, 112, 123, 134, 144, 154, 139, 115, 105, 118, 123, 115, 110, 98, 96, 92, 97, 93, 100, 117, 
    121, 119, 100, 92, 96, 98, 105, 109, 113, 117, 122, 138, 153, 152, 152, 144, 129, 108, 95, 97, 109, 127, 124, 114, 111, 97, 92, 93, 102, 112, 
    107, 105, 87, 72, 84, 97, 101, 92, 94, 109, 127, 145, 150, 146, 130, 104, 95, 105, 103, 93, 103, 133, 131, 130, 118, 106, 97, 98, 104, 108, 
    107, 111, 108, 90, 79, 89, 107, 108, 100, 100, 114, 125, 127, 122, 107, 101, 109, 115, 108, 110, 126, 148, 150, 144, 115, 102, 95, 97, 109, 110, 
    108, 117, 117, 106, 87, 79, 91, 123, 134, 120, 115, 107, 83, 69, 72, 99, 127, 130, 127, 134, 142, 148, 144, 135, 114, 102, 96, 97, 106, 104, 
    111, 122, 123, 115, 104, 80, 71, 93, 120, 122, 108, 95, 82, 70, 68, 89, 111, 118, 121, 130, 133, 128, 110, 115, 122, 112, 103, 103, 101, 97, 
    110, 117, 123, 126, 120, 97, 71, 69, 90, 101, 88, 82, 94, 113, 119, 113, 112, 105, 90, 84, 87, 101, 110, 128, 129, 119, 115, 108, 95, 85, 
    89, 97, 105, 118, 120, 116, 91, 87, 95, 95, 88, 85, 77, 78, 90, 103, 104, 93, 83, 70, 62, 65, 81, 113, 121, 116, 108, 105, 96, 82, 
    104, 106, 103, 108, 115, 117, 98, 79, 84, 91, 96, 95, 83, 71, 62, 61, 65, 78, 89, 91, 80, 66, 53, 66, 99, 113, 114, 112, 114, 114, 
    119, 118, 111, 102, 101, 104, 101, 68, 48, 61, 87, 103, 89, 81, 74, 61, 57, 58, 58, 66, 75, 80, 63, 49, 63, 91, 116, 117, 124, 130, 
    104, 107, 104, 100, 95, 106, 110, 104, 76, 53, 48, 64, 67, 63, 67, 78, 80, 65, 54, 49, 53, 71, 83, 75, 57, 85, 103, 113, 108, 102, 
    94, 93, 97, 111, 119, 132, 123, 117, 100, 66, 37, 32, 62, 72, 60, 60, 65, 75, 83, 87, 83, 73, 70, 84, 97, 104, 111, 118, 104, 95, 
    90, 93, 101, 116, 128, 129, 130, 110, 107, 90, 73, 54, 59, 69, 65, 59, 52, 51, 50, 59, 76, 83, 76, 73, 97, 116, 139, 135, 115, 87, 
    93, 106, 129, 134, 125, 118, 127, 112, 109, 113, 105, 87, 54, 40, 45, 53, 62, 58, 56, 62, 72, 77, 77, 75, 83, 91, 99, 110, 116, 96, 
    109, 122, 134, 120, 116, 114, 117, 131, 124, 113, 104, 107, 80, 50, 47, 47, 54, 61, 67, 65, 67, 72, 78, 81, 84, 83, 76, 81, 88, 103, 
    115, 124, 118, 106, 113, 111, 105, 107, 112, 102, 87, 80, 82, 64, 56, 54, 51, 61, 76, 75, 75, 79, 81, 81, 90, 101, 96, 89, 89, 116, 
    103, 96, 95, 103, 113, 117, 115, 96, 94, 105, 97, 74, 70, 72, 69, 61, 58, 61, 65, 72, 70, 64, 69, 78, 91, 98, 97, 104, 125, 142, 
    73, 47, 41, 74, 101, 112, 120, 120, 109, 111, 105, 85, 72, 72, 76, 70, 65, 64, 63, 58, 58, 59, 71, 91, 106, 105, 106, 122, 140, 141, 
    75, 72, 77, 88, 100, 106, 110, 123, 126, 105, 84, 74, 74, 73, 77, 80, 71, 64, 62, 56, 50, 54, 74, 94, 106, 120, 138, 147, 140, 140, 
    140, 157, 151, 127, 109, 113, 121, 121, 122, 115, 103, 89, 83, 90, 102, 116, 105, 82, 60, 58, 59, 69, 72, 79, 85, 115, 145, 154, 145, 148, 
    144, 171, 185, 169, 144, 122, 119, 124, 123, 125, 138, 142, 129, 116, 121, 124, 109, 90, 67, 61, 70, 72, 64, 75, 97, 118, 137, 143, 148, 156, 
    117, 145, 182, 196, 186, 149, 118, 112, 124, 131, 134, 139, 140, 121, 99, 83, 76, 75, 73, 70, 67, 69, 83, 100, 117, 128, 136, 125, 138, 129, 
    108, 121, 144, 176, 191, 170, 135, 113, 109, 119, 130, 133, 138, 133, 115, 95, 85, 82, 81, 76, 73, 76, 89, 112, 121, 122, 129, 138, 124, 88, 
    121, 118, 116, 127, 171, 189, 168, 136, 111, 103, 109, 118, 131, 139, 140, 136, 122, 107, 98, 90, 97, 107, 106, 98, 87, 94, 105, 121, 118, 119, 
    143, 149, 133, 112, 140, 185, 200, 183, 155, 132, 110, 102, 111, 113, 100, 95, 106, 121, 130, 130, 136, 122, 95, 68, 54, 59, 60, 73, 99, 122, 
    
    -- channel=74
    17, 16, 23, 29, 21, 28, 44, 43, 47, 60, 52, 34, 31, 36, 44, 39, 30, 45, 51, 40, 30, 34, 33, 4, 0, 29, 61, 44, 29, 26, 
    17, 21, 13, 22, 22, 36, 41, 38, 45, 59, 56, 52, 57, 55, 54, 39, 19, 25, 34, 29, 26, 32, 30, 2, 0, 7, 21, 4, 0, 17, 
    10, 12, 1, 23, 30, 41, 39, 37, 46, 64, 67, 71, 67, 49, 32, 28, 24, 18, 20, 25, 29, 32, 22, 0, 0, 0, 0, 0, 3, 7, 
    27, 27, 20, 33, 44, 44, 46, 48, 48, 62, 58, 50, 32, 19, 13, 22, 38, 39, 44, 55, 47, 24, 15, 0, 0, 0, 0, 12, 7, 0, 
    49, 60, 68, 43, 41, 36, 48, 59, 53, 50, 25, 1, 0, 2, 23, 54, 63, 44, 43, 66, 47, 12, 7, 0, 0, 0, 0, 1, 0, 10, 
    52, 57, 56, 27, 28, 31, 40, 55, 58, 37, 0, 0, 0, 23, 60, 89, 80, 48, 19, 35, 25, 4, 4, 0, 0, 0, 0, 0, 7, 36, 
    39, 34, 8, 0, 0, 28, 32, 25, 33, 21, 0, 0, 20, 46, 74, 61, 28, 25, 20, 0, 0, 0, 0, 0, 7, 0, 0, 6, 18, 44, 
    24, 31, 5, 0, 0, 4, 36, 20, 0, 0, 0, 8, 32, 58, 55, 8, 0, 0, 3, 0, 0, 0, 0, 8, 6, 5, 4, 11, 27, 53, 
    25, 40, 28, 0, 0, 0, 20, 46, 24, 0, 0, 7, 11, 22, 9, 0, 0, 0, 0, 0, 0, 16, 31, 25, 0, 5, 8, 10, 25, 51, 
    28, 49, 40, 14, 0, 0, 0, 23, 30, 7, 14, 13, 0, 0, 0, 0, 0, 0, 0, 2, 19, 20, 9, 0, 0, 13, 11, 4, 16, 40, 
    39, 59, 51, 32, 16, 0, 0, 0, 0, 0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 8, 7, 9, 0, 0, 0, 19, 25, 8, 9, 31, 
    23, 37, 41, 37, 34, 6, 0, 0, 0, 0, 0, 0, 0, 4, 21, 27, 17, 0, 0, 0, 0, 0, 0, 0, 7, 10, 16, 8, 3, 11, 
    5, 16, 20, 25, 32, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 4, 4, 7, 14, 
    21, 31, 27, 20, 21, 27, 0, 0, 0, 0, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 11, 12, 12, 35, 55, 
    28, 29, 30, 13, 1, 4, 6, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 20, 37, 52, 
    17, 6, 7, 14, 12, 17, 19, 10, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 8, 25, 15, 25, 
    9, 0, 0, 13, 36, 51, 32, 24, 9, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 38, 40, 46, 21, 2, 
    2, 1, 13, 30, 42, 50, 37, 16, 6, 13, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 31, 60, 51, 43, 3, 
    7, 22, 44, 43, 37, 38, 41, 25, 33, 16, 36, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 16, 20, 8, 
    21, 41, 44, 16, 21, 30, 29, 25, 37, 28, 0, 26, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 7, 2, 0, 0, 
    28, 36, 28, 1, 11, 27, 24, 8, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 10, 0, 7, 
    12, 0, 0, 0, 0, 7, 30, 16, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 15, 27, 
    0, 0, 0, 0, 0, 0, 0, 18, 23, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 27, 24, 24, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 26, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 9, 51, 53, 25, 24, 
    45, 61, 60, 12, 0, 0, 0, 0, 0, 0, 23, 6, 0, 1, 17, 48, 47, 12, 0, 0, 0, 0, 0, 0, 0, 18, 53, 55, 28, 38, 
    41, 58, 92, 76, 23, 0, 0, 0, 0, 0, 3, 26, 17, 12, 19, 25, 26, 9, 0, 0, 0, 0, 0, 0, 5, 44, 50, 32, 32, 36, 
    23, 39, 82, 101, 76, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 40, 51, 42, 25, 25, 0, 
    11, 19, 39, 62, 83, 50, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 32, 40, 37, 26, 15, 0, 
    25, 30, 26, 20, 55, 76, 48, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 29, 26, 26, 38, 41, 25, 0, 0, 0, 0, 0, 0, 0, 
    61, 65, 37, 10, 33, 69, 82, 50, 20, 5, 0, 0, 0, 0, 0, 0, 0, 0, 32, 45, 50, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=75
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=76
    77, 49, 36, 66, 78, 83, 100, 88, 41, 35, 73, 89, 84, 78, 98, 129, 133, 134, 142, 136, 104, 88, 145, 165, 75, 55, 92, 82, 83, 88, 
    97, 65, 58, 95, 91, 96, 107, 82, 35, 43, 84, 102, 95, 76, 102, 123, 111, 104, 126, 135, 97, 85, 154, 173, 66, 30, 71, 85, 93, 81, 
    104, 83, 83, 110, 97, 107, 112, 75, 33, 48, 74, 93, 81, 63, 99, 125, 109, 97, 118, 132, 97, 88, 156, 177, 76, 48, 95, 118, 107, 69, 
    131, 104, 106, 112, 104, 115, 114, 71, 31, 39, 53, 69, 68, 72, 100, 125, 126, 120, 126, 132, 105, 97, 159, 190, 116, 92, 129, 145, 119, 92, 
    141, 118, 122, 107, 106, 105, 104, 65, 28, 32, 54, 70, 86, 100, 111, 121, 125, 117, 94, 119, 118, 108, 164, 210, 152, 118, 140, 153, 146, 133, 
    102, 98, 111, 107, 105, 86, 84, 50, 33, 60, 93, 110, 127, 121, 102, 108, 131, 101, 46, 101, 127, 118, 181, 223, 172, 133, 148, 167, 153, 110, 
    67, 87, 104, 105, 103, 83, 68, 26, 41, 104, 130, 144, 146, 100, 61, 75, 121, 90, 51, 102, 121, 134, 190, 230, 192, 157, 166, 179, 127, 56, 
    68, 115, 145, 125, 95, 85, 75, 31, 60, 123, 139, 153, 119, 58, 49, 83, 103, 90, 99, 128, 134, 159, 188, 230, 193, 173, 174, 178, 100, 31, 
    84, 142, 188, 170, 110, 80, 83, 80, 115, 136, 142, 129, 64, 37, 80, 128, 120, 123, 141, 156, 166, 163, 190, 229, 183, 172, 179, 167, 74, 21, 
    83, 147, 197, 201, 147, 86, 61, 101, 155, 150, 148, 112, 44, 49, 99, 133, 146, 154, 162, 179, 167, 128, 176, 216, 178, 177, 184, 153, 55, 12, 
    74, 141, 195, 209, 191, 118, 60, 97, 136, 135, 138, 107, 88, 124, 137, 139, 147, 150, 150, 157, 130, 118, 174, 200, 177, 185, 189, 154, 50, 0, 
    60, 122, 172, 201, 212, 169, 123, 124, 120, 125, 125, 93, 95, 141, 163, 160, 145, 137, 129, 113, 99, 121, 171, 198, 173, 174, 190, 161, 50, 8, 
    65, 108, 145, 177, 201, 208, 181, 156, 135, 128, 118, 98, 87, 101, 115, 122, 124, 126, 129, 111, 109, 111, 135, 170, 157, 167, 189, 157, 73, 59, 
    97, 124, 146, 152, 185, 211, 189, 143, 120, 107, 117, 126, 121, 113, 100, 95, 95, 104, 118, 122, 133, 134, 130, 126, 136, 165, 184, 158, 103, 98, 
    109, 132, 151, 144, 172, 194, 194, 169, 125, 70, 84, 131, 132, 128, 137, 129, 107, 96, 94, 94, 117, 156, 162, 133, 123, 142, 173, 140, 76, 94, 
    106, 127, 149, 165, 173, 193, 192, 207, 179, 83, 59, 110, 129, 132, 135, 136, 144, 138, 135, 120, 116, 134, 168, 184, 133, 137, 151, 111, 50, 100, 
    123, 134, 156, 170, 173, 191, 178, 189, 199, 142, 106, 103, 135, 150, 134, 133, 136, 141, 152, 150, 142, 132, 151, 167, 157, 149, 142, 119, 70, 102, 
    148, 158, 168, 145, 153, 159, 172, 162, 178, 191, 176, 123, 123, 140, 148, 153, 137, 138, 139, 132, 143, 147, 145, 129, 133, 107, 129, 135, 103, 123, 
    167, 163, 159, 133, 129, 135, 169, 166, 153, 181, 194, 164, 139, 137, 152, 152, 158, 167, 151, 127, 139, 146, 139, 128, 91, 70, 92, 102, 132, 181, 
    160, 135, 141, 121, 103, 133, 146, 156, 151, 142, 150, 179, 180, 169, 165, 152, 162, 174, 160, 137, 141, 145, 136, 126, 95, 93, 87, 102, 155, 188, 
    122, 123, 143, 115, 101, 132, 133, 124, 151, 134, 122, 154, 192, 190, 174, 168, 161, 159, 156, 146, 141, 140, 128, 118, 109, 100, 111, 164, 179, 180, 
    93, 113, 132, 118, 105, 120, 152, 143, 149, 152, 148, 161, 186, 192, 184, 178, 165, 155, 137, 136, 137, 132, 127, 127, 109, 92, 138, 188, 187, 188, 
    117, 149, 144, 131, 111, 110, 152, 178, 149, 143, 161, 184, 182, 182, 183, 168, 165, 156, 136, 138, 139, 133, 138, 132, 113, 125, 161, 175, 185, 189, 
    199, 234, 216, 184, 146, 133, 150, 162, 147, 140, 160, 179, 179, 179, 174, 166, 170, 159, 137, 151, 151, 136, 128, 116, 111, 128, 157, 178, 191, 194, 
    223, 257, 270, 247, 198, 170, 168, 150, 143, 164, 188, 192, 184, 181, 161, 160, 180, 176, 146, 165, 160, 139, 112, 115, 104, 87, 132, 182, 195, 177, 
    158, 186, 251, 279, 251, 209, 183, 167, 153, 161, 186, 196, 191, 155, 115, 119, 161, 182, 165, 155, 155, 143, 122, 123, 95, 62, 125, 174, 169, 149, 
    103, 98, 168, 240, 269, 243, 213, 191, 168, 160, 163, 169, 175, 141, 98, 86, 131, 173, 169, 153, 156, 137, 133, 120, 71, 65, 142, 144, 138, 129, 
    87, 48, 69, 152, 229, 262, 251, 218, 183, 171, 167, 169, 172, 171, 161, 132, 146, 165, 155, 158, 165, 143, 122, 89, 49, 94, 123, 135, 187, 139, 
    97, 61, 40, 72, 164, 243, 273, 259, 226, 193, 179, 183, 177, 176, 173, 159, 158, 165, 162, 169, 172, 147, 115, 71, 52, 86, 76, 149, 217, 174, 
    93, 98, 77, 48, 92, 178, 252, 280, 271, 246, 220, 202, 183, 175, 160, 130, 110, 132, 146, 142, 138, 128, 126, 109, 96, 99, 108, 165, 197, 178, 
    
    -- channel=77
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 50, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 74, 37, 0, 0, 25, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 84, 57, 16, 28, 50, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 77, 70, 40, 51, 53, 0, 
    0, 0, 0, 15, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 58, 63, 51, 61, 45, 0, 
    0, 0, 0, 45, 37, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 49, 57, 58, 59, 26, 0, 
    0, 0, 0, 50, 52, 28, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 50, 52, 58, 57, 14, 0, 
    0, 0, 0, 39, 56, 43, 0, 0, 0, 0, 3, 14, 16, 13, 31, 29, 12, 3, 0, 0, 0, 0, 0, 20, 53, 47, 45, 52, 10, 0, 
    0, 0, 0, 23, 39, 54, 47, 22, 3, 5, 16, 11, 6, 8, 32, 38, 24, 17, 19, 17, 10, 0, 6, 22, 39, 27, 28, 45, 5, 0, 
    0, 0, 0, 15, 24, 46, 75, 62, 40, 23, 22, 18, 12, 10, 19, 16, 23, 33, 43, 50, 48, 37, 35, 37, 31, 18, 32, 44, 15, 0, 
    0, 0, 0, 6, 17, 32, 71, 56, 46, 46, 22, 15, 35, 38, 38, 40, 39, 35, 31, 45, 52, 59, 77, 67, 48, 19, 36, 52, 18, 0, 
    0, 0, 0, 1, 22, 36, 72, 86, 72, 68, 22, 0, 30, 50, 68, 75, 62, 49, 42, 39, 51, 73, 92, 98, 87, 44, 31, 42, 0, 0, 
    0, 0, 0, 24, 39, 47, 52, 80, 85, 67, 46, 24, 48, 70, 77, 75, 79, 84, 91, 86, 69, 66, 82, 116, 107, 69, 35, 12, 0, 0, 
    0, 0, 15, 29, 28, 19, 27, 38, 77, 75, 91, 90, 70, 81, 88, 81, 81, 80, 76, 84, 76, 72, 81, 86, 99, 67, 32, 0, 0, 0, 
    12, 34, 36, 15, 3, 0, 0, 11, 49, 82, 86, 103, 79, 68, 96, 105, 100, 100, 108, 99, 76, 72, 81, 73, 65, 20, 0, 0, 0, 0, 
    43, 40, 9, 0, 0, 0, 0, 19, 9, 52, 65, 71, 93, 98, 112, 120, 115, 114, 121, 107, 78, 74, 81, 75, 39, 2, 0, 0, 0, 4, 
    46, 0, 0, 0, 0, 0, 0, 1, 0, 0, 30, 37, 75, 120, 135, 128, 129, 130, 118, 106, 93, 83, 78, 67, 40, 22, 0, 0, 0, 29, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 31, 70, 119, 140, 140, 134, 128, 111, 90, 76, 74, 67, 57, 37, 13, 0, 15, 38, 32, 
    0, 0, 0, 0, 0, 0, 0, 5, 19, 23, 12, 38, 81, 116, 133, 140, 134, 125, 101, 81, 79, 81, 75, 61, 36, 1, 1, 27, 29, 11, 
    6, 33, 63, 54, 4, 0, 0, 15, 23, 4, 16, 47, 86, 110, 120, 125, 121, 117, 106, 83, 88, 100, 85, 58, 32, 14, 3, 14, 7, 0, 
    66, 96, 109, 89, 48, 8, 0, 0, 9, 0, 19, 71, 90, 109, 118, 114, 104, 108, 105, 101, 109, 119, 86, 41, 29, 13, 0, 0, 0, 3, 
    41, 52, 63, 86, 76, 44, 17, 0, 0, 9, 35, 75, 94, 98, 94, 67, 58, 83, 102, 119, 119, 104, 76, 56, 42, 0, 0, 0, 0, 0, 
    0, 0, 0, 29, 67, 60, 38, 20, 0, 0, 1, 19, 41, 42, 20, 2, 6, 54, 106, 108, 108, 101, 86, 70, 46, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 47, 60, 52, 28, 0, 0, 0, 0, 1, 0, 0, 20, 58, 98, 105, 98, 99, 86, 56, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 56, 73, 58, 29, 1, 0, 0, 0, 8, 20, 32, 57, 79, 90, 101, 99, 62, 11, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 13, 70, 86, 71, 47, 23, 7, 0, 0, 6, 18, 25, 61, 84, 81, 58, 16, 0, 0, 0, 0, 0, 0, 42, 
    0, 0, 0, 0, 0, 0, 0, 12, 64, 80, 82, 69, 47, 26, 15, 17, 12, 0, 9, 9, 0, 0, 1, 25, 28, 9, 6, 14, 40, 39, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    73, 68, 75, 76, 59, 38, 15, 10, 25, 37, 47, 60, 59, 48, 46, 48, 50, 41, 39, 46, 48, 47, 62, 89, 94, 64, 41, 61, 67, 51, 
    63, 65, 83, 68, 50, 28, 15, 16, 34, 41, 36, 36, 31, 32, 40, 53, 62, 58, 50, 50, 53, 53, 63, 94, 107, 95, 85, 93, 77, 51, 
    68, 75, 83, 56, 42, 24, 17, 20, 38, 36, 29, 20, 28, 47, 59, 63, 65, 66, 57, 50, 54, 58, 70, 104, 130, 122, 100, 82, 61, 67, 
    56, 63, 60, 43, 29, 17, 15, 19, 38, 40, 46, 46, 64, 74, 64, 46, 35, 33, 27, 32, 47, 64, 77, 108, 127, 103, 71, 56, 63, 93, 
    17, 33, 26, 42, 32, 23, 16, 17, 41, 63, 82, 93, 92, 73, 43, 17, 16, 22, 22, 30, 52, 69, 84, 102, 109, 85, 61, 63, 68, 56, 
    12, 32, 42, 59, 50, 43, 31, 27, 49, 81, 94, 94, 75, 42, 10, 0, 20, 35, 60, 60, 66, 78, 84, 96, 96, 84, 71, 67, 44, 21, 
    36, 57, 80, 86, 68, 61, 57, 67, 78, 82, 77, 69, 42, 25, 28, 47, 56, 65, 87, 98, 99, 93, 83, 87, 76, 72, 69, 53, 32, 30, 
    52, 55, 75, 88, 80, 72, 69, 97, 108, 89, 78, 57, 34, 44, 74, 103, 90, 93, 107, 110, 111, 82, 80, 74, 75, 63, 60, 40, 27, 35, 
    45, 38, 39, 63, 76, 74, 67, 80, 88, 88, 83, 69, 76, 90, 99, 92, 92, 97, 106, 106, 85, 50, 62, 72, 86, 64, 48, 33, 33, 42, 
    44, 29, 26, 37, 68, 78, 79, 73, 56, 72, 89, 107, 132, 143, 128, 104, 90, 86, 83, 80, 62, 63, 84, 96, 88, 56, 37, 42, 53, 53, 
    41, 23, 16, 21, 42, 76, 112, 111, 84, 96, 130, 144, 138, 120, 115, 110, 96, 98, 102, 90, 95, 100, 105, 111, 85, 45, 30, 49, 68, 69, 
    60, 41, 23, 17, 18, 57, 108, 127, 132, 143, 171, 178, 145, 109, 93, 92, 99, 121, 147, 147, 155, 133, 109, 98, 73, 45, 37, 51, 81, 99, 
    80, 63, 49, 29, 26, 31, 73, 113, 141, 151, 174, 193, 194, 177, 158, 144, 140, 148, 154, 162, 170, 171, 155, 120, 87, 59, 46, 53, 79, 90, 
    59, 51, 48, 41, 39, 30, 63, 137, 172, 166, 148, 158, 183, 192, 203, 210, 200, 182, 166, 152, 150, 166, 179, 166, 129, 74, 41, 40, 41, 44, 
    46, 46, 43, 58, 53, 49, 58, 137, 188, 183, 156, 143, 168, 188, 191, 196, 208, 216, 220, 202, 180, 154, 148, 175, 162, 113, 45, 26, 34, 55, 
    64, 62, 58, 54, 45, 36, 37, 74, 143, 174, 189, 179, 180, 189, 184, 182, 186, 194, 202, 207, 193, 168, 145, 134, 150, 122, 67, 42, 71, 78, 
    74, 71, 68, 38, 24, 6, 33, 50, 99, 155, 178, 195, 172, 161, 179, 189, 188, 183, 174, 175, 179, 177, 159, 123, 121, 79, 50, 46, 67, 80, 
    68, 63, 49, 35, 22, 20, 33, 64, 69, 104, 122, 166, 180, 165, 175, 182, 192, 199, 198, 181, 169, 167, 162, 155, 107, 73, 29, 32, 55, 86, 
    47, 32, 27, 34, 30, 43, 29, 52, 52, 58, 87, 117, 170, 190, 175, 177, 178, 176, 174, 175, 169, 168, 164, 159, 130, 104, 66, 55, 64, 58, 
    21, 32, 43, 57, 50, 48, 38, 34, 56, 49, 84, 106, 133, 171, 172, 172, 170, 165, 157, 164, 169, 166, 159, 153, 142, 98, 81, 86, 70, 41, 
    30, 56, 68, 82, 69, 45, 55, 57, 66, 73, 87, 128, 139, 154, 169, 170, 160, 157, 151, 150, 158, 170, 172, 171, 149, 99, 81, 63, 44, 25, 
    77, 112, 136, 131, 101, 66, 46, 62, 53, 62, 75, 119, 148, 160, 165, 160, 153, 145, 155, 168, 176, 184, 190, 183, 163, 137, 92, 36, 17, 11, 
    133, 173, 190, 176, 149, 112, 68, 43, 45, 46, 78, 109, 142, 169, 172, 162, 147, 143, 158, 174, 185, 191, 181, 165, 157, 138, 72, 24, 15, 16, 
    95, 108, 136, 155, 168, 149, 112, 70, 62, 67, 79, 120, 149, 168, 167, 142, 132, 146, 163, 178, 182, 183, 172, 165, 158, 113, 46, 10, 19, 13, 
    15, 17, 49, 104, 146, 155, 135, 114, 94, 82, 63, 78, 127, 133, 117, 88, 95, 134, 170, 168, 170, 167, 180, 177, 153, 101, 44, 9, 10, 4, 
    20, 7, 2, 32, 92, 131, 142, 144, 126, 96, 68, 59, 88, 110, 98, 81, 98, 136, 166, 159, 165, 171, 177, 157, 125, 85, 46, 17, 9, 29, 
    55, 36, 0, 0, 34, 99, 137, 150, 145, 127, 106, 99, 98, 122, 131, 127, 138, 150, 154, 164, 163, 174, 163, 123, 88, 78, 34, 32, 59, 93, 
    74, 75, 49, 29, 23, 58, 113, 144, 153, 148, 132, 119, 110, 109, 107, 109, 117, 142, 149, 150, 155, 154, 137, 110, 96, 66, 26, 65, 102, 133, 
    58, 79, 84, 71, 37, 25, 60, 109, 136, 147, 148, 136, 119, 108, 104, 104, 101, 107, 114, 107, 95, 100, 115, 132, 138, 98, 99, 105, 107, 111, 
    24, 44, 74, 91, 53, 21, 19, 50, 84, 107, 124, 136, 133, 140, 166, 180, 170, 130, 81, 66, 73, 101, 131, 150, 147, 138, 140, 117, 112, 100, 
    
    -- channel=80
    214, 163, 161, 178, 188, 181, 187, 198, 200, 196, 189, 186, 176, 160, 146, 140, 129, 95, 68, 67, 79, 85, 82, 84, 79, 79, 83, 97, 89, 71, 
    211, 201, 213, 214, 199, 183, 199, 205, 207, 209, 203, 198, 194, 181, 166, 163, 139, 103, 64, 55, 70, 81, 86, 86, 86, 95, 99, 103, 93, 82, 
    212, 221, 228, 225, 202, 194, 210, 210, 218, 218, 216, 214, 204, 191, 188, 186, 170, 122, 73, 53, 64, 79, 87, 88, 99, 111, 112, 107, 95, 88, 
    218, 224, 221, 227, 209, 209, 219, 218, 225, 227, 225, 227, 217, 202, 203, 199, 194, 154, 101, 74, 78, 97, 100, 96, 110, 116, 120, 112, 100, 102, 
    224, 206, 208, 227, 214, 219, 228, 225, 231, 237, 239, 233, 228, 215, 205, 207, 207, 189, 149, 116, 112, 122, 110, 95, 103, 111, 111, 110, 107, 109, 
    223, 179, 207, 225, 218, 222, 228, 231, 237, 243, 243, 235, 232, 221, 207, 208, 214, 211, 193, 159, 153, 148, 131, 108, 101, 103, 99, 105, 113, 113, 
    200, 179, 208, 221, 224, 223, 226, 233, 239, 245, 239, 236, 232, 220, 203, 194, 200, 206, 212, 202, 192, 175, 156, 119, 104, 100, 99, 108, 113, 116, 
    182, 184, 202, 220, 228, 226, 229, 234, 243, 246, 241, 235, 223, 216, 203, 194, 190, 192, 200, 208, 196, 180, 167, 127, 99, 96, 100, 109, 111, 116, 
    173, 171, 199, 219, 227, 236, 232, 241, 248, 245, 229, 218, 206, 201, 201, 204, 187, 175, 178, 196, 190, 185, 168, 123, 85, 97, 104, 105, 111, 115, 
    135, 149, 199, 209, 219, 238, 236, 237, 245, 243, 227, 213, 203, 188, 190, 206, 192, 166, 162, 181, 175, 167, 149, 95, 78, 98, 103, 102, 107, 111, 
    86, 153, 222, 216, 232, 248, 241, 239, 240, 231, 217, 212, 208, 173, 167, 175, 159, 149, 146, 160, 162, 149, 118, 68, 65, 85, 89, 93, 99, 109, 
    54, 155, 213, 203, 230, 243, 237, 234, 218, 207, 215, 231, 224, 184, 163, 166, 153, 155, 154, 156, 155, 126, 80, 45, 52, 76, 85, 88, 94, 102, 
    59, 153, 190, 215, 244, 240, 230, 229, 208, 206, 229, 242, 221, 192, 177, 153, 157, 175, 166, 177, 156, 113, 74, 41, 47, 69, 83, 90, 90, 94, 
    89, 129, 162, 215, 243, 232, 227, 217, 207, 225, 255, 254, 232, 207, 206, 183, 187, 198, 192, 196, 164, 122, 73, 42, 47, 67, 93, 104, 95, 83, 
    123, 114, 138, 200, 234, 220, 213, 205, 217, 242, 263, 250, 233, 216, 219, 220, 218, 215, 218, 210, 177, 132, 67, 41, 41, 65, 110, 121, 106, 76, 
    140, 121, 144, 203, 235, 225, 205, 194, 213, 245, 234, 233, 239, 224, 219, 216, 210, 211, 206, 191, 168, 115, 53, 28, 28, 60, 119, 142, 116, 74, 
    154, 138, 145, 197, 230, 223, 189, 171, 198, 249, 216, 222, 234, 211, 187, 192, 176, 177, 164, 149, 132, 78, 34, 19, 20, 69, 122, 161, 131, 76, 
    160, 148, 146, 191, 226, 234, 184, 146, 171, 220, 200, 211, 229, 201, 185, 199, 176, 147, 120, 98, 81, 45, 26, 20, 24, 72, 126, 168, 152, 86, 
    173, 152, 153, 190, 220, 227, 179, 103, 100, 146, 174, 205, 207, 155, 165, 187, 169, 125, 74, 47, 40, 30, 34, 28, 31, 70, 130, 180, 176, 105, 
    174, 151, 148, 179, 211, 212, 177, 76, 28, 82, 114, 139, 142, 118, 147, 180, 158, 105, 50, 21, 20, 30, 47, 45, 43, 72, 125, 184, 196, 125, 
    180, 164, 152, 174, 201, 201, 172, 77, 15, 49, 67, 79, 88, 91, 114, 149, 128, 76, 35, 17, 18, 23, 39, 42, 47, 66, 116, 169, 204, 145, 
    187, 162, 150, 171, 190, 195, 166, 97, 63, 50, 46, 59, 78, 79, 92, 92, 60, 34, 11, 0, 0, 0, 10, 27, 43, 59, 100, 148, 191, 158, 
    176, 153, 156, 171, 180, 187, 179, 152, 129, 86, 78, 77, 83, 88, 93, 69, 26, 2, 0, 0, 0, 0, 0, 14, 32, 59, 82, 112, 160, 162, 
    170, 160, 170, 167, 163, 167, 187, 202, 181, 135, 131, 126, 116, 123, 112, 70, 27, 0, 0, 0, 0, 0, 0, 0, 10, 50, 63, 65, 115, 144, 
    164, 167, 183, 178, 163, 164, 188, 193, 177, 152, 137, 136, 135, 146, 132, 97, 61, 39, 25, 12, 5, 0, 0, 3, 21, 53, 52, 56, 89, 130, 
    162, 170, 168, 170, 174, 163, 159, 173, 173, 171, 146, 130, 133, 158, 152, 129, 96, 79, 68, 57, 48, 37, 40, 51, 61, 69, 60, 63, 86, 105, 
    158, 159, 148, 165, 183, 166, 132, 142, 162, 139, 133, 141, 148, 169, 167, 148, 122, 109, 103, 97, 94, 87, 93, 105, 100, 95, 90, 90, 111, 98, 
    151, 148, 138, 171, 181, 169, 148, 145, 162, 142, 143, 154, 157, 169, 171, 155, 135, 128, 125, 120, 125, 129, 138, 144, 139, 132, 129, 125, 121, 110, 
    165, 155, 154, 178, 175, 163, 158, 164, 158, 152, 173, 176, 165, 163, 161, 153, 148, 143, 134, 132, 141, 151, 159, 163, 160, 152, 152, 137, 115, 116, 
    166, 171, 176, 171, 156, 151, 159, 169, 167, 159, 174, 174, 168, 159, 148, 144, 149, 146, 139, 141, 152, 163, 166, 172, 168, 161, 158, 148, 136, 140, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    32, 40, 59, 52, 39, 39, 44, 50, 44, 47, 52, 49, 46, 48, 55, 43, 21, 14, 20, 25, 27, 30, 32, 38, 36, 38, 39, 26, 16, 25, 
    27, 45, 41, 38, 43, 44, 41, 43, 43, 48, 52, 54, 59, 56, 58, 55, 32, 22, 20, 21, 24, 27, 30, 36, 43, 46, 38, 28, 22, 27, 
    20, 32, 18, 28, 46, 52, 45, 46, 49, 46, 50, 51, 54, 58, 58, 60, 47, 31, 31, 29, 28, 28, 29, 30, 34, 34, 31, 31, 31, 31, 
    17, 24, 16, 23, 43, 51, 44, 47, 48, 45, 48, 46, 46, 53, 53, 53, 59, 42, 41, 48, 44, 42, 43, 41, 38, 32, 29, 30, 38, 40, 
    13, 21, 24, 27, 40, 47, 44, 43, 43, 44, 49, 47, 48, 52, 54, 51, 55, 50, 44, 57, 58, 43, 40, 41, 38, 34, 30, 29, 34, 38, 
    9, 13, 31, 25, 35, 43, 44, 45, 42, 40, 51, 52, 49, 47, 54, 55, 52, 50, 43, 45, 55, 34, 31, 34, 28, 33, 33, 32, 32, 31, 
    5, 24, 29, 23, 35, 38, 41, 44, 40, 39, 48, 50, 44, 40, 43, 44, 44, 46, 47, 41, 52, 41, 33, 34, 31, 35, 43, 41, 34, 33, 
    9, 33, 23, 31, 38, 38, 41, 37, 38, 44, 48, 43, 38, 42, 42, 41, 38, 40, 44, 41, 44, 41, 25, 29, 31, 34, 40, 38, 32, 34, 
    15, 20, 28, 35, 35, 41, 44, 44, 40, 39, 39, 26, 22, 37, 40, 37, 34, 40, 41, 39, 36, 28, 1, 15, 25, 30, 27, 26, 29, 32, 
    11, 21, 29, 26, 28, 37, 41, 39, 39, 35, 32, 19, 13, 22, 17, 10, 20, 37, 41, 37, 31, 17, 0, 1, 25, 29, 27, 28, 29, 30, 
    29, 45, 37, 38, 39, 36, 37, 23, 29, 35, 36, 14, 4, 3, 0, 0, 0, 20, 31, 26, 24, 13, 2, 6, 23, 21, 27, 31, 31, 32, 
    51, 41, 24, 33, 36, 27, 24, 16, 25, 39, 41, 8, 0, 1, 8, 12, 3, 22, 31, 12, 11, 3, 3, 15, 21, 21, 26, 30, 30, 30, 
    58, 36, 17, 25, 15, 12, 14, 19, 32, 41, 32, 5, 0, 13, 13, 37, 42, 32, 31, 15, 5, 4, 8, 14, 22, 28, 32, 33, 28, 26, 
    47, 36, 31, 28, 12, 15, 13, 12, 32, 37, 22, 16, 33, 41, 16, 13, 27, 12, 12, 10, 1, 10, 11, 14, 23, 32, 37, 34, 28, 24, 
    36, 41, 48, 26, 9, 10, 18, 12, 22, 19, 7, 9, 38, 49, 22, 5, 4, 1, 1, 0, 0, 3, 0, 7, 17, 31, 36, 23, 25, 22, 
    40, 54, 59, 33, 13, 7, 23, 25, 5, 0, 0, 0, 17, 35, 17, 0, 0, 5, 0, 0, 0, 0, 0, 0, 18, 35, 33, 7, 8, 23, 
    43, 47, 49, 30, 12, 2, 12, 30, 0, 2, 12, 10, 3, 19, 8, 4, 0, 0, 0, 0, 0, 0, 1, 14, 33, 48, 34, 8, 0, 17, 
    40, 44, 39, 18, 5, 0, 0, 30, 0, 0, 36, 26, 1, 25, 32, 43, 24, 0, 0, 0, 0, 11, 25, 32, 39, 53, 39, 9, 0, 4, 
    40, 48, 58, 25, 0, 0, 0, 14, 0, 0, 10, 5, 0, 28, 40, 30, 41, 17, 10, 7, 17, 35, 32, 30, 33, 47, 46, 10, 0, 0, 
    37, 45, 60, 29, 0, 0, 0, 0, 22, 0, 0, 0, 0, 29, 28, 0, 3, 15, 21, 13, 9, 22, 20, 28, 38, 49, 49, 10, 0, 0, 
    36, 39, 48, 29, 0, 0, 0, 0, 46, 39, 3, 0, 0, 28, 33, 0, 0, 0, 11, 15, 1, 6, 10, 19, 38, 48, 49, 9, 0, 0, 
    31, 34, 51, 39, 0, 0, 10, 29, 48, 47, 50, 47, 39, 35, 30, 4, 0, 0, 0, 7, 2, 6, 8, 8, 22, 33, 46, 21, 0, 0, 
    30, 37, 48, 41, 14, 1, 24, 47, 50, 37, 53, 59, 57, 45, 27, 7, 10, 13, 8, 7, 2, 3, 10, 17, 21, 24, 38, 34, 0, 0, 
    44, 52, 40, 32, 29, 8, 9, 23, 45, 52, 53, 48, 48, 47, 33, 26, 30, 29, 26, 19, 11, 8, 10, 20, 27, 19, 20, 29, 15, 0, 
    45, 57, 44, 33, 43, 31, 4, 0, 9, 30, 20, 37, 42, 46, 46, 38, 35, 35, 34, 32, 31, 34, 30, 30, 36, 19, 20, 45, 37, 13, 
    34, 37, 40, 32, 34, 35, 33, 9, 0, 21, 14, 32, 43, 41, 40, 39, 35, 39, 41, 42, 42, 51, 53, 48, 49, 38, 41, 53, 33, 35, 
    31, 31, 39, 33, 23, 20, 39, 38, 4, 20, 44, 52, 49, 36, 37, 44, 42, 40, 42, 44, 45, 55, 56, 48, 47, 50, 52, 47, 22, 19, 
    31, 34, 48, 47, 31, 35, 44, 49, 36, 31, 47, 52, 48, 38, 36, 41, 45, 38, 38, 41, 50, 56, 53, 44, 45, 46, 43, 46, 37, 31, 
    45, 45, 54, 49, 37, 45, 53, 43, 40, 53, 49, 43, 42, 32, 29, 33, 41, 36, 38, 45, 49, 50, 48, 42, 44, 40, 36, 38, 46, 49, 
    54, 50, 40, 25, 28, 33, 41, 35, 29, 32, 32, 35, 38, 31, 29, 31, 37, 38, 44, 50, 46, 46, 46, 40, 38, 40, 37, 42, 52, 47, 
    
    -- channel=83
    110, 103, 93, 92, 89, 93, 95, 90, 90, 80, 72, 70, 64, 53, 56, 65, 53, 28, 17, 27, 33, 34, 27, 24, 33, 42, 51, 57, 47, 35, 
    143, 133, 122, 103, 89, 97, 101, 103, 101, 90, 82, 74, 65, 64, 65, 60, 39, 9, 3, 18, 32, 40, 44, 48, 50, 50, 51, 49, 44, 44, 
    151, 143, 136, 110, 96, 102, 107, 111, 107, 104, 101, 89, 73, 70, 69, 64, 47, 14, 0, 8, 25, 33, 42, 52, 61, 63, 55, 43, 46, 54, 
    146, 137, 138, 121, 107, 110, 115, 113, 116, 117, 106, 99, 84, 69, 77, 82, 73, 51, 20, 21, 42, 41, 36, 46, 57, 61, 60, 53, 49, 57, 
    138, 131, 144, 130, 115, 115, 119, 121, 126, 123, 112, 110, 98, 75, 75, 90, 95, 93, 73, 60, 69, 61, 43, 39, 43, 46, 53, 59, 58, 62, 
    131, 136, 143, 136, 125, 120, 126, 132, 135, 130, 118, 115, 110, 91, 75, 87, 104, 113, 107, 80, 70, 65, 48, 40, 35, 29, 39, 54, 61, 66, 
    138, 135, 136, 137, 128, 127, 131, 136, 135, 128, 117, 111, 110, 98, 81, 84, 95, 102, 108, 92, 79, 80, 56, 36, 33, 32, 41, 52, 60, 65, 
    137, 122, 138, 138, 133, 126, 125, 135, 132, 126, 121, 114, 106, 100, 95, 89, 85, 91, 103, 104, 99, 97, 68, 38, 41, 48, 48, 55, 60, 62, 
    111, 128, 144, 141, 139, 129, 126, 138, 140, 130, 120, 123, 126, 129, 135, 115, 85, 78, 92, 100, 105, 108, 75, 38, 39, 45, 48, 55, 60, 64, 
    87, 129, 129, 130, 139, 143, 141, 137, 127, 126, 143, 168, 169, 162, 170, 151, 102, 78, 89, 101, 97, 85, 51, 31, 34, 37, 41, 48, 58, 64, 
    76, 128, 134, 147, 162, 158, 150, 133, 120, 137, 186, 215, 190, 155, 147, 135, 104, 87, 99, 107, 91, 60, 33, 20, 25, 32, 31, 38, 51, 58, 
    68, 137, 163, 173, 174, 170, 160, 134, 127, 157, 203, 219, 200, 154, 113, 114, 123, 114, 124, 125, 94, 58, 21, 0, 13, 26, 28, 36, 46, 48, 
    57, 116, 162, 188, 195, 189, 171, 151, 157, 185, 201, 193, 182, 179, 159, 146, 161, 159, 159, 146, 102, 59, 24, 8, 14, 25, 32, 33, 38, 39, 
    43, 85, 152, 193, 198, 184, 178, 178, 188, 208, 213, 189, 173, 191, 215, 211, 206, 214, 199, 166, 125, 71, 34, 17, 18, 40, 54, 44, 35, 32, 
    58, 76, 135, 189, 195, 167, 164, 192, 216, 233, 235, 204, 172, 187, 220, 230, 230, 230, 223, 204, 148, 76, 30, 7, 19, 62, 91, 71, 37, 28, 
    77, 81, 135, 188, 199, 170, 149, 187, 229, 214, 203, 205, 184, 178, 192, 204, 207, 203, 204, 183, 121, 51, 3, 0, 14, 65, 115, 107, 49, 21, 
    94, 98, 141, 193, 211, 175, 127, 166, 207, 181, 187, 211, 177, 130, 132, 149, 152, 136, 118, 96, 58, 13, 0, 0, 8, 67, 126, 137, 76, 15, 
    82, 88, 148, 206, 225, 193, 114, 117, 185, 193, 187, 189, 148, 124, 135, 121, 101, 69, 43, 28, 11, 2, 0, 0, 12, 70, 137, 166, 107, 19, 
    87, 92, 145, 213, 240, 211, 102, 39, 115, 165, 161, 163, 139, 135, 159, 129, 73, 32, 10, 11, 11, 9, 0, 0, 10, 69, 154, 202, 143, 36, 
    110, 99, 132, 199, 227, 197, 95, 0, 4, 76, 97, 102, 87, 79, 123, 133, 71, 15, 0, 2, 6, 10, 9, 0, 9, 69, 153, 217, 180, 62, 
    114, 98, 126, 178, 196, 160, 84, 6, 0, 0, 19, 39, 38, 33, 56, 67, 44, 3, 0, 0, 0, 0, 10, 10, 10, 49, 128, 203, 190, 83, 
    112, 101, 115, 150, 171, 143, 100, 61, 26, 3, 2, 17, 35, 41, 20, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 30, 87, 163, 179, 98, 
    104, 113, 115, 127, 152, 167, 149, 87, 51, 52, 50, 44, 45, 37, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 26, 39, 99, 154, 115, 
    104, 117, 119, 109, 130, 170, 168, 122, 92, 88, 75, 66, 59, 55, 44, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 34, 101, 121, 
    100, 103, 122, 122, 112, 124, 154, 159, 120, 91, 71, 71, 89, 85, 65, 41, 20, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 21, 60, 94, 
    100, 101, 117, 135, 119, 87, 105, 141, 115, 87, 85, 86, 104, 103, 80, 59, 48, 43, 39, 29, 13, 12, 23, 19, 14, 23, 32, 55, 54, 44, 
    96, 86, 105, 128, 121, 93, 75, 103, 104, 81, 85, 88, 104, 114, 93, 71, 74, 75, 63, 53, 50, 55, 63, 60, 53, 49, 49, 55, 61, 57, 
    91, 89, 105, 115, 108, 100, 95, 89, 97, 109, 101, 90, 98, 108, 101, 84, 79, 73, 65, 67, 69, 75, 85, 87, 80, 73, 61, 44, 63, 92, 
    108, 116, 114, 114, 113, 105, 108, 112, 109, 112, 114, 102, 91, 90, 91, 83, 73, 69, 68, 71, 76, 83, 96, 99, 92, 87, 74, 62, 67, 87, 
    116, 125, 117, 102, 94, 98, 105, 111, 111, 109, 106, 96, 82, 70, 69, 73, 75, 76, 71, 75, 87, 91, 103, 108, 99, 92, 90, 83, 82, 92, 
    
    -- channel=84
    0, 0, 0, 0, 14, 11, 0, 0, 8, 5, 7, 23, 24, 10, 0, 6, 28, 32, 20, 15, 11, 0, 0, 0, 0, 0, 0, 11, 20, 0, 
    0, 0, 0, 6, 22, 11, 15, 17, 6, 3, 0, 0, 3, 1, 0, 0, 23, 36, 38, 29, 23, 8, 0, 0, 0, 0, 0, 25, 30, 0, 
    9, 2, 31, 29, 7, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 2, 0, 1, 11, 19, 25, 32, 22, 3, 0, 6, 15, 10, 0, 
    27, 47, 48, 28, 3, 0, 0, 0, 2, 10, 4, 12, 18, 20, 20, 2, 0, 0, 0, 0, 0, 0, 0, 12, 27, 32, 22, 5, 0, 0, 
    35, 38, 14, 7, 0, 4, 18, 9, 4, 11, 17, 12, 6, 8, 11, 19, 6, 0, 0, 0, 0, 0, 0, 0, 15, 40, 37, 17, 0, 0, 
    63, 25, 0, 19, 11, 7, 7, 4, 6, 13, 12, 11, 11, 6, 0, 7, 24, 6, 0, 0, 0, 17, 22, 18, 37, 47, 42, 28, 19, 12, 
    51, 3, 11, 38, 23, 16, 9, 9, 22, 34, 31, 25, 41, 45, 27, 22, 37, 37, 25, 12, 0, 0, 10, 16, 27, 11, 0, 2, 13, 15, 
    33, 0, 19, 15, 10, 16, 26, 35, 27, 18, 22, 27, 38, 36, 22, 22, 48, 59, 41, 23, 0, 0, 0, 12, 7, 0, 0, 0, 8, 13, 
    64, 23, 2, 1, 6, 7, 7, 8, 14, 12, 16, 23, 18, 0, 0, 0, 11, 36, 46, 47, 32, 26, 62, 48, 20, 18, 31, 29, 20, 13, 
    98, 21, 24, 52, 32, 7, 0, 0, 28, 35, 3, 0, 0, 0, 0, 0, 3, 4, 15, 38, 50, 83, 127, 78, 21, 26, 36, 32, 25, 19, 
    38, 0, 0, 0, 0, 0, 10, 34, 51, 26, 0, 0, 0, 33, 103, 142, 92, 25, 0, 11, 40, 82, 97, 55, 21, 35, 23, 14, 16, 22, 
    0, 0, 0, 0, 0, 0, 17, 44, 34, 0, 0, 14, 54, 34, 38, 73, 47, 0, 0, 4, 38, 68, 56, 20, 23, 36, 25, 14, 19, 29, 
    0, 29, 57, 5, 25, 35, 20, 13, 0, 0, 0, 72, 80, 1, 0, 0, 0, 0, 0, 0, 34, 44, 34, 5, 0, 0, 0, 3, 20, 37, 
    0, 36, 33, 5, 30, 37, 35, 0, 0, 0, 0, 14, 2, 0, 0, 0, 0, 0, 0, 0, 4, 5, 3, 0, 0, 0, 0, 0, 13, 29, 
    0, 1, 0, 7, 36, 48, 45, 15, 0, 0, 4, 0, 0, 0, 0, 7, 13, 18, 2, 0, 0, 25, 39, 33, 10, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 27, 36, 35, 7, 6, 64, 94, 67, 41, 39, 71, 78, 65, 66, 78, 91, 113, 127, 101, 67, 19, 0, 0, 0, 6, 21, 
    4, 0, 0, 0, 1, 30, 48, 23, 47, 90, 68, 31, 71, 105, 132, 143, 130, 140, 177, 220, 234, 171, 74, 20, 0, 0, 0, 0, 23, 17, 
    38, 37, 0, 0, 0, 27, 73, 71, 82, 46, 0, 0, 82, 52, 0, 11, 89, 152, 171, 178, 141, 54, 0, 0, 0, 0, 0, 0, 15, 28, 
    24, 0, 0, 0, 15, 30, 85, 113, 149, 134, 43, 86, 128, 34, 0, 0, 1, 85, 76, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    2, 0, 0, 4, 44, 89, 140, 117, 115, 221, 228, 200, 174, 114, 109, 145, 96, 64, 40, 17, 9, 0, 10, 0, 0, 0, 0, 0, 25, 23, 
    19, 30, 22, 32, 66, 114, 134, 35, 0, 33, 149, 169, 143, 88, 99, 184, 190, 117, 50, 41, 68, 67, 49, 4, 0, 0, 16, 38, 65, 56, 
    48, 31, 9, 27, 61, 69, 25, 0, 0, 0, 0, 0, 0, 0, 28, 124, 159, 130, 78, 37, 40, 52, 65, 66, 27, 16, 38, 69, 79, 59, 
    69, 17, 0, 22, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 61, 40, 28, 33, 23, 24, 20, 26, 50, 33, 22, 51, 81, 87, 39, 
    28, 1, 15, 36, 43, 25, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 28, 72, 83, 108, 82, 
    0, 0, 27, 18, 0, 50, 94, 63, 0, 0, 25, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 21, 0, 16, 93, 
    28, 48, 41, 10, 0, 20, 66, 87, 73, 68, 83, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    34, 62, 50, 41, 61, 55, 18, 33, 90, 29, 0, 0, 0, 27, 28, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 5, 
    44, 20, 0, 18, 56, 35, 0, 0, 15, 1, 0, 0, 0, 28, 32, 9, 0, 11, 22, 0, 0, 0, 0, 0, 0, 0, 0, 10, 19, 0, 
    15, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 18, 23, 50, 62, 46, 26, 30, 22, 1, 0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 
    0, 0, 8, 63, 72, 50, 27, 33, 41, 28, 37, 40, 37, 60, 73, 64, 35, 11, 0, 0, 1, 3, 3, 11, 16, 15, 7, 0, 0, 0, 
    
    -- channel=85
    43, 46, 52, 76, 88, 87, 86, 84, 85, 87, 92, 94, 88, 83, 83, 79, 73, 75, 82, 83, 76, 66, 65, 62, 66, 68, 75, 68, 65, 62, 
    58, 58, 66, 83, 90, 95, 89, 89, 88, 83, 84, 89, 86, 81, 85, 78, 78, 79, 88, 92, 85, 75, 62, 53, 54, 58, 74, 76, 71, 67, 
    80, 79, 84, 82, 88, 87, 81, 90, 85, 83, 85, 85, 87, 88, 86, 83, 67, 62, 72, 86, 89, 88, 85, 83, 77, 71, 71, 73, 72, 70, 
    84, 87, 92, 82, 88, 87, 85, 88, 86, 89, 91, 90, 94, 101, 95, 89, 59, 38, 41, 54, 65, 66, 72, 87, 87, 84, 74, 67, 69, 69, 
    72, 82, 87, 76, 85, 90, 91, 91, 85, 92, 92, 89, 85, 91, 102, 101, 80, 46, 31, 39, 53, 58, 63, 77, 87, 90, 85, 76, 71, 70, 
    66, 90, 82, 83, 87, 86, 89, 88, 84, 89, 93, 92, 84, 82, 92, 98, 95, 76, 57, 67, 74, 81, 81, 84, 91, 93, 94, 88, 80, 79, 
    75, 85, 83, 92, 90, 91, 90, 88, 93, 96, 100, 99, 97, 94, 93, 99, 101, 99, 87, 81, 74, 76, 73, 81, 81, 79, 80, 79, 80, 80, 
    79, 76, 85, 84, 85, 94, 96, 96, 94, 94, 95, 89, 93, 88, 86, 90, 102, 107, 102, 83, 71, 64, 62, 71, 77, 73, 71, 73, 79, 78, 
    85, 88, 81, 77, 85, 84, 87, 90, 94, 94, 88, 77, 74, 61, 56, 58, 81, 101, 109, 94, 90, 80, 75, 76, 92, 88, 86, 86, 81, 79, 
    110, 106, 89, 94, 95, 83, 80, 88, 102, 99, 70, 48, 50, 58, 55, 53, 64, 82, 95, 89, 96, 101, 87, 92, 94, 88, 89, 89, 85, 82, 
    114, 89, 60, 70, 72, 74, 81, 91, 96, 90, 59, 37, 39, 80, 103, 98, 93, 82, 79, 77, 81, 83, 79, 91, 92, 89, 86, 84, 86, 85, 
    103, 85, 59, 59, 54, 65, 80, 82, 78, 77, 68, 60, 56, 58, 71, 76, 78, 66, 63, 69, 69, 68, 70, 80, 90, 93, 88, 85, 87, 87, 
    92, 98, 100, 81, 71, 70, 69, 59, 60, 64, 72, 79, 76, 46, 7, 5, 15, 16, 37, 47, 57, 62, 60, 68, 74, 79, 81, 79, 85, 88, 
    76, 96, 103, 78, 68, 77, 68, 55, 52, 50, 49, 60, 64, 55, 21, 16, 15, 22, 30, 28, 42, 43, 50, 61, 66, 67, 62, 65, 75, 84, 
    65, 83, 93, 81, 68, 79, 78, 70, 57, 53, 47, 54, 60, 66, 57, 51, 52, 55, 42, 33, 39, 44, 67, 73, 77, 75, 50, 49, 61, 79, 
    56, 60, 76, 74, 62, 68, 77, 75, 82, 80, 88, 82, 77, 91, 91, 80, 80, 81, 83, 82, 75, 81, 89, 88, 90, 88, 64, 44, 51, 75, 
    70, 65, 67, 60, 53, 58, 79, 86, 96, 74, 90, 82, 86, 102, 127, 117, 116, 117, 130, 137, 117, 103, 86, 74, 85, 83, 74, 40, 42, 64, 
    86, 90, 88, 60, 47, 45, 81, 103, 94, 61, 66, 72, 72, 66, 70, 79, 101, 115, 120, 117, 95, 76, 61, 55, 75, 81, 66, 31, 27, 53, 
    67, 79, 83, 65, 50, 42, 64, 122, 138, 114, 94, 92, 83, 80, 46, 42, 61, 80, 80, 68, 57, 55, 55, 66, 82, 90, 69, 28, 10, 35, 
    61, 70, 78, 74, 66, 69, 59, 99, 157, 170, 157, 133, 122, 137, 127, 101, 75, 71, 75, 75, 75, 74, 67, 66, 82, 95, 83, 46, 13, 25, 
    71, 80, 92, 85, 76, 82, 55, 46, 73, 103, 135, 135, 124, 125, 141, 134, 114, 94, 87, 90, 99, 102, 85, 71, 73, 100, 101, 79, 33, 32, 
    73, 77, 87, 82, 74, 58, 35, 33, 20, 28, 46, 62, 66, 85, 99, 110, 123, 110, 94, 84, 88, 101, 108, 102, 90, 104, 114, 102, 54, 37, 
    84, 76, 74, 79, 67, 38, 26, 41, 40, 48, 33, 36, 50, 68, 68, 69, 75, 80, 78, 77, 73, 79, 97, 100, 99, 98, 115, 122, 78, 35, 
    87, 85, 72, 79, 83, 72, 50, 38, 36, 50, 52, 60, 70, 65, 48, 34, 32, 43, 53, 63, 65, 65, 70, 77, 92, 91, 107, 136, 115, 61, 
    81, 85, 73, 61, 75, 105, 96, 74, 69, 73, 82, 74, 70, 55, 43, 35, 33, 32, 33, 36, 38, 41, 44, 61, 80, 79, 80, 83, 104, 92, 
    89, 91, 86, 70, 58, 80, 106, 91, 89, 89, 97, 84, 74, 61, 60, 53, 46, 32, 27, 25, 24, 24, 25, 34, 46, 50, 54, 50, 58, 78, 
    84, 88, 100, 94, 79, 71, 86, 94, 77, 69, 70, 75, 82, 76, 69, 60, 55, 49, 46, 46, 43, 40, 38, 34, 37, 42, 60, 81, 63, 61, 
    78, 69, 86, 81, 79, 71, 66, 68, 62, 69, 63, 70, 83, 84, 73, 67, 70, 74, 72, 70, 64, 63, 60, 57, 54, 58, 69, 77, 70, 63, 
    70, 60, 65, 67, 70, 67, 67, 56, 52, 64, 69, 80, 90, 97, 93, 88, 83, 81, 81, 79, 77, 78, 74, 71, 67, 71, 68, 66, 67, 73, 
    68, 72, 76, 90, 95, 92, 86, 84, 85, 92, 87, 86, 89, 97, 103, 100, 87, 77, 75, 78, 81, 80, 80, 76, 76, 73, 67, 62, 67, 78, 
    
    -- channel=86
    2, 0, 0, 44, 73, 72, 71, 68, 69, 68, 79, 81, 75, 69, 65, 65, 57, 58, 65, 67, 57, 42, 39, 34, 29, 30, 51, 55, 46, 35, 
    15, 10, 34, 65, 75, 82, 79, 73, 70, 64, 64, 70, 68, 60, 62, 58, 68, 70, 77, 78, 67, 53, 33, 12, 10, 25, 56, 67, 60, 44, 
    62, 63, 75, 69, 64, 66, 61, 68, 69, 64, 58, 61, 69, 68, 72, 64, 46, 41, 46, 63, 71, 77, 75, 71, 63, 56, 60, 61, 51, 43, 
    81, 84, 86, 63, 63, 67, 66, 73, 72, 71, 75, 76, 82, 92, 83, 69, 25, 0, 0, 0, 18, 34, 52, 75, 81, 80, 64, 47, 44, 47, 
    70, 72, 65, 49, 64, 76, 79, 77, 71, 78, 76, 75, 68, 77, 85, 88, 62, 9, 0, 0, 0, 21, 36, 62, 82, 90, 81, 62, 53, 51, 
    65, 72, 58, 63, 71, 74, 73, 72, 69, 75, 75, 81, 71, 66, 74, 88, 87, 56, 22, 35, 54, 73, 71, 75, 93, 95, 93, 82, 70, 67, 
    58, 62, 70, 83, 78, 76, 75, 80, 84, 89, 97, 103, 99, 94, 90, 96, 103, 102, 79, 72, 55, 53, 54, 67, 72, 62, 59, 63, 68, 69, 
    59, 61, 71, 67, 67, 81, 91, 95, 88, 85, 90, 95, 97, 87, 80, 87, 106, 114, 103, 74, 45, 36, 43, 53, 53, 43, 48, 56, 67, 67, 
    89, 76, 58, 58, 67, 69, 75, 74, 73, 79, 89, 81, 65, 37, 27, 31, 67, 97, 115, 101, 87, 77, 79, 66, 74, 76, 82, 79, 72, 67, 
    115, 91, 84, 97, 89, 64, 58, 74, 93, 97, 61, 22, 15, 30, 40, 31, 41, 66, 92, 92, 104, 123, 113, 89, 77, 79, 81, 80, 74, 71, 
    88, 64, 43, 42, 39, 52, 71, 93, 98, 76, 22, 0, 14, 81, 130, 129, 104, 70, 67, 72, 87, 109, 85, 75, 74, 77, 72, 71, 74, 76, 
    54, 58, 26, 19, 28, 52, 72, 78, 67, 49, 46, 58, 52, 59, 85, 71, 59, 34, 32, 55, 66, 71, 61, 63, 74, 76, 71, 69, 76, 83, 
    52, 100, 101, 78, 68, 63, 64, 43, 22, 31, 71, 92, 75, 18, 0, 0, 0, 0, 0, 22, 47, 54, 43, 40, 42, 46, 52, 60, 77, 84, 
    65, 100, 100, 73, 66, 73, 61, 30, 11, 24, 40, 41, 35, 25, 0, 0, 0, 0, 0, 2, 16, 17, 20, 29, 29, 22, 21, 34, 58, 75, 
    52, 64, 79, 79, 70, 87, 76, 55, 33, 35, 26, 31, 40, 56, 51, 46, 45, 46, 30, 6, 15, 27, 55, 60, 48, 28, 4, 18, 38, 65, 
    35, 33, 54, 69, 59, 67, 70, 63, 75, 95, 111, 97, 83, 100, 116, 104, 97, 96, 96, 100, 108, 104, 101, 82, 59, 53, 31, 23, 32, 56, 
    57, 46, 52, 49, 40, 54, 82, 83, 118, 97, 90, 76, 100, 140, 177, 154, 160, 168, 196, 217, 183, 130, 77, 43, 43, 45, 48, 19, 25, 43, 
    99, 95, 83, 57, 42, 38, 91, 119, 120, 47, 28, 72, 100, 67, 60, 65, 120, 166, 174, 166, 107, 50, 18, 6, 31, 38, 36, 7, 5, 28, 
    73, 65, 67, 61, 46, 31, 83, 156, 173, 143, 115, 126, 102, 56, 18, 25, 58, 93, 81, 48, 11, 4, 20, 36, 55, 60, 39, 2, 0, 0, 
    46, 54, 74, 83, 77, 82, 89, 131, 192, 230, 233, 199, 166, 174, 170, 145, 105, 80, 61, 52, 53, 54, 50, 41, 49, 66, 70, 33, 0, 0, 
    75, 86, 101, 101, 97, 108, 65, 14, 39, 105, 165, 167, 149, 152, 182, 191, 158, 111, 83, 84, 96, 96, 71, 41, 39, 83, 107, 90, 33, 11, 
    86, 81, 90, 95, 88, 61, 0, 0, 0, 0, 0, 13, 17, 49, 103, 149, 154, 118, 87, 68, 72, 91, 99, 95, 77, 103, 125, 122, 62, 19, 
    96, 71, 72, 86, 70, 6, 0, 0, 6, 6, 0, 0, 0, 48, 72, 65, 54, 51, 49, 49, 46, 54, 78, 86, 77, 88, 128, 146, 90, 19, 
    78, 73, 80, 95, 81, 52, 26, 16, 0, 1, 20, 46, 64, 54, 22, 0, 0, 0, 5, 24, 27, 21, 28, 31, 56, 88, 122, 162, 138, 60, 
    74, 91, 80, 61, 71, 115, 107, 68, 35, 54, 85, 68, 50, 26, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 65, 54, 60, 103, 91, 
    97, 106, 92, 62, 53, 93, 115, 102, 107, 93, 96, 65, 54, 47, 47, 32, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 75, 
    95, 106, 108, 106, 91, 76, 89, 98, 88, 60, 43, 50, 75, 77, 68, 46, 25, 13, 12, 9, 0, 0, 0, 0, 0, 0, 14, 62, 62, 40, 
    94, 64, 73, 88, 93, 65, 48, 65, 47, 35, 35, 55, 80, 88, 75, 57, 55, 70, 68, 53, 35, 34, 35, 30, 24, 27, 50, 77, 54, 19, 
    57, 27, 47, 65, 66, 54, 49, 38, 25, 37, 56, 74, 93, 110, 104, 95, 85, 82, 72, 64, 64, 67, 63, 61, 54, 59, 57, 45, 37, 50, 
    45, 56, 84, 111, 115, 107, 96, 89, 85, 97, 97, 96, 99, 111, 115, 110, 84, 64, 59, 63, 70, 71, 71, 71, 71, 69, 53, 38, 42, 66, 
    
    -- channel=87
    97, 120, 105, 89, 77, 70, 72, 73, 79, 81, 78, 79, 81, 79, 78, 81, 86, 88, 82, 76, 73, 75, 77, 77, 83, 80, 68, 66, 72, 76, 
    99, 103, 95, 91, 80, 73, 73, 77, 81, 79, 79, 78, 75, 78, 77, 78, 81, 83, 83, 81, 78, 75, 76, 76, 74, 65, 62, 64, 69, 72, 
    90, 89, 97, 93, 86, 80, 79, 81, 78, 79, 83, 81, 76, 75, 72, 73, 81, 84, 85, 84, 79, 71, 68, 65, 61, 59, 61, 64, 71, 74, 
    84, 86, 99, 97, 89, 83, 83, 78, 76, 83, 81, 79, 80, 73, 74, 82, 83, 91, 87, 85, 83, 70, 59, 57, 56, 56, 62, 68, 67, 65, 
    83, 88, 105, 97, 85, 81, 82, 80, 78, 83, 83, 81, 79, 74, 76, 84, 81, 89, 93, 87, 81, 72, 61, 53, 51, 54, 60, 66, 64, 61, 
    82, 98, 99, 94, 87, 78, 81, 83, 81, 84, 81, 76, 74, 75, 74, 75, 77, 83, 88, 77, 66, 72, 66, 59, 56, 55, 60, 62, 61, 60, 
    91, 100, 89, 93, 86, 83, 82, 80, 81, 81, 73, 64, 65, 70, 72, 72, 70, 68, 71, 70, 66, 82, 77, 68, 65, 64, 64, 62, 60, 59, 
    98, 84, 89, 90, 86, 85, 80, 83, 81, 75, 68, 61, 61, 63, 68, 69, 66, 66, 65, 68, 73, 83, 80, 75, 76, 74, 65, 61, 62, 58, 
    81, 87, 90, 83, 86, 85, 81, 86, 90, 82, 66, 62, 67, 66, 70, 71, 68, 64, 60, 58, 66, 78, 83, 79, 81, 70, 65, 66, 64, 60, 
    85, 98, 77, 75, 85, 89, 88, 84, 86, 84, 79, 78, 78, 67, 67, 76, 76, 66, 59, 55, 59, 67, 77, 85, 85, 71, 71, 71, 68, 62, 
    104, 94, 70, 79, 89, 87, 81, 79, 82, 98, 101, 92, 74, 60, 61, 73, 81, 73, 65, 57, 56, 60, 79, 91, 85, 82, 77, 71, 68, 60, 
    98, 90, 85, 85, 75, 75, 78, 80, 86, 98, 92, 81, 79, 69, 55, 71, 95, 83, 74, 69, 61, 69, 79, 80, 84, 88, 83, 75, 68, 59, 
    77, 71, 79, 75, 72, 78, 78, 79, 90, 91, 77, 77, 87, 87, 79, 75, 89, 81, 76, 75, 68, 72, 77, 84, 90, 93, 87, 75, 67, 61, 
    57, 59, 76, 73, 72, 74, 78, 86, 87, 80, 76, 84, 86, 79, 78, 76, 72, 80, 79, 71, 78, 77, 80, 87, 90, 95, 88, 75, 69, 66, 
    56, 61, 66, 69, 69, 67, 72, 86, 82, 78, 83, 85, 70, 60, 62, 63, 68, 74, 72, 78, 79, 73, 80, 83, 91, 97, 88, 74, 68, 72, 
    56, 48, 54, 64, 67, 71, 72, 82, 87, 72, 66, 69, 60, 56, 59, 61, 66, 64, 70, 71, 66, 71, 81, 87, 97, 92, 81, 76, 68, 74, 
    49, 46, 48, 58, 67, 73, 69, 75, 83, 63, 72, 74, 59, 45, 58, 67, 63, 53, 54, 59, 71, 84, 91, 96, 95, 87, 76, 74, 78, 73, 
    34, 38, 54, 58, 59, 71, 71, 62, 85, 85, 81, 62, 47, 51, 71, 65, 60, 51, 56, 71, 84, 95, 94, 90, 90, 83, 75, 71, 82, 77, 
    33, 43, 55, 59, 62, 73, 70, 50, 81, 86, 59, 56, 64, 68, 65, 48, 43, 58, 70, 84, 88, 85, 80, 77, 80, 77, 76, 75, 81, 82, 
    43, 45, 42, 51, 61, 70, 74, 56, 64, 80, 66, 60, 61, 40, 34, 46, 45, 58, 76, 89, 83, 73, 74, 73, 76, 77, 69, 70, 86, 88, 
    34, 34, 40, 50, 59, 70, 82, 89, 77, 68, 76, 78, 69, 40, 31, 44, 63, 77, 78, 84, 87, 84, 86, 83, 75, 67, 60, 66, 84, 93, 
    31, 34, 37, 45, 66, 79, 93, 108, 90, 74, 77, 80, 78, 66, 49, 49, 75, 96, 98, 96, 96, 90, 92, 90, 77, 66, 56, 64, 81, 94, 
    34, 39, 32, 41, 67, 88, 100, 87, 69, 78, 76, 70, 63, 52, 49, 73, 93, 102, 105, 101, 99, 98, 97, 93, 89, 79, 58, 60, 80, 89, 
    43, 40, 30, 36, 64, 86, 79, 71, 74, 76, 55, 48, 45, 48, 68, 86, 94, 98, 97, 98, 102, 110, 110, 102, 94, 77, 62, 60, 72, 88, 
    41, 27, 31, 45, 51, 61, 73, 90, 86, 70, 49, 39, 47, 51, 59, 72, 81, 89, 94, 98, 102, 106, 112, 106, 90, 80, 79, 69, 64, 78, 
    34, 32, 37, 47, 47, 45, 58, 80, 72, 66, 73, 58, 48, 42, 48, 58, 70, 79, 89, 94, 95, 97, 100, 94, 85, 93, 93, 79, 64, 54, 
    32, 29, 36, 40, 43, 54, 50, 59, 73, 65, 66, 53, 40, 37, 41, 47, 63, 68, 65, 69, 79, 82, 79, 78, 82, 84, 76, 65, 64, 69, 
    32, 35, 38, 32, 35, 49, 53, 45, 56, 71, 56, 40, 37, 35, 38, 46, 53, 49, 45, 55, 61, 60, 59, 62, 65, 67, 64, 54, 64, 80, 
    46, 49, 35, 27, 38, 40, 41, 49, 53, 49, 42, 41, 40, 39, 42, 47, 46, 45, 46, 50, 50, 49, 50, 50, 49, 53, 58, 64, 65, 55, 
    44, 40, 30, 29, 33, 33, 32, 43, 51, 48, 40, 38, 43, 46, 49, 52, 52, 53, 48, 45, 49, 47, 47, 46, 43, 45, 55, 58, 53, 47, 
    
    -- channel=88
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 27, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 32, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 38, 34, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 53, 37, 10, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 57, 35, 6, 0, 0, 0, 0, 48, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 37, 23, 4, 0, 0, 0, 0, 78, 26, 
    0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 14, 0, 0, 0, 0, 0, 99, 76, 
    0, 0, 0, 0, 0, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 5, 1, 4, 0, 6, 3, 0, 0, 0, 0, 112, 121, 
    0, 0, 0, 0, 0, 0, 102, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 8, 0, 0, 0, 0, 5, 0, 0, 0, 0, 96, 144, 
    0, 0, 0, 0, 0, 0, 73, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 135, 
    0, 0, 0, 0, 0, 0, 18, 10, 6, 14, 0, 0, 0, 0, 0, 0, 0, 0, 17, 10, 22, 0, 0, 0, 0, 0, 0, 0, 0, 110, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 41, 21, 27, 29, 44, 38, 0, 0, 0, 0, 0, 0, 0, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 50, 43, 42, 43, 51, 45, 27, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 23, 31, 37, 42, 51, 32, 18, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=89
    77, 70, 60, 74, 80, 75, 72, 75, 83, 84, 87, 90, 90, 89, 91, 96, 97, 95, 88, 83, 80, 79, 81, 84, 85, 77, 73, 74, 75, 72, 
    72, 66, 73, 86, 87, 86, 82, 85, 84, 80, 81, 84, 85, 84, 83, 85, 97, 100, 98, 91, 83, 75, 67, 60, 57, 60, 72, 80, 81, 77, 
    80, 80, 87, 85, 84, 83, 81, 84, 80, 80, 78, 76, 78, 77, 77, 85, 93, 95, 93, 92, 90, 85, 80, 72, 67, 67, 72, 79, 79, 72, 
    87, 94, 99, 88, 84, 81, 80, 81, 80, 80, 81, 84, 86, 86, 82, 82, 76, 74, 72, 76, 79, 75, 77, 80, 77, 77, 75, 73, 71, 70, 
    81, 92, 94, 81, 81, 84, 85, 84, 80, 83, 87, 87, 82, 86, 88, 88, 79, 69, 60, 57, 61, 61, 61, 65, 72, 78, 78, 73, 67, 67, 
    84, 95, 85, 84, 82, 81, 85, 84, 79, 83, 85, 81, 74, 79, 83, 88, 88, 77, 65, 61, 69, 81, 78, 75, 80, 83, 85, 81, 74, 71, 
    94, 90, 86, 93, 87, 84, 83, 83, 83, 84, 86, 81, 79, 82, 82, 83, 81, 82, 79, 80, 81, 89, 82, 79, 81, 80, 78, 75, 75, 73, 
    85, 80, 90, 88, 84, 88, 90, 91, 86, 85, 85, 76, 75, 79, 81, 81, 85, 87, 82, 75, 68, 70, 72, 75, 77, 69, 64, 67, 72, 71, 
    89, 91, 82, 76, 81, 85, 90, 90, 86, 81, 78, 70, 63, 55, 54, 57, 73, 83, 83, 77, 79, 82, 85, 81, 84, 79, 80, 79, 75, 73, 
    111, 98, 79, 86, 89, 84, 79, 79, 90, 97, 87, 64, 50, 46, 46, 51, 64, 73, 77, 75, 83, 98, 104, 98, 91, 88, 91, 87, 80, 74, 
    110, 86, 78, 86, 80, 75, 75, 83, 97, 100, 76, 47, 44, 72, 88, 88, 85, 72, 65, 64, 75, 96, 105, 98, 88, 87, 86, 83, 79, 76, 
    88, 73, 59, 51, 49, 65, 77, 82, 89, 88, 75, 68, 76, 84, 97, 107, 102, 76, 65, 65, 70, 83, 86, 87, 95, 96, 92, 85, 79, 77, 
    77, 89, 89, 74, 71, 74, 75, 75, 76, 72, 77, 90, 97, 73, 41, 33, 41, 40, 50, 60, 72, 82, 84, 86, 89, 89, 89, 82, 81, 80, 
    70, 94, 96, 77, 74, 78, 76, 68, 58, 58, 68, 81, 84, 68, 38, 23, 26, 36, 42, 49, 66, 69, 73, 78, 79, 79, 75, 72, 77, 81, 
    74, 81, 78, 73, 69, 78, 83, 77, 61, 59, 55, 54, 55, 61, 58, 58, 63, 65, 59, 55, 57, 63, 81, 86, 88, 79, 61, 61, 70, 80, 
    59, 58, 68, 74, 70, 78, 85, 83, 77, 72, 77, 73, 66, 74, 82, 82, 83, 81, 81, 77, 80, 94, 106, 106, 98, 84, 67, 60, 66, 80, 
    57, 49, 55, 60, 55, 63, 81, 85, 91, 89, 99, 81, 71, 87, 114, 108, 103, 101, 112, 126, 129, 126, 115, 102, 94, 84, 76, 63, 67, 75, 
    64, 70, 74, 60, 50, 60, 90, 96, 98, 75, 61, 59, 73, 86, 94, 89, 105, 118, 128, 134, 122, 106, 89, 78, 79, 77, 72, 56, 59, 72, 
    63, 72, 76, 66, 53, 55, 83, 107, 118, 91, 67, 76, 78, 59, 33, 33, 64, 97, 104, 96, 76, 64, 69, 76, 81, 82, 73, 52, 50, 68, 
    48, 51, 63, 72, 67, 74, 91, 111, 145, 150, 128, 109, 97, 88, 81, 75, 69, 82, 90, 85, 74, 71, 78, 82, 85, 86, 77, 60, 54, 62, 
    51, 61, 78, 82, 80, 94, 99, 91, 101, 129, 150, 137, 113, 99, 110, 117, 109, 97, 95, 104, 108, 102, 90, 76, 71, 83, 87, 81, 72, 72, 
    56, 62, 72, 80, 85, 85, 79, 62, 48, 60, 81, 91, 83, 76, 84, 110, 129, 124, 111, 105, 107, 110, 107, 96, 83, 92, 97, 99, 88, 78, 
    64, 56, 57, 75, 82, 67, 49, 49, 57, 62, 44, 41, 46, 60, 82, 106, 113, 116, 112, 104, 101, 104, 111, 109, 101, 94, 96, 107, 96, 72, 
    68, 57, 55, 75, 86, 70, 48, 53, 55, 52, 43, 48, 55, 65, 75, 75, 74, 82, 88, 95, 101, 103, 103, 96, 91, 87, 97, 114, 106, 76, 
    52, 54, 59, 65, 77, 94, 91, 79, 53, 47, 56, 57, 55, 51, 55, 58, 61, 68, 73, 79, 85, 90, 90, 86, 91, 96, 96, 94, 105, 96, 
    60, 60, 57, 52, 53, 79, 102, 102, 94, 93, 95, 67, 49, 45, 57, 60, 61, 59, 58, 57, 59, 61, 61, 65, 77, 82, 71, 56, 66, 84, 
    62, 65, 70, 68, 65, 70, 80, 90, 85, 74, 70, 60, 58, 56, 60, 63, 61, 54, 51, 57, 59, 54, 50, 52, 56, 56, 61, 71, 74, 73, 
    63, 60, 63, 63, 70, 70, 64, 69, 74, 64, 47, 50, 60, 58, 57, 57, 58, 61, 62, 64, 60, 56, 56, 57, 57, 58, 67, 81, 84, 65, 
    65, 48, 43, 48, 54, 49, 49, 50, 48, 47, 51, 62, 68, 68, 67, 69, 69, 71, 67, 61, 60, 60, 59, 58, 57, 61, 65, 67, 61, 54, 
    46, 43, 47, 57, 59, 56, 57, 64, 62, 59, 58, 65, 72, 80, 84, 82, 74, 65, 58, 58, 64, 63, 62, 59, 58, 61, 63, 62, 58, 62, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 19, 16, 7, 0, 0, 0, 0, 0, 0, 1, 5, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 29, 29, 16, 5, 0, 0, 0, 0, 0, 1, 10, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 18, 11, 10, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 3, 1, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 26, 15, 3, 6, 5, 0, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 2, 0, 0, 0, 0, 2, 23, 32, 20, 13, 7, 2, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 23, 29, 26, 18, 12, 5, 2, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 20, 26, 17, 7, 1, 0, 4, 7, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 19, 14, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 36, 30, 4, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 32, 58, 57, 42, 12, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 18, 21, 17, 40, 63, 74, 74, 59, 45, 26, 5, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 14, 24, 0, 0, 0, 0, 0, 0, 0, 0, 35, 56, 68, 59, 44, 24, 18, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 29, 80, 41, 0, 0, 0, 0, 0, 0, 0, 12, 40, 36, 14, 6, 8, 18, 24, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 41, 81, 106, 87, 58, 33, 22, 21, 12, 0, 8, 33, 45, 34, 25, 20, 15, 14, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 19, 11, 34, 76, 77, 53, 26, 25, 41, 53, 49, 42, 53, 61, 57, 45, 20, 2, 4, 12, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 41, 74, 81, 70, 61, 61, 62, 63, 54, 32, 20, 17, 25, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 31, 46, 55, 62, 64, 66, 63, 60, 55, 43, 22, 19, 36, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 32, 48, 58, 61, 54, 38, 34, 26, 33, 47, 46, 20, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 16, 23, 24, 15, 20, 29, 24, 11, 6, 22, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=92
    19, 35, 53, 60, 53, 51, 54, 51, 44, 42, 42, 38, 30, 25, 40, 44, 29, 22, 31, 36, 29, 18, 17, 13, 21, 31, 48, 35, 22, 22, 
    65, 76, 69, 59, 54, 66, 62, 59, 52, 43, 36, 33, 25, 21, 31, 28, 16, 8, 26, 40, 38, 30, 19, 13, 20, 27, 40, 35, 28, 28, 
    103, 100, 86, 58, 56, 65, 57, 65, 57, 49, 47, 37, 27, 29, 30, 22, 0, 0, 6, 33, 41, 40, 39, 44, 43, 37, 32, 25, 28, 35, 
    107, 104, 95, 65, 66, 69, 65, 69, 63, 64, 61, 47, 40, 42, 38, 33, 2, 0, 0, 9, 26, 20, 22, 42, 47, 43, 31, 22, 30, 38, 
    91, 96, 100, 73, 71, 75, 75, 75, 71, 72, 63, 52, 41, 36, 49, 53, 36, 8, 0, 7, 27, 15, 11, 27, 36, 39, 38, 35, 35, 39, 
    78, 107, 104, 84, 79, 74, 78, 80, 78, 73, 64, 60, 47, 35, 45, 57, 60, 49, 31, 35, 42, 33, 24, 28, 32, 31, 41, 45, 43, 47, 
    84, 113, 102, 95, 84, 81, 86, 85, 86, 76, 70, 65, 60, 50, 49, 60, 69, 69, 57, 41, 35, 33, 20, 24, 21, 18, 32, 38, 43, 47, 
    99, 97, 98, 91, 83, 86, 90, 91, 83, 72, 70, 62, 62, 54, 53, 58, 67, 70, 68, 45, 44, 42, 20, 19, 25, 28, 32, 35, 42, 44, 
    96, 99, 100, 89, 88, 79, 80, 86, 87, 78, 73, 66, 68, 62, 60, 49, 51, 62, 75, 61, 73, 70, 37, 26, 47, 47, 44, 47, 45, 44, 
    96, 118, 100, 99, 99, 83, 81, 89, 95, 89, 82, 83, 90, 101, 100, 71, 46, 52, 69, 65, 80, 77, 39, 38, 53, 42, 42, 48, 47, 47, 
    107, 114, 73, 87, 98, 95, 95, 93, 89, 98, 113, 121, 109, 124, 138, 113, 77, 65, 72, 68, 66, 47, 21, 43, 50, 40, 37, 39, 46, 48, 
    114, 115, 85, 102, 103, 99, 102, 85, 82, 113, 152, 152, 120, 97, 87, 88, 84, 75, 83, 79, 56, 25, 14, 31, 44, 43, 37, 38, 45, 44, 
    105, 121, 134, 140, 125, 118, 105, 77, 94, 132, 152, 139, 118, 86, 42, 52, 72, 71, 90, 79, 51, 25, 12, 21, 33, 36, 34, 35, 40, 39, 
    65, 95, 143, 140, 124, 124, 111, 96, 118, 137, 124, 103, 100, 111, 92, 106, 109, 110, 112, 75, 50, 20, 12, 22, 30, 39, 33, 26, 29, 34, 
    28, 73, 133, 142, 121, 117, 119, 131, 147, 149, 128, 103, 97, 127, 141, 148, 149, 153, 131, 97, 64, 26, 28, 28, 41, 63, 48, 26, 18, 32, 
    18, 53, 118, 137, 118, 101, 113, 148, 175, 162, 155, 133, 114, 138, 153, 150, 153, 155, 151, 134, 81, 41, 31, 26, 54, 87, 81, 41, 13, 29, 
    35, 60, 111, 129, 122, 95, 103, 156, 178, 126, 143, 139, 115, 118, 136, 142, 145, 139, 145, 131, 73, 33, 11, 9, 50, 89, 104, 58, 17, 19, 
    45, 74, 129, 141, 135, 96, 86, 149, 162, 106, 130, 131, 84, 68, 77, 84, 94, 87, 81, 63, 23, 5, 0, 0, 44, 89, 111, 75, 22, 10, 
    26, 61, 127, 154, 150, 106, 52, 111, 170, 156, 148, 127, 72, 85, 74, 45, 27, 18, 18, 10, 0, 4, 0, 6, 45, 96, 127, 105, 28, 0, 
    30, 59, 116, 157, 162, 127, 28, 37, 131, 169, 163, 124, 85, 120, 131, 87, 24, 0, 9, 24, 27, 28, 6, 2, 36, 98, 146, 140, 53, 0, 
    49, 62, 112, 150, 147, 111, 9, 0, 24, 62, 96, 91, 66, 76, 103, 85, 45, 12, 12, 28, 39, 45, 25, 9, 28, 90, 148, 165, 80, 7, 
    49, 52, 94, 126, 123, 73, 3, 0, 0, 0, 0, 16, 18, 36, 43, 31, 36, 26, 15, 14, 18, 33, 43, 41, 39, 74, 127, 162, 93, 14, 
    50, 56, 73, 100, 104, 67, 37, 24, 0, 0, 0, 0, 10, 25, 3, 0, 0, 3, 6, 9, 3, 8, 30, 36, 47, 54, 91, 139, 106, 21, 
    52, 69, 63, 74, 102, 116, 93, 35, 10, 25, 23, 22, 29, 17, 0, 0, 0, 0, 0, 0, 0, 0, 4, 16, 48, 38, 51, 110, 120, 57, 
    55, 67, 60, 54, 82, 127, 129, 82, 61, 58, 43, 30, 33, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 36, 15, 15, 49, 88, 83, 
    63, 65, 71, 67, 58, 70, 110, 111, 89, 68, 59, 52, 57, 36, 20, 6, 2, 0, 0, 0, 0, 0, 0, 0, 3, 0, 10, 33, 41, 49, 
    57, 56, 84, 90, 64, 40, 69, 92, 64, 42, 42, 56, 68, 52, 29, 15, 21, 21, 16, 9, 1, 8, 13, 4, 1, 6, 27, 59, 31, 25, 
    44, 37, 73, 71, 53, 38, 47, 57, 39, 52, 46, 48, 60, 57, 36, 27, 38, 39, 29, 26, 24, 34, 36, 29, 25, 28, 32, 35, 28, 44, 
    40, 43, 59, 50, 43, 40, 51, 42, 38, 58, 53, 51, 58, 61, 52, 47, 43, 33, 30, 36, 38, 46, 48, 44, 39, 42, 29, 17, 34, 62, 
    52, 67, 65, 61, 63, 64, 67, 66, 70, 78, 61, 52, 50, 52, 56, 53, 41, 30, 32, 40, 47, 50, 58, 52, 48, 44, 32, 28, 43, 62, 
    
    -- channel=93
    0, 0, 0, 4, 3, 3, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 12, 20, 11, 0, 0, 10, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 38, 32, 14, 0, 0, 8, 10, 7, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    46, 34, 20, 16, 5, 4, 14, 14, 15, 16, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 23, 17, 23, 15, 15, 17, 18, 22, 23, 13, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 16, 27, 32, 23, 19, 19, 24, 29, 27, 20, 16, 16, 3, 0, 0, 1, 5, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 16, 31, 28, 23, 23, 25, 31, 36, 30, 23, 23, 27, 13, 4, 4, 11, 14, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 21, 24, 25, 25, 25, 26, 26, 27, 25, 25, 27, 28, 11, 6, 10, 12, 9, 13, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 12, 29, 35, 32, 23, 18, 20, 30, 32, 33, 36, 37, 29, 32, 34, 19, 5, 12, 19, 20, 19, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 44, 35, 27, 29, 29, 35, 34, 18, 17, 42, 72, 75, 71, 67, 34, 5, 8, 22, 24, 23, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 16, 32, 47, 46, 40, 24, 5, 33, 85, 105, 94, 84, 63, 30, 10, 12, 32, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 48, 56, 74, 70, 62, 45, 17, 19, 70, 104, 95, 52, 28, 6, 0, 14, 23, 42, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 21, 44, 69, 91, 78, 64, 44, 27, 49, 91, 87, 60, 42, 31, 32, 32, 44, 53, 55, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 67, 88, 82, 63, 55, 59, 79, 87, 67, 45, 53, 78, 101, 97, 96, 91, 73, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 73, 92, 80, 59, 58, 83, 109, 112, 93, 76, 73, 99, 119, 115, 110, 102, 90, 67, 23, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 27, 69, 84, 73, 52, 48, 102, 128, 107, 93, 94, 88, 92, 98, 99, 101, 102, 101, 70, 12, 0, 0, 0, 0, 6, 20, 3, 0, 
    24, 20, 39, 79, 99, 86, 59, 43, 84, 91, 56, 82, 109, 72, 55, 57, 63, 75, 63, 46, 3, 0, 0, 0, 0, 0, 10, 34, 18, 0, 
    35, 20, 36, 86, 114, 95, 63, 33, 40, 75, 69, 94, 84, 19, 4, 34, 24, 16, 0, 0, 0, 0, 0, 0, 0, 0, 10, 51, 42, 0, 
    21, 9, 31, 87, 125, 114, 64, 21, 10, 61, 85, 87, 65, 40, 48, 71, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 70, 67, 0, 
    40, 33, 42, 83, 121, 116, 45, 0, 0, 0, 39, 43, 35, 34, 56, 72, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 84, 87, 16, 
    56, 40, 39, 68, 97, 84, 6, 0, 0, 0, 0, 0, 0, 0, 3, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 74, 85, 27, 
    53, 33, 35, 52, 68, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 39, 60, 27, 
    40, 29, 44, 51, 41, 32, 25, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 27, 20, 
    26, 39, 50, 44, 39, 50, 60, 39, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 13, 
    34, 42, 40, 30, 33, 46, 48, 51, 55, 34, 27, 10, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    44, 48, 42, 48, 48, 29, 23, 21, 38, 18, 0, 6, 26, 35, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 39, 33, 51, 58, 24, 6, 19, 19, 0, 0, 13, 31, 41, 27, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 21, 29, 44, 40, 18, 8, 11, 12, 11, 22, 32, 32, 42, 32, 18, 12, 14, 2, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    14, 28, 45, 53, 41, 34, 34, 30, 29, 33, 41, 37, 31, 37, 28, 20, 12, 3, 0, 0, 6, 11, 17, 23, 20, 14, 3, 0, 0, 10, 
    32, 54, 64, 63, 46, 38, 42, 45, 45, 45, 45, 33, 21, 17, 7, 2, 2, 2, 5, 7, 14, 19, 26, 34, 34, 23, 11, 3, 7, 20, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    292, 286, 292, 295, 299, 305, 308, 313, 314, 312, 309, 306, 295, 279, 259, 231, 202, 175, 168, 176, 186, 193, 186, 186, 189, 195, 193, 190, 180, 175, 
    295, 297, 301, 300, 299, 292, 299, 312, 321, 324, 330, 330, 326, 315, 303, 280, 234, 188, 158, 161, 178, 194, 206, 220, 224, 221, 205, 192, 182, 185, 
    271, 280, 286, 303, 311, 306, 315, 322, 328, 333, 342, 346, 344, 337, 328, 321, 280, 221, 172, 158, 172, 184, 193, 203, 216, 221, 214, 205, 201, 200, 
    254, 256, 269, 301, 312, 317, 324, 325, 332, 333, 337, 342, 339, 330, 339, 341, 329, 271, 220, 204, 210, 218, 215, 212, 217, 218, 220, 220, 215, 211, 
    246, 247, 269, 301, 312, 317, 321, 324, 328, 333, 341, 347, 347, 335, 335, 339, 332, 305, 275, 267, 262, 256, 245, 231, 224, 218, 217, 220, 220, 221, 
    234, 236, 268, 294, 306, 316, 323, 321, 326, 338, 353, 353, 352, 342, 331, 330, 324, 316, 306, 289, 276, 255, 241, 227, 213, 211, 209, 212, 216, 217, 
    229, 232, 263, 281, 300, 312, 317, 319, 323, 340, 349, 346, 338, 328, 316, 309, 306, 309, 317, 306, 301, 280, 253, 228, 215, 221, 223, 221, 219, 218, 
    221, 241, 261, 286, 306, 308, 308, 310, 326, 350, 346, 330, 318, 315, 302, 287, 282, 294, 314, 319, 311, 289, 256, 225, 220, 226, 227, 225, 219, 220, 
    206, 238, 268, 292, 306, 316, 315, 322, 338, 348, 324, 297, 288, 301, 299, 289, 277, 283, 291, 295, 279, 254, 216, 201, 197, 204, 203, 206, 213, 220, 
    189, 229, 259, 270, 292, 321, 324, 325, 322, 316, 290, 267, 254, 250, 250, 262, 268, 272, 272, 273, 248, 209, 169, 165, 179, 193, 195, 198, 210, 217, 
    182, 242, 278, 287, 304, 312, 306, 296, 293, 290, 271, 241, 218, 187, 165, 173, 207, 236, 245, 248, 227, 184, 157, 144, 165, 185, 194, 200, 207, 213, 
    189, 248, 289, 298, 302, 296, 285, 278, 278, 275, 241, 203, 196, 182, 163, 169, 189, 218, 224, 220, 209, 181, 150, 132, 145, 171, 188, 197, 202, 206, 
    184, 212, 236, 253, 261, 262, 262, 269, 271, 260, 228, 208, 214, 236, 240, 244, 243, 238, 228, 212, 193, 168, 142, 130, 144, 177, 195, 197, 194, 196, 
    188, 200, 217, 246, 251, 247, 248, 262, 266, 257, 253, 264, 271, 262, 255, 236, 234, 231, 219, 220, 202, 177, 150, 132, 148, 188, 213, 209, 191, 186, 
    221, 212, 220, 239, 248, 234, 231, 233, 246, 252, 271, 292, 299, 267, 232, 205, 202, 199, 208, 220, 203, 173, 129, 114, 137, 186, 224, 216, 191, 173, 
    258, 242, 233, 236, 247, 238, 222, 217, 218, 213, 221, 253, 273, 251, 212, 197, 193, 192, 192, 178, 154, 126, 95, 96, 127, 172, 214, 208, 183, 162, 
    275, 253, 239, 243, 249, 237, 206, 193, 181, 205, 218, 247, 249, 219, 189, 183, 175, 163, 134, 102, 95, 94, 101, 111, 136, 178, 203, 205, 171, 151, 
    262, 237, 221, 222, 228, 229, 182, 153, 161, 231, 253, 246, 234, 244, 242, 240, 195, 145, 112, 94, 113, 133, 139, 141, 153, 191, 205, 206, 170, 141, 
    273, 253, 226, 206, 204, 218, 169, 111, 108, 156, 201, 206, 227, 257, 286, 286, 248, 176, 136, 134, 158, 170, 160, 145, 153, 186, 207, 201, 176, 146, 
    291, 265, 232, 193, 177, 180, 155, 92, 61, 60, 89, 134, 177, 192, 214, 223, 223, 187, 142, 121, 127, 147, 157, 155, 166, 185, 193, 187, 171, 154, 
    278, 254, 223, 187, 169, 165, 168, 153, 123, 95, 70, 96, 145, 181, 184, 169, 159, 146, 122, 97, 87, 107, 141, 166, 178, 178, 173, 164, 163, 155, 
    271, 262, 236, 200, 179, 192, 224, 227, 211, 188, 169, 171, 200, 216, 189, 138, 100, 89, 85, 83, 76, 79, 103, 127, 156, 162, 164, 156, 167, 169, 
    268, 272, 258, 217, 194, 232, 275, 264, 248, 233, 243, 246, 249, 222, 183, 135, 99, 84, 76, 72, 65, 62, 72, 103, 141, 160, 157, 157, 172, 191, 
    283, 285, 266, 227, 206, 219, 255, 277, 288, 275, 269, 257, 246, 239, 215, 179, 151, 125, 105, 84, 71, 66, 75, 112, 136, 146, 143, 138, 151, 179, 
    290, 285, 276, 255, 226, 195, 205, 240, 264, 257, 246, 260, 271, 276, 253, 218, 186, 161, 145, 132, 119, 111, 117, 130, 134, 145, 161, 168, 159, 161, 
    271, 268, 270, 273, 256, 219, 200, 194, 193, 211, 215, 246, 269, 281, 266, 240, 216, 206, 198, 190, 187, 190, 193, 186, 182, 192, 204, 214, 183, 173, 
    251, 243, 247, 252, 252, 241, 220, 208, 197, 226, 251, 258, 264, 279, 274, 258, 242, 234, 226, 224, 232, 242, 243, 242, 240, 241, 231, 204, 191, 200, 
    245, 252, 259, 263, 258, 263, 256, 235, 240, 253, 276, 278, 275, 281, 284, 271, 254, 239, 239, 249, 263, 268, 269, 267, 263, 259, 245, 218, 218, 231, 
    274, 287, 285, 287, 284, 288, 283, 274, 275, 280, 290, 286, 273, 264, 264, 260, 255, 253, 258, 268, 276, 279, 282, 279, 275, 264, 258, 254, 245, 242, 
    302, 296, 279, 260, 256, 263, 266, 262, 256, 263, 282, 282, 264, 242, 241, 247, 262, 269, 269, 275, 278, 281, 283, 282, 275, 267, 269, 267, 259, 250, 
    
    -- channel=96
    285, 299, 301, 303, 318, 327, 322, 316, 309, 291, 272, 261, 259, 257, 241, 221, 198, 176, 183, 171, 157, 144, 112, 78, 50, 39, 37, 62, 86, 88, 
    316, 316, 306, 295, 298, 292, 280, 269, 260, 245, 229, 220, 219, 219, 205, 190, 175, 162, 147, 143, 143, 127, 98, 71, 33, 5, 16, 58, 94, 94, 
    299, 291, 280, 267, 259, 246, 232, 221, 211, 200, 188, 180, 181, 183, 173, 164, 153, 148, 138, 129, 126, 116, 100, 65, 16, 0, 16, 67, 99, 99, 
    250, 241, 230, 223, 211, 200, 191, 181, 173, 166, 158, 153, 155, 158, 153, 149, 142, 144, 138, 120, 104, 110, 98, 60, 30, 22, 45, 92, 110, 106, 
    194, 188, 185, 176, 169, 162, 159, 152, 149, 145, 141, 140, 144, 148, 148, 145, 141, 145, 136, 102, 86, 87, 62, 43, 57, 53, 81, 111, 117, 109, 
    153, 148, 144, 138, 139, 139, 140, 137, 137, 137, 137, 139, 142, 148, 151, 152, 148, 154, 138, 98, 85, 57, 21, 36, 67, 80, 105, 121, 123, 113, 
    121, 122, 122, 124, 128, 128, 131, 132, 135, 139, 141, 143, 149, 159, 164, 170, 163, 161, 137, 100, 76, 22, 0, 38, 85, 107, 121, 123, 120, 110, 
    109, 116, 120, 123, 127, 127, 129, 132, 136, 144, 150, 156, 163, 166, 166, 167, 160, 153, 131, 100, 60, 12, 11, 53, 105, 123, 120, 118, 112, 105, 
    110, 117, 123, 124, 128, 128, 131, 131, 134, 139, 146, 151, 154, 162, 169, 180, 186, 191, 176, 144, 68, 25, 25, 52, 106, 121, 116, 112, 105, 100, 
    114, 120, 125, 127, 129, 128, 131, 131, 127, 129, 138, 146, 166, 191, 200, 202, 196, 189, 190, 160, 109, 92, 57, 28, 66, 88, 114, 108, 99, 93, 
    120, 123, 127, 128, 130, 129, 130, 126, 122, 125, 135, 132, 141, 145, 136, 131, 128, 127, 141, 120, 128, 163, 94, 24, 14, 45, 87, 107, 93, 88, 
    127, 126, 128, 128, 129, 130, 125, 120, 110, 110, 106, 93, 99, 109, 94, 87, 84, 81, 68, 64, 157, 226, 143, 46, 0, 0, 50, 81, 81, 79, 
    131, 129, 130, 128, 126, 125, 113, 101, 94, 97, 87, 80, 86, 75, 39, 21, 15, 20, 0, 25, 163, 233, 189, 94, 0, 0, 12, 38, 52, 67, 
    131, 131, 132, 126, 125, 118, 107, 86, 94, 84, 68, 50, 55, 33, 0, 0, 8, 28, 21, 91, 178, 210, 207, 135, 23, 0, 0, 5, 31, 72, 
    130, 130, 130, 117, 111, 104, 94, 92, 78, 68, 37, 39, 56, 46, 46, 70, 99, 110, 121, 175, 204, 198, 202, 124, 18, 0, 0, 0, 37, 97, 
    127, 127, 120, 98, 77, 71, 69, 62, 50, 35, 15, 27, 40, 30, 86, 139, 148, 170, 201, 219, 209, 207, 169, 69, 24, 15, 0, 3, 77, 135, 
    124, 120, 112, 91, 77, 51, 42, 29, 41, 11, 0, 10, 16, 24, 136, 205, 213, 224, 230, 229, 235, 236, 154, 45, 37, 51, 38, 56, 116, 160, 
    118, 117, 108, 118, 92, 17, 0, 13, 25, 0, 0, 0, 0, 37, 173, 221, 212, 207, 211, 218, 235, 223, 153, 83, 68, 80, 84, 109, 133, 163, 
    111, 101, 115, 170, 114, 22, 0, 4, 2, 0, 0, 0, 0, 43, 166, 192, 177, 170, 169, 145, 144, 160, 151, 127, 118, 124, 133, 137, 127, 144, 
    90, 66, 131, 175, 114, 32, 0, 1, 0, 0, 0, 0, 0, 53, 160, 176, 157, 161, 124, 64, 55, 89, 116, 146, 153, 144, 132, 120, 115, 94, 
    56, 50, 110, 102, 83, 43, 0, 2, 0, 0, 0, 0, 0, 71, 161, 168, 162, 159, 58, 4, 0, 10, 54, 109, 142, 130, 111, 107, 79, 32, 
    50, 63, 57, 38, 64, 52, 10, 0, 0, 0, 0, 0, 18, 89, 172, 171, 183, 121, 0, 0, 0, 0, 0, 63, 118, 113, 99, 84, 26, 0, 
    56, 51, 0, 0, 45, 60, 19, 0, 0, 0, 0, 31, 43, 117, 172, 175, 179, 74, 0, 0, 0, 0, 0, 14, 75, 97, 94, 41, 0, 0, 
    44, 26, 0, 0, 39, 66, 16, 0, 0, 0, 16, 38, 53, 131, 167, 177, 163, 55, 0, 0, 0, 0, 0, 0, 41, 89, 72, 2, 0, 0, 
    26, 10, 1, 0, 37, 67, 25, 0, 0, 32, 71, 80, 108, 159, 173, 180, 154, 51, 0, 16, 27, 12, 0, 0, 14, 68, 35, 0, 0, 0, 
    18, 5, 0, 0, 28, 52, 5, 0, 0, 15, 45, 56, 78, 102, 106, 121, 107, 31, 0, 14, 18, 6, 0, 0, 0, 22, 0, 0, 0, 0, 
    23, 7, 0, 0, 5, 16, 0, 0, 0, 0, 20, 30, 37, 44, 46, 55, 47, 0, 0, 18, 38, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 20, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 27, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 27, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=97
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=98
    148, 139, 131, 130, 131, 129, 129, 127, 123, 118, 114, 112, 111, 107, 102, 99, 107, 103, 65, 54, 83, 68, 68, 43, 16, 1, 9, 40, 65, 72, 
    136, 131, 125, 121, 123, 120, 120, 119, 114, 109, 105, 103, 103, 100, 95, 93, 97, 93, 79, 77, 78, 73, 67, 35, 3, 0, 27, 53, 73, 77, 
    121, 120, 115, 109, 111, 111, 110, 108, 103, 99, 95, 95, 95, 94, 90, 88, 90, 87, 83, 81, 73, 64, 64, 40, 14, 24, 45, 65, 75, 79, 
    99, 97, 93, 88, 92, 101, 100, 97, 94, 90, 90, 90, 91, 91, 88, 86, 88, 87, 87, 86, 58, 35, 33, 31, 33, 43, 55, 72, 72, 74, 
    75, 74, 78, 77, 84, 91, 91, 91, 92, 90, 90, 92, 92, 94, 93, 90, 89, 88, 91, 84, 38, 0, 0, 4, 44, 53, 62, 72, 72, 66, 
    72, 73, 80, 83, 88, 87, 88, 90, 95, 95, 94, 97, 98, 100, 95, 93, 92, 86, 88, 76, 22, 0, 0, 6, 42, 63, 66, 69, 71, 68, 
    82, 87, 91, 91, 91, 90, 91, 92, 97, 99, 96, 95, 95, 101, 96, 94, 91, 81, 81, 61, 4, 0, 14, 43, 60, 76, 73, 70, 74, 75, 
    86, 91, 95, 94, 93, 92, 93, 93, 96, 100, 96, 92, 83, 85, 87, 81, 79, 71, 68, 47, 0, 0, 32, 56, 71, 81, 78, 74, 75, 76, 
    87, 91, 95, 94, 94, 93, 93, 91, 92, 93, 83, 77, 61, 61, 72, 73, 81, 82, 71, 52, 5, 0, 16, 24, 44, 64, 72, 74, 73, 72, 
    89, 92, 95, 93, 92, 93, 91, 90, 88, 85, 74, 67, 57, 57, 65, 55, 49, 33, 14, 16, 4, 0, 4, 0, 1, 24, 61, 71, 70, 69, 
    93, 93, 94, 93, 91, 91, 89, 87, 86, 83, 73, 54, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 22, 63, 69, 67, 
    96, 93, 94, 95, 90, 88, 84, 86, 77, 57, 38, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 13, 0, 0, 21, 55, 63, 
    96, 93, 93, 93, 87, 85, 80, 77, 58, 31, 7, 0, 0, 0, 0, 0, 0, 0, 27, 37, 0, 0, 0, 0, 25, 14, 0, 0, 23, 50, 
    94, 93, 92, 88, 83, 77, 78, 57, 37, 4, 5, 6, 0, 0, 0, 17, 23, 34, 64, 52, 0, 0, 0, 0, 1, 27, 4, 0, 9, 42, 
    93, 92, 89, 83, 69, 49, 49, 37, 0, 0, 6, 10, 0, 0, 22, 62, 73, 57, 53, 14, 0, 0, 0, 0, 0, 18, 23, 17, 15, 26, 
    91, 90, 82, 67, 43, 7, 0, 0, 0, 0, 0, 0, 0, 3, 20, 31, 26, 10, 0, 0, 0, 0, 0, 0, 0, 11, 47, 45, 18, 0, 
    89, 89, 83, 58, 36, 4, 0, 0, 0, 0, 0, 0, 12, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 41, 28, 51, 47, 0, 0, 
    88, 91, 84, 48, 15, 0, 0, 0, 0, 0, 3, 0, 30, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 41, 20, 11, 2, 0, 0, 
    94, 93, 66, 17, 0, 0, 0, 0, 0, 0, 6, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    100, 79, 23, 0, 0, 0, 0, 0, 0, 1, 14, 10, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    95, 52, 0, 0, 0, 0, 0, 0, 0, 14, 20, 25, 41, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    90, 39, 0, 0, 0, 0, 0, 0, 0, 21, 11, 4, 16, 0, 0, 0, 0, 0, 0, 0, 0, 17, 18, 0, 0, 0, 0, 0, 0, 0, 
    80, 25, 0, 20, 0, 0, 0, 0, 8, 22, 10, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 30, 0, 0, 0, 0, 0, 0, 24, 
    67, 24, 0, 14, 0, 0, 0, 0, 12, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 22, 0, 0, 0, 0, 10, 22, 
    60, 33, 0, 0, 0, 0, 0, 11, 26, 19, 7, 12, 10, 0, 0, 0, 0, 0, 3, 0, 0, 0, 11, 31, 0, 0, 0, 0, 11, 18, 
    56, 42, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 8, 14, 
    53, 44, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 1, 9, 12, 
    47, 42, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 4, 8, 9, 12, 
    35, 26, 14, 2, 0, 0, 1, 4, 1, 0, 1, 3, 5, 4, 3, 4, 5, 15, 14, 0, 0, 0, 0, 3, 8, 7, 9, 9, 10, 10, 
    26, 20, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 10, 16, 7, 0, 0, 0, 7, 7, 7, 8, 10, 11, 7, 
    
    -- channel=99
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 29, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 49, 33, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 26, 26, 25, 25, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 3, 0, 0, 0, 8, 11, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 25, 28, 41, 69, 99, 104, 84, 69, 39, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 96, 128, 151, 181, 214, 240, 225, 200, 186, 111, 20, 2, 7, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 64, 133, 188, 206, 204, 206, 211, 217, 236, 288, 315, 212, 46, 0, 9, 35, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 63, 101, 131, 153, 150, 126, 119, 112, 97, 142, 277, 382, 331, 141, 0, 0, 22, 35, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 42, 55, 70, 105, 111, 74, 33, 25, 22, 16, 99, 254, 375, 395, 258, 61, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 20, 34, 50, 72, 87, 79, 42, 0, 0, 32, 92, 195, 302, 380, 412, 333, 146, 11, 0, 0, 4, 8, 0, 
    0, 0, 0, 0, 1, 32, 40, 42, 63, 65, 63, 72, 74, 89, 113, 143, 206, 277, 318, 366, 411, 390, 287, 161, 53, 0, 0, 45, 100, 55, 
    0, 0, 0, 0, 6, 52, 71, 92, 79, 38, 40, 52, 90, 198, 295, 328, 348, 371, 393, 418, 406, 298, 163, 98, 50, 7, 35, 130, 193, 134, 
    0, 0, 0, 5, 15, 46, 89, 92, 55, 20, 17, 34, 108, 262, 368, 397, 402, 413, 428, 432, 380, 260, 130, 54, 67, 107, 140, 191, 243, 195, 
    0, 0, 67, 103, 63, 39, 56, 57, 29, 0, 7, 45, 117, 259, 373, 397, 395, 407, 414, 413, 401, 323, 195, 139, 169, 207, 220, 235, 258, 204, 
    0, 70, 198, 201, 118, 54, 47, 39, 0, 0, 0, 40, 133, 270, 365, 381, 384, 369, 321, 299, 336, 357, 313, 270, 265, 275, 281, 270, 232, 149, 
    0, 137, 247, 254, 174, 75, 41, 13, 0, 0, 0, 29, 147, 287, 359, 374, 358, 270, 165, 133, 177, 274, 347, 347, 324, 302, 281, 241, 155, 68, 
    7, 89, 177, 234, 188, 94, 34, 0, 0, 0, 21, 78, 169, 293, 357, 366, 299, 165, 82, 44, 34, 117, 258, 329, 309, 273, 238, 155, 64, 15, 
    0, 22, 91, 175, 186, 109, 28, 0, 0, 6, 82, 134, 205, 310, 369, 354, 246, 116, 46, 12, 0, 11, 124, 249, 277, 248, 169, 73, 15, 0, 
    0, 23, 59, 120, 176, 114, 23, 0, 0, 38, 98, 163, 260, 343, 373, 337, 218, 88, 29, 21, 19, 0, 39, 172, 251, 215, 118, 31, 0, 0, 
    0, 25, 62, 113, 171, 121, 25, 0, 33, 84, 129, 190, 270, 334, 360, 324, 206, 82, 51, 52, 25, 0, 3, 105, 208, 181, 80, 0, 0, 0, 
    0, 15, 65, 117, 166, 133, 58, 57, 114, 181, 223, 251, 296, 343, 361, 326, 205, 81, 73, 97, 74, 24, 0, 44, 135, 126, 38, 0, 0, 0, 
    0, 11, 64, 113, 157, 141, 90, 94, 143, 199, 234, 243, 262, 286, 290, 265, 172, 75, 78, 111, 85, 27, 0, 0, 42, 44, 0, 0, 0, 0, 
    0, 5, 43, 74, 92, 79, 47, 40, 63, 94, 118, 130, 137, 142, 142, 138, 99, 53, 59, 82, 78, 38, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 17, 19, 16, 1, 0, 0, 3, 9, 14, 18, 20, 16, 12, 5, 7, 40, 67, 69, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 3, 14, 30, 39, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 34, 65, 90, 99, 95, 70, 38, 34, 43, 48, 47, 39, 32, 24, 10, 0, 0, 0, 9, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=100
    0, 11, 41, 57, 76, 95, 101, 106, 110, 105, 98, 93, 92, 95, 89, 77, 77, 93, 117, 124, 69, 49, 38, 30, 53, 89, 73, 35, 23, 16, 
    72, 80, 73, 69, 91, 110, 108, 108, 109, 100, 91, 85, 84, 87, 82, 71, 66, 62, 48, 42, 45, 31, 27, 55, 74, 48, 5, 8, 23, 21, 
    88, 77, 66, 71, 91, 101, 97, 94, 93, 88, 80, 73, 71, 72, 66, 57, 51, 46, 40, 20, 0, 0, 23, 49, 38, 0, 0, 0, 14, 20, 
    73, 89, 106, 113, 107, 91, 86, 81, 77, 71, 63, 56, 57, 57, 48, 40, 32, 29, 28, 0, 0, 0, 12, 15, 0, 0, 0, 0, 1, 16, 
    112, 122, 129, 113, 93, 77, 73, 65, 56, 48, 40, 35, 35, 33, 27, 22, 19, 20, 10, 0, 0, 55, 68, 7, 0, 0, 0, 0, 21, 30, 
    111, 99, 79, 57, 49, 51, 48, 41, 33, 28, 26, 22, 20, 14, 11, 10, 6, 3, 0, 0, 72, 149, 111, 38, 0, 0, 9, 50, 54, 45, 
    51, 42, 35, 31, 29, 29, 28, 24, 22, 20, 18, 8, 0, 0, 0, 0, 0, 0, 0, 26, 90, 102, 37, 9, 14, 14, 39, 50, 49, 37, 
    22, 25, 24, 28, 30, 28, 27, 24, 22, 10, 0, 0, 0, 0, 6, 16, 21, 22, 25, 39, 36, 0, 0, 0, 16, 40, 38, 34, 35, 32, 
    20, 27, 28, 30, 32, 33, 34, 30, 26, 13, 10, 12, 17, 22, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 37, 41, 35, 33, 33, 
    21, 27, 28, 29, 31, 32, 37, 33, 30, 30, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 51, 15, 15, 32, 33, 36, 
    23, 27, 28, 28, 29, 30, 34, 30, 12, 0, 0, 0, 0, 0, 0, 42, 115, 193, 216, 56, 0, 0, 0, 37, 79, 35, 4, 20, 33, 35, 
    25, 29, 30, 29, 30, 32, 35, 7, 0, 0, 0, 24, 118, 247, 325, 341, 342, 347, 278, 91, 0, 0, 0, 0, 17, 42, 67, 48, 39, 36, 
    26, 28, 31, 31, 38, 42, 25, 0, 0, 43, 115, 142, 166, 194, 193, 158, 122, 69, 0, 0, 0, 16, 0, 0, 0, 13, 84, 96, 50, 41, 
    30, 29, 32, 28, 16, 0, 0, 0, 46, 97, 69, 21, 31, 45, 1, 0, 0, 0, 0, 0, 0, 11, 28, 0, 0, 0, 24, 31, 0, 0, 
    35, 33, 32, 17, 0, 0, 0, 0, 25, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 183, 194, 38, 0, 0, 0, 0, 0, 
    34, 34, 32, 25, 32, 50, 48, 13, 23, 31, 56, 82, 30, 0, 0, 0, 0, 0, 0, 0, 31, 178, 304, 243, 88, 0, 0, 0, 0, 0, 
    37, 30, 0, 0, 5, 63, 84, 65, 85, 100, 52, 47, 0, 0, 0, 0, 21, 60, 56, 24, 46, 136, 141, 3, 0, 0, 0, 0, 0, 23, 
    35, 0, 0, 0, 0, 8, 23, 59, 102, 79, 0, 0, 0, 0, 0, 99, 85, 59, 43, 39, 24, 0, 0, 0, 0, 0, 0, 0, 2, 98, 
    3, 0, 0, 0, 0, 2, 2, 42, 71, 37, 10, 0, 0, 0, 0, 48, 20, 54, 167, 254, 218, 77, 0, 0, 0, 0, 0, 5, 63, 164, 
    0, 0, 0, 44, 66, 0, 0, 50, 65, 12, 0, 0, 0, 0, 0, 18, 42, 186, 327, 350, 320, 256, 118, 0, 0, 16, 40, 86, 178, 225, 
    0, 44, 210, 243, 111, 15, 7, 51, 44, 0, 0, 0, 0, 0, 0, 17, 110, 252, 236, 110, 93, 152, 175, 130, 96, 92, 120, 199, 245, 176, 
    21, 96, 186, 133, 63, 31, 29, 42, 0, 0, 0, 0, 0, 0, 0, 11, 138, 198, 75, 0, 0, 19, 71, 134, 110, 85, 135, 200, 157, 27, 
    37, 39, 0, 0, 0, 38, 31, 16, 0, 0, 0, 0, 0, 0, 0, 42, 142, 114, 0, 0, 0, 10, 10, 45, 49, 49, 123, 132, 29, 0, 
    43, 21, 0, 0, 0, 62, 37, 0, 0, 0, 0, 0, 0, 0, 46, 78, 131, 64, 0, 0, 0, 0, 3, 4, 53, 104, 144, 92, 8, 0, 
    29, 10, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 4, 30, 87, 37, 0, 0, 0, 0, 0, 1, 82, 168, 158, 69, 18, 22, 
    9, 0, 0, 0, 0, 49, 0, 0, 0, 0, 10, 26, 54, 120, 143, 159, 164, 61, 0, 0, 27, 25, 23, 29, 114, 193, 133, 35, 7, 9, 
    0, 0, 21, 42, 97, 163, 141, 115, 163, 234, 295, 323, 329, 342, 347, 341, 296, 127, 0, 26, 80, 65, 39, 40, 75, 123, 71, 6, 0, 0, 
    0, 0, 38, 93, 123, 125, 80, 66, 88, 108, 128, 144, 156, 167, 172, 173, 162, 94, 30, 18, 0, 27, 28, 20, 10, 17, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 81, 85, 81, 59, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 58, 13, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=101
    146, 156, 163, 175, 183, 184, 186, 186, 181, 176, 172, 173, 172, 165, 159, 156, 154, 152, 142, 145, 129, 124, 110, 96, 86, 93, 109, 113, 107, 102, 
    177, 173, 167, 175, 179, 182, 181, 178, 172, 165, 160, 160, 161, 156, 150, 146, 141, 129, 125, 125, 122, 117, 111, 91, 70, 76, 97, 112, 108, 105, 
    170, 162, 155, 160, 166, 169, 167, 164, 159, 152, 148, 147, 148, 144, 139, 134, 133, 126, 121, 111, 97, 92, 85, 73, 66, 60, 87, 104, 104, 104, 
    157, 159, 161, 159, 161, 157, 153, 151, 147, 141, 136, 136, 137, 134, 129, 124, 124, 122, 116, 92, 72, 53, 51, 66, 65, 63, 85, 94, 98, 101, 
    158, 161, 159, 154, 150, 146, 140, 139, 135, 129, 125, 125, 126, 124, 122, 118, 117, 117, 111, 97, 77, 61, 62, 70, 62, 78, 92, 102, 106, 106, 
    150, 144, 137, 134, 131, 132, 127, 126, 125, 122, 119, 117, 117, 115, 115, 115, 110, 107, 108, 102, 81, 85, 96, 85, 80, 98, 109, 118, 118, 112, 
    127, 124, 122, 121, 119, 120, 117, 119, 121, 120, 118, 112, 107, 101, 101, 103, 104, 101, 104, 90, 64, 74, 89, 98, 104, 110, 117, 122, 118, 112, 
    117, 118, 119, 120, 118, 119, 116, 118, 120, 114, 110, 104, 100, 104, 106, 108, 110, 105, 97, 65, 34, 38, 61, 96, 111, 113, 116, 117, 115, 111, 
    116, 119, 120, 121, 121, 122, 119, 120, 120, 116, 113, 104, 104, 105, 89, 67, 38, 10, 5, 0, 0, 16, 53, 93, 99, 108, 115, 115, 114, 111, 
    117, 119, 119, 120, 120, 123, 121, 121, 124, 121, 100, 65, 33, 9, 0, 0, 0, 0, 0, 0, 0, 0, 52, 107, 90, 96, 99, 109, 113, 112, 
    119, 118, 118, 118, 119, 121, 120, 119, 106, 82, 50, 30, 19, 28, 48, 73, 100, 119, 80, 16, 0, 0, 7, 80, 104, 89, 85, 93, 110, 112, 
    120, 119, 117, 117, 119, 119, 118, 101, 83, 68, 65, 80, 103, 131, 159, 169, 175, 166, 127, 88, 1, 0, 0, 15, 93, 101, 92, 90, 106, 112, 
    118, 119, 118, 119, 119, 115, 108, 93, 89, 89, 101, 106, 95, 91, 111, 111, 99, 62, 40, 37, 0, 0, 0, 0, 41, 102, 100, 100, 105, 111, 
    118, 119, 120, 117, 97, 89, 83, 91, 80, 83, 74, 64, 42, 35, 44, 48, 14, 0, 0, 0, 0, 0, 0, 0, 6, 62, 79, 71, 68, 80, 
    120, 120, 117, 109, 81, 62, 61, 46, 57, 55, 61, 54, 21, 0, 0, 0, 0, 0, 0, 0, 0, 26, 32, 24, 39, 40, 43, 23, 4, 24, 
    120, 119, 113, 106, 102, 90, 68, 46, 49, 63, 92, 89, 31, 0, 0, 0, 0, 0, 0, 0, 16, 54, 78, 102, 64, 23, 1, 0, 0, 0, 
    120, 115, 89, 69, 64, 81, 75, 73, 58, 77, 77, 70, 44, 29, 0, 0, 10, 14, 6, 0, 0, 1, 25, 44, 11, 0, 0, 0, 0, 8, 
    116, 78, 36, 0, 0, 43, 64, 68, 63, 71, 55, 31, 31, 44, 24, 22, 19, 17, 14, 9, 0, 0, 0, 0, 0, 0, 0, 1, 29, 33, 
    94, 35, 0, 0, 0, 27, 54, 55, 58, 74, 77, 55, 47, 39, 10, 0, 2, 33, 72, 108, 81, 0, 0, 0, 0, 0, 0, 15, 52, 58, 
    88, 67, 26, 0, 0, 13, 53, 55, 64, 67, 65, 58, 53, 37, 3, 0, 29, 68, 116, 167, 179, 120, 42, 0, 0, 4, 20, 52, 78, 85, 
    115, 128, 104, 72, 21, 12, 49, 54, 64, 39, 14, 0, 12, 16, 0, 7, 47, 52, 84, 86, 113, 141, 110, 57, 23, 29, 62, 83, 94, 95, 
    119, 94, 100, 77, 25, 18, 41, 52, 51, 33, 19, 0, 0, 0, 0, 8, 22, 32, 62, 44, 51, 101, 112, 83, 34, 34, 60, 71, 81, 74, 
    101, 44, 43, 35, 16, 15, 33, 46, 35, 33, 34, 16, 20, 0, 0, 7, 2, 26, 43, 37, 43, 67, 97, 76, 34, 25, 37, 57, 69, 66, 
    95, 51, 37, 36, 24, 17, 29, 39, 22, 12, 5, 8, 25, 11, 12, 8, 0, 24, 30, 22, 24, 45, 83, 85, 62, 38, 41, 68, 79, 81, 
    89, 61, 43, 43, 21, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 31, 9, 3, 17, 64, 92, 92, 64, 60, 77, 84, 86, 
    82, 58, 41, 39, 34, 14, 13, 23, 31, 35, 30, 40, 52, 61, 65, 46, 26, 33, 56, 40, 35, 34, 63, 100, 113, 89, 76, 74, 76, 79, 
    77, 74, 63, 75, 83, 82, 92, 106, 126, 148, 157, 162, 162, 163, 165, 145, 103, 72, 64, 59, 47, 56, 56, 88, 97, 88, 77, 70, 70, 71, 
    70, 71, 72, 89, 86, 79, 78, 78, 88, 96, 101, 106, 109, 111, 114, 113, 99, 100, 72, 48, 39, 43, 52, 70, 70, 68, 67, 66, 63, 64, 
    71, 55, 36, 27, 15, 6, 6, 14, 25, 27, 24, 27, 32, 35, 40, 45, 50, 73, 87, 84, 75, 63, 66, 63, 60, 60, 60, 60, 58, 60, 
    64, 37, 0, 0, 0, 0, 0, 1, 10, 7, 3, 3, 5, 6, 8, 13, 20, 31, 47, 58, 59, 56, 56, 52, 50, 50, 51, 51, 53, 57, 
    
    -- channel=102
    136, 165, 183, 200, 214, 224, 229, 232, 227, 219, 212, 208, 206, 199, 189, 181, 189, 208, 176, 168, 144, 126, 116, 106, 107, 104, 91, 87, 92, 93, 
    214, 210, 197, 202, 214, 227, 228, 226, 219, 207, 197, 192, 191, 186, 177, 167, 164, 150, 130, 131, 127, 117, 115, 110, 74, 52, 53, 79, 98, 101, 
    211, 193, 179, 190, 202, 211, 209, 205, 199, 188, 178, 174, 172, 168, 159, 149, 145, 136, 124, 112, 95, 84, 86, 76, 40, 15, 34, 70, 99, 101, 
    187, 193, 206, 206, 201, 194, 189, 183, 176, 166, 156, 153, 154, 149, 140, 130, 125, 124, 115, 76, 51, 41, 46, 39, 27, 16, 31, 59, 88, 95, 
    204, 210, 208, 191, 180, 174, 167, 159, 150, 141, 133, 131, 133, 128, 122, 115, 115, 115, 104, 82, 86, 74, 53, 34, 13, 21, 47, 83, 102, 105, 
    183, 171, 157, 146, 144, 144, 139, 134, 129, 126, 124, 121, 120, 115, 114, 110, 106, 101, 93, 117, 131, 112, 81, 50, 36, 59, 103, 129, 126, 115, 
    134, 130, 127, 126, 125, 124, 121, 121, 122, 124, 122, 115, 108, 93, 91, 88, 87, 87, 96, 120, 100, 68, 58, 59, 80, 106, 124, 129, 123, 114, 
    115, 121, 124, 128, 126, 125, 123, 123, 124, 116, 103, 88, 90, 91, 102, 111, 116, 111, 111, 90, 27, 0, 0, 51, 102, 121, 120, 118, 117, 112, 
    116, 124, 128, 131, 131, 131, 131, 129, 128, 119, 117, 109, 112, 109, 95, 55, 0, 0, 0, 0, 0, 0, 0, 56, 92, 106, 114, 115, 115, 112, 
    119, 126, 128, 129, 130, 132, 133, 130, 133, 136, 120, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 94, 87, 78, 78, 102, 114, 114, 
    124, 128, 127, 126, 127, 129, 130, 127, 115, 80, 15, 0, 0, 0, 33, 90, 154, 206, 153, 3, 0, 0, 0, 66, 89, 69, 68, 79, 107, 110, 
    128, 129, 127, 126, 127, 129, 127, 103, 68, 41, 52, 106, 173, 234, 284, 297, 303, 292, 208, 96, 0, 0, 0, 0, 65, 83, 93, 86, 100, 107, 
    127, 128, 128, 131, 134, 133, 113, 82, 84, 120, 159, 164, 153, 147, 151, 131, 118, 58, 0, 0, 0, 0, 0, 0, 0, 79, 99, 102, 96, 102, 
    127, 129, 130, 129, 110, 89, 62, 97, 117, 117, 71, 49, 34, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 57, 41, 23, 38, 
    131, 132, 128, 117, 74, 41, 41, 56, 53, 23, 28, 37, 4, 0, 0, 0, 0, 0, 0, 0, 0, 37, 75, 39, 14, 0, 0, 0, 0, 0, 
    131, 133, 126, 122, 116, 102, 83, 30, 26, 46, 89, 101, 1, 0, 0, 0, 0, 0, 0, 0, 28, 132, 175, 135, 59, 0, 0, 0, 0, 0, 
    134, 128, 91, 73, 73, 90, 72, 74, 66, 78, 68, 62, 0, 0, 0, 0, 38, 51, 29, 5, 33, 46, 19, 10, 0, 0, 0, 0, 0, 0, 
    131, 75, 0, 0, 0, 22, 52, 76, 60, 54, 20, 0, 0, 16, 50, 63, 51, 32, 23, 23, 0, 0, 0, 0, 0, 0, 0, 0, 22, 38, 
    93, 0, 0, 0, 0, 0, 29, 45, 40, 49, 50, 29, 12, 26, 21, 10, 1, 52, 139, 205, 145, 0, 0, 0, 0, 0, 0, 4, 67, 90, 
    70, 40, 36, 8, 0, 0, 23, 43, 42, 36, 39, 31, 11, 19, 4, 0, 45, 151, 244, 293, 282, 189, 70, 0, 0, 0, 23, 72, 136, 133, 
    123, 210, 215, 138, 27, 0, 27, 33, 30, 0, 0, 0, 0, 0, 0, 5, 99, 135, 127, 93, 142, 187, 165, 105, 57, 57, 92, 146, 157, 100, 
    159, 192, 162, 88, 16, 0, 17, 22, 5, 0, 0, 0, 0, 0, 0, 10, 70, 43, 30, 4, 33, 110, 141, 136, 65, 46, 98, 114, 78, 30, 
    136, 63, 16, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 25, 25, 2, 5, 0, 1, 48, 97, 89, 39, 32, 56, 48, 23, 16, 
    118, 53, 11, 5, 9, 0, 0, 0, 0, 0, 0, 0, 0, 13, 27, 30, 4, 0, 0, 0, 0, 12, 66, 79, 76, 65, 51, 43, 43, 53, 
    98, 63, 30, 21, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 86, 122, 102, 65, 55, 58, 65, 
    78, 48, 23, 15, 15, 0, 0, 0, 0, 10, 23, 53, 85, 107, 119, 98, 55, 14, 21, 10, 20, 11, 44, 99, 148, 125, 71, 43, 44, 50, 
    66, 62, 62, 83, 109, 111, 112, 138, 187, 235, 262, 276, 283, 287, 289, 251, 166, 73, 54, 57, 45, 36, 26, 81, 107, 86, 48, 29, 31, 34, 
    48, 69, 84, 115, 117, 92, 74, 77, 96, 113, 125, 135, 142, 147, 152, 146, 110, 86, 59, 38, 4, 14, 25, 40, 37, 30, 25, 22, 18, 19, 
    55, 45, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 44, 72, 80, 86, 64, 40, 19, 14, 13, 13, 12, 6, 12, 
    48, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 38, 45, 24, 9, 0, 0, 0, 0, 0, 1, 11, 
    
    -- channel=103
    32, 29, 27, 29, 31, 30, 29, 29, 27, 26, 25, 26, 29, 31, 31, 32, 22, 10, 30, 59, 48, 50, 42, 36, 44, 68, 92, 77, 53, 47, 
    18, 25, 27, 26, 22, 17, 11, 7, 7, 9, 12, 15, 19, 22, 24, 27, 24, 24, 36, 45, 45, 41, 38, 45, 68, 90, 95, 72, 45, 39, 
    12, 22, 22, 17, 10, 5, 0, 0, 0, 3, 8, 11, 13, 17, 22, 26, 27, 27, 35, 34, 32, 40, 49, 65, 87, 91, 85, 58, 35, 33, 
    14, 15, 7, 4, 5, 0, 0, 0, 4, 8, 10, 11, 12, 18, 25, 28, 30, 30, 33, 28, 30, 40, 55, 83, 90, 84, 78, 52, 36, 30, 
    13, 6, 4, 7, 7, 2, 1, 9, 13, 14, 13, 12, 13, 19, 30, 30, 29, 32, 31, 24, 30, 50, 74, 93, 92, 86, 68, 48, 37, 30, 
    20, 17, 13, 13, 9, 9, 9, 16, 18, 16, 13, 8, 9, 15, 25, 29, 31, 34, 33, 20, 30, 74, 104, 107, 85, 68, 48, 38, 36, 36, 
    23, 17, 13, 14, 11, 13, 12, 17, 15, 12, 8, 4, 10, 18, 24, 31, 37, 35, 30, 22, 48, 96, 108, 99, 66, 41, 36, 35, 35, 35, 
    19, 12, 8, 9, 8, 10, 8, 11, 10, 6, 10, 17, 23, 22, 20, 23, 26, 27, 26, 31, 68, 109, 104, 79, 44, 33, 35, 35, 34, 32, 
    14, 7, 4, 5, 3, 5, 3, 7, 5, 4, 14, 22, 30, 23, 15, 25, 32, 35, 39, 49, 85, 107, 92, 70, 46, 40, 39, 37, 36, 31, 
    9, 3, 0, 4, 4, 4, 4, 7, 4, 0, 4, 18, 41, 45, 44, 56, 57, 49, 42, 50, 83, 90, 83, 80, 66, 60, 48, 40, 36, 31, 
    5, 1, 0, 4, 4, 6, 7, 8, 1, 1, 24, 48, 56, 52, 45, 41, 30, 23, 38, 71, 88, 77, 73, 80, 93, 82, 53, 41, 39, 35, 
    3, 1, 0, 2, 3, 7, 11, 5, 10, 25, 34, 26, 22, 29, 35, 42, 44, 39, 51, 74, 79, 79, 83, 78, 92, 84, 69, 46, 46, 41, 
    2, 3, 0, 0, 1, 4, 8, 11, 23, 19, 18, 30, 47, 60, 75, 84, 84, 78, 80, 66, 43, 64, 81, 78, 90, 86, 78, 65, 58, 54, 
    2, 3, 0, 0, 0, 6, 15, 15, 17, 40, 64, 69, 71, 90, 99, 97, 100, 104, 97, 53, 23, 46, 75, 78, 85, 88, 83, 87, 80, 71, 
    0, 0, 0, 0, 10, 24, 21, 19, 53, 85, 80, 71, 73, 94, 111, 108, 110, 110, 68, 30, 36, 44, 52, 75, 85, 72, 82, 99, 99, 74, 
    0, 0, 0, 3, 20, 40, 40, 58, 86, 80, 86, 84, 89, 112, 117, 92, 69, 43, 27, 34, 44, 31, 35, 72, 70, 54, 79, 98, 80, 64, 
    0, 0, 0, 11, 28, 55, 75, 80, 79, 92, 95, 95, 96, 95, 58, 32, 27, 25, 34, 38, 28, 34, 68, 61, 44, 62, 72, 61, 49, 64, 
    0, 0, 12, 38, 50, 70, 73, 78, 90, 105, 99, 104, 80, 50, 29, 31, 34, 39, 41, 36, 42, 62, 63, 53, 50, 51, 45, 36, 47, 69, 
    0, 0, 31, 33, 53, 75, 78, 88, 95, 100, 95, 92, 70, 46, 36, 42, 45, 43, 31, 31, 48, 64, 56, 46, 40, 38, 46, 53, 55, 66, 
    0, 6, 11, 28, 75, 83, 83, 89, 99, 101, 88, 84, 74, 59, 43, 45, 47, 29, 22, 45, 57, 61, 59, 42, 40, 50, 56, 60, 56, 72, 
    0, 0, 0, 58, 88, 85, 86, 93, 107, 103, 102, 95, 71, 56, 47, 49, 45, 35, 72, 91, 69, 56, 61, 49, 37, 44, 62, 60, 66, 101, 
    0, 0, 31, 80, 93, 88, 90, 101, 107, 104, 105, 86, 59, 49, 49, 50, 52, 75, 110, 98, 88, 66, 50, 52, 46, 58, 63, 69, 103, 111, 
    0, 27, 71, 67, 85, 85, 89, 107, 107, 94, 79, 68, 68, 56, 45, 50, 68, 92, 94, 86, 101, 90, 60, 61, 63, 60, 69, 95, 112, 100, 
    10, 42, 72, 62, 78, 88, 93, 105, 103, 86, 74, 73, 64, 43, 42, 55, 81, 94, 94, 91, 88, 89, 75, 64, 68, 64, 80, 104, 103, 90, 
    24, 39, 62, 63, 74, 86, 92, 102, 98, 86, 79, 67, 50, 46, 51, 63, 83, 85, 86, 86, 85, 90, 83, 68, 71, 76, 91, 101, 96, 89, 
    36, 41, 59, 63, 76, 91, 95, 95, 85, 73, 65, 51, 43, 48, 46, 53, 73, 78, 84, 83, 80, 80, 87, 76, 78, 90, 104, 104, 97, 92, 
    43, 44, 57, 63, 71, 83, 87, 75, 64, 57, 54, 53, 52, 51, 50, 61, 87, 88, 76, 65, 77, 93, 100, 90, 87, 107, 118, 109, 101, 97, 
    49, 39, 47, 66, 76, 92, 96, 90, 89, 87, 84, 83, 83, 83, 80, 84, 99, 102, 89, 76, 84, 96, 96, 107, 107, 113, 114, 111, 109, 105, 
    49, 46, 55, 78, 100, 114, 111, 103, 106, 107, 106, 108, 107, 105, 102, 104, 108, 97, 85, 91, 80, 84, 108, 115, 113, 112, 113, 114, 114, 111, 
    50, 53, 71, 92, 100, 99, 95, 94, 102, 105, 104, 106, 106, 105, 104, 105, 108, 104, 88, 79, 87, 105, 117, 115, 112, 112, 112, 113, 112, 109, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 36, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 44, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 31, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 86, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 98, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 87, 85, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 100, 94, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 95, 115, 170, 79, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 50, 231, 205, 40, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 21, 0, 18, 40, 0, 0, 0, 197, 285, 161, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 118, 85, 21, 38, 63, 0, 0, 0, 116, 268, 260, 105, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 81, 129, 98, 22, 7, 17, 0, 0, 11, 72, 206, 287, 160, 62, 27, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 35, 0, 5, 70, 74, 58, 38, 2, 1, 0, 13, 56, 98, 184, 194, 131, 98, 40, 0, 0, 32, 
    0, 0, 0, 0, 0, 0, 0, 21, 82, 65, 1, 15, 10, 0, 0, 26, 6, 9, 25, 47, 78, 162, 181, 79, 44, 81, 14, 0, 0, 99, 
    0, 0, 0, 0, 10, 2, 16, 55, 100, 91, 29, 43, 0, 0, 0, 28, 22, 23, 32, 40, 105, 207, 180, 40, 0, 41, 13, 0, 0, 119, 
    0, 0, 0, 11, 135, 81, 34, 76, 115, 82, 26, 41, 0, 0, 0, 65, 50, 37, 34, 30, 74, 187, 178, 53, 11, 32, 37, 29, 31, 120, 
    0, 0, 0, 97, 222, 136, 53, 93, 125, 63, 23, 14, 0, 0, 17, 79, 59, 73, 81, 26, 0, 50, 123, 87, 60, 66, 68, 68, 78, 129, 
    0, 0, 0, 128, 241, 170, 75, 104, 111, 56, 38, 19, 0, 0, 43, 72, 84, 158, 147, 49, 0, 0, 1, 82, 101, 99, 84, 93, 126, 117, 
    0, 0, 0, 68, 185, 181, 104, 113, 93, 37, 32, 49, 0, 0, 53, 70, 149, 229, 151, 79, 39, 0, 0, 26, 115, 105, 99, 138, 135, 72, 
    0, 0, 47, 0, 116, 192, 127, 110, 72, 13, 8, 46, 0, 0, 62, 94, 217, 235, 104, 69, 82, 17, 0, 0, 95, 119, 150, 161, 100, 24, 
    0, 29, 83, 0, 71, 204, 145, 93, 54, 18, 21, 31, 0, 0, 68, 121, 249, 209, 66, 76, 87, 80, 0, 0, 50, 143, 189, 149, 47, 0, 
    0, 7, 67, 8, 55, 204, 158, 70, 34, 34, 57, 31, 0, 9, 68, 131, 254, 179, 43, 88, 104, 102, 24, 0, 1, 156, 198, 111, 11, 0, 
    0, 0, 52, 25, 53, 193, 160, 61, 27, 43, 81, 61, 9, 45, 74, 137, 259, 173, 23, 70, 127, 133, 74, 0, 0, 148, 178, 79, 8, 0, 
    0, 0, 42, 39, 53, 161, 136, 50, 20, 20, 46, 49, 25, 44, 53, 103, 217, 157, 17, 45, 120, 135, 99, 10, 0, 114, 130, 64, 24, 5, 
    0, 0, 27, 43, 60, 119, 101, 51, 35, 27, 32, 37, 35, 42, 45, 64, 134, 92, 17, 58, 101, 128, 114, 62, 33, 79, 85, 57, 41, 20, 
    0, 6, 37, 62, 73, 98, 94, 82, 74, 68, 70, 69, 68, 71, 72, 69, 82, 39, 0, 56, 88, 128, 114, 73, 56, 64, 59, 50, 44, 28, 
    0, 18, 64, 86, 89, 93, 115, 117, 93, 86, 91, 90, 89, 86, 86, 81, 76, 51, 0, 28, 83, 106, 98, 66, 60, 59, 55, 49, 40, 32, 
    0, 17, 62, 98, 110, 112, 142, 143, 105, 101, 104, 101, 101, 97, 98, 96, 91, 85, 61, 54, 92, 108, 82, 62, 62, 65, 60, 51, 43, 41, 
    
    -- channel=105
    73, 82, 84, 88, 95, 100, 101, 102, 100, 97, 94, 93, 95, 95, 92, 91, 91, 104, 109, 117, 100, 92, 86, 70, 80, 96, 93, 84, 82, 80, 
    88, 94, 90, 88, 91, 93, 89, 87, 86, 84, 82, 82, 85, 87, 86, 85, 83, 82, 86, 90, 84, 80, 88, 88, 98, 103, 89, 82, 79, 77, 
    82, 81, 75, 73, 77, 80, 76, 74, 75, 74, 74, 73, 77, 80, 80, 79, 79, 75, 79, 79, 68, 64, 79, 91, 98, 84, 73, 70, 70, 69, 
    69, 69, 71, 74, 75, 71, 69, 71, 73, 73, 71, 69, 72, 76, 77, 75, 77, 75, 76, 69, 49, 36, 55, 80, 84, 70, 66, 66, 65, 62, 
    79, 83, 85, 81, 74, 68, 67, 72, 74, 71, 66, 64, 69, 73, 75, 72, 74, 72, 69, 66, 56, 57, 67, 73, 72, 69, 64, 68, 70, 69, 
    91, 86, 78, 73, 68, 68, 68, 69, 69, 66, 61, 58, 61, 65, 69, 66, 68, 67, 68, 77, 87, 109, 111, 96, 80, 76, 77, 80, 84, 80, 
    74, 69, 65, 66, 62, 64, 63, 63, 62, 61, 59, 53, 49, 50, 58, 60, 63, 61, 68, 85, 98, 115, 108, 94, 83, 83, 86, 82, 81, 77, 
    60, 60, 59, 63, 59, 61, 60, 59, 58, 56, 56, 53, 46, 43, 51, 58, 62, 61, 70, 79, 83, 85, 67, 64, 66, 71, 77, 76, 75, 73, 
    58, 59, 58, 60, 58, 60, 59, 58, 56, 52, 54, 57, 55, 51, 49, 44, 32, 15, 21, 28, 40, 49, 46, 55, 54, 57, 69, 75, 73, 71, 
    58, 57, 56, 59, 57, 59, 61, 60, 59, 59, 61, 56, 33, 8, 0, 0, 0, 0, 0, 0, 0, 20, 60, 87, 67, 56, 57, 72, 73, 72, 
    57, 56, 55, 58, 58, 60, 62, 61, 55, 48, 37, 15, 0, 0, 0, 9, 33, 58, 64, 32, 0, 0, 43, 104, 104, 66, 48, 57, 70, 72, 
    56, 55, 54, 56, 60, 61, 62, 56, 44, 26, 19, 34, 69, 111, 145, 169, 184, 187, 167, 112, 32, 0, 10, 59, 105, 90, 64, 51, 63, 72, 
    56, 56, 54, 54, 60, 61, 58, 48, 42, 52, 87, 116, 126, 138, 152, 147, 138, 116, 85, 50, 16, 0, 0, 19, 74, 104, 95, 79, 70, 74, 
    55, 56, 55, 55, 52, 46, 41, 48, 60, 89, 95, 89, 80, 80, 83, 81, 69, 35, 2, 0, 0, 8, 0, 4, 47, 89, 104, 90, 67, 62, 
    55, 55, 56, 57, 42, 23, 24, 44, 72, 72, 63, 65, 66, 56, 31, 3, 0, 0, 0, 0, 6, 31, 51, 61, 64, 70, 85, 63, 25, 18, 
    54, 53, 56, 62, 60, 53, 53, 55, 65, 75, 95, 98, 71, 20, 0, 0, 0, 0, 0, 2, 25, 63, 115, 128, 86, 62, 52, 25, 0, 0, 
    53, 53, 52, 61, 71, 93, 95, 85, 88, 114, 117, 115, 79, 30, 0, 0, 10, 25, 29, 21, 29, 62, 85, 69, 35, 12, 0, 0, 1, 17, 
    56, 42, 23, 14, 25, 64, 85, 97, 105, 112, 95, 78, 49, 37, 37, 48, 48, 41, 31, 23, 8, 0, 0, 0, 0, 0, 0, 9, 38, 46, 
    50, 16, 0, 0, 18, 59, 80, 90, 97, 105, 98, 81, 54, 38, 34, 35, 29, 35, 57, 85, 68, 10, 0, 0, 0, 0, 19, 36, 59, 76, 
    43, 15, 0, 13, 42, 50, 75, 89, 101, 104, 100, 95, 72, 48, 30, 27, 38, 71, 132, 182, 176, 120, 53, 5, 8, 27, 41, 61, 89, 114, 
    59, 70, 88, 101, 69, 53, 80, 96, 106, 88, 68, 48, 36, 35, 30, 32, 61, 99, 142, 139, 143, 149, 117, 66, 43, 55, 76, 100, 128, 133, 
    78, 104, 137, 124, 77, 59, 78, 94, 94, 71, 45, 17, 14, 21, 20, 34, 67, 94, 101, 75, 85, 113, 119, 103, 71, 67, 88, 116, 130, 105, 
    79, 78, 77, 64, 58, 57, 78, 93, 80, 63, 59, 52, 42, 20, 14, 35, 61, 79, 80, 80, 87, 94, 103, 96, 65, 55, 80, 104, 100, 82, 
    78, 69, 60, 57, 59, 61, 74, 82, 64, 47, 46, 45, 37, 29, 37, 49, 63, 69, 64, 57, 60, 80, 98, 95, 79, 68, 85, 99, 95, 90, 
    79, 76, 73, 68, 60, 59, 60, 56, 33, 11, 0, 4, 16, 32, 37, 38, 51, 61, 62, 51, 47, 60, 86, 100, 107, 101, 103, 105, 100, 97, 
    75, 73, 73, 67, 65, 58, 49, 42, 31, 22, 17, 22, 36, 51, 54, 56, 66, 68, 72, 56, 52, 61, 88, 110, 128, 128, 118, 104, 96, 93, 
    71, 75, 78, 85, 99, 108, 111, 116, 133, 151, 162, 166, 166, 167, 167, 158, 138, 103, 88, 88, 93, 98, 99, 116, 133, 136, 119, 101, 96, 94, 
    63, 75, 93, 114, 128, 134, 131, 131, 140, 147, 152, 156, 160, 161, 161, 160, 150, 126, 94, 78, 72, 78, 91, 108, 109, 110, 106, 101, 98, 93, 
    60, 65, 71, 80, 78, 65, 56, 60, 71, 71, 70, 72, 77, 81, 84, 88, 94, 103, 106, 97, 86, 93, 107, 103, 99, 98, 99, 99, 95, 91, 
    64, 58, 43, 26, 18, 19, 32, 47, 57, 55, 51, 51, 52, 53, 53, 57, 65, 73, 82, 95, 104, 106, 101, 94, 91, 91, 91, 91, 90, 90, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 35, 47, 36, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 55, 52, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 50, 32, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 25, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 19, 30, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 76, 77, 33, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 49, 73, 52, 14, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 38, 31, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 69, 83, 47, 0, 0, 0, 43, 72, 30, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 52, 94, 135, 154, 156, 163, 160, 108, 11, 0, 0, 0, 64, 70, 32, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 47, 76, 86, 92, 105, 108, 98, 78, 60, 18, 0, 0, 0, 0, 17, 72, 73, 42, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 40, 44, 43, 41, 48, 47, 38, 24, 0, 0, 0, 0, 0, 0, 0, 0, 40, 70, 59, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 23, 26, 29, 31, 14, 0, 0, 0, 0, 0, 0, 0, 0, 21, 56, 39, 23, 55, 32, 0, 0, 
    0, 0, 0, 0, 13, 30, 32, 23, 30, 37, 66, 73, 63, 3, 0, 0, 0, 0, 0, 0, 0, 17, 75, 104, 74, 29, 8, 0, 0, 0, 
    0, 0, 0, 0, 6, 50, 71, 65, 63, 82, 82, 73, 53, 22, 0, 0, 0, 0, 0, 0, 0, 0, 11, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 39, 69, 71, 72, 90, 77, 56, 27, 18, 4, 12, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 30, 62, 64, 66, 81, 86, 85, 63, 29, 3, 5, 1, 5, 43, 99, 102, 36, 0, 0, 0, 0, 0, 0, 15, 34, 
    0, 0, 0, 0, 12, 21, 51, 64, 75, 78, 76, 78, 69, 39, 3, 0, 8, 45, 120, 172, 177, 159, 84, 0, 0, 3, 17, 28, 59, 83, 
    7, 53, 100, 127, 62, 24, 49, 62, 79, 66, 42, 11, 6, 13, 2, 0, 21, 66, 117, 101, 96, 132, 147, 85, 36, 39, 50, 74, 102, 97, 
    26, 68, 109, 121, 64, 25, 48, 65, 69, 55, 38, 14, 6, 0, 0, 0, 15, 57, 83, 55, 61, 81, 114, 119, 60, 39, 53, 79, 93, 60, 
    31, 51, 57, 52, 45, 24, 42, 64, 56, 44, 44, 43, 30, 0, 0, 0, 12, 45, 54, 40, 50, 65, 86, 105, 63, 26, 43, 69, 62, 35, 
    37, 54, 53, 49, 48, 34, 46, 59, 47, 27, 19, 22, 22, 9, 16, 14, 15, 37, 45, 30, 27, 46, 72, 94, 84, 51, 57, 70, 57, 46, 
    37, 55, 62, 61, 52, 32, 25, 24, 1, 0, 0, 0, 0, 0, 0, 0, 0, 28, 48, 26, 3, 18, 51, 85, 105, 88, 82, 78, 62, 56, 
    30, 50, 58, 54, 55, 49, 42, 41, 43, 48, 48, 48, 53, 68, 75, 71, 59, 52, 58, 53, 49, 45, 64, 85, 119, 122, 102, 78, 64, 59, 
    20, 42, 68, 81, 97, 111, 119, 124, 140, 160, 175, 182, 182, 182, 182, 174, 151, 108, 74, 56, 70, 64, 62, 84, 102, 110, 94, 74, 66, 61, 
    11, 29, 60, 94, 108, 109, 97, 96, 107, 113, 117, 123, 126, 129, 130, 128, 121, 109, 93, 68, 41, 49, 58, 77, 77, 77, 72, 68, 65, 58, 
    17, 31, 41, 45, 40, 27, 17, 28, 48, 50, 43, 40, 43, 48, 51, 53, 55, 66, 82, 100, 88, 78, 79, 69, 66, 65, 64, 63, 60, 53, 
    25, 30, 21, 3, 0, 0, 14, 31, 41, 37, 32, 26, 22, 21, 22, 23, 27, 37, 50, 64, 72, 70, 66, 59, 56, 56, 57, 56, 53, 51, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 16, 6, 4, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 10, 9, 6, 6, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 6, 5, 5, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 4, 3, 2, 2, 0, 0, 
    
    -- channel=108
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 35, 19, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 41, 53, 57, 29, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 9, 22, 37, 29, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 23, 22, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 12, 29, 52, 76, 53, 24, 32, 17, 35, 53, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 92, 117, 142, 178, 212, 237, 200, 184, 144, 27, 4, 35, 60, 41, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 72, 138, 185, 203, 215, 217, 212, 197, 200, 277, 258, 95, 0, 0, 56, 77, 35, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 28, 67, 103, 138, 133, 103, 93, 90, 71, 41, 110, 250, 272, 178, 40, 0, 7, 73, 58, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 21, 46, 55, 67, 84, 56, 22, 9, 22, 9, 6, 122, 231, 262, 245, 123, 0, 0, 27, 36, 25, 4, 0, 
    0, 0, 0, 0, 0, 0, 9, 25, 40, 48, 65, 73, 41, 15, 0, 3, 25, 90, 188, 238, 267, 278, 178, 60, 13, 0, 4, 31, 30, 0, 
    0, 0, 0, 0, 24, 60, 63, 57, 66, 63, 94, 91, 67, 92, 101, 111, 159, 220, 253, 267, 283, 236, 128, 86, 33, 0, 1, 84, 93, 14, 
    0, 0, 0, 0, 22, 76, 98, 108, 69, 62, 74, 70, 112, 231, 265, 273, 295, 299, 292, 287, 243, 120, 31, 32, 8, 0, 52, 140, 157, 63, 
    0, 0, 0, 0, 1, 52, 92, 87, 44, 38, 47, 48, 138, 275, 301, 293, 287, 290, 294, 291, 214, 81, 4, 15, 50, 80, 131, 169, 191, 99, 
    0, 0, 78, 50, 21, 45, 76, 52, 20, 23, 57, 77, 170, 268, 271, 260, 266, 285, 293, 308, 287, 198, 115, 109, 144, 171, 185, 186, 190, 98, 
    0, 105, 184, 123, 62, 44, 66, 33, 7, 11, 39, 78, 186, 268, 258, 254, 273, 247, 214, 240, 290, 294, 257, 217, 209, 211, 206, 197, 155, 67, 
    31, 167, 215, 193, 104, 54, 55, 13, 2, 1, 22, 57, 173, 255, 251, 260, 241, 132, 89, 92, 141, 236, 293, 272, 229, 211, 208, 165, 86, 35, 
    35, 75, 136, 184, 119, 65, 35, 3, 0, 28, 76, 98, 185, 244, 243, 252, 158, 48, 50, 35, 37, 123, 225, 254, 208, 188, 156, 76, 28, 12, 
    2, 0, 63, 140, 121, 64, 19, 6, 11, 66, 119, 143, 225, 257, 253, 233, 97, 36, 43, 31, 25, 54, 144, 203, 192, 158, 81, 22, 10, 9, 
    0, 12, 65, 137, 133, 64, 16, 19, 39, 82, 106, 153, 245, 263, 264, 212, 81, 44, 47, 33, 20, 19, 90, 175, 200, 135, 46, 17, 17, 17, 
    0, 29, 70, 138, 135, 62, 16, 35, 69, 98, 104, 157, 223, 239, 245, 189, 76, 50, 72, 56, 25, 5, 48, 141, 184, 111, 32, 15, 14, 15, 
    0, 25, 63, 124, 138, 79, 55, 92, 145, 185, 195, 222, 247, 260, 265, 207, 92, 58, 101, 98, 64, 21, 27, 97, 135, 76, 21, 6, 4, 9, 
    0, 27, 65, 121, 139, 105, 105, 135, 177, 214, 229, 239, 246, 247, 246, 205, 111, 77, 101, 101, 68, 37, 12, 44, 58, 32, 10, 0, 1, 10, 
    0, 14, 42, 85, 83, 62, 58, 62, 76, 88, 93, 100, 104, 105, 103, 92, 57, 77, 88, 73, 51, 26, 0, 3, 2, 0, 0, 0, 2, 12, 
    2, 1, 5, 18, 18, 14, 7, 0, 10, 13, 12, 12, 12, 9, 6, 4, 0, 35, 73, 88, 71, 22, 0, 0, 0, 0, 0, 0, 6, 19, 
    15, 13, 14, 25, 41, 51, 36, 22, 31, 37, 35, 31, 25, 17, 11, 5, 0, 6, 34, 57, 42, 13, 0, 0, 0, 0, 0, 3, 15, 24, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 36, 67, 112, 150, 151, 103, 62, 54, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 110, 167, 186, 194, 210, 211, 180, 146, 153, 145, 36, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 66, 102, 133, 137, 102, 64, 53, 35, 17, 77, 186, 210, 99, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 44, 41, 35, 34, 7, 0, 0, 0, 0, 0, 68, 217, 248, 162, 41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 1, 0, 0, 0, 0, 0, 14, 153, 253, 272, 226, 107, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 82, 175, 242, 273, 294, 245, 108, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 17, 26, 25, 20, 0, 0, 0, 0, 0, 94, 181, 225, 263, 281, 283, 298, 262, 137, 20, 0, 0, 0, 0, 72, 96, 
    0, 0, 0, 0, 0, 0, 0, 22, 4, 0, 0, 0, 0, 69, 225, 298, 296, 288, 283, 284, 265, 185, 48, 0, 0, 0, 23, 88, 144, 138, 
    0, 0, 0, 22, 37, 0, 0, 0, 0, 0, 0, 0, 0, 105, 237, 274, 257, 260, 275, 281, 255, 194, 106, 46, 64, 110, 140, 151, 164, 142, 
    0, 0, 72, 138, 95, 1, 0, 0, 0, 0, 0, 0, 13, 120, 228, 247, 246, 273, 276, 245, 227, 218, 207, 182, 174, 183, 181, 169, 163, 110, 
    0, 47, 172, 191, 115, 20, 0, 0, 0, 0, 0, 0, 4, 121, 225, 238, 256, 244, 150, 72, 87, 131, 191, 232, 227, 205, 182, 172, 125, 26, 
    0, 80, 142, 121, 92, 35, 0, 0, 0, 0, 0, 0, 32, 134, 219, 237, 237, 140, 0, 0, 0, 18, 100, 199, 219, 183, 162, 118, 23, 0, 
    0, 0, 16, 19, 59, 50, 0, 0, 0, 0, 0, 29, 81, 158, 224, 238, 191, 62, 0, 0, 0, 0, 13, 102, 158, 152, 114, 28, 0, 0, 
    0, 0, 0, 3, 56, 56, 0, 0, 0, 0, 0, 44, 103, 190, 246, 236, 159, 25, 0, 0, 0, 0, 0, 29, 116, 140, 74, 0, 0, 0, 
    0, 0, 0, 16, 59, 59, 0, 0, 0, 0, 20, 61, 127, 207, 236, 213, 138, 18, 0, 0, 0, 0, 0, 0, 82, 118, 39, 0, 0, 0, 
    0, 0, 0, 17, 51, 48, 0, 0, 0, 26, 73, 111, 154, 199, 215, 200, 135, 25, 0, 0, 0, 0, 0, 0, 30, 61, 0, 0, 0, 0, 
    0, 0, 0, 17, 55, 58, 16, 10, 62, 123, 164, 183, 198, 213, 217, 192, 119, 20, 0, 27, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 32, 24, 0, 0, 13, 40, 60, 70, 79, 84, 85, 72, 27, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=111
    632, 631, 626, 629, 639, 642, 636, 623, 607, 583, 562, 551, 544, 534, 514, 494, 457, 377, 347, 350, 364, 353, 322, 247, 143, 112, 163, 251, 299, 307, 
    641, 625, 611, 605, 606, 602, 591, 578, 560, 537, 515, 506, 500, 491, 473, 455, 433, 404, 376, 374, 377, 351, 281, 180, 97, 86, 169, 269, 320, 323, 
    607, 591, 574, 560, 558, 551, 537, 520, 503, 482, 464, 458, 456, 449, 434, 421, 407, 399, 381, 366, 358, 322, 237, 158, 113, 128, 209, 298, 337, 336, 
    534, 516, 496, 489, 493, 495, 480, 464, 450, 436, 425, 423, 424, 419, 409, 404, 395, 395, 390, 361, 313, 256, 203, 169, 154, 188, 256, 324, 344, 339, 
    428, 422, 421, 427, 436, 440, 431, 422, 416, 411, 408, 410, 412, 410, 406, 404, 397, 397, 393, 329, 208, 130, 125, 156, 198, 241, 297, 333, 338, 333, 
    374, 382, 395, 400, 407, 407, 406, 406, 408, 407, 409, 416, 419, 416, 411, 410, 402, 403, 383, 266, 113, 28, 57, 146, 235, 279, 311, 332, 334, 329, 
    371, 382, 390, 391, 395, 396, 397, 403, 410, 414, 416, 421, 426, 428, 422, 419, 410, 404, 354, 218, 85, 29, 84, 193, 277, 319, 332, 345, 348, 339, 
    375, 388, 395, 394, 397, 398, 398, 404, 413, 422, 421, 413, 415, 423, 414, 401, 386, 368, 305, 188, 96, 76, 154, 255, 326, 350, 349, 349, 350, 340, 
    379, 392, 400, 398, 401, 401, 398, 401, 408, 412, 394, 363, 354, 367, 373, 375, 384, 382, 316, 213, 122, 97, 153, 236, 304, 336, 338, 337, 338, 332, 
    387, 397, 402, 399, 401, 401, 397, 397, 395, 376, 343, 321, 328, 351, 365, 361, 350, 323, 260, 206, 155, 123, 116, 130, 198, 272, 319, 324, 324, 321, 
    398, 401, 402, 399, 399, 397, 393, 387, 373, 351, 327, 289, 254, 220, 186, 140, 88, 33, 21, 56, 111, 144, 116, 67, 90, 174, 266, 303, 307, 310, 
    403, 402, 402, 401, 394, 390, 382, 372, 347, 300, 227, 132, 42, 0, 0, 0, 0, 0, 0, 0, 36, 118, 128, 90, 41, 87, 164, 242, 278, 294, 
    404, 402, 403, 402, 386, 373, 363, 338, 266, 172, 93, 35, 0, 0, 0, 0, 7, 22, 38, 27, 36, 79, 117, 118, 60, 37, 75, 146, 222, 263, 
    403, 402, 402, 392, 375, 361, 335, 253, 161, 106, 96, 77, 53, 41, 51, 78, 103, 142, 134, 79, 37, 42, 76, 97, 91, 48, 44, 88, 177, 246, 
    400, 401, 394, 367, 338, 311, 261, 172, 119, 107, 112, 90, 69, 86, 143, 194, 224, 212, 144, 78, 33, 4, 0, 35, 76, 88, 64, 100, 175, 241, 
    397, 396, 375, 308, 226, 167, 124, 106, 63, 58, 44, 33, 56, 123, 202, 231, 201, 137, 80, 46, 15, 0, 0, 20, 80, 112, 118, 120, 156, 207, 
    392, 383, 350, 257, 142, 63, 35, 14, 9, 0, 6, 9, 48, 65, 80, 62, 29, 14, 20, 31, 24, 44, 84, 116, 162, 169, 155, 107, 100, 147, 
    383, 371, 337, 237, 125, 42, 7, 0, 7, 8, 26, 36, 42, 18, 0, 0, 0, 0, 11, 22, 67, 140, 199, 212, 189, 156, 107, 68, 50, 91, 
    374, 354, 285, 182, 79, 28, 9, 9, 21, 25, 15, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 55, 136, 151, 106, 63, 42, 36, 18, 45, 
    350, 251, 135, 66, 24, 27, 15, 17, 26, 31, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 23, 1, 0, 0, 0, 17, 
    281, 89, 0, 0, 0, 18, 12, 25, 30, 48, 53, 45, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 
    222, 50, 0, 0, 0, 12, 19, 33, 41, 53, 45, 40, 21, 13, 12, 0, 0, 0, 10, 35, 17, 0, 0, 0, 0, 0, 0, 0, 21, 84, 
    215, 107, 22, 0, 0, 8, 27, 37, 48, 34, 0, 0, 0, 9, 8, 0, 4, 22, 32, 42, 38, 5, 0, 0, 0, 0, 0, 22, 71, 115, 
    202, 105, 31, 0, 0, 4, 25, 37, 45, 29, 14, 11, 0, 0, 0, 0, 12, 28, 49, 54, 51, 35, 0, 0, 0, 0, 0, 37, 81, 110, 
    181, 89, 24, 0, 0, 5, 35, 49, 60, 63, 71, 55, 24, 5, 0, 8, 21, 27, 39, 53, 66, 59, 23, 0, 0, 0, 0, 35, 74, 97, 
    175, 102, 38, 0, 0, 0, 22, 21, 7, 0, 0, 0, 0, 0, 0, 0, 0, 11, 19, 26, 26, 39, 21, 0, 0, 0, 0, 39, 68, 85, 
    181, 119, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 16, 25, 0, 0, 0, 16, 43, 57, 68, 
    192, 129, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 42, 33, 39, 28, 31, 34, 41, 48, 52, 61, 
    178, 134, 77, 37, 34, 48, 50, 40, 27, 27, 31, 34, 35, 35, 36, 39, 42, 20, 10, 0, 0, 16, 29, 44, 48, 48, 49, 51, 55, 59, 
    149, 122, 89, 68, 57, 45, 30, 20, 16, 18, 23, 33, 43, 51, 54, 58, 59, 49, 25, 4, 1, 20, 38, 50, 53, 51, 51, 52, 52, 54, 
    
    -- channel=112
    69, 68, 66, 65, 63, 67, 76, 82, 99, 115, 118, 109, 93, 75, 61, 55, 50, 47, 46, 43, 33, 26, 21, 14, 8, 3, 2, 4, 5, 1, 
    70, 69, 67, 66, 63, 69, 76, 78, 107, 123, 128, 128, 121, 104, 81, 63, 51, 44, 48, 46, 37, 32, 29, 26, 25, 22, 21, 23, 22, 19, 
    68, 67, 66, 64, 64, 75, 70, 74, 112, 122, 125, 135, 137, 129, 111, 85, 61, 47, 54, 56, 55, 52, 50, 50, 46, 43, 44, 45, 45, 41, 
    65, 64, 65, 63, 66, 75, 61, 81, 116, 126, 130, 140, 151, 151, 137, 112, 83, 67, 72, 77, 76, 75, 74, 75, 71, 67, 67, 65, 60, 54, 
    62, 61, 63, 60, 58, 59, 55, 83, 117, 124, 131, 138, 151, 160, 158, 144, 111, 89, 88, 96, 97, 97, 97, 95, 83, 76, 73, 70, 65, 59, 
    60, 59, 60, 58, 53, 47, 55, 83, 112, 121, 128, 137, 145, 155, 164, 163, 144, 120, 110, 114, 118, 117, 112, 96, 81, 77, 75, 72, 69, 64, 
    61, 62, 64, 72, 70, 62, 65, 85, 116, 125, 135, 146, 149, 157, 171, 174, 168, 151, 138, 128, 128, 131, 124, 102, 82, 78, 76, 74, 74, 74, 
    73, 79, 90, 101, 103, 102, 81, 85, 111, 120, 133, 149, 155, 168, 177, 181, 181, 170, 159, 151, 150, 154, 139, 113, 94, 90, 91, 92, 94, 95, 
    100, 109, 121, 132, 145, 146, 93, 84, 104, 110, 125, 151, 164, 179, 181, 179, 187, 188, 180, 172, 169, 166, 155, 130, 114, 112, 114, 113, 112, 111, 
    128, 140, 151, 163, 181, 162, 94, 81, 105, 109, 124, 151, 171, 179, 181, 178, 183, 190, 193, 187, 183, 177, 165, 146, 128, 125, 130, 128, 126, 122, 
    157, 165, 171, 174, 188, 152, 90, 77, 110, 115, 133, 162, 177, 180, 176, 173, 174, 184, 189, 190, 188, 180, 169, 153, 141, 135, 139, 136, 127, 117, 
    164, 166, 167, 166, 176, 152, 91, 70, 92, 114, 140, 173, 179, 181, 174, 167, 165, 176, 179, 183, 187, 178, 167, 157, 148, 137, 132, 128, 116, 103, 
    155, 157, 158, 158, 164, 164, 121, 87, 84, 104, 122, 154, 175, 175, 173, 166, 168, 174, 175, 180, 185, 178, 162, 160, 150, 133, 118, 113, 101, 87, 
    148, 150, 152, 156, 163, 172, 156, 117, 104, 100, 101, 134, 176, 177, 175, 173, 176, 182, 179, 182, 185, 179, 163, 161, 151, 132, 108, 97, 87, 80, 
    149, 154, 159, 165, 171, 173, 167, 147, 148, 114, 101, 129, 164, 173, 172, 174, 179, 184, 184, 184, 184, 179, 168, 158, 150, 135, 112, 98, 91, 83, 
    159, 164, 169, 178, 193, 195, 188, 185, 202, 169, 120, 148, 162, 182, 181, 175, 182, 184, 188, 186, 183, 181, 174, 159, 150, 139, 117, 101, 97, 89, 
    171, 182, 196, 211, 233, 240, 211, 206, 215, 219, 177, 175, 164, 192, 189, 176, 176, 180, 184, 184, 184, 184, 180, 163, 150, 138, 119, 102, 97, 89, 
    202, 218, 229, 238, 253, 273, 249, 235, 236, 229, 212, 186, 164, 194, 198, 179, 173, 176, 181, 182, 187, 189, 187, 168, 150, 135, 117, 96, 84, 74, 
    234, 246, 255, 261, 265, 264, 267, 236, 218, 212, 228, 190, 165, 193, 201, 183, 176, 177, 180, 183, 189, 194, 189, 172, 149, 134, 110, 85, 66, 60, 
    264, 277, 288, 289, 262, 214, 234, 216, 184, 191, 220, 191, 159, 181, 191, 181, 182, 182, 180, 184, 189, 193, 185, 169, 145, 128, 107, 86, 68, 61, 
    287, 286, 288, 291, 239, 181, 197, 193, 168, 174, 187, 175, 151, 155, 160, 159, 178, 181, 176, 176, 182, 187, 183, 170, 144, 123, 111, 99, 85, 68, 
    273, 256, 246, 243, 189, 151, 158, 158, 157, 155, 154, 148, 138, 131, 126, 126, 146, 163, 164, 165, 173, 178, 177, 163, 138, 116, 116, 116, 100, 79, 
    225, 210, 198, 184, 149, 130, 139, 137, 135, 135, 129, 125, 124, 123, 105, 107, 131, 151, 155, 153, 160, 172, 178, 169, 144, 113, 112, 122, 113, 93, 
    180, 162, 140, 123, 117, 117, 127, 130, 122, 119, 121, 117, 129, 137, 111, 96, 111, 133, 145, 150, 166, 178, 181, 174, 149, 123, 109, 119, 119, 106, 
    121, 110, 107, 108, 110, 110, 110, 114, 114, 103, 94, 100, 121, 136, 131, 119, 120, 133, 143, 152, 173, 181, 180, 178, 157, 131, 113, 110, 118, 116, 
    96, 98, 103, 106, 107, 109, 110, 109, 108, 103, 99, 105, 112, 120, 132, 132, 127, 130, 133, 143, 167, 177, 175, 173, 165, 139, 116, 104, 110, 117, 
    94, 94, 96, 104, 109, 110, 106, 100, 94, 92, 102, 106, 101, 104, 126, 126, 117, 117, 116, 126, 146, 158, 161, 160, 155, 136, 113, 101, 100, 106, 
    91, 93, 96, 100, 102, 101, 95, 86, 79, 80, 103, 117, 105, 103, 114, 111, 105, 103, 102, 106, 117, 127, 133, 136, 134, 120, 101, 94, 92, 91, 
    87, 86, 87, 88, 89, 88, 82, 76, 75, 80, 103, 118, 110, 116, 108, 100, 96, 91, 93, 92, 93, 100, 109, 113, 111, 102, 90, 86, 85, 79, 
    74, 73, 73, 71, 74, 76, 75, 74, 74, 80, 101, 114, 111, 115, 101, 93, 90, 86, 88, 87, 83, 86, 92, 93, 93, 90, 82, 78, 75, 71, 
    
    -- channel=113
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=114
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 4, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 10, 14, 13, 12, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 7, 10, 12, 14, 15, 14, 15, 13, 10, 9, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 2, 5, 5, 5, 8, 11, 14, 12, 11, 11, 8, 5, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 5, 4, 11, 15, 12, 6, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 11, 19, 24, 20, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 
    0, 0, 0, 0, 0, 5, 18, 3, 0, 0, 5, 10, 12, 16, 18, 16, 20, 17, 0, 0, 0, 0, 0, 0, 0, 2, 1, 3, 8, 14, 
    0, 2, 6, 7, 0, 0, 13, 10, 4, 4, 6, 12, 14, 13, 15, 13, 13, 19, 15, 1, 0, 0, 0, 6, 7, 8, 11, 14, 18, 22, 
    11, 11, 8, 4, 0, 0, 0, 7, 5, 5, 0, 0, 0, 0, 3, 12, 11, 12, 15, 13, 6, 0, 0, 3, 9, 12, 19, 20, 21, 21, 
    4, 0, 0, 0, 0, 0, 0, 6, 7, 12, 4, 0, 0, 0, 0, 5, 6, 8, 12, 16, 13, 10, 0, 0, 6, 11, 19, 19, 16, 14, 
    0, 0, 0, 0, 0, 0, 0, 11, 7, 17, 20, 0, 0, 0, 0, 1, 1, 3, 10, 15, 12, 13, 8, 5, 12, 12, 14, 14, 10, 6, 
    0, 0, 0, 0, 0, 0, 0, 15, 0, 2, 13, 0, 0, 0, 0, 0, 0, 0, 3, 11, 9, 10, 12, 5, 12, 13, 6, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 27, 9, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 5, 4, 6, 13, 5, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 25, 14, 3, 0, 0, 0, 8, 11, 3, 0, 0, 0, 1, 4, 12, 10, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 37, 23, 8, 11, 13, 9, 0, 0, 0, 0, 0, 3, 8, 12, 0, 0, 9, 5, 9, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 23, 27, 0, 11, 17, 8, 0, 0, 0, 0, 0, 2, 4, 9, 2, 0, 8, 11, 12, 11, 
    0, 0, 0, 0, 0, 0, 7, 14, 0, 0, 0, 11, 0, 0, 11, 7, 0, 0, 0, 0, 0, 0, 1, 4, 4, 0, 2, 5, 3, 9, 
    0, 3, 3, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 7, 8, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 19, 24, 29, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 4, 6, 9, 27, 33, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 16, 14, 21, 32, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 22, 20, 14, 24, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 7, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 2, 16, 23, 26, 14, 14, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 25, 17, 0, 0, 6, 10, 1, 6, 4, 0, 0, 0, 0, 15, 30, 30, 22, 10, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 14, 6, 0, 0, 0, 3, 0, 2, 0, 0, 0, 0, 0, 0, 24, 32, 31, 17, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 1, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 8, 27, 32, 27, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 9, 9, 22, 18, 8, 2, 9, 8, 4, 0, 0, 0, 0, 0, 0, 5, 22, 33, 33, 21, 
    0, 0, 0, 0, 0, 0, 5, 14, 26, 32, 21, 9, 16, 20, 19, 18, 24, 22, 16, 15, 4, 0, 0, 0, 3, 10, 25, 35, 34, 29, 
    0, 0, 0, 5, 13, 16, 23, 27, 36, 37, 23, 12, 13, 19, 19, 29, 35, 33, 27, 26, 28, 20, 16, 14, 15, 21, 32, 36, 32, 30, 
    0, 3, 14, 23, 30, 29, 27, 27, 35, 39, 26, 18, 14, 18, 25, 34, 37, 38, 33, 30, 33, 32, 30, 30, 29, 31, 34, 35, 31, 29, 
    
    -- channel=115
    115, 111, 104, 103, 110, 117, 115, 109, 105, 108, 110, 105, 97, 90, 88, 82, 73, 67, 62, 53, 47, 39, 29, 21, 13, 8, 7, 7, 4, 3, 
    113, 110, 103, 101, 107, 97, 88, 99, 97, 95, 106, 108, 96, 84, 79, 73, 67, 62, 55, 46, 39, 33, 29, 26, 25, 27, 30, 32, 30, 28, 
    111, 110, 103, 100, 100, 80, 72, 88, 84, 71, 76, 90, 89, 77, 69, 62, 59, 59, 58, 55, 51, 52, 53, 54, 55, 58, 60, 60, 56, 50, 
    107, 106, 102, 94, 90, 79, 63, 61, 62, 52, 46, 56, 66, 62, 58, 58, 65, 78, 86, 87, 84, 83, 83, 81, 80, 83, 82, 75, 65, 54, 
    98, 98, 97, 86, 69, 56, 45, 44, 46, 39, 33, 31, 32, 39, 49, 62, 80, 101, 111, 112, 107, 106, 105, 96, 90, 87, 80, 70, 58, 45, 
    90, 90, 90, 76, 44, 20, 25, 33, 28, 25, 22, 18, 21, 30, 40, 50, 67, 95, 116, 121, 122, 118, 105, 93, 86, 82, 77, 66, 54, 42, 
    88, 89, 93, 92, 73, 31, 6, 14, 20, 26, 29, 29, 31, 34, 40, 42, 45, 67, 96, 112, 117, 109, 98, 92, 90, 85, 77, 66, 55, 48, 
    104, 119, 136, 155, 142, 67, 8, 7, 22, 42, 56, 60, 60, 51, 42, 44, 46, 47, 62, 81, 96, 104, 99, 93, 95, 89, 80, 74, 68, 65, 
    159, 180, 199, 215, 186, 96, 25, 11, 18, 43, 75, 93, 96, 79, 54, 44, 46, 46, 45, 53, 68, 84, 94, 95, 99, 100, 93, 87, 82, 76, 
    212, 227, 239, 248, 210, 111, 34, 20, 20, 36, 76, 101, 106, 93, 67, 52, 49, 47, 42, 41, 46, 59, 78, 91, 101, 107, 101, 96, 91, 85, 
    242, 250, 254, 256, 226, 124, 37, 37, 49, 53, 85, 101, 99, 95, 76, 62, 63, 55, 45, 43, 39, 42, 61, 81, 93, 105, 108, 104, 97, 87, 
    247, 247, 244, 243, 233, 154, 52, 34, 63, 76, 97, 113, 100, 85, 77, 72, 76, 69, 55, 50, 43, 36, 55, 76, 83, 96, 105, 102, 92, 78, 
    233, 234, 232, 232, 232, 197, 103, 45, 49, 59, 77, 99, 93, 74, 72, 78, 89, 88, 72, 60, 48, 37, 47, 71, 79, 83, 93, 92, 79, 65, 
    222, 224, 227, 233, 237, 229, 183, 113, 52, 27, 51, 81, 84, 73, 73, 85, 105, 109, 92, 71, 52, 39, 39, 61, 75, 70, 75, 76, 71, 66, 
    221, 228, 237, 243, 236, 215, 209, 188, 122, 69, 71, 93, 87, 71, 71, 91, 112, 119, 105, 78, 57, 45, 38, 51, 69, 64, 65, 77, 78, 70, 
    231, 240, 247, 254, 250, 217, 206, 237, 228, 165, 118, 118, 118, 89, 74, 87, 110, 121, 110, 87, 66, 53, 44, 46, 64, 71, 74, 79, 68, 45, 
    246, 262, 284, 312, 333, 298, 246, 259, 266, 231, 178, 146, 150, 114, 80, 84, 104, 117, 111, 95, 78, 64, 52, 46, 60, 72, 67, 58, 37, 13, 
    304, 334, 364, 388, 404, 390, 309, 262, 276, 268, 217, 152, 146, 132, 92, 84, 101, 113, 113, 104, 92, 77, 61, 49, 55, 58, 41, 26, 13, 0, 
    385, 404, 417, 409, 392, 396, 343, 248, 232, 254, 221, 149, 130, 133, 100, 88, 100, 110, 113, 111, 103, 86, 66, 50, 48, 48, 31, 12, 1, 0, 
    432, 444, 445, 387, 303, 283, 270, 215, 186, 191, 180, 138, 108, 111, 100, 91, 101, 109, 112, 111, 99, 81, 61, 46, 44, 51, 39, 15, 2, 0, 
    458, 458, 436, 344, 227, 183, 182, 163, 135, 118, 111, 100, 83, 77, 76, 82, 93, 99, 101, 96, 85, 74, 63, 50, 44, 53, 56, 32, 10, 1, 
    429, 399, 358, 299, 221, 170, 146, 108, 76, 59, 54, 62, 70, 60, 43, 48, 63, 72, 78, 84, 90, 85, 72, 52, 38, 46, 65, 54, 22, 5, 
    327, 293, 271, 255, 213, 171, 149, 107, 59, 31, 25, 49, 86, 75, 32, 27, 45, 60, 74, 91, 100, 98, 86, 61, 37, 36, 54, 66, 42, 13, 
    242, 226, 206, 185, 165, 152, 152, 141, 95, 53, 42, 59, 85, 89, 63, 37, 43, 60, 80, 107, 121, 117, 105, 76, 44, 29, 38, 61, 61, 30, 
    172, 157, 149, 145, 146, 146, 141, 136, 121, 89, 60, 48, 58, 77, 75, 55, 52, 68, 95, 132, 142, 123, 106, 91, 61, 34, 28, 43, 63, 48, 
    122, 125, 132, 136, 133, 125, 113, 97, 86, 84, 69, 45, 44, 63, 69, 54, 49, 62, 86, 120, 135, 119, 94, 82, 70, 44, 22, 25, 46, 55, 
    114, 117, 116, 112, 103, 87, 68, 51, 46, 60, 69, 50, 36, 50, 55, 41, 33, 38, 49, 73, 97, 100, 85, 72, 57, 35, 18, 14, 23, 42, 
    104, 96, 84, 71, 59, 44, 30, 21, 22, 40, 61, 61, 51, 41, 31, 20, 11, 15, 20, 28, 48, 65, 65, 52, 35, 18, 7, 5, 7, 17, 
    73, 56, 40, 32, 27, 19, 9, 1, 8, 32, 54, 60, 50, 34, 21, 7, 0, 3, 9, 5, 11, 22, 28, 25, 17, 3, 0, 0, 0, 0, 
    31, 20, 11, 7, 5, 1, 0, 0, 2, 23, 43, 52, 44, 27, 11, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0, 
    
    -- channel=116
    1, 4, 5, 3, 0, 7, 24, 25, 19, 15, 0, 0, 0, 5, 8, 4, 2, 1, 5, 11, 12, 14, 14, 11, 5, 0, 0, 0, 0, 0, 
    2, 4, 5, 0, 0, 27, 48, 25, 1, 2, 2, 0, 0, 0, 0, 9, 13, 11, 11, 15, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 2, 30, 26, 3, 11, 24, 31, 36, 20, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 8, 6, 7, 15, 26, 0, 0, 42, 43, 30, 37, 47, 35, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    13, 12, 13, 19, 42, 63, 34, 8, 26, 16, 2, 4, 15, 16, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 29, 34, 32, 
    7, 5, 9, 23, 45, 59, 46, 27, 15, 12, 12, 13, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 25, 21, 21, 27, 23, 15, 7, 
    0, 0, 0, 0, 0, 0, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 13, 32, 24, 4, 3, 14, 17, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 18, 16, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 78, 34, 0, 0, 0, 0, 0, 6, 13, 1, 0, 0, 0, 0, 0, 0, 13, 20, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 43, 58, 4, 0, 0, 0, 0, 0, 3, 22, 11, 0, 0, 0, 0, 0, 0, 3, 5, 1, 0, 5, 6, 5, 11, 21, 
    13, 24, 32, 37, 40, 30, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 12, 24, 27, 39, 51, 
    37, 40, 38, 29, 15, 0, 0, 0, 15, 66, 64, 51, 41, 14, 0, 0, 0, 0, 0, 0, 3, 5, 0, 0, 8, 19, 40, 53, 61, 60, 
    26, 21, 9, 0, 0, 0, 0, 0, 0, 27, 57, 38, 36, 22, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 18, 25, 45, 56, 40, 13, 
    0, 0, 0, 0, 0, 32, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 4, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 2, 11, 40, 75, 83, 
    0, 0, 0, 0, 0, 0, 0, 0, 40, 12, 0, 8, 11, 27, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 51, 72, 78, 49, 
    0, 0, 0, 0, 68, 105, 99, 60, 65, 78, 68, 58, 8, 37, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 33, 28, 22, 9, 
    0, 0, 0, 98, 211, 259, 262, 190, 85, 92, 125, 101, 17, 37, 42, 0, 0, 0, 0, 0, 6, 19, 22, 15, 7, 0, 0, 0, 0, 3, 
    6, 21, 55, 136, 162, 128, 145, 143, 97, 105, 124, 93, 50, 71, 82, 35, 8, 9, 14, 22, 28, 21, 7, 0, 0, 0, 0, 0, 0, 5, 
    81, 141, 197, 208, 104, 0, 0, 32, 77, 103, 90, 55, 22, 30, 64, 80, 74, 61, 44, 25, 8, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    229, 242, 225, 178, 94, 24, 32, 29, 16, 35, 36, 5, 0, 0, 0, 4, 32, 25, 5, 0, 0, 0, 0, 1, 13, 12, 10, 13, 0, 0, 
    220, 166, 116, 90, 82, 71, 51, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 24, 8, 0, 
    94, 75, 67, 55, 40, 21, 5, 6, 12, 0, 0, 0, 20, 33, 11, 0, 0, 0, 0, 0, 0, 0, 6, 11, 0, 0, 4, 18, 22, 11, 
    54, 46, 29, 8, 0, 6, 36, 71, 92, 73, 33, 23, 40, 34, 13, 1, 0, 1, 7, 15, 34, 36, 25, 23, 26, 19, 13, 19, 27, 30, 
    17, 2, 0, 12, 43, 73, 94, 96, 73, 31, 6, 0, 0, 0, 22, 39, 27, 26, 44, 67, 88, 69, 30, 16, 30, 46, 38, 26, 26, 35, 
    0, 16, 50, 78, 92, 90, 77, 56, 24, 0, 0, 5, 0, 0, 28, 48, 40, 35, 38, 45, 63, 64, 46, 38, 44, 47, 36, 26, 29, 36, 
    58, 83, 92, 83, 60, 38, 22, 15, 9, 3, 12, 17, 11, 23, 38, 28, 20, 12, 11, 17, 27, 45, 61, 64, 52, 35, 24, 26, 32, 35, 
    98, 84, 61, 36, 22, 19, 14, 14, 12, 6, 19, 24, 22, 30, 34, 26, 21, 11, 12, 17, 15, 21, 35, 40, 33, 25, 22, 27, 32, 30, 
    
    -- channel=117
    44, 44, 47, 50, 52, 54, 54, 61, 68, 66, 61, 55, 56, 56, 52, 47, 48, 51, 56, 56, 57, 58, 58, 59, 57, 56, 54, 49, 46, 43, 
    45, 44, 47, 48, 54, 63, 63, 69, 66, 72, 71, 60, 56, 60, 61, 58, 54, 57, 58, 60, 60, 56, 52, 47, 42, 38, 36, 32, 32, 33, 
    45, 43, 44, 49, 55, 55, 65, 76, 73, 86, 97, 91, 80, 72, 69, 65, 56, 54, 49, 47, 42, 37, 33, 30, 29, 28, 29, 31, 34, 40, 
    50, 48, 47, 54, 58, 49, 66, 78, 86, 93, 101, 106, 105, 99, 88, 69, 47, 34, 29, 27, 29, 28, 30, 33, 37, 40, 43, 48, 53, 58, 
    53, 53, 50, 58, 70, 73, 80, 84, 86, 89, 91, 98, 101, 101, 99, 83, 62, 39, 30, 33, 41, 43, 46, 47, 54, 58, 61, 64, 68, 68, 
    52, 53, 53, 55, 64, 82, 92, 93, 91, 95, 98, 99, 99, 97, 95, 97, 96, 82, 64, 53, 54, 61, 60, 59, 60, 60, 61, 62, 63, 63, 
    50, 47, 42, 29, 23, 42, 68, 89, 86, 83, 81, 79, 84, 93, 98, 101, 102, 105, 93, 80, 70, 68, 67, 61, 54, 50, 53, 57, 57, 56, 
    29, 19, 7, 0, 0, 10, 50, 79, 79, 71, 60, 53, 59, 72, 92, 101, 98, 100, 102, 98, 90, 77, 67, 58, 53, 50, 50, 51, 52, 53, 
    0, 0, 0, 0, 8, 21, 59, 79, 85, 87, 79, 63, 59, 64, 81, 95, 98, 99, 103, 104, 103, 95, 80, 68, 57, 52, 50, 50, 53, 56, 
    0, 2, 9, 17, 20, 34, 62, 73, 76, 87, 88, 85, 77, 76, 82, 89, 92, 95, 99, 103, 106, 105, 98, 86, 72, 62, 57, 58, 60, 63, 
    21, 27, 32, 35, 15, 25, 50, 65, 55, 61, 65, 72, 79, 81, 84, 81, 83, 84, 93, 97, 100, 101, 97, 94, 85, 75, 67, 63, 64, 67, 
    37, 39, 41, 42, 19, 10, 41, 68, 70, 66, 64, 61, 70, 76, 84, 82, 78, 75, 85, 93, 95, 96, 94, 92, 87, 82, 75, 69, 70, 74, 
    46, 45, 43, 39, 25, 0, 2, 38, 83, 99, 105, 98, 86, 85, 86, 83, 73, 69, 76, 88, 93, 94, 100, 95, 92, 89, 84, 77, 75, 75, 
    44, 41, 35, 30, 27, 8, 0, 0, 31, 73, 97, 98, 84, 88, 85, 78, 66, 60, 67, 80, 89, 93, 102, 97, 94, 92, 89, 78, 67, 60, 
    32, 28, 24, 25, 35, 49, 35, 16, 0, 4, 33, 47, 58, 74, 86, 84, 73, 66, 69, 78, 85, 90, 96, 95, 88, 82, 73, 65, 55, 57, 
    27, 25, 25, 20, 14, 31, 38, 25, 0, 0, 15, 25, 46, 59, 79, 90, 81, 76, 74, 76, 81, 86, 90, 93, 85, 75, 65, 64, 69, 83, 
    20, 13, 0, 0, 0, 0, 0, 12, 15, 0, 24, 33, 55, 55, 72, 84, 81, 75, 72, 72, 75, 81, 85, 91, 86, 82, 84, 92, 95, 97, 
    0, 0, 0, 0, 0, 0, 0, 24, 50, 37, 26, 46, 69, 70, 71, 80, 79, 75, 73, 72, 72, 77, 81, 89, 90, 90, 95, 101, 96, 86, 
    0, 0, 0, 11, 38, 42, 29, 50, 72, 86, 52, 63, 78, 79, 73, 78, 77, 74, 73, 73, 74, 78, 82, 88, 90, 83, 85, 85, 83, 78, 
    0, 0, 4, 45, 92, 138, 113, 94, 96, 110, 92, 88, 91, 87, 82, 80, 76, 73, 73, 77, 83, 86, 90, 91, 89, 76, 70, 71, 75, 75, 
    2, 8, 19, 26, 58, 98, 100, 99, 112, 122, 115, 103, 101, 101, 102, 98, 87, 85, 86, 87, 87, 84, 82, 81, 85, 79, 66, 65, 70, 77, 
    36, 61, 71, 42, 32, 29, 38, 68, 101, 122, 117, 100, 82, 81, 100, 115, 114, 106, 100, 89, 77, 73, 73, 78, 85, 90, 76, 64, 67, 77, 
    93, 99, 91, 65, 50, 47, 41, 43, 62, 85, 97, 91, 73, 49, 58, 83, 96, 93, 87, 76, 66, 64, 68, 78, 86, 98, 90, 70, 64, 70, 
    96, 81, 71, 68, 65, 64, 54, 32, 17, 25, 49, 74, 80, 62, 52, 57, 68, 72, 68, 60, 55, 61, 68, 68, 78, 88, 97, 84, 67, 65, 
    71, 68, 66, 64, 59, 53, 53, 53, 43, 34, 51, 77, 90, 84, 71, 68, 73, 77, 72, 62, 52, 62, 79, 80, 77, 80, 91, 94, 80, 67, 
    66, 63, 58, 54, 55, 61, 74, 88, 90, 79, 72, 77, 87, 88, 80, 76, 80, 87, 94, 91, 77, 75, 86, 94, 91, 90, 90, 97, 93, 75, 
    57, 55, 58, 66, 79, 90, 98, 99, 93, 85, 69, 61, 65, 79, 82, 85, 88, 93, 106, 113, 103, 88, 83, 89, 95, 100, 98, 96, 97, 87, 
    57, 69, 82, 93, 98, 99, 97, 93, 86, 82, 72, 63, 67, 76, 83, 90, 91, 90, 95, 101, 101, 96, 91, 91, 95, 101, 101, 96, 95, 95, 
    83, 94, 99, 98, 92, 87, 85, 88, 89, 89, 80, 71, 80, 81, 90, 90, 86, 86, 84, 85, 91, 99, 100, 98, 95, 97, 100, 98, 94, 95, 
    99, 98, 93, 91, 89, 86, 86, 87, 91, 93, 86, 77, 81, 83, 94, 93, 91, 90, 86, 84, 86, 91, 93, 94, 92, 92, 97, 98, 94, 90, 
    
    -- channel=118
    12, 13, 16, 18, 22, 30, 33, 37, 36, 28, 18, 10, 15, 21, 20, 15, 15, 17, 22, 24, 26, 26, 25, 24, 20, 16, 12, 5, 0, 0, 
    13, 12, 15, 13, 24, 48, 46, 38, 23, 25, 22, 10, 4, 9, 19, 26, 26, 27, 27, 27, 25, 20, 10, 0, 0, 0, 0, 0, 0, 0, 
    13, 10, 10, 12, 27, 38, 29, 32, 32, 48, 61, 53, 34, 19, 17, 23, 22, 21, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 17, 15, 23, 32, 17, 20, 40, 55, 56, 61, 65, 60, 49, 32, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 23, 32, 
    23, 23, 20, 32, 52, 52, 52, 47, 38, 34, 32, 42, 47, 44, 34, 15, 0, 0, 0, 0, 0, 0, 5, 14, 26, 36, 43, 48, 51, 49, 
    20, 20, 21, 32, 51, 65, 58, 48, 36, 36, 41, 43, 39, 30, 29, 36, 44, 42, 33, 20, 14, 23, 34, 42, 44, 43, 41, 37, 33, 29, 
    13, 8, 1, 0, 0, 0, 9, 35, 25, 13, 9, 4, 8, 22, 34, 46, 55, 64, 59, 44, 30, 33, 37, 33, 28, 19, 18, 19, 17, 14, 
    0, 0, 0, 0, 0, 0, 0, 18, 7, 0, 0, 0, 0, 0, 24, 37, 37, 45, 52, 54, 47, 30, 21, 15, 18, 15, 12, 9, 6, 5, 
    0, 0, 0, 0, 0, 0, 9, 19, 25, 26, 15, 0, 0, 0, 10, 29, 35, 34, 40, 45, 50, 44, 33, 25, 18, 13, 7, 7, 11, 18, 
    0, 0, 0, 0, 8, 10, 13, 17, 21, 28, 31, 32, 25, 23, 16, 22, 30, 30, 33, 39, 48, 54, 53, 43, 32, 27, 25, 29, 33, 38, 
    0, 5, 15, 23, 3, 0, 0, 7, 0, 0, 0, 14, 24, 23, 21, 15, 18, 20, 27, 32, 39, 44, 43, 44, 44, 51, 48, 43, 47, 52, 
    26, 34, 38, 40, 0, 0, 0, 21, 20, 0, 0, 0, 6, 9, 19, 15, 15, 14, 22, 30, 34, 37, 29, 36, 46, 59, 64, 61, 66, 71, 
    43, 43, 39, 31, 0, 0, 0, 0, 48, 82, 88, 66, 44, 31, 23, 17, 10, 5, 9, 23, 31, 33, 36, 39, 54, 64, 77, 76, 74, 69, 
    31, 26, 17, 5, 0, 0, 0, 0, 0, 51, 75, 66, 39, 31, 19, 10, 0, 0, 0, 12, 24, 27, 40, 42, 54, 61, 75, 71, 51, 29, 
    3, 0, 0, 0, 12, 35, 0, 0, 0, 0, 0, 0, 0, 10, 23, 23, 16, 6, 6, 13, 19, 21, 32, 37, 39, 40, 37, 28, 11, 14, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 19, 40, 33, 25, 16, 12, 12, 13, 22, 31, 28, 20, 9, 18, 40, 73, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 14, 32, 28, 20, 12, 5, 4, 8, 15, 26, 25, 30, 45, 77, 101, 104, 
    0, 0, 0, 0, 0, 0, 0, 0, 33, 1, 0, 13, 38, 32, 18, 24, 24, 17, 10, 4, 0, 4, 8, 20, 29, 50, 76, 98, 93, 70, 
    0, 0, 0, 11, 66, 68, 46, 54, 69, 76, 45, 45, 42, 41, 22, 18, 17, 12, 9, 7, 6, 9, 14, 22, 34, 42, 52, 57, 58, 52, 
    0, 0, 12, 91, 162, 220, 179, 120, 91, 114, 94, 65, 53, 54, 41, 24, 14, 10, 11, 17, 27, 32, 34, 32, 34, 22, 20, 28, 44, 51, 
    8, 19, 43, 76, 95, 122, 110, 87, 98, 119, 107, 75, 73, 84, 78, 60, 38, 33, 37, 45, 46, 34, 21, 16, 26, 24, 18, 23, 36, 50, 
    67, 118, 149, 95, 22, 0, 0, 39, 81, 101, 87, 60, 44, 53, 74, 96, 93, 75, 62, 46, 24, 8, 6, 17, 36, 47, 37, 30, 33, 46, 
    185, 192, 159, 87, 40, 30, 25, 21, 20, 37, 47, 31, 7, 0, 16, 42, 54, 42, 26, 12, 4, 1, 7, 23, 40, 65, 64, 44, 30, 34, 
    154, 108, 79, 74, 74, 69, 37, 0, 0, 0, 0, 0, 20, 9, 0, 0, 0, 1, 0, 0, 0, 0, 4, 8, 22, 49, 76, 61, 37, 30, 
    72, 68, 67, 59, 41, 25, 21, 20, 5, 0, 1, 38, 66, 49, 18, 6, 9, 13, 2, 0, 0, 3, 21, 19, 25, 36, 63, 73, 56, 40, 
    62, 54, 34, 18, 18, 34, 61, 91, 97, 70, 52, 55, 61, 53, 32, 21, 24, 33, 45, 53, 45, 32, 35, 40, 42, 49, 62, 80, 75, 53, 
    27, 19, 24, 41, 67, 89, 105, 106, 88, 61, 35, 26, 23, 39, 45, 51, 53, 59, 83, 99, 87, 56, 33, 35, 52, 68, 75, 79, 84, 70, 
    22, 47, 75, 96, 105, 101, 90, 78, 61, 54, 44, 28, 22, 43, 61, 72, 71, 68, 75, 83, 81, 67, 55, 57, 66, 73, 78, 79, 85, 85, 
    79, 100, 106, 97, 79, 65, 58, 62, 65, 68, 61, 44, 50, 58, 67, 67, 64, 58, 53, 59, 69, 82, 88, 85, 74, 70, 76, 82, 83, 86, 
    108, 97, 80, 70, 66, 65, 63, 64, 68, 73, 71, 56, 61, 60, 70, 73, 69, 65, 62, 62, 64, 73, 78, 78, 72, 70, 77, 82, 80, 77, 
    
    -- channel=119
    113, 114, 114, 112, 106, 100, 102, 113, 133, 149, 153, 142, 131, 121, 117, 115, 114, 115, 119, 117, 115, 115, 115, 117, 117, 115, 112, 112, 113, 115, 
    113, 114, 115, 114, 110, 103, 107, 131, 149, 161, 169, 164, 155, 148, 139, 124, 113, 112, 117, 120, 119, 116, 118, 120, 119, 116, 113, 112, 112, 111, 
    113, 114, 116, 115, 111, 109, 121, 147, 160, 171, 179, 183, 185, 180, 167, 146, 124, 116, 119, 124, 122, 121, 121, 122, 119, 113, 106, 103, 103, 102, 
    114, 115, 116, 115, 113, 121, 133, 147, 168, 186, 193, 199, 209, 212, 202, 176, 142, 125, 122, 125, 124, 119, 117, 114, 109, 104, 98, 96, 97, 96, 
    116, 116, 117, 115, 112, 122, 136, 157, 188, 207, 213, 216, 220, 227, 225, 204, 170, 138, 121, 117, 119, 115, 112, 106, 100, 95, 92, 94, 97, 98, 
    119, 119, 119, 114, 106, 116, 147, 182, 207, 221, 223, 223, 228, 233, 227, 210, 185, 157, 134, 123, 127, 127, 116, 103, 93, 91, 95, 100, 103, 106, 
    121, 121, 119, 115, 116, 125, 148, 191, 220, 228, 225, 225, 227, 225, 222, 215, 199, 183, 167, 156, 152, 144, 130, 113, 98, 94, 100, 105, 107, 107, 
    120, 121, 121, 123, 127, 125, 145, 195, 224, 229, 221, 216, 216, 215, 217, 224, 223, 211, 198, 189, 183, 178, 160, 128, 105, 96, 100, 105, 107, 108, 
    117, 115, 113, 111, 112, 118, 151, 192, 211, 211, 207, 205, 207, 212, 220, 228, 231, 232, 227, 220, 214, 205, 186, 148, 115, 102, 101, 102, 102, 100, 
    102, 97, 94, 93, 103, 121, 152, 182, 195, 197, 200, 201, 203, 214, 225, 230, 230, 234, 239, 237, 230, 221, 206, 172, 132, 106, 94, 92, 92, 93, 
    87, 84, 85, 89, 105, 124, 137, 170, 191, 196, 196, 201, 205, 223, 231, 226, 224, 224, 231, 235, 233, 228, 219, 189, 143, 108, 90, 86, 86, 86, 
    84, 83, 82, 87, 103, 121, 122, 144, 172, 185, 190, 204, 214, 224, 233, 223, 214, 212, 219, 226, 231, 232, 228, 202, 153, 115, 92, 83, 82, 84, 
    84, 83, 84, 87, 97, 114, 113, 116, 143, 159, 175, 197, 213, 221, 228, 219, 209, 209, 214, 221, 230, 235, 229, 209, 169, 127, 101, 87, 87, 90, 
    93, 91, 88, 90, 96, 108, 116, 111, 113, 128, 158, 183, 201, 217, 222, 216, 211, 212, 215, 222, 231, 238, 231, 213, 187, 148, 119, 102, 98, 102, 
    101, 97, 94, 93, 93, 96, 110, 122, 115, 126, 146, 164, 179, 197, 209, 212, 210, 212, 217, 224, 233, 241, 235, 218, 201, 170, 139, 122, 112, 106, 
    105, 99, 92, 87, 88, 96, 104, 126, 139, 136, 123, 129, 156, 176, 197, 208, 211, 214, 219, 226, 234, 241, 239, 225, 211, 189, 158, 131, 105, 93, 
    97, 91, 85, 85, 94, 106, 108, 122, 129, 117, 116, 110, 147, 166, 190, 210, 214, 218, 222, 228, 234, 240, 242, 233, 218, 197, 160, 121, 92, 86, 
    90, 87, 82, 74, 71, 86, 93, 96, 129, 127, 119, 108, 135, 168, 193, 213, 219, 220, 224, 227, 231, 239, 244, 239, 222, 195, 150, 112, 92, 92, 
    77, 66, 54, 45, 44, 70, 102, 104, 128, 140, 133, 128, 145, 182, 199, 215, 221, 222, 224, 225, 227, 236, 243, 243, 223, 190, 147, 110, 91, 87, 
    46, 39, 40, 46, 51, 81, 119, 144, 154, 149, 154, 174, 175, 187, 201, 212, 221, 224, 221, 217, 219, 228, 239, 240, 219, 183, 142, 105, 87, 84, 
    43, 42, 45, 59, 76, 109, 145, 177, 181, 175, 188, 207, 196, 181, 187, 201, 213, 220, 216, 207, 206, 220, 235, 232, 207, 169, 132, 104, 89, 87, 
    49, 45, 47, 77, 112, 129, 145, 161, 180, 203, 220, 221, 198, 168, 163, 181, 203, 215, 213, 203, 204, 217, 224, 216, 186, 149, 122, 107, 94, 91, 
    52, 55, 69, 97, 111, 108, 122, 139, 166, 202, 222, 217, 196, 164, 144, 162, 199, 217, 219, 208, 200, 204, 208, 200, 173, 139, 113, 107, 102, 95, 
    85, 100, 103, 96, 89, 92, 109, 133, 148, 166, 191, 193, 179, 167, 165, 170, 196, 217, 216, 202, 193, 200, 207, 196, 169, 136, 110, 106, 107, 100, 
    108, 105, 101, 100, 103, 108, 109, 114, 126, 136, 145, 149, 154, 169, 180, 183, 199, 216, 213, 200, 192, 198, 209, 209, 181, 141, 114, 103, 107, 106, 
    102, 105, 111, 117, 116, 111, 106, 101, 102, 112, 119, 123, 145, 169, 182, 186, 197, 209, 202, 189, 189, 204, 215, 214, 194, 156, 118, 102, 103, 109, 
    114, 115, 113, 113, 114, 112, 107, 103, 103, 108, 116, 122, 133, 152, 163, 169, 176, 182, 176, 171, 185, 204, 214, 211, 190, 155, 120, 103, 97, 103, 
    113, 107, 104, 107, 111, 111, 110, 107, 104, 101, 107, 120, 132, 135, 132, 137, 141, 148, 151, 154, 169, 185, 188, 182, 167, 143, 115, 98, 92, 94, 
    104, 100, 100, 105, 110, 110, 106, 101, 95, 94, 100, 115, 125, 121, 118, 113, 111, 121, 129, 134, 140, 146, 144, 141, 137, 125, 106, 93, 88, 89, 
    99, 101, 103, 102, 99, 97, 97, 98, 95, 93, 96, 107, 115, 113, 109, 99, 99, 106, 110, 112, 114, 114, 111, 110, 110, 105, 97, 91, 90, 91, 
    
    -- channel=120
    36, 41, 40, 25, 17, 25, 29, 14, 0, 0, 0, 5, 21, 24, 28, 37, 40, 35, 35, 43, 43, 49, 52, 50, 50, 46, 41, 46, 53, 48, 
    37, 41, 43, 24, 17, 41, 21, 0, 0, 0, 0, 0, 2, 6, 8, 24, 33, 31, 31, 35, 33, 36, 38, 37, 38, 35, 33, 37, 42, 37, 
    37, 38, 44, 26, 19, 56, 15, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 20, 22, 25, 22, 20, 22, 22, 21, 20, 22, 26, 30, 28, 
    35, 34, 40, 31, 21, 45, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 12, 10, 4, 5, 9, 6, 6, 14, 18, 21, 22, 
    35, 31, 34, 38, 35, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 4, 3, 5, 13, 16, 15, 16, 
    33, 30, 29, 46, 57, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 14, 18, 15, 11, 7, 
    28, 25, 26, 40, 63, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 15, 5, 0, 0, 
    19, 15, 16, 17, 53, 94, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 3, 2, 0, 55, 115, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 72, 137, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 71, 152, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 3, 44, 136, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 3, 6, 4, 16, 81, 112, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    5, 3, 1, 0, 0, 24, 66, 63, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 
    0, 0, 0, 0, 0, 9, 0, 11, 72, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 37, 0, 0, 27, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 59, 25, 0, 0, 8, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 81, 0, 0, 0, 23, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 53, 41, 0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 69, 51, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 114, 106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 14, 24, 78, 85, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 30, 29, 35, 40, 4, 7, 34, 11, 0, 0, 0, 0, 2, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 29, 30, 23, 18, 9, 0, 14, 31, 7, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 16, 17, 15, 9, 2, 0, 0, 2, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=121
    89, 90, 91, 91, 88, 86, 89, 101, 116, 124, 120, 110, 107, 103, 100, 95, 93, 95, 99, 100, 101, 102, 103, 104, 102, 100, 97, 96, 94, 90, 
    91, 92, 93, 92, 92, 96, 104, 118, 124, 132, 131, 122, 118, 119, 115, 107, 100, 99, 103, 105, 104, 102, 102, 100, 94, 88, 82, 78, 76, 74, 
    90, 90, 90, 90, 93, 101, 112, 123, 128, 144, 153, 150, 143, 138, 132, 123, 109, 102, 98, 98, 94, 89, 84, 80, 74, 69, 65, 66, 69, 73, 
    95, 93, 92, 94, 98, 100, 110, 127, 148, 163, 172, 178, 179, 172, 159, 136, 109, 91, 82, 78, 72, 70, 70, 72, 72, 71, 71, 75, 80, 84, 
    99, 99, 96, 98, 105, 111, 122, 140, 159, 167, 169, 175, 183, 187, 179, 153, 117, 88, 76, 74, 76, 78, 81, 82, 82, 80, 82, 88, 94, 98, 
    100, 100, 98, 97, 106, 125, 144, 159, 166, 173, 175, 177, 179, 177, 170, 163, 149, 127, 109, 100, 100, 100, 96, 93, 90, 89, 92, 95, 96, 97, 
    99, 97, 93, 83, 82, 98, 129, 166, 177, 175, 170, 167, 167, 167, 167, 169, 169, 164, 148, 132, 124, 119, 113, 100, 88, 84, 88, 90, 91, 90, 
    86, 79, 69, 52, 44, 61, 111, 159, 168, 156, 142, 136, 138, 148, 163, 174, 173, 171, 169, 164, 157, 144, 124, 99, 84, 81, 86, 88, 87, 85, 
    54, 43, 36, 32, 44, 73, 120, 153, 162, 155, 145, 135, 133, 141, 157, 172, 177, 178, 179, 180, 177, 165, 140, 110, 89, 82, 81, 79, 78, 78, 
    34, 35, 41, 50, 69, 94, 123, 145, 154, 158, 159, 154, 150, 155, 163, 170, 173, 176, 181, 184, 186, 182, 165, 133, 100, 84, 77, 77, 79, 82, 
    51, 57, 63, 70, 72, 86, 106, 131, 134, 136, 144, 153, 162, 169, 170, 165, 163, 163, 172, 177, 181, 183, 172, 146, 114, 95, 83, 79, 80, 82, 
    65, 67, 72, 78, 72, 72, 89, 118, 128, 123, 128, 141, 156, 166, 173, 163, 154, 152, 160, 168, 175, 182, 173, 150, 119, 101, 88, 81, 82, 88, 
    75, 75, 76, 77, 70, 58, 64, 93, 131, 144, 152, 159, 164, 169, 172, 164, 153, 148, 153, 163, 174, 182, 177, 158, 132, 110, 100, 94, 94, 98, 
    81, 77, 73, 69, 65, 53, 38, 45, 86, 135, 162, 169, 167, 170, 166, 159, 149, 144, 149, 161, 174, 181, 180, 168, 150, 128, 117, 107, 101, 97, 
    76, 69, 64, 61, 65, 74, 66, 54, 48, 76, 99, 114, 127, 145, 158, 158, 151, 147, 151, 161, 174, 179, 179, 171, 157, 136, 120, 106, 92, 86, 
    67, 61, 57, 56, 62, 81, 88, 82, 54, 34, 52, 74, 105, 125, 152, 167, 163, 160, 159, 164, 171, 176, 178, 173, 160, 139, 113, 94, 86, 95, 
    60, 54, 46, 33, 18, 20, 40, 52, 56, 43, 64, 75, 102, 115, 146, 166, 165, 161, 160, 161, 166, 172, 176, 175, 164, 146, 121, 108, 107, 115, 
    33, 17, 1, 0, 0, 0, 17, 58, 91, 75, 71, 81, 109, 130, 149, 166, 166, 162, 161, 160, 162, 170, 177, 178, 168, 152, 132, 121, 113, 106, 
    0, 0, 0, 8, 35, 54, 65, 88, 118, 119, 98, 106, 127, 147, 155, 165, 167, 164, 163, 161, 162, 169, 177, 180, 169, 148, 125, 105, 95, 91, 
    0, 3, 20, 58, 104, 149, 155, 151, 146, 149, 148, 149, 147, 154, 159, 161, 164, 163, 160, 158, 164, 175, 183, 182, 166, 134, 105, 87, 84, 88, 
    21, 24, 34, 67, 113, 156, 174, 173, 165, 173, 188, 183, 166, 158, 159, 163, 164, 165, 161, 159, 165, 174, 178, 172, 154, 123, 96, 83, 83, 88, 
    43, 58, 76, 87, 90, 86, 104, 134, 167, 193, 200, 186, 158, 144, 152, 169, 178, 179, 173, 163, 158, 156, 155, 152, 140, 121, 100, 87, 84, 89, 
    101, 122, 128, 113, 89, 78, 89, 110, 142, 172, 181, 166, 136, 110, 123, 157, 179, 181, 170, 152, 140, 140, 145, 146, 136, 123, 106, 94, 86, 87, 
    144, 131, 111, 98, 95, 102, 103, 94, 93, 113, 133, 137, 131, 119, 115, 125, 146, 157, 149, 137, 132, 137, 140, 134, 125, 117, 114, 103, 91, 85, 
    113, 105, 104, 104, 102, 95, 89, 86, 83, 84, 97, 118, 139, 144, 135, 137, 152, 159, 149, 134, 127, 139, 152, 144, 125, 110, 110, 109, 101, 92, 
    105, 108, 105, 97, 92, 92, 100, 111, 119, 116, 114, 125, 143, 148, 142, 146, 159, 165, 158, 150, 147, 156, 165, 163, 142, 118, 108, 111, 110, 101, 
    101, 95, 93, 99, 109, 116, 124, 128, 126, 116, 102, 102, 116, 133, 139, 147, 154, 159, 164, 170, 174, 172, 168, 163, 147, 127, 114, 111, 112, 108, 
    90, 95, 105, 120, 129, 131, 126, 117, 106, 100, 99, 101, 106, 112, 122, 134, 139, 143, 148, 159, 168, 166, 157, 151, 143, 129, 114, 105, 107, 109, 
    105, 115, 123, 127, 124, 116, 106, 102, 99, 100, 104, 106, 111, 111, 114, 113, 115, 120, 123, 129, 138, 144, 143, 140, 132, 120, 109, 103, 103, 107, 
    124, 124, 117, 110, 103, 100, 100, 101, 99, 101, 106, 105, 109, 107, 106, 104, 106, 108, 109, 112, 114, 117, 117, 116, 111, 106, 105, 103, 102, 103, 
    
    -- channel=122
    32, 33, 32, 33, 33, 32, 35, 33, 25, 20, 16, 11, 18, 32, 39, 37, 36, 37, 39, 42, 48, 50, 52, 53, 53, 51, 48, 44, 40, 37, 
    32, 33, 32, 31, 33, 35, 44, 41, 15, 11, 16, 8, 2, 11, 28, 38, 42, 42, 39, 40, 44, 43, 40, 35, 30, 25, 20, 18, 16, 16, 
    33, 32, 31, 29, 33, 34, 36, 34, 17, 18, 26, 28, 18, 8, 13, 26, 37, 39, 29, 22, 16, 13, 8, 4, 3, 3, 2, 4, 8, 13, 
    38, 38, 34, 32, 36, 35, 27, 25, 28, 26, 24, 25, 25, 18, 14, 17, 15, 10, 0, 0, 0, 0, 0, 0, 0, 5, 8, 14, 21, 27, 
    40, 41, 39, 36, 43, 54, 50, 30, 24, 19, 13, 10, 11, 9, 2, 4, 8, 2, 0, 0, 0, 0, 0, 5, 15, 22, 26, 29, 33, 35, 
    38, 38, 38, 38, 43, 53, 57, 42, 24, 21, 18, 14, 9, 0, 0, 0, 6, 22, 23, 10, 3, 3, 11, 22, 26, 27, 28, 26, 23, 22, 
    35, 32, 26, 16, 2, 0, 17, 33, 23, 13, 2, 0, 0, 0, 0, 0, 0, 12, 28, 25, 12, 6, 8, 19, 20, 15, 15, 14, 12, 8, 
    14, 2, 0, 0, 0, 0, 0, 21, 17, 8, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 14, 7, 1, 1, 7, 4, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13, 20, 19, 24, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 22, 13, 20, 21, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 23, 1, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 1, 
    0, 0, 3, 7, 1, 0, 0, 23, 28, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 10, 20, 
    10, 10, 8, 6, 0, 0, 0, 0, 26, 44, 42, 26, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 19, 21, 27, 32, 
    10, 7, 1, 0, 0, 0, 0, 0, 0, 18, 47, 28, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 10, 28, 33, 29, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 11, 8, 13, 15, 6, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 1, 9, 5, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 7, 9, 7, 20, 29, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 0, 0, 6, 15, 20, 33, 35, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 13, 13, 15, 20, 14, 
    0, 0, 0, 0, 16, 79, 76, 47, 23, 23, 23, 20, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 9, 8, 0, 0, 5, 11, 
    0, 0, 0, 0, 3, 39, 43, 40, 35, 37, 41, 35, 24, 23, 28, 17, 2, 1, 3, 3, 2, 0, 0, 0, 0, 4, 0, 0, 0, 10, 
    0, 5, 32, 34, 9, 0, 0, 0, 25, 45, 44, 36, 25, 15, 24, 44, 39, 27, 22, 13, 0, 0, 0, 0, 0, 5, 1, 0, 0, 3, 
    57, 70, 69, 53, 29, 9, 11, 8, 3, 17, 28, 24, 12, 0, 0, 16, 29, 18, 11, 4, 0, 0, 0, 0, 0, 9, 7, 0, 0, 0, 
    78, 63, 48, 42, 41, 36, 24, 9, 0, 0, 0, 0, 1, 6, 7, 0, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 0, 0, 
    48, 44, 42, 37, 29, 19, 10, 8, 10, 3, 0, 5, 21, 22, 13, 5, 9, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 0, 
    40, 38, 29, 17, 9, 9, 18, 31, 42, 40, 24, 13, 26, 27, 13, 8, 12, 18, 21, 26, 20, 7, 3, 1, 0, 0, 0, 7, 12, 9, 
    24, 18, 13, 15, 22, 31, 40, 42, 38, 27, 12, 1, 3, 9, 11, 19, 22, 27, 35, 47, 51, 33, 13, 3, 0, 5, 8, 8, 12, 17, 
    11, 17, 28, 38, 42, 40, 35, 28, 22, 14, 4, 0, 0, 1, 8, 20, 23, 27, 30, 35, 42, 39, 25, 17, 12, 12, 11, 9, 13, 19, 
    33, 42, 45, 41, 32, 21, 14, 12, 12, 14, 10, 4, 2, 2, 8, 9, 9, 13, 14, 17, 23, 30, 30, 28, 20, 12, 9, 11, 15, 19, 
    53, 45, 35, 24, 17, 15, 14, 12, 11, 13, 11, 7, 5, 0, 6, 6, 7, 8, 9, 11, 14, 16, 16, 17, 13, 8, 9, 15, 19, 20, 
    
    -- channel=123
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=124
    108, 104, 102, 103, 109, 113, 113, 113, 117, 114, 105, 95, 93, 91, 84, 78, 76, 77, 76, 68, 64, 59, 52, 46, 39, 34, 32, 26, 19, 15, 
    107, 102, 99, 100, 108, 107, 104, 111, 108, 111, 113, 102, 89, 84, 83, 78, 73, 74, 70, 62, 57, 50, 42, 36, 30, 27, 27, 24, 22, 23, 
    106, 102, 96, 100, 104, 83, 90, 114, 105, 108, 122, 120, 103, 88, 80, 70, 64, 67, 61, 53, 46, 40, 38, 36, 36, 38, 40, 40, 40, 41, 
    107, 105, 97, 101, 98, 69, 87, 106, 99, 97, 105, 114, 112, 100, 86, 66, 55, 58, 59, 56, 54, 53, 56, 57, 60, 64, 64, 63, 60, 57, 
    103, 104, 97, 94, 91, 80, 91, 92, 87, 83, 83, 90, 91, 89, 88, 79, 76, 76, 78, 82, 85, 84, 83, 77, 81, 83, 79, 73, 65, 56, 
    96, 98, 94, 81, 65, 67, 85, 91, 82, 83, 82, 79, 78, 81, 83, 88, 101, 111, 108, 105, 104, 104, 93, 81, 82, 80, 74, 65, 54, 44, 
    91, 91, 87, 64, 34, 29, 55, 79, 76, 76, 73, 68, 73, 82, 86, 86, 91, 111, 118, 117, 115, 105, 88, 76, 72, 68, 64, 57, 48, 39, 
    83, 84, 83, 74, 54, 21, 35, 66, 73, 79, 75, 69, 74, 77, 84, 85, 82, 91, 105, 116, 118, 105, 86, 74, 71, 65, 59, 53, 48, 43, 
    90, 101, 112, 128, 106, 41, 45, 66, 78, 102, 110, 103, 100, 86, 83, 87, 87, 87, 93, 101, 111, 112, 97, 84, 75, 66, 59, 55, 55, 54, 
    132, 147, 163, 178, 127, 52, 54, 66, 69, 100, 124, 132, 126, 107, 93, 90, 89, 87, 88, 90, 100, 110, 108, 98, 87, 77, 68, 66, 66, 65, 
    173, 182, 190, 195, 126, 52, 49, 70, 62, 84, 111, 123, 125, 116, 102, 94, 91, 86, 85, 85, 88, 96, 103, 102, 96, 89, 79, 74, 73, 71, 
    188, 189, 189, 191, 138, 58, 44, 75, 89, 101, 120, 117, 114, 110, 105, 102, 100, 89, 88, 89, 84, 87, 98, 102, 94, 93, 88, 82, 80, 75, 
    187, 183, 179, 178, 153, 77, 31, 49, 97, 121, 142, 140, 120, 108, 104, 109, 107, 97, 93, 93, 85, 82, 102, 107, 97, 95, 95, 86, 79, 69, 
    175, 172, 168, 167, 163, 120, 56, 33, 44, 72, 114, 127, 108, 104, 104, 111, 113, 107, 100, 97, 87, 82, 99, 107, 99, 94, 92, 79, 65, 55, 
    164, 163, 165, 170, 172, 162, 133, 95, 23, 16, 64, 90, 84, 90, 105, 120, 128, 124, 113, 101, 90, 85, 90, 102, 96, 84, 74, 66, 57, 55, 
    166, 169, 174, 175, 161, 145, 155, 148, 83, 46, 73, 85, 88, 84, 102, 126, 136, 136, 122, 105, 95, 90, 87, 98, 96, 81, 72, 70, 63, 60, 
    173, 175, 176, 175, 159, 120, 144, 177, 157, 111, 105, 102, 115, 91, 94, 118, 133, 136, 124, 110, 100, 96, 89, 95, 98, 91, 87, 80, 59, 39, 
    175, 182, 196, 214, 223, 179, 168, 199, 205, 177, 120, 113, 135, 110, 96, 113, 131, 135, 129, 119, 109, 102, 92, 94, 99, 91, 76, 58, 32, 13, 
    211, 232, 257, 279, 295, 283, 220, 200, 206, 223, 147, 119, 135, 122, 100, 112, 128, 132, 130, 126, 119, 109, 97, 93, 94, 73, 48, 25, 11, 5, 
    272, 285, 295, 280, 273, 304, 248, 198, 194, 217, 163, 129, 133, 122, 109, 116, 125, 128, 128, 127, 124, 111, 100, 91, 84, 63, 34, 14, 7, 5, 
    302, 307, 296, 219, 175, 203, 188, 173, 179, 178, 149, 128, 127, 119, 120, 127, 128, 130, 130, 126, 115, 103, 92, 80, 75, 67, 42, 17, 7, 8, 
    315, 318, 293, 190, 133, 127, 120, 124, 135, 135, 121, 114, 102, 88, 102, 126, 134, 131, 127, 117, 105, 99, 88, 75, 67, 71, 58, 28, 10, 10, 
    300, 277, 243, 188, 157, 144, 120, 90, 80, 85, 93, 103, 100, 63, 53, 82, 107, 111, 112, 111, 110, 107, 93, 73, 58, 67, 68, 44, 18, 9, 
    229, 201, 181, 167, 153, 141, 122, 87, 53, 41, 61, 98, 115, 79, 50, 60, 82, 95, 107, 117, 120, 119, 105, 70, 47, 49, 63, 58, 34, 14, 
    161, 154, 146, 138, 126, 118, 116, 108, 83, 60, 65, 93, 107, 98, 79, 78, 91, 106, 123, 139, 133, 127, 121, 93, 57, 38, 48, 61, 54, 27, 
    127, 123, 119, 116, 114, 112, 114, 112, 102, 86, 73, 69, 83, 97, 90, 81, 91, 110, 139, 162, 152, 134, 125, 112, 78, 51, 38, 51, 61, 41, 
    103, 102, 107, 112, 112, 105, 93, 76, 67, 72, 61, 44, 52, 78, 79, 71, 79, 93, 121, 147, 146, 129, 114, 107, 84, 57, 37, 37, 51, 50, 
    96, 99, 101, 99, 89, 72, 54, 40, 40, 59, 62, 47, 52, 61, 53, 49, 52, 59, 72, 91, 105, 108, 101, 90, 68, 46, 32, 26, 33, 45, 
    93, 86, 73, 61, 48, 34, 25, 21, 32, 56, 61, 54, 60, 45, 34, 25, 21, 29, 34, 41, 57, 72, 73, 62, 44, 29, 22, 19, 18, 29, 
    67, 50, 35, 29, 25, 19, 17, 16, 28, 50, 55, 54, 51, 32, 26, 14, 10, 19, 20, 19, 26, 34, 33, 29, 21, 13, 12, 14, 12, 14, 
    
    -- channel=125
    1, 0, 0, 0, 0, 12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 28, 50, 72, 81, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 94, 106, 115, 100, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    112, 121, 124, 123, 98, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 6, 3, 
    120, 123, 119, 114, 96, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 11, 1, 
    111, 109, 106, 99, 93, 57, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    91, 92, 92, 93, 98, 89, 46, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    77, 84, 92, 103, 112, 107, 77, 49, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    85, 98, 108, 112, 105, 90, 58, 44, 62, 29, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    98, 107, 116, 131, 140, 130, 117, 91, 105, 90, 60, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    124, 149, 184, 222, 245, 227, 193, 146, 111, 107, 85, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    215, 246, 274, 298, 289, 257, 212, 147, 83, 89, 77, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    287, 297, 301, 292, 231, 165, 125, 71, 33, 37, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    304, 309, 303, 244, 133, 36, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    306, 299, 263, 183, 92, 27, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    235, 190, 148, 114, 87, 64, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    107, 86, 79, 74, 59, 41, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 43, 35, 26, 20, 18, 20, 20, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 4, 2, 5, 11, 15, 14, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=127
    47, 46, 48, 54, 56, 53, 51, 59, 77, 95, 105, 102, 86, 71, 63, 60, 58, 58, 56, 55, 51, 47, 47, 47, 51, 56, 60, 64, 69, 75, 
    46, 46, 48, 56, 57, 46, 49, 66, 93, 109, 117, 120, 117, 105, 89, 73, 63, 58, 61, 65, 65, 66, 70, 75, 83, 90, 95, 98, 100, 101, 
    46, 48, 51, 58, 57, 53, 65, 80, 102, 109, 112, 117, 126, 131, 123, 103, 82, 71, 79, 90, 101, 107, 112, 116, 119, 120, 118, 115, 111, 106, 
    42, 43, 49, 53, 56, 68, 76, 85, 99, 111, 118, 123, 130, 141, 148, 140, 125, 110, 113, 123, 134, 136, 134, 130, 124, 119, 114, 108, 102, 97, 
    42, 42, 47, 50, 50, 57, 65, 91, 112, 131, 144, 148, 153, 163, 174, 174, 158, 142, 129, 125, 124, 129, 125, 119, 109, 100, 94, 93, 94, 95, 
    47, 47, 51, 53, 53, 53, 66, 87, 115, 133, 144, 154, 168, 187, 200, 195, 166, 137, 116, 111, 116, 122, 119, 111, 99, 90, 90, 98, 109, 118, 
    55, 58, 65, 84, 105, 107, 100, 97, 117, 140, 155, 170, 181, 192, 204, 202, 185, 155, 127, 117, 122, 127, 130, 124, 113, 107, 110, 120, 133, 145, 
    80, 91, 107, 135, 151, 143, 126, 116, 130, 152, 171, 187, 193, 195, 201, 208, 207, 188, 164, 142, 139, 148, 153, 149, 137, 133, 138, 150, 162, 173, 
    124, 132, 138, 140, 128, 123, 115, 118, 121, 128, 140, 163, 174, 183, 194, 202, 206, 202, 193, 181, 170, 165, 164, 161, 161, 167, 176, 183, 185, 185, 
    131, 124, 114, 102, 94, 101, 105, 116, 119, 119, 122, 132, 139, 151, 175, 191, 197, 203, 207, 205, 192, 172, 163, 164, 176, 188, 194, 190, 184, 178, 
    101, 94, 84, 74, 87, 98, 108, 116, 136, 147, 147, 136, 133, 138, 158, 179, 187, 195, 206, 213, 202, 181, 170, 174, 184, 190, 192, 185, 173, 160, 
    79, 76, 71, 62, 85, 105, 112, 105, 115, 136, 148, 150, 145, 150, 156, 171, 174, 181, 192, 204, 200, 184, 180, 182, 190, 186, 176, 163, 144, 128, 
    63, 66, 68, 69, 89, 125, 136, 129, 97, 86, 96, 119, 133, 151, 165, 168, 165, 167, 178, 189, 193, 184, 177, 176, 175, 170, 149, 130, 113, 106, 
    64, 73, 81, 90, 102, 135, 167, 177, 139, 94, 86, 110, 141, 159, 177, 175, 167, 161, 167, 178, 186, 187, 176, 168, 157, 150, 129, 113, 111, 119, 
    83, 95, 103, 107, 104, 103, 132, 158, 181, 170, 162, 162, 175, 182, 183, 173, 156, 148, 154, 167, 180, 187, 178, 166, 153, 146, 139, 136, 142, 147, 
    102, 110, 113, 114, 117, 112, 124, 149, 198, 210, 188, 181, 180, 194, 182, 159, 141, 131, 142, 159, 175, 183, 179, 166, 156, 153, 161, 161, 158, 145, 
    111, 121, 135, 152, 177, 186, 176, 168, 169, 200, 170, 172, 169, 190, 185, 158, 138, 128, 139, 157, 171, 178, 176, 164, 155, 148, 150, 148, 145, 145, 
    147, 167, 178, 176, 176, 189, 162, 144, 127, 160, 165, 154, 150, 170, 179, 159, 135, 126, 135, 151, 166, 172, 174, 163, 152, 140, 139, 146, 157, 167, 
    174, 169, 151, 114, 81, 85, 95, 96, 104, 114, 139, 134, 149, 162, 176, 163, 140, 130, 137, 150, 162, 168, 169, 161, 150, 151, 160, 176, 181, 179, 
    131, 118, 101, 59, 19, 0, 18, 51, 87, 90, 111, 118, 141, 156, 165, 163, 152, 143, 146, 154, 158, 159, 159, 156, 155, 171, 186, 197, 192, 182, 
    92, 87, 76, 58, 45, 30, 43, 60, 77, 86, 98, 112, 120, 128, 133, 142, 147, 143, 144, 148, 152, 159, 164, 169, 170, 183, 196, 202, 199, 189, 
    54, 26, 10, 42, 81, 111, 110, 92, 80, 85, 103, 119, 126, 123, 113, 104, 111, 120, 130, 144, 158, 169, 176, 179, 180, 186, 197, 202, 203, 194, 
    0, 0, 0, 29, 62, 84, 92, 95, 102, 103, 114, 131, 145, 143, 128, 114, 108, 121, 138, 149, 153, 159, 173, 184, 191, 187, 191, 199, 205, 202, 
    0, 0, 22, 36, 45, 55, 81, 112, 132, 141, 144, 145, 141, 144, 141, 138, 134, 139, 150, 151, 145, 147, 167, 194, 212, 204, 192, 196, 202, 203, 
    31, 36, 39, 50, 68, 86, 101, 115, 126, 134, 142, 132, 121, 126, 134, 133, 127, 129, 140, 139, 133, 132, 150, 183, 208, 221, 205, 193, 193, 195, 
    52, 57, 71, 87, 100, 106, 104, 98, 97, 110, 124, 130, 123, 122, 134, 135, 127, 120, 115, 104, 99, 107, 127, 155, 188, 211, 211, 195, 186, 187, 
    84, 95, 101, 102, 101, 102, 106, 115, 128, 143, 157, 159, 152, 142, 145, 143, 134, 122, 103, 83, 77, 94, 123, 145, 169, 194, 207, 201, 188, 180, 
    105, 105, 100, 98, 105, 120, 139, 158, 171, 171, 170, 169, 168, 163, 169, 167, 158, 146, 130, 112, 101, 109, 128, 142, 161, 188, 207, 210, 194, 175, 
    96, 99, 109, 126, 147, 165, 178, 185, 188, 180, 171, 171, 169, 180, 194, 200, 194, 184, 174, 160, 147, 141, 146, 155, 173, 194, 209, 211, 198, 177, 
    99, 120, 146, 170, 184, 187, 187, 186, 189, 187, 179, 176, 175, 192, 205, 214, 212, 203, 196, 188, 182, 178, 181, 188, 197, 204, 207, 203, 193, 179, 
    
    -- channel=128
    0, 0, 0, 94, 202, 234, 208, 193, 197, 211, 218, 224, 231, 226, 222, 222, 214, 183, 127, 93, 88, 149, 237, 259, 262, 266, 265, 266, 265, 262, 
    0, 0, 0, 70, 185, 230, 194, 171, 184, 194, 203, 208, 223, 228, 226, 226, 219, 199, 149, 94, 88, 176, 255, 266, 269, 271, 272, 273, 273, 270, 
    0, 0, 0, 45, 159, 215, 176, 153, 177, 190, 187, 183, 193, 205, 218, 226, 226, 217, 178, 113, 110, 205, 266, 274, 277, 275, 274, 274, 272, 268, 
    0, 0, 0, 24, 132, 197, 165, 149, 172, 196, 188, 168, 163, 174, 190, 208, 212, 205, 173, 133, 148, 224, 260, 269, 272, 273, 273, 276, 276, 271, 
    0, 0, 0, 7, 107, 188, 177, 157, 173, 205, 198, 163, 142, 137, 154, 175, 174, 171, 153, 144, 190, 240, 253, 264, 270, 268, 271, 275, 273, 271, 
    8, 0, 0, 12, 114, 205, 198, 160, 171, 210, 210, 179, 148, 128, 135, 141, 136, 135, 132, 152, 211, 239, 235, 254, 273, 268, 272, 277, 268, 270, 
    94, 69, 47, 60, 150, 219, 208, 161, 159, 199, 214, 199, 168, 152, 146, 125, 119, 118, 120, 159, 221, 241, 230, 255, 269, 266, 271, 265, 257, 264, 
    173, 139, 111, 141, 208, 243, 217, 157, 147, 185, 207, 208, 193, 180, 157, 125, 106, 116, 120, 156, 223, 241, 246, 279, 287, 291, 291, 262, 248, 259, 
    240, 208, 187, 214, 245, 252, 221, 149, 144, 184, 204, 209, 209, 193, 164, 127, 112, 119, 122, 147, 212, 238, 261, 294, 303, 309, 301, 266, 246, 257, 
    254, 240, 233, 242, 256, 261, 222, 159, 159, 189, 202, 205, 206, 186, 155, 115, 113, 126, 120, 145, 200, 235, 267, 300, 311, 321, 308, 277, 252, 253, 
    258, 247, 239, 245, 260, 262, 216, 175, 175, 188, 194, 198, 198, 182, 145, 119, 126, 142, 125, 150, 193, 222, 263, 302, 315, 325, 317, 292, 267, 258, 
    268, 257, 247, 245, 257, 246, 210, 195, 180, 177, 174, 178, 187, 170, 137, 130, 153, 153, 136, 158, 183, 207, 259, 299, 312, 319, 321, 302, 283, 266, 
    275, 263, 252, 247, 248, 221, 208, 221, 197, 190, 178, 177, 187, 164, 133, 133, 174, 166, 154, 170, 187, 212, 259, 301, 310, 313, 317, 310, 290, 267, 
    277, 261, 249, 250, 237, 196, 201, 232, 208, 187, 171, 177, 181, 165, 145, 159, 184, 180, 173, 171, 191, 210, 250, 288, 308, 311, 313, 316, 287, 272, 
    275, 256, 236, 241, 224, 179, 188, 227, 222, 203, 187, 189, 185, 167, 144, 163, 175, 184, 179, 174, 195, 199, 215, 234, 268, 297, 313, 312, 283, 283, 
    275, 252, 222, 223, 221, 180, 190, 224, 233, 225, 216, 205, 184, 176, 176, 164, 166, 186, 188, 181, 205, 217, 194, 191, 215, 251, 283, 281, 273, 295, 
    282, 252, 217, 208, 220, 196, 195, 222, 228, 221, 227, 225, 204, 192, 202, 169, 152, 177, 187, 173, 202, 223, 179, 160, 181, 214, 245, 244, 245, 282, 
    290, 258, 220, 205, 222, 222, 212, 222, 222, 221, 230, 232, 216, 208, 212, 185, 158, 177, 179, 181, 213, 215, 185, 167, 159, 180, 213, 217, 218, 248, 
    292, 267, 229, 214, 226, 233, 232, 228, 226, 225, 226, 228, 218, 219, 219, 214, 193, 189, 180, 193, 207, 194, 186, 190, 170, 175, 198, 197, 191, 212, 
    288, 274, 242, 224, 227, 236, 244, 238, 232, 231, 226, 210, 204, 218, 211, 216, 220, 200, 194, 204, 191, 172, 180, 188, 180, 188, 197, 188, 177, 181, 
    284, 278, 251, 223, 220, 238, 245, 246, 244, 245, 235, 204, 198, 213, 212, 220, 234, 216, 209, 197, 167, 162, 178, 185, 189, 199, 196, 176, 168, 166, 
    280, 279, 260, 225, 209, 234, 247, 249, 253, 259, 242, 209, 206, 218, 217, 220, 230, 225, 216, 180, 154, 168, 183, 186, 194, 206, 191, 174, 171, 164, 
    278, 279, 269, 230, 206, 228, 246, 248, 249, 246, 229, 200, 212, 228, 222, 221, 223, 224, 206, 164, 154, 175, 184, 177, 189, 204, 189, 181, 169, 157, 
    277, 277, 274, 238, 213, 225, 241, 246, 242, 229, 193, 176, 216, 237, 227, 223, 223, 217, 188, 159, 157, 179, 180, 168, 183, 193, 186, 178, 165, 154, 
    277, 276, 273, 245, 220, 224, 240, 245, 245, 223, 164, 154, 215, 238, 224, 219, 218, 201, 176, 154, 158, 175, 171, 158, 169, 173, 170, 167, 169, 167, 
    277, 274, 270, 248, 222, 221, 240, 248, 251, 219, 157, 160, 221, 228, 212, 208, 199, 181, 165, 140, 152, 170, 162, 155, 158, 152, 150, 159, 170, 171, 
    274, 268, 265, 245, 214, 211, 237, 251, 251, 223, 178, 188, 219, 213, 199, 195, 183, 169, 148, 129, 152, 164, 157, 156, 152, 138, 136, 154, 170, 174, 
    262, 254, 254, 241, 203, 193, 227, 247, 245, 229, 214, 218, 215, 197, 185, 181, 166, 156, 127, 124, 149, 153, 153, 156, 151, 136, 136, 151, 167, 172, 
    244, 235, 247, 239, 195, 176, 208, 239, 240, 232, 228, 219, 193, 168, 164, 164, 155, 139, 114, 131, 145, 147, 152, 160, 151, 140, 142, 152, 160, 167, 
    217, 207, 229, 229, 184, 156, 184, 224, 230, 222, 216, 197, 161, 135, 132, 137, 139, 119, 115, 132, 136, 138, 152, 157, 146, 141, 142, 147, 153, 162, 
    
    -- channel=129
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=130
    0, 4, 40, 36, 8, 12, 1, 0, 0, 4, 5, 5, 8, 10, 9, 3, 0, 0, 8, 19, 19, 22, 13, 8, 15, 14, 14, 11, 11, 14, 
    1, 1, 32, 42, 7, 5, 1, 0, 0, 0, 3, 0, 0, 8, 11, 5, 0, 0, 0, 21, 40, 25, 0, 0, 4, 5, 8, 8, 9, 12, 
    3, 0, 21, 44, 12, 3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 40, 17, 0, 0, 0, 0, 2, 3, 3, 4, 
    5, 2, 12, 39, 18, 5, 21, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 5, 6, 31, 27, 11, 30, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 14, 19, 39, 44, 16, 15, 14, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 51, 54, 53, 41, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 1, 3, 0, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 33, 54, 48, 9, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 8, 0, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 15, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 8, 0, 0, 0, 32, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 9, 0, 6, 0, 0, 0, 10, 27, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 10, 16, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 5, 0, 2, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 17, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 25, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 7, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 0, 0, 3, 9, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 0, 0, 0, 0, 0, 4, 8, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 4, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=131
    0, 0, 25, 143, 207, 201, 196, 196, 192, 188, 194, 200, 199, 198, 209, 223, 215, 165, 96, 83, 150, 225, 256, 255, 249, 245, 245, 244, 238, 232, 
    0, 0, 4, 117, 198, 198, 201, 222, 224, 205, 202, 217, 226, 231, 239, 255, 263, 222, 133, 99, 172, 256, 284, 277, 267, 262, 260, 259, 253, 246, 
    0, 0, 0, 86, 174, 183, 198, 243, 267, 245, 213, 218, 230, 240, 252, 262, 262, 232, 171, 148, 210, 287, 311, 302, 292, 283, 277, 272, 265, 257, 
    0, 0, 0, 54, 145, 168, 188, 250, 300, 291, 231, 194, 194, 209, 232, 244, 236, 214, 188, 195, 247, 302, 325, 323, 316, 308, 303, 297, 290, 282, 
    0, 0, 0, 30, 132, 181, 193, 250, 317, 320, 258, 188, 156, 163, 183, 196, 195, 192, 207, 242, 279, 307, 327, 339, 338, 337, 339, 333, 326, 321, 
    0, 0, 0, 67, 176, 221, 212, 247, 312, 332, 293, 221, 174, 160, 150, 152, 163, 172, 219, 281, 309, 313, 335, 362, 367, 369, 365, 352, 348, 353, 
    75, 48, 87, 166, 227, 242, 219, 233, 294, 332, 323, 278, 228, 195, 167, 151, 157, 168, 210, 283, 319, 325, 358, 387, 391, 384, 358, 336, 345, 366, 
    203, 166, 186, 231, 271, 265, 212, 208, 272, 320, 326, 314, 281, 236, 196, 162, 161, 173, 202, 270, 317, 337, 367, 397, 401, 379, 343, 314, 323, 359, 
    286, 263, 258, 285, 305, 272, 212, 204, 256, 304, 319, 318, 297, 252, 195, 168, 171, 176, 203, 258, 308, 343, 376, 404, 406, 375, 328, 294, 294, 336, 
    304, 294, 299, 315, 313, 274, 228, 228, 268, 304, 315, 308, 278, 231, 189, 174, 178, 184, 205, 251, 291, 335, 386, 411, 409, 383, 332, 290, 281, 304, 
    315, 303, 302, 313, 311, 281, 246, 246, 279, 301, 301, 291, 261, 217, 189, 197, 207, 203, 220, 254, 279, 322, 383, 414, 414, 396, 351, 300, 280, 284, 
    314, 305, 299, 298, 288, 276, 259, 245, 257, 265, 267, 278, 261, 223, 211, 231, 238, 232, 240, 253, 277, 321, 376, 410, 418, 411, 380, 328, 292, 293, 
    310, 300, 296, 280, 246, 254, 274, 261, 252, 254, 270, 282, 261, 228, 228, 250, 257, 251, 252, 264, 285, 325, 375, 405, 417, 421, 410, 363, 321, 326, 
    310, 299, 295, 275, 222, 226, 285, 303, 292, 281, 278, 280, 266, 232, 232, 263, 269, 252, 262, 283, 281, 306, 355, 391, 409, 420, 417, 382, 353, 355, 
    306, 292, 287, 279, 226, 209, 281, 323, 314, 300, 287, 283, 286, 268, 229, 229, 261, 249, 245, 270, 269, 251, 270, 326, 378, 404, 397, 376, 369, 373, 
    298, 271, 266, 275, 249, 221, 275, 331, 328, 324, 323, 296, 284, 287, 239, 195, 233, 246, 221, 251, 269, 211, 177, 227, 302, 345, 346, 340, 359, 381, 
    304, 262, 252, 275, 286, 260, 273, 331, 354, 354, 353, 335, 309, 294, 260, 193, 189, 227, 220, 243, 265, 226, 165, 148, 201, 262, 285, 290, 322, 367, 
    322, 280, 265, 287, 307, 304, 295, 315, 342, 356, 369, 366, 343, 319, 286, 222, 181, 208, 232, 243, 247, 231, 201, 163, 164, 212, 237, 237, 263, 315, 
    339, 306, 286, 300, 319, 324, 316, 308, 318, 333, 341, 350, 356, 339, 320, 292, 231, 220, 248, 238, 218, 206, 204, 201, 202, 219, 222, 205, 206, 245, 
    348, 322, 296, 304, 324, 326, 327, 326, 324, 321, 303, 300, 327, 336, 334, 333, 293, 252, 242, 221, 201, 196, 207, 223, 228, 225, 214, 202, 198, 200, 
    354, 336, 300, 295, 326, 337, 334, 340, 344, 326, 290, 272, 291, 312, 316, 326, 320, 278, 227, 195, 193, 205, 219, 235, 239, 229, 213, 200, 190, 174, 
    352, 343, 306, 288, 322, 353, 354, 351, 351, 337, 303, 275, 285, 303, 303, 309, 309, 272, 211, 179, 193, 215, 226, 240, 253, 239, 217, 197, 175, 162, 
    344, 341, 313, 288, 314, 353, 365, 361, 348, 319, 291, 283, 295, 305, 304, 304, 292, 252, 203, 181, 193, 215, 222, 238, 254, 244, 221, 198, 181, 171, 
    337, 329, 311, 290, 308, 346, 359, 355, 328, 262, 232, 269, 301, 304, 298, 292, 275, 238, 198, 179, 194, 210, 212, 221, 236, 234, 212, 199, 190, 171, 
    331, 315, 298, 282, 299, 340, 356, 346, 303, 219, 184, 241, 291, 289, 276, 266, 249, 219, 183, 174, 191, 202, 199, 199, 201, 199, 198, 198, 188, 176, 
    325, 305, 280, 263, 284, 333, 358, 345, 306, 238, 196, 229, 267, 263, 247, 234, 217, 189, 162, 164, 182, 188, 186, 182, 170, 166, 179, 194, 200, 196, 
    315, 293, 268, 245, 262, 322, 358, 347, 321, 285, 247, 237, 242, 236, 219, 205, 190, 158, 142, 157, 174, 181, 179, 173, 159, 148, 161, 192, 210, 203, 
    295, 280, 259, 229, 242, 306, 351, 349, 327, 304, 277, 254, 231, 212, 201, 185, 160, 134, 132, 150, 165, 175, 178, 170, 154, 150, 166, 186, 198, 195, 
    266, 264, 257, 222, 220, 282, 339, 347, 329, 309, 283, 242, 199, 179, 176, 166, 141, 124, 131, 144, 157, 171, 179, 172, 163, 163, 167, 173, 183, 189, 
    229, 234, 241, 213, 190, 244, 315, 333, 321, 300, 255, 192, 145, 128, 137, 142, 128, 124, 130, 140, 152, 166, 174, 173, 168, 157, 154, 166, 183, 192, 
    
    -- channel=132
    0, 0, 0, 0, 9, 11, 15, 9, 8, 21, 24, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 34, 52, 30, 0, 0, 0, 12, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 40, 70, 28, 0, 0, 0, 0, 25, 38, 17, 0, 0, 10, 46, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 8, 
    0, 0, 0, 0, 33, 61, 13, 0, 0, 0, 0, 43, 100, 109, 89, 74, 79, 83, 31, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 31, 62, 78, 98, 125, 129, 99, 11, 0, 0, 0, 22, 11, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 7, 0, 0, 0, 21, 73, 84, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 0, 
    0, 0, 0, 0, 0, 0, 29, 29, 22, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 0, 0, 0, 0, 29, 55, 35, 0, 
    0, 0, 0, 0, 0, 13, 57, 37, 23, 33, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 13, 31, 71, 72, 37, 16, 
    0, 0, 0, 0, 0, 25, 40, 0, 0, 6, 26, 23, 26, 40, 48, 27, 6, 5, 0, 0, 8, 0, 0, 0, 0, 13, 35, 27, 11, 18, 
    0, 0, 0, 0, 0, 32, 23, 0, 0, 0, 0, 22, 61, 95, 79, 15, 0, 0, 0, 0, 10, 8, 0, 0, 0, 16, 21, 6, 4, 16, 
    1, 0, 0, 5, 25, 37, 2, 0, 0, 9, 32, 47, 58, 61, 27, 0, 0, 0, 0, 0, 1, 0, 0, 6, 9, 10, 9, 0, 0, 8, 
    11, 18, 12, 26, 66, 55, 0, 0, 47, 99, 91, 62, 48, 17, 0, 0, 0, 0, 0, 0, 7, 0, 0, 5, 8, 0, 0, 0, 0, 0, 
    8, 17, 12, 34, 82, 61, 0, 0, 0, 9, 0, 0, 11, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 3, 0, 0, 0, 0, 
    15, 15, 6, 25, 62, 22, 0, 0, 0, 0, 0, 0, 4, 0, 0, 5, 11, 3, 0, 0, 0, 0, 26, 24, 13, 6, 17, 28, 0, 0, 
    26, 36, 31, 33, 45, 0, 0, 0, 0, 5, 2, 20, 33, 0, 0, 14, 47, 14, 4, 20, 36, 88, 159, 162, 83, 32, 48, 64, 15, 0, 
    27, 49, 58, 45, 26, 0, 0, 17, 0, 0, 0, 0, 0, 0, 22, 45, 51, 44, 17, 10, 30, 55, 116, 176, 183, 145, 128, 94, 22, 0, 
    17, 22, 17, 3, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 13, 29, 11, 53, 32, 0, 4, 16, 0, 0, 83, 154, 160, 119, 56, 30, 
    7, 0, 0, 0, 0, 0, 0, 0, 40, 31, 19, 3, 0, 0, 0, 0, 0, 11, 13, 0, 33, 66, 4, 0, 0, 4, 48, 65, 82, 104, 
    2, 0, 0, 0, 0, 1, 1, 0, 16, 47, 72, 81, 49, 6, 0, 0, 0, 0, 0, 0, 58, 72, 27, 0, 0, 0, 0, 33, 50, 90, 
    3, 1, 0, 0, 9, 8, 12, 0, 0, 0, 45, 74, 68, 52, 13, 0, 0, 0, 0, 58, 72, 25, 0, 0, 0, 0, 39, 46, 24, 36, 
    11, 7, 11, 9, 5, 0, 0, 0, 0, 0, 24, 28, 22, 39, 38, 39, 46, 23, 40, 89, 45, 0, 0, 0, 0, 20, 40, 29, 27, 57, 
    16, 15, 18, 4, 0, 0, 0, 0, 0, 21, 20, 0, 0, 0, 6, 15, 37, 58, 79, 59, 0, 0, 0, 0, 0, 11, 7, 6, 29, 49, 
    17, 21, 26, 0, 0, 1, 15, 13, 27, 67, 72, 8, 0, 0, 0, 1, 21, 57, 66, 13, 0, 0, 25, 17, 10, 16, 13, 15, 14, 0, 
    19, 25, 35, 8, 0, 2, 26, 39, 78, 148, 151, 70, 9, 14, 26, 33, 54, 69, 53, 4, 0, 18, 35, 28, 43, 63, 47, 30, 18, 7, 
    19, 27, 40, 28, 0, 0, 10, 20, 67, 123, 90, 21, 25, 48, 52, 61, 76, 78, 56, 21, 10, 30, 36, 33, 63, 93, 65, 25, 5, 8, 
    22, 30, 40, 36, 14, 2, 4, 10, 30, 17, 0, 0, 20, 74, 69, 75, 80, 80, 67, 31, 13, 34, 35, 37, 58, 65, 45, 17, 0, 0, 
    33, 35, 40, 35, 11, 0, 7, 18, 18, 0, 0, 0, 40, 77, 61, 62, 71, 79, 57, 13, 6, 25, 18, 20, 36, 25, 4, 0, 2, 3, 
    59, 47, 36, 35, 17, 0, 11, 26, 19, 0, 0, 22, 64, 56, 44, 49, 62, 69, 30, 0, 13, 23, 8, 10, 18, 0, 0, 0, 20, 41, 
    79, 48, 28, 29, 22, 13, 24, 30, 20, 8, 28, 76, 98, 79, 60, 57, 63, 45, 0, 0, 22, 15, 8, 13, 2, 0, 0, 17, 37, 33, 
    87, 59, 49, 53, 37, 25, 40, 43, 40, 46, 83, 127, 144, 128, 103, 84, 57, 14, 0, 6, 19, 3, 9, 18, 13, 12, 28, 29, 10, 0, 
    
    -- channel=133
    56, 74, 102, 102, 79, 58, 51, 44, 56, 69, 70, 64, 58, 58, 52, 36, 13, 3, 30, 52, 64, 53, 36, 44, 47, 49, 51, 53, 55, 57, 
    57, 67, 98, 111, 96, 69, 51, 31, 23, 46, 57, 57, 46, 40, 39, 34, 23, 5, 5, 23, 47, 40, 34, 44, 47, 50, 52, 53, 52, 53, 
    58, 60, 90, 112, 106, 78, 55, 28, 1, 12, 39, 60, 62, 52, 46, 44, 45, 35, 19, 19, 34, 26, 27, 32, 35, 40, 44, 47, 49, 52, 
    57, 56, 80, 110, 108, 81, 63, 34, 5, 0, 22, 61, 89, 92, 85, 75, 70, 50, 28, 24, 39, 38, 41, 34, 30, 28, 30, 31, 33, 36, 
    59, 58, 71, 96, 90, 63, 49, 33, 18, 0, 7, 39, 67, 88, 97, 93, 90, 65, 31, 18, 21, 33, 40, 34, 26, 23, 22, 20, 19, 17, 
    40, 55, 41, 46, 41, 34, 38, 37, 29, 6, 0, 0, 17, 43, 61, 73, 75, 61, 42, 26, 14, 18, 17, 8, 0, 3, 14, 22, 27, 19, 
    0, 0, 0, 0, 6, 30, 54, 60, 46, 20, 0, 0, 0, 5, 18, 38, 41, 44, 51, 45, 31, 25, 25, 9, 5, 16, 28, 42, 43, 30, 
    0, 0, 0, 0, 15, 37, 50, 64, 58, 36, 18, 3, 0, 4, 19, 30, 39, 41, 51, 53, 32, 27, 29, 17, 22, 33, 38, 55, 59, 44, 
    2, 0, 7, 15, 27, 34, 31, 44, 41, 31, 27, 26, 24, 28, 32, 42, 47, 45, 49, 53, 37, 33, 24, 14, 17, 20, 29, 45, 60, 58, 
    23, 26, 29, 30, 32, 29, 26, 29, 20, 16, 20, 31, 39, 49, 41, 39, 35, 33, 41, 45, 46, 48, 35, 19, 17, 15, 24, 39, 56, 67, 
    31, 31, 37, 42, 40, 27, 30, 34, 30, 30, 33, 34, 35, 34, 30, 23, 18, 11, 29, 31, 37, 48, 40, 22, 17, 11, 14, 30, 47, 59, 
    39, 40, 42, 55, 57, 41, 39, 41, 59, 63, 56, 45, 30, 15, 10, 11, 6, 8, 27, 29, 34, 43, 36, 25, 16, 7, 0, 10, 23, 33, 
    38, 40, 39, 54, 64, 60, 41, 14, 25, 26, 26, 22, 20, 31, 29, 27, 14, 24, 25, 24, 31, 37, 36, 26, 20, 11, 0, 0, 5, 18, 
    38, 39, 39, 38, 52, 61, 38, 2, 0, 0, 8, 13, 8, 16, 40, 38, 25, 31, 26, 26, 29, 53, 55, 39, 26, 22, 21, 7, 11, 18, 
    43, 49, 52, 36, 40, 58, 44, 20, 15, 17, 25, 29, 17, 2, 34, 46, 44, 39, 43, 47, 50, 93, 117, 103, 64, 41, 37, 29, 30, 25, 
    42, 54, 66, 47, 25, 44, 40, 24, 7, 3, 3, 5, 14, 17, 28, 60, 65, 52, 47, 48, 43, 54, 109, 139, 124, 96, 69, 55, 46, 32, 
    28, 40, 50, 45, 18, 20, 30, 25, 8, 0, 0, 0, 0, 6, 7, 44, 68, 62, 46, 47, 38, 15, 36, 76, 107, 111, 94, 83, 73, 50, 
    18, 20, 25, 31, 21, 13, 22, 33, 39, 33, 18, 0, 0, 0, 0, 8, 49, 49, 44, 48, 50, 46, 37, 33, 49, 63, 63, 76, 96, 88, 
    18, 19, 26, 29, 30, 28, 20, 27, 38, 46, 51, 40, 26, 6, 0, 0, 0, 18, 40, 46, 55, 67, 57, 34, 31, 36, 42, 56, 80, 98, 
    21, 21, 34, 36, 33, 32, 23, 18, 15, 25, 42, 55, 54, 32, 17, 0, 0, 13, 43, 54, 56, 60, 47, 34, 36, 43, 50, 53, 58, 74, 
    26, 22, 31, 37, 33, 18, 15, 16, 15, 15, 24, 43, 48, 43, 41, 37, 25, 37, 52, 60, 58, 49, 40, 39, 41, 45, 46, 55, 60, 69, 
    32, 25, 28, 34, 37, 18, 9, 12, 19, 15, 14, 21, 27, 31, 30, 33, 35, 47, 50, 56, 54, 45, 42, 40, 39, 32, 36, 48, 54, 59, 
    37, 33, 28, 34, 38, 28, 21, 21, 28, 40, 37, 33, 26, 25, 28, 27, 36, 41, 43, 50, 51, 50, 50, 51, 44, 34, 42, 41, 42, 42, 
    37, 43, 35, 40, 39, 31, 28, 31, 49, 71, 82, 71, 42, 35, 42, 44, 47, 45, 48, 52, 57, 54, 53, 63, 60, 56, 53, 48, 48, 50, 
    37, 45, 46, 52, 47, 33, 22, 26, 35, 51, 76, 76, 51, 47, 55, 59, 56, 56, 56, 60, 62, 57, 55, 66, 71, 73, 63, 53, 45, 45, 
    37, 45, 51, 60, 58, 39, 21, 20, 11, 3, 24, 45, 47, 58, 67, 66, 65, 68, 63, 69, 63, 57, 59, 63, 65, 72, 69, 54, 40, 33, 
    40, 46, 52, 60, 59, 45, 26, 19, 12, 4, 16, 32, 49, 63, 66, 65, 69, 69, 65, 70, 58, 53, 55, 54, 55, 59, 62, 56, 47, 44, 
    51, 50, 52, 59, 62, 51, 31, 20, 21, 27, 36, 42, 54, 61, 62, 61, 69, 63, 67, 66, 58, 56, 52, 49, 48, 51, 54, 57, 57, 57, 
    63, 60, 49, 55, 66, 60, 40, 24, 21, 28, 42, 56, 70, 78, 72, 67, 65, 57, 66, 60, 61, 58, 55, 45, 43, 47, 54, 61, 62, 54, 
    74, 78, 64, 60, 71, 71, 55, 35, 33, 42, 56, 73, 96, 105, 95, 81, 60, 58, 60, 58, 60, 59, 55, 50, 55, 58, 62, 60, 55, 47, 
    
    -- channel=134
    20, 41, 69, 79, 65, 50, 48, 37, 44, 53, 58, 50, 41, 37, 28, 7, 0, 0, 0, 25, 19, 11, 5, 20, 25, 27, 29, 32, 34, 38, 
    20, 32, 67, 90, 95, 75, 52, 18, 0, 22, 40, 44, 24, 11, 9, 2, 0, 0, 0, 0, 0, 0, 7, 26, 35, 39, 38, 38, 37, 39, 
    22, 25, 59, 89, 109, 88, 54, 16, 0, 0, 17, 50, 58, 45, 33, 30, 40, 36, 0, 0, 0, 0, 0, 9, 16, 23, 30, 36, 41, 44, 
    20, 18, 49, 85, 107, 85, 59, 28, 0, 0, 9, 67, 114, 119, 108, 96, 93, 66, 9, 0, 0, 19, 29, 17, 10, 7, 9, 11, 14, 19, 
    23, 23, 41, 66, 68, 39, 27, 23, 11, 0, 0, 36, 76, 105, 124, 129, 127, 77, 5, 0, 0, 17, 32, 23, 11, 4, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 9, 30, 34, 4, 0, 0, 0, 16, 63, 86, 88, 59, 13, 0, 0, 0, 0, 0, 0, 0, 0, 8, 12, 0, 
    0, 0, 0, 0, 0, 0, 49, 68, 64, 21, 0, 0, 0, 0, 0, 12, 17, 22, 30, 39, 33, 8, 0, 0, 0, 9, 36, 49, 40, 19, 
    0, 0, 0, 0, 0, 22, 51, 70, 67, 43, 15, 0, 0, 0, 0, 6, 18, 21, 40, 53, 27, 0, 6, 11, 21, 39, 48, 58, 53, 38, 
    0, 0, 0, 0, 0, 19, 18, 24, 28, 33, 29, 23, 20, 27, 36, 32, 31, 33, 37, 50, 25, 9, 6, 0, 2, 12, 13, 26, 47, 51, 
    0, 0, 4, 7, 11, 18, 0, 0, 0, 4, 14, 34, 53, 70, 46, 23, 11, 13, 21, 37, 40, 36, 26, 7, 4, 0, 0, 7, 34, 58, 
    10, 13, 19, 29, 32, 13, 0, 4, 19, 33, 41, 49, 48, 37, 12, 0, 0, 0, 0, 16, 30, 36, 33, 16, 7, 0, 0, 0, 15, 41, 
    23, 26, 28, 51, 59, 31, 20, 32, 75, 97, 85, 57, 29, 0, 0, 0, 0, 0, 0, 20, 24, 27, 24, 17, 5, 0, 0, 0, 0, 0, 
    20, 25, 24, 56, 76, 54, 32, 0, 16, 16, 4, 2, 10, 21, 9, 11, 0, 0, 9, 9, 6, 15, 24, 17, 12, 0, 0, 0, 0, 0, 
    20, 24, 22, 38, 57, 51, 31, 0, 0, 0, 0, 0, 3, 7, 19, 27, 18, 14, 2, 1, 10, 45, 60, 45, 23, 13, 13, 0, 0, 0, 
    28, 38, 47, 33, 39, 48, 45, 16, 1, 8, 27, 30, 6, 0, 17, 43, 47, 31, 26, 45, 59, 120, 167, 159, 93, 48, 48, 27, 8, 0, 
    30, 49, 69, 48, 19, 31, 38, 31, 2, 0, 0, 0, 0, 0, 31, 66, 63, 54, 44, 43, 41, 69, 145, 187, 180, 146, 108, 67, 33, 13, 
    10, 21, 35, 30, 0, 1, 23, 23, 0, 0, 0, 0, 0, 0, 0, 33, 57, 69, 39, 25, 25, 0, 12, 74, 135, 160, 134, 101, 78, 50, 
    0, 0, 0, 0, 0, 0, 15, 31, 43, 41, 19, 0, 0, 0, 0, 0, 21, 37, 28, 30, 52, 35, 7, 9, 35, 58, 66, 84, 116, 116, 
    0, 0, 0, 5, 17, 14, 15, 24, 38, 60, 75, 59, 35, 0, 0, 0, 0, 0, 11, 42, 67, 69, 49, 12, 0, 6, 30, 60, 100, 126, 
    0, 0, 13, 24, 27, 27, 13, 2, 0, 15, 54, 73, 73, 37, 5, 0, 0, 0, 31, 66, 63, 48, 29, 9, 10, 34, 55, 53, 53, 84, 
    8, 0, 16, 26, 22, 6, 0, 0, 0, 7, 21, 39, 52, 49, 50, 46, 21, 31, 64, 72, 47, 24, 17, 21, 32, 43, 42, 43, 53, 81, 
    17, 7, 12, 17, 24, 5, 0, 0, 13, 12, 0, 0, 7, 19, 29, 36, 33, 53, 62, 48, 28, 22, 30, 30, 28, 19, 18, 35, 53, 58, 
    24, 16, 11, 11, 24, 27, 20, 21, 37, 55, 44, 27, 9, 11, 19, 21, 34, 50, 39, 25, 25, 39, 47, 43, 38, 24, 29, 32, 27, 13, 
    24, 28, 18, 16, 22, 33, 35, 40, 76, 122, 124, 91, 44, 30, 42, 49, 58, 51, 39, 32, 44, 50, 52, 63, 67, 62, 56, 39, 29, 33, 
    21, 31, 29, 33, 34, 29, 21, 26, 58, 84, 89, 82, 60, 54, 65, 75, 71, 63, 54, 50, 54, 53, 51, 71, 87, 91, 67, 42, 30, 30, 
    21, 29, 35, 43, 44, 33, 15, 14, 6, 0, 0, 23, 57, 72, 80, 83, 78, 79, 64, 61, 56, 55, 54, 65, 74, 76, 62, 42, 19, 2, 
    28, 32, 34, 40, 45, 38, 20, 15, 0, 0, 0, 24, 63, 74, 76, 74, 75, 79, 59, 54, 47, 44, 43, 45, 46, 47, 48, 38, 28, 27, 
    49, 41, 34, 38, 46, 47, 29, 17, 7, 1, 25, 49, 61, 61, 63, 62, 76, 65, 48, 48, 47, 44, 37, 34, 31, 27, 28, 39, 52, 58, 
    65, 48, 28, 32, 51, 60, 46, 23, 13, 17, 40, 66, 86, 90, 81, 73, 69, 43, 41, 43, 50, 43, 39, 30, 19, 15, 33, 57, 62, 47, 
    74, 70, 48, 46, 63, 74, 66, 42, 34, 46, 77, 106, 127, 133, 117, 94, 57, 33, 36, 44, 45, 42, 43, 34, 35, 47, 62, 55, 39, 25, 
    
    -- channel=135
    96, 97, 85, 91, 93, 80, 70, 68, 80, 91, 91, 89, 88, 88, 90, 89, 85, 81, 74, 77, 90, 87, 79, 80, 78, 81, 85, 86, 83, 82, 
    97, 98, 85, 87, 93, 78, 65, 61, 71, 82, 84, 87, 86, 88, 89, 88, 86, 81, 72, 74, 85, 82, 78, 78, 75, 78, 84, 85, 82, 80, 
    96, 97, 88, 86, 95, 80, 63, 53, 61, 75, 74, 80, 81, 79, 82, 80, 71, 68, 79, 85, 83, 80, 83, 82, 79, 79, 80, 79, 76, 74, 
    96, 96, 90, 86, 98, 87, 62, 44, 49, 64, 64, 62, 68, 71, 76, 74, 66, 66, 80, 88, 84, 83, 92, 90, 84, 81, 79, 77, 75, 74, 
    95, 95, 90, 85, 100, 101, 69, 42, 43, 52, 59, 61, 63, 67, 70, 68, 67, 71, 83, 81, 77, 83, 91, 87, 81, 78, 81, 82, 82, 82, 
    100, 98, 95, 98, 111, 111, 78, 45, 36, 45, 61, 67, 71, 74, 66, 65, 73, 72, 76, 75, 73, 83, 83, 73, 67, 69, 74, 80, 85, 86, 
    108, 111, 119, 120, 101, 97, 84, 54, 39, 44, 62, 71, 72, 70, 68, 70, 75, 71, 61, 59, 70, 83, 82, 65, 56, 63, 68, 78, 90, 89, 
    126, 120, 116, 94, 86, 103, 91, 61, 50, 48, 53, 63, 67, 63, 71, 70, 69, 68, 55, 54, 74, 89, 80, 61, 60, 70, 85, 99, 103, 96, 
    119, 117, 97, 87, 100, 107, 95, 72, 52, 46, 50, 56, 59, 61, 61, 65, 72, 67, 60, 60, 78, 95, 84, 73, 81, 93, 110, 122, 114, 106, 
    102, 99, 94, 97, 103, 105, 99, 82, 56, 49, 51, 52, 53, 58, 66, 71, 70, 68, 62, 61, 72, 90, 91, 84, 89, 108, 126, 134, 131, 118, 
    103, 97, 93, 98, 104, 107, 99, 77, 58, 51, 49, 50, 55, 63, 70, 74, 71, 66, 63, 59, 67, 82, 90, 87, 93, 111, 129, 138, 141, 133, 
    107, 105, 99, 101, 103, 102, 91, 67, 58, 53, 49, 58, 65, 66, 68, 67, 66, 66, 65, 56, 68, 82, 86, 88, 94, 105, 120, 132, 137, 140, 
    113, 110, 101, 98, 89, 88, 84, 64, 62, 61, 66, 66, 61, 64, 63, 56, 60, 73, 67, 62, 74, 82, 85, 89, 92, 97, 107, 117, 123, 135, 
    117, 113, 98, 89, 76, 65, 71, 72, 76, 71, 65, 56, 55, 53, 53, 59, 68, 76, 76, 79, 73, 77, 85, 87, 89, 90, 96, 104, 116, 121, 
    118, 114, 95, 80, 66, 41, 50, 61, 65, 62, 55, 53, 65, 66, 53, 49, 75, 82, 75, 76, 71, 75, 79, 86, 87, 87, 90, 102, 118, 116, 
    120, 113, 96, 75, 59, 32, 35, 56, 56, 59, 68, 60, 56, 62, 56, 50, 78, 89, 67, 70, 81, 74, 73, 87, 92, 89, 92, 104, 117, 119, 
    125, 118, 100, 77, 61, 38, 30, 57, 70, 63, 59, 58, 54, 51, 63, 70, 70, 86, 75, 74, 84, 88, 89, 73, 75, 87, 99, 107, 109, 112, 
    130, 127, 107, 82, 60, 48, 44, 57, 67, 57, 55, 57, 51, 51, 65, 77, 70, 79, 80, 70, 72, 87, 98, 81, 69, 82, 92, 92, 94, 99, 
    128, 128, 107, 84, 66, 60, 62, 64, 65, 59, 54, 53, 56, 53, 61, 82, 76, 71, 82, 66, 66, 78, 82, 81, 78, 77, 78, 78, 75, 82, 
    120, 119, 103, 86, 75, 65, 70, 78, 73, 68, 61, 55, 61, 61, 61, 72, 76, 66, 68, 65, 74, 81, 77, 76, 73, 65, 67, 76, 81, 77, 
    113, 115, 104, 86, 80, 71, 67, 73, 74, 70, 68, 66, 66, 62, 53, 57, 71, 70, 64, 71, 86, 85, 73, 69, 64, 64, 71, 79, 79, 75, 
    110, 114, 110, 91, 79, 69, 62, 57, 61, 67, 73, 68, 68, 67, 54, 55, 66, 71, 71, 82, 89, 81, 70, 65, 68, 71, 75, 77, 72, 78, 
    110, 117, 119, 100, 79, 63, 57, 54, 55, 58, 59, 61, 65, 67, 61, 60, 65, 69, 79, 89, 83, 76, 70, 67, 69, 70, 75, 75, 79, 87, 
    113, 120, 126, 113, 87, 64, 53, 53, 55, 45, 39, 55, 63, 67, 64, 62, 65, 71, 84, 83, 78, 76, 72, 67, 66, 70, 72, 76, 85, 82, 
    116, 124, 133, 126, 99, 75, 60, 58, 57, 44, 37, 48, 61, 69, 66, 64, 68, 77, 81, 79, 80, 79, 76, 68, 64, 70, 76, 81, 78, 77, 
    118, 129, 137, 135, 113, 86, 70, 66, 67, 61, 41, 40, 56, 71, 72, 69, 73, 79, 80, 83, 81, 79, 77, 74, 69, 75, 82, 81, 80, 84, 
    117, 128, 140, 142, 119, 90, 73, 69, 74, 75, 52, 37, 55, 76, 74, 72, 78, 81, 83, 89, 81, 81, 80, 78, 80, 81, 78, 80, 82, 79, 
    116, 127, 140, 144, 123, 90, 70, 70, 74, 73, 58, 54, 70, 79, 77, 75, 77, 83, 92, 89, 81, 83, 82, 81, 82, 84, 83, 78, 75, 75, 
    118, 129, 142, 146, 122, 89, 68, 68, 72, 72, 72, 73, 77, 77, 75, 74, 79, 88, 94, 85, 82, 83, 83, 82, 85, 87, 81, 74, 75, 80, 
    126, 132, 143, 150, 121, 86, 70, 66, 70, 72, 72, 71, 78, 78, 76, 80, 83, 91, 90, 84, 86, 84, 81, 82, 87, 81, 75, 78, 83, 84, 
    
    -- channel=136
    63, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    61, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 108, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 55, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 17, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    58, 59, 0, 0, 0, 0, 0, 0, 0, 41, 52, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    54, 57, 27, 0, 0, 0, 0, 0, 0, 39, 89, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    74, 53, 13, 0, 0, 0, 0, 0, 0, 21, 77, 86, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    103, 64, 0, 0, 0, 0, 0, 0, 0, 0, 36, 65, 48, 21, 32, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    61, 35, 0, 0, 0, 0, 21, 0, 0, 0, 1, 18, 32, 39, 51, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 15, 43, 60, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 14, 0, 0, 0, 0, 2, 23, 46, 47, 13, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 33, 53, 33, 0, 6, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 44, 12, 0, 18, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 4, 11, 0, 0, 40, 42, 0, 0, 24, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 11, 17, 0, 0, 44, 61, 0, 0, 11, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 8, 5, 8, 11, 21, 43, 31, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 3, 14, 41, 16, 10, 59, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 45, 39, 19, 59, 50, 0, 0, 0, 0, 0, 24, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 33, 37, 52, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 27, 38, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 2, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=137
    88, 93, 93, 89, 81, 70, 64, 59, 66, 74, 75, 70, 68, 70, 68, 56, 43, 43, 63, 79, 76, 56, 46, 52, 54, 59, 62, 64, 64, 65, 
    88, 92, 94, 95, 95, 82, 68, 52, 46, 61, 70, 71, 63, 62, 62, 57, 45, 34, 41, 55, 59, 48, 47, 53, 55, 61, 65, 65, 64, 64, 
    89, 90, 93, 96, 104, 91, 69, 45, 29, 39, 53, 65, 64, 60, 59, 58, 58, 58, 57, 47, 41, 40, 47, 51, 52, 55, 58, 57, 57, 57, 
    88, 88, 91, 97, 108, 96, 72, 45, 26, 25, 41, 69, 90, 92, 87, 77, 72, 69, 62, 48, 45, 52, 61, 54, 48, 46, 46, 47, 48, 50, 
    89, 88, 90, 96, 101, 84, 60, 43, 31, 24, 36, 60, 84, 99, 103, 97, 95, 83, 62, 43, 46, 65, 74, 63, 50, 45, 41, 39, 39, 38, 
    82, 91, 84, 78, 69, 58, 49, 41, 35, 29, 30, 37, 50, 65, 79, 91, 94, 81, 61, 41, 39, 51, 51, 39, 30, 33, 40, 47, 53, 47, 
    36, 54, 48, 31, 26, 54, 71, 61, 49, 37, 25, 15, 17, 31, 49, 63, 67, 63, 57, 52, 56, 58, 45, 23, 20, 31, 49, 70, 75, 62, 
    0, 0, 2, 14, 43, 75, 85, 78, 64, 47, 35, 25, 20, 26, 41, 47, 53, 54, 55, 60, 63, 62, 51, 38, 46, 62, 80, 96, 91, 74, 
    47, 31, 29, 43, 62, 73, 74, 66, 53, 48, 46, 42, 40, 46, 56, 64, 65, 61, 60, 62, 62, 61, 50, 43, 50, 65, 81, 95, 98, 90, 
    65, 62, 61, 64, 67, 73, 70, 52, 35, 35, 39, 44, 53, 67, 69, 64, 57, 57, 56, 58, 66, 73, 63, 48, 53, 66, 80, 91, 100, 102, 
    69, 66, 69, 75, 77, 74, 65, 49, 39, 39, 43, 49, 59, 68, 65, 51, 43, 40, 46, 47, 60, 73, 69, 56, 59, 66, 76, 89, 101, 107, 
    79, 78, 77, 86, 90, 80, 66, 56, 66, 70, 68, 63, 53, 44, 39, 31, 30, 34, 40, 43, 56, 66, 63, 60, 60, 59, 60, 72, 84, 91, 
    81, 80, 75, 83, 91, 86, 68, 49, 63, 68, 63, 51, 46, 47, 37, 35, 39, 48, 48, 52, 58, 62, 64, 63, 62, 55, 50, 56, 65, 71, 
    82, 78, 68, 68, 74, 72, 61, 33, 23, 19, 23, 27, 35, 45, 52, 55, 58, 62, 57, 52, 49, 65, 73, 69, 64, 58, 57, 59, 65, 65, 
    87, 84, 71, 56, 52, 52, 53, 40, 34, 35, 42, 50, 45, 28, 35, 54, 71, 68, 64, 66, 68, 94, 114, 110, 85, 69, 72, 78, 78, 70, 
    89, 93, 86, 59, 38, 39, 47, 47, 41, 42, 41, 38, 40, 36, 44, 70, 86, 79, 69, 75, 77, 92, 136, 153, 132, 106, 98, 97, 90, 79, 
    85, 89, 83, 59, 27, 20, 35, 47, 34, 16, 9, 12, 19, 28, 41, 65, 78, 84, 68, 61, 58, 55, 75, 102, 129, 137, 127, 115, 101, 87, 
    79, 75, 64, 47, 26, 22, 36, 51, 55, 43, 31, 19, 12, 18, 26, 42, 62, 75, 68, 58, 65, 69, 61, 56, 72, 93, 99, 105, 112, 108, 
    77, 69, 58, 48, 40, 39, 45, 55, 65, 67, 66, 57, 43, 29, 25, 21, 30, 44, 56, 54, 72, 83, 75, 60, 51, 51, 61, 77, 99, 117, 
    74, 71, 69, 63, 55, 52, 53, 51, 47, 51, 64, 74, 69, 51, 36, 20, 15, 27, 52, 70, 81, 78, 64, 52, 45, 50, 66, 75, 78, 90, 
    74, 72, 72, 67, 58, 46, 42, 42, 41, 42, 56, 70, 69, 62, 57, 53, 48, 49, 65, 84, 83, 66, 54, 52, 52, 61, 70, 73, 72, 82, 
    76, 75, 75, 68, 58, 40, 29, 31, 41, 44, 47, 51, 51, 52, 51, 55, 59, 66, 76, 85, 76, 61, 57, 56, 56, 56, 61, 67, 75, 86, 
    80, 81, 80, 70, 60, 46, 35, 33, 41, 49, 49, 49, 43, 44, 46, 47, 54, 65, 75, 74, 65, 64, 65, 62, 57, 53, 59, 63, 69, 69, 
    82, 89, 89, 79, 64, 52, 45, 46, 56, 70, 79, 76, 57, 52, 56, 58, 64, 70, 73, 70, 70, 72, 72, 71, 69, 69, 70, 70, 69, 65, 
    84, 95, 100, 95, 77, 58, 46, 48, 57, 71, 81, 79, 65, 63, 68, 73, 76, 79, 77, 77, 78, 76, 73, 75, 80, 86, 82, 73, 68, 72, 
    85, 97, 107, 109, 93, 66, 46, 45, 41, 31, 29, 45, 62, 75, 80, 81, 83, 87, 84, 85, 80, 78, 77, 78, 83, 91, 86, 73, 63, 58, 
    88, 98, 109, 113, 99, 71, 48, 46, 38, 16, 5, 27, 64, 83, 83, 83, 87, 91, 90, 87, 78, 77, 76, 76, 79, 80, 79, 73, 65, 60, 
    95, 100, 108, 115, 102, 74, 52, 48, 46, 38, 38, 54, 74, 80, 79, 77, 85, 90, 89, 81, 75, 75, 72, 71, 73, 74, 72, 69, 71, 74, 
    107, 107, 106, 114, 106, 80, 59, 51, 49, 51, 60, 71, 82, 85, 82, 81, 87, 87, 85, 78, 80, 79, 74, 70, 70, 68, 67, 74, 80, 79, 
    117, 117, 113, 117, 109, 87, 69, 56, 54, 58, 69, 89, 107, 110, 102, 94, 85, 82, 77, 78, 80, 76, 73, 72, 72, 70, 77, 81, 77, 69, 
    
    -- channel=138
    62, 56, 43, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 58, 47, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 61, 51, 31, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 60, 54, 36, 14, 0, 0, 2, 0, 0, 0, 0, 19, 23, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 62, 58, 42, 12, 0, 0, 0, 0, 0, 0, 0, 9, 24, 26, 28, 29, 18, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 50, 46, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 30, 16, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 21, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 3, 0, 0, 35, 46, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 9, 58, 63, 25, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 22, 43, 25, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 6, 0, 0, 0, 0, 3, 10, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 3, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 4, 0, 0, 0, 25, 12, 0, 0, 0, 0, 5, 29, 41, 38, 25, 11, 4, 0, 0, 1, 0, 0, 0, 0, 0, 1, 2, 0, 0, 
    
    -- channel=139
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=140
    9, 30, 111, 170, 157, 129, 125, 127, 137, 144, 142, 137, 130, 133, 138, 130, 95, 50, 50, 76, 140, 178, 161, 154, 150, 149, 152, 150, 145, 141, 
    10, 18, 94, 173, 173, 135, 132, 140, 139, 145, 152, 155, 146, 146, 155, 160, 143, 89, 39, 59, 154, 192, 179, 174, 168, 166, 166, 164, 156, 151, 
    12, 11, 73, 162, 172, 131, 138, 161, 154, 145, 151, 171, 174, 173, 175, 180, 175, 127, 65, 86, 176, 205, 197, 188, 180, 176, 175, 173, 167, 162, 
    11, 9, 54, 142, 161, 123, 142, 177, 185, 160, 148, 163, 183, 194, 200, 195, 179, 135, 95, 132, 207, 228, 226, 212, 201, 193, 189, 183, 177, 172, 
    11, 11, 36, 115, 147, 123, 137, 182, 212, 184, 141, 129, 138, 163, 184, 184, 170, 141, 129, 168, 210, 227, 236, 232, 224, 218, 216, 209, 200, 192, 
    0, 7, 15, 87, 142, 138, 139, 185, 224, 200, 146, 103, 97, 119, 130, 139, 140, 137, 165, 207, 212, 214, 226, 231, 225, 231, 238, 234, 233, 228, 
    0, 0, 18, 110, 162, 161, 157, 194, 228, 215, 173, 122, 105, 105, 93, 103, 111, 126, 182, 230, 225, 222, 248, 249, 246, 253, 246, 243, 251, 254, 
    34, 19, 88, 163, 190, 173, 146, 179, 224, 228, 207, 175, 151, 126, 105, 106, 116, 130, 177, 227, 223, 233, 265, 265, 267, 260, 234, 235, 254, 268, 
    151, 141, 175, 200, 207, 170, 122, 154, 202, 218, 218, 209, 187, 154, 120, 118, 132, 134, 170, 218, 227, 251, 268, 267, 267, 242, 212, 214, 241, 270, 
    196, 197, 211, 222, 215, 165, 126, 157, 189, 203, 211, 210, 190, 158, 119, 123, 128, 129, 164, 205, 230, 266, 282, 279, 274, 242, 212, 207, 226, 259, 
    211, 206, 218, 232, 219, 165, 147, 177, 201, 210, 214, 202, 171, 133, 116, 129, 131, 124, 163, 192, 216, 261, 289, 288, 280, 251, 218, 206, 214, 236, 
    219, 212, 216, 228, 213, 179, 169, 182, 209, 215, 211, 198, 163, 121, 121, 148, 144, 140, 173, 188, 207, 255, 284, 289, 282, 262, 227, 206, 203, 216, 
    217, 209, 209, 205, 184, 189, 183, 159, 169, 169, 182, 187, 161, 144, 159, 181, 162, 168, 179, 182, 207, 253, 280, 285, 285, 277, 252, 217, 204, 225, 
    218, 208, 206, 176, 143, 180, 194, 167, 159, 155, 180, 186, 157, 139, 174, 195, 174, 174, 182, 191, 205, 252, 283, 284, 284, 289, 280, 237, 229, 250, 
    220, 212, 212, 167, 121, 167, 208, 204, 199, 197, 200, 196, 175, 146, 164, 184, 186, 171, 187, 208, 204, 241, 281, 300, 296, 296, 282, 251, 259, 267, 
    213, 205, 211, 179, 122, 155, 209, 219, 203, 198, 193, 181, 183, 179, 154, 163, 191, 172, 169, 193, 184, 162, 200, 266, 304, 304, 272, 256, 273, 275, 
    201, 183, 191, 188, 147, 155, 198, 225, 216, 212, 199, 177, 179, 184, 137, 133, 175, 169, 152, 184, 174, 110, 104, 156, 227, 262, 246, 249, 277, 281, 
    201, 174, 179, 196, 185, 177, 197, 227, 248, 254, 244, 218, 199, 188, 144, 114, 146, 154, 156, 186, 175, 139, 112, 102, 137, 180, 187, 207, 256, 282, 
    217, 191, 197, 213, 214, 210, 204, 214, 235, 250, 258, 250, 236, 206, 171, 128, 124, 137, 170, 176, 155, 152, 141, 114, 126, 153, 153, 160, 196, 241, 
    233, 210, 212, 224, 226, 223, 213, 209, 212, 219, 222, 235, 246, 225, 214, 188, 148, 152, 175, 160, 138, 144, 142, 136, 151, 160, 149, 143, 152, 181, 
    243, 220, 208, 219, 231, 219, 214, 219, 223, 207, 184, 202, 223, 223, 230, 230, 196, 182, 163, 140, 136, 146, 149, 159, 165, 156, 139, 141, 145, 147, 
    250, 229, 203, 210, 237, 231, 223, 226, 231, 206, 174, 179, 197, 204, 208, 214, 205, 184, 137, 122, 144, 155, 159, 168, 169, 147, 135, 137, 130, 120, 
    250, 238, 203, 205, 239, 246, 242, 240, 232, 211, 187, 190, 197, 199, 200, 201, 196, 163, 119, 124, 150, 160, 160, 176, 176, 151, 145, 130, 114, 107, 
    246, 242, 209, 210, 235, 247, 247, 246, 228, 195, 191, 215, 211, 203, 206, 203, 189, 149, 123, 134, 156, 157, 154, 178, 181, 166, 150, 132, 125, 120, 
    240, 235, 215, 216, 234, 244, 239, 234, 192, 129, 149, 208, 211, 201, 200, 196, 175, 146, 127, 138, 155, 149, 147, 164, 167, 162, 147, 139, 128, 117, 
    234, 226, 211, 211, 233, 247, 240, 227, 163, 87, 110, 178, 192, 189, 188, 176, 158, 140, 121, 138, 149, 140, 142, 145, 136, 138, 145, 143, 129, 117, 
    228, 216, 201, 199, 223, 250, 249, 227, 179, 129, 139, 165, 170, 172, 165, 152, 143, 121, 111, 136, 138, 130, 133, 126, 113, 116, 134, 146, 145, 136, 
    223, 211, 195, 185, 212, 250, 252, 229, 204, 187, 183, 168, 158, 154, 147, 134, 124, 98, 109, 131, 130, 130, 129, 117, 104, 109, 128, 147, 152, 144, 
    213, 210, 190, 171, 199, 245, 254, 232, 214, 205, 192, 169, 151, 148, 140, 125, 104, 87, 114, 123, 125, 131, 132, 116, 105, 115, 131, 142, 144, 135, 
    200, 212, 197, 166, 178, 231, 253, 234, 220, 211, 187, 152, 138, 140, 137, 122, 92, 94, 114, 114, 121, 132, 131, 119, 121, 125, 128, 130, 135, 132, 
    
    -- channel=141
    0, 0, 0, 0, 72, 93, 85, 85, 87, 79, 72, 78, 80, 76, 80, 90, 87, 65, 32, 0, 5, 72, 125, 127, 118, 115, 112, 111, 110, 105, 
    0, 0, 0, 0, 62, 92, 83, 97, 109, 103, 85, 85, 94, 94, 99, 114, 127, 115, 63, 4, 18, 99, 150, 147, 137, 131, 124, 121, 120, 114, 
    0, 0, 0, 0, 39, 78, 76, 106, 140, 136, 117, 107, 115, 118, 121, 132, 140, 125, 73, 27, 57, 133, 166, 160, 152, 145, 140, 138, 136, 132, 
    0, 0, 0, 0, 10, 54, 70, 111, 164, 174, 148, 113, 101, 102, 113, 130, 133, 109, 69, 58, 103, 160, 175, 173, 172, 166, 160, 158, 153, 147, 
    0, 0, 0, 0, 0, 40, 73, 115, 176, 199, 166, 112, 68, 61, 80, 97, 97, 86, 66, 91, 135, 161, 163, 176, 186, 188, 188, 188, 182, 173, 
    0, 0, 0, 0, 3, 79, 104, 125, 178, 205, 172, 119, 71, 55, 62, 60, 54, 62, 76, 124, 170, 172, 164, 192, 210, 212, 219, 209, 194, 193, 
    0, 0, 0, 0, 84, 124, 121, 121, 159, 200, 190, 153, 118, 94, 71, 54, 45, 60, 89, 137, 175, 177, 185, 227, 251, 245, 230, 201, 177, 191, 
    61, 27, 36, 88, 132, 132, 105, 92, 131, 188, 199, 186, 164, 139, 108, 74, 62, 73, 93, 131, 158, 171, 194, 232, 245, 231, 197, 160, 151, 176, 
    126, 115, 116, 136, 150, 139, 96, 75, 117, 173, 190, 191, 183, 159, 111, 75, 64, 77, 89, 122, 154, 171, 199, 231, 235, 212, 171, 128, 125, 153, 
    145, 143, 143, 151, 159, 139, 97, 85, 130, 176, 188, 192, 180, 144, 93, 64, 69, 78, 89, 117, 149, 166, 199, 233, 236, 208, 167, 123, 109, 130, 
    153, 152, 150, 154, 157, 134, 110, 114, 152, 185, 191, 178, 156, 115, 76, 66, 89, 94, 100, 127, 144, 159, 193, 230, 234, 211, 172, 131, 103, 104, 
    149, 147, 141, 147, 147, 121, 120, 135, 151, 161, 156, 153, 147, 115, 87, 104, 124, 121, 124, 141, 141, 157, 194, 227, 235, 222, 193, 158, 117, 99, 
    145, 139, 136, 139, 130, 100, 115, 135, 122, 117, 122, 141, 153, 138, 114, 130, 147, 135, 125, 135, 141, 157, 193, 222, 233, 232, 221, 196, 151, 131, 
    146, 139, 141, 138, 123, 92, 117, 165, 154, 151, 162, 168, 154, 132, 122, 127, 141, 135, 121, 136, 157, 166, 183, 211, 227, 236, 241, 215, 176, 167, 
    149, 138, 144, 145, 133, 109, 127, 189, 195, 180, 172, 170, 156, 145, 148, 131, 116, 128, 126, 128, 152, 159, 155, 164, 198, 228, 233, 207, 177, 183, 
    146, 127, 126, 139, 135, 129, 140, 184, 190, 176, 173, 172, 161, 162, 150, 117, 87, 109, 114, 101, 123, 108, 77, 85, 136, 189, 195, 173, 161, 182, 
    142, 116, 103, 130, 153, 156, 163, 184, 201, 207, 206, 201, 185, 175, 149, 109, 77, 87, 104, 104, 129, 107, 51, 42, 66, 106, 131, 132, 141, 173, 
    146, 121, 109, 138, 176, 178, 178, 188, 200, 219, 233, 229, 217, 202, 166, 116, 88, 72, 93, 119, 133, 112, 76, 60, 51, 66, 91, 102, 119, 148, 
    158, 142, 136, 151, 185, 193, 180, 176, 176, 191, 211, 215, 216, 209, 182, 146, 122, 98, 109, 134, 121, 91, 77, 76, 76, 93, 107, 95, 88, 106, 
    169, 157, 151, 153, 173, 187, 180, 172, 173, 183, 186, 174, 182, 198, 199, 193, 174, 147, 134, 126, 90, 73, 80, 96, 111, 122, 113, 89, 78, 87, 
    175, 167, 157, 148, 161, 184, 190, 189, 192, 192, 170, 143, 148, 173, 184, 194, 187, 168, 138, 95, 63, 74, 100, 115, 125, 124, 102, 87, 87, 80, 
    177, 167, 157, 145, 157, 197, 211, 211, 210, 201, 170, 141, 145, 163, 170, 175, 176, 161, 116, 65, 55, 88, 111, 115, 125, 123, 102, 88, 77, 54, 
    172, 163, 151, 140, 153, 202, 226, 228, 224, 216, 175, 149, 162, 172, 172, 173, 173, 146, 97, 60, 67, 98, 110, 115, 128, 130, 113, 90, 69, 55, 
    166, 157, 141, 134, 148, 193, 221, 223, 223, 197, 140, 124, 163, 177, 169, 169, 161, 130, 90, 65, 75, 94, 99, 107, 121, 124, 105, 87, 77, 71, 
    160, 145, 128, 120, 134, 176, 208, 212, 196, 147, 87, 93, 155, 170, 153, 148, 136, 110, 80, 62, 70, 88, 88, 93, 103, 95, 80, 78, 75, 64, 
    156, 135, 112, 99, 113, 159, 201, 209, 184, 129, 90, 108, 150, 148, 130, 122, 107, 89, 62, 48, 64, 77, 77, 76, 73, 61, 60, 69, 78, 77, 
    151, 126, 101, 83, 93, 144, 198, 210, 191, 159, 147, 146, 142, 119, 103, 94, 84, 62, 36, 34, 58, 67, 66, 65, 58, 43, 45, 66, 87, 94, 
    139, 112, 92, 75, 81, 131, 195, 209, 194, 178, 169, 152, 125, 96, 86, 83, 68, 37, 19, 33, 57, 61, 64, 64, 51, 37, 47, 72, 88, 89, 
    113, 94, 81, 71, 73, 112, 182, 206, 190, 176, 167, 145, 107, 80, 71, 68, 49, 19, 15, 35, 48, 52, 64, 62, 50, 48, 61, 70, 72, 69, 
    83, 74, 72, 64, 63, 88, 158, 197, 190, 181, 161, 117, 68, 41, 38, 43, 29, 16, 23, 37, 40, 50, 63, 63, 61, 61, 56, 52, 58, 71, 
    
    -- channel=142
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=143
    46, 55, 97, 166, 223, 235, 204, 182, 186, 207, 222, 232, 238, 233, 225, 223, 223, 199, 144, 117, 136, 184, 233, 254, 264, 262, 260, 263, 266, 267, 
    46, 53, 80, 143, 196, 211, 180, 152, 154, 168, 181, 189, 208, 213, 204, 199, 200, 189, 158, 148, 155, 186, 219, 234, 243, 243, 246, 252, 257, 260, 
    47, 51, 67, 122, 176, 198, 169, 130, 133, 143, 152, 149, 159, 175, 182, 183, 175, 163, 156, 159, 163, 183, 201, 217, 227, 232, 237, 241, 244, 247, 
    51, 51, 57, 104, 163, 196, 170, 122, 112, 124, 122, 110, 100, 112, 129, 143, 145, 143, 149, 152, 142, 148, 162, 184, 200, 210, 218, 223, 226, 228, 
    55, 51, 52, 89, 158, 206, 186, 132, 98, 106, 112, 107, 99, 97, 97, 101, 103, 117, 135, 141, 133, 127, 132, 149, 159, 169, 179, 188, 198, 205, 
    91, 69, 81, 124, 188, 216, 189, 134, 92, 97, 118, 133, 142, 129, 111, 99, 94, 105, 120, 121, 127, 131, 143, 155, 159, 154, 149, 147, 152, 166, 
    196, 172, 179, 183, 192, 185, 153, 108, 79, 92, 123, 152, 165, 156, 139, 124, 119, 116, 110, 100, 105, 127, 143, 150, 149, 135, 120, 118, 125, 140, 
    239, 248, 225, 183, 163, 156, 137, 101, 76, 80, 103, 130, 145, 148, 137, 120, 117, 112, 100, 93, 108, 133, 140, 138, 129, 121, 116, 113, 122, 128, 
    185, 192, 175, 159, 151, 157, 155, 126, 99, 87, 93, 106, 116, 117, 106, 102, 98, 99, 95, 90, 112, 132, 145, 147, 142, 144, 147, 141, 133, 128, 
    158, 152, 146, 142, 148, 159, 167, 147, 125, 107, 101, 99, 98, 90, 94, 96, 104, 101, 96, 91, 102, 117, 132, 139, 142, 152, 157, 157, 143, 129, 
    155, 149, 141, 134, 140, 163, 167, 147, 117, 97, 90, 90, 98, 102, 106, 111, 114, 116, 104, 99, 100, 113, 121, 127, 132, 149, 159, 163, 153, 137, 
    153, 146, 141, 133, 136, 159, 160, 134, 88, 60, 61, 82, 103, 120, 127, 127, 118, 117, 102, 95, 99, 113, 126, 125, 130, 146, 164, 167, 164, 158, 
    157, 153, 154, 144, 146, 156, 154, 148, 114, 96, 96, 102, 106, 103, 106, 103, 108, 98, 94, 97, 106, 118, 131, 132, 131, 140, 157, 161, 167, 166, 
    156, 156, 162, 169, 175, 172, 158, 162, 154, 145, 125, 109, 102, 99, 101, 94, 100, 98, 105, 107, 112, 114, 120, 132, 135, 136, 136, 143, 151, 152, 
    146, 143, 149, 178, 193, 182, 151, 133, 126, 109, 93, 88, 93, 113, 109, 104, 100, 111, 114, 98, 99, 84, 73, 79, 109, 124, 119, 126, 132, 141, 
    140, 132, 129, 165, 197, 184, 146, 113, 113, 117, 114, 106, 100, 104, 101, 103, 109, 118, 123, 117, 117, 112, 86, 61, 58, 75, 94, 110, 126, 140, 
    146, 142, 137, 159, 199, 187, 150, 115, 121, 135, 139, 136, 121, 109, 121, 118, 125, 126, 138, 143, 146, 175, 169, 135, 87, 65, 83, 99, 114, 132, 
    154, 158, 160, 159, 177, 174, 141, 112, 94, 94, 104, 113, 119, 117, 134, 142, 145, 144, 146, 146, 144, 167, 190, 183, 156, 134, 128, 120, 105, 105, 
    152, 157, 153, 141, 144, 148, 133, 117, 101, 84, 73, 77, 87, 104, 133, 166, 174, 180, 155, 143, 141, 150, 170, 182, 181, 174, 163, 144, 120, 104, 
    143, 145, 133, 121, 120, 127, 133, 132, 133, 117, 91, 76, 76, 96, 113, 144, 169, 179, 152, 133, 139, 156, 172, 179, 172, 161, 150, 148, 146, 128, 
    136, 139, 126, 116, 118, 132, 144, 145, 138, 130, 122, 104, 98, 103, 97, 101, 129, 143, 140, 131, 144, 160, 169, 161, 152, 148, 148, 148, 144, 128, 
    130, 135, 129, 122, 117, 130, 141, 143, 133, 136, 146, 140, 137, 133, 121, 113, 123, 130, 139, 146, 153, 157, 151, 146, 148, 155, 159, 149, 139, 134, 
    128, 133, 133, 129, 117, 114, 120, 124, 123, 127, 138, 142, 148, 149, 141, 135, 134, 137, 151, 158, 158, 149, 139, 138, 142, 154, 154, 151, 153, 159, 
    128, 130, 136, 132, 121, 107, 104, 106, 105, 100, 108, 117, 136, 147, 141, 135, 131, 141, 150, 153, 148, 141, 134, 125, 126, 132, 137, 149, 152, 151, 
    130, 131, 137, 129, 121, 111, 109, 112, 115, 128, 134, 130, 134, 139, 138, 132, 132, 137, 140, 143, 139, 139, 134, 121, 114, 112, 129, 144, 150, 150, 
    132, 135, 137, 130, 118, 110, 113, 119, 149, 192, 205, 175, 143, 135, 138, 135, 135, 131, 133, 134, 137, 136, 133, 123, 118, 119, 130, 143, 159, 167, 
    132, 136, 141, 135, 118, 106, 106, 115, 152, 200, 212, 181, 148, 139, 143, 144, 137, 129, 134, 135, 140, 141, 138, 136, 135, 134, 138, 146, 152, 154, 
    124, 133, 142, 137, 116, 97, 96, 109, 132, 157, 161, 156, 147, 149, 154, 151, 137, 135, 138, 139, 141, 140, 143, 145, 144, 147, 148, 145, 139, 135, 
    114, 126, 143, 141, 113, 85, 83, 102, 119, 131, 136, 133, 132, 138, 143, 143, 136, 141, 138, 140, 136, 140, 143, 147, 153, 155, 147, 135, 132, 138, 
    103, 110, 130, 133, 108, 79, 72, 94, 109, 114, 109, 105, 103, 106, 116, 122, 134, 142, 137, 137, 136, 140, 141, 146, 146, 139, 132, 133, 142, 151, 
    
    -- channel=144
    263, 263, 256, 256, 256, 253, 226, 199, 184, 179, 176, 180, 193, 194, 204, 226, 240, 265, 273, 274, 269, 268, 265, 270, 265, 255, 255, 259, 244, 223, 
    273, 273, 271, 265, 269, 254, 213, 168, 159, 162, 146, 165, 170, 172, 198, 215, 229, 259, 269, 276, 269, 260, 261, 272, 269, 272, 273, 271, 246, 240, 
    274, 273, 274, 274, 274, 247, 174, 100, 96, 92, 82, 103, 95, 100, 127, 129, 152, 183, 213, 244, 250, 242, 252, 273, 273, 283, 287, 269, 255, 256, 
    277, 276, 276, 275, 278, 256, 161, 55, 34, 30, 32, 47, 35, 46, 55, 51, 74, 93, 131, 188, 213, 230, 254, 272, 274, 280, 278, 259, 253, 263, 
    277, 276, 275, 272, 270, 244, 153, 44, 0, 12, 23, 29, 18, 23, 26, 20, 27, 34, 58, 122, 177, 212, 255, 268, 271, 273, 257, 244, 240, 252, 
    277, 276, 272, 269, 254, 217, 153, 48, 2, 46, 76, 69, 51, 34, 24, 22, 13, 14, 28, 60, 145, 199, 233, 260, 269, 264, 260, 240, 227, 233, 
    277, 275, 275, 269, 241, 197, 154, 36, 0, 53, 91, 89, 77, 46, 33, 39, 40, 33, 38, 50, 107, 174, 214, 251, 263, 257, 259, 241, 208, 208, 
    276, 275, 277, 260, 215, 176, 123, 18, 5, 64, 84, 99, 88, 39, 22, 28, 44, 46, 47, 60, 95, 130, 185, 242, 259, 267, 273, 263, 227, 211, 
    272, 275, 275, 244, 194, 132, 82, 0, 0, 30, 20, 43, 49, 15, 9, 16, 28, 40, 35, 43, 77, 102, 152, 209, 244, 267, 282, 263, 240, 233, 
    259, 270, 273, 253, 187, 105, 61, 0, 0, 3, 1, 11, 13, 0, 0, 3, 9, 16, 10, 19, 46, 64, 108, 173, 222, 261, 278, 262, 252, 257, 
    242, 257, 264, 248, 165, 94, 60, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 6, 22, 37, 51, 83, 139, 205, 260, 277, 276, 276, 277, 
    221, 233, 245, 216, 160, 116, 74, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 1, 24, 50, 52, 57, 69, 103, 168, 228, 251, 261, 274, 277, 
    208, 223, 223, 182, 151, 136, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 27, 25, 28, 43, 80, 134, 175, 198, 220, 253, 277, 
    206, 211, 181, 137, 124, 138, 107, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 25, 52, 79, 106, 158, 217, 268, 
    208, 195, 153, 104, 103, 127, 128, 67, 0, 0, 11, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 33, 86, 180, 256, 
    221, 200, 146, 79, 91, 131, 132, 37, 1, 4, 20, 18, 21, 13, 28, 17, 5, 13, 15, 13, 35, 35, 12, 5, 0, 7, 34, 63, 153, 236, 
    205, 184, 127, 65, 85, 139, 100, 0, 0, 20, 26, 28, 24, 24, 51, 29, 41, 56, 40, 56, 84, 65, 55, 44, 33, 49, 50, 54, 118, 203, 
    213, 191, 128, 64, 85, 127, 51, 0, 0, 19, 28, 27, 16, 27, 31, 32, 66, 61, 39, 61, 89, 62, 50, 55, 55, 79, 62, 40, 83, 175, 
    220, 194, 125, 44, 62, 88, 21, 0, 0, 0, 2, 0, 0, 5, 2, 28, 75, 71, 53, 61, 66, 60, 59, 54, 74, 86, 49, 15, 44, 144, 
    215, 200, 137, 41, 45, 50, 12, 0, 0, 0, 0, 0, 0, 0, 0, 10, 19, 4, 0, 3, 1, 2, 2, 7, 30, 34, 13, 9, 42, 129, 
    207, 199, 143, 42, 24, 39, 11, 0, 0, 0, 0, 0, 0, 12, 22, 0, 3, 31, 48, 31, 22, 31, 42, 60, 58, 8, 4, 32, 47, 114, 
    191, 188, 133, 43, 15, 34, 23, 18, 1, 0, 0, 0, 0, 9, 24, 0, 0, 35, 67, 38, 35, 41, 53, 90, 54, 0, 0, 28, 21, 95, 
    166, 171, 118, 23, 17, 22, 30, 49, 18, 0, 0, 0, 0, 11, 12, 0, 0, 30, 57, 46, 58, 56, 67, 112, 40, 0, 11, 20, 0, 75, 
    138, 152, 112, 34, 21, 33, 46, 67, 27, 0, 0, 0, 0, 0, 0, 0, 0, 20, 69, 114, 130, 123, 113, 118, 28, 0, 0, 0, 0, 64, 
    120, 134, 108, 60, 35, 40, 64, 74, 27, 10, 0, 0, 0, 0, 0, 0, 0, 0, 34, 111, 132, 124, 121, 84, 1, 0, 0, 0, 0, 57, 
    113, 120, 112, 80, 59, 54, 66, 67, 19, 17, 8, 0, 0, 0, 0, 0, 0, 0, 47, 115, 133, 125, 140, 97, 0, 0, 0, 0, 0, 49, 
    115, 121, 123, 107, 78, 57, 65, 52, 11, 21, 15, 0, 0, 0, 0, 0, 0, 0, 28, 68, 79, 92, 117, 84, 0, 0, 0, 0, 0, 46, 
    105, 110, 109, 98, 82, 55, 59, 33, 8, 17, 12, 0, 0, 0, 0, 0, 0, 0, 1, 7, 17, 40, 78, 53, 0, 0, 0, 0, 0, 46, 
    95, 88, 85, 83, 88, 70, 43, 9, 4, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 26, 58, 39, 0, 0, 0, 0, 0, 64, 
    88, 86, 88, 85, 88, 78, 41, 0, 0, 5, 2, 0, 0, 0, 0, 0, 0, 0, 8, 15, 20, 28, 44, 42, 8, 0, 0, 0, 21, 91, 
    
    -- channel=145
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=146
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 11, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 11, 11, 27, 19, 15, 24, 12, 18, 19, 1, 0, 0, 0, 0, 
    0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 23, 29, 17, 0, 6, 26, 40, 39, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 3, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 6, 25, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 15, 7, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 24, 9, 
    0, 0, 0, 0, 24, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 26, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 5, 4, 14, 34, 0, 0, 0, 0, 0, 0, 0, 4, 7, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 5, 1, 0, 8, 0, 0, 0, 0, 0, 0, 0, 9, 14, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 10, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 8, 8, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 18, 19, 20, 21, 0, 
    
    -- channel=147
    398, 392, 385, 392, 393, 349, 301, 297, 304, 302, 308, 318, 333, 350, 363, 379, 393, 407, 410, 403, 389, 388, 401, 400, 384, 361, 350, 343, 329, 329, 
    423, 423, 422, 422, 414, 362, 293, 275, 284, 290, 297, 298, 312, 337, 350, 371, 390, 394, 394, 388, 376, 378, 396, 408, 406, 386, 357, 351, 358, 357, 
    443, 441, 441, 440, 427, 357, 264, 235, 239, 239, 255, 246, 242, 259, 269, 293, 318, 324, 337, 343, 351, 371, 390, 397, 399, 386, 352, 345, 365, 374, 
    450, 449, 449, 446, 423, 346, 233, 196, 210, 214, 229, 226, 217, 220, 217, 220, 236, 241, 263, 297, 329, 370, 393, 390, 387, 367, 331, 315, 342, 379, 
    449, 448, 449, 440, 419, 356, 237, 185, 221, 250, 258, 261, 261, 261, 250, 235, 230, 226, 223, 265, 320, 367, 401, 398, 373, 343, 309, 283, 308, 367, 
    448, 449, 445, 421, 399, 365, 272, 210, 263, 319, 336, 325, 314, 309, 304, 293, 280, 274, 264, 260, 298, 343, 389, 399, 368, 343, 317, 282, 281, 332, 
    448, 449, 440, 409, 388, 357, 278, 229, 276, 324, 354, 351, 317, 309, 314, 319, 317, 306, 319, 304, 277, 308, 363, 384, 382, 372, 340, 288, 255, 292, 
    447, 448, 440, 408, 370, 327, 257, 221, 252, 285, 317, 339, 314, 297, 301, 306, 319, 312, 316, 337, 312, 300, 337, 387, 406, 398, 360, 312, 290, 303, 
    444, 447, 438, 386, 318, 287, 238, 214, 251, 268, 265, 288, 288, 277, 283, 290, 300, 301, 302, 328, 328, 317, 343, 387, 412, 425, 410, 379, 366, 365, 
    431, 444, 432, 369, 307, 272, 216, 178, 207, 240, 237, 245, 252, 252, 258, 263, 260, 265, 272, 296, 314, 304, 311, 359, 416, 445, 448, 436, 422, 424, 
    411, 430, 414, 372, 320, 267, 197, 135, 153, 209, 227, 234, 230, 222, 220, 220, 219, 231, 244, 254, 267, 268, 279, 339, 410, 443, 450, 449, 449, 450, 
    376, 391, 368, 328, 298, 270, 201, 154, 167, 202, 232, 246, 234, 210, 199, 204, 219, 243, 257, 235, 218, 233, 262, 306, 360, 403, 427, 442, 449, 449, 
    351, 350, 318, 276, 251, 250, 226, 209, 204, 208, 225, 240, 239, 204, 185, 193, 210, 227, 232, 206, 175, 175, 200, 239, 289, 329, 365, 412, 442, 449, 
    345, 303, 250, 228, 229, 257, 245, 213, 213, 203, 175, 168, 177, 174, 159, 156, 163, 169, 170, 162, 143, 136, 152, 175, 206, 232, 270, 354, 425, 447, 
    316, 254, 185, 187, 239, 271, 235, 194, 184, 174, 156, 143, 141, 145, 126, 98, 90, 86, 85, 97, 94, 83, 85, 96, 141, 195, 223, 295, 398, 445, 
    312, 262, 178, 168, 222, 234, 196, 175, 173, 189, 195, 184, 166, 158, 119, 83, 86, 92, 112, 142, 120, 87, 82, 100, 159, 211, 240, 282, 370, 435, 
    327, 269, 186, 175, 204, 171, 128, 141, 176, 186, 191, 206, 212, 202, 180, 182, 187, 185, 205, 235, 221, 187, 175, 185, 216, 240, 247, 251, 325, 417, 
    340, 275, 187, 174, 197, 143, 84, 99, 145, 147, 128, 149, 175, 180, 219, 250, 234, 224, 232, 253, 266, 243, 224, 243, 258, 233, 199, 207, 291, 399, 
    354, 284, 170, 130, 157, 136, 81, 67, 95, 127, 110, 92, 98, 137, 180, 214, 223, 214, 219, 225, 220, 212, 210, 235, 249, 208, 164, 176, 257, 378, 
    359, 300, 179, 106, 117, 125, 86, 55, 59, 89, 97, 95, 105, 110, 111, 160, 194, 177, 164, 166, 165, 166, 179, 171, 174, 186, 171, 173, 240, 366, 
    356, 308, 200, 123, 108, 109, 90, 61, 37, 40, 75, 118, 153, 152, 99, 89, 151, 186, 169, 161, 160, 176, 209, 183, 142, 173, 208, 190, 223, 351, 
    351, 294, 183, 133, 126, 119, 123, 94, 43, 21, 43, 88, 144, 151, 85, 64, 144, 204, 189, 185, 189, 203, 249, 201, 105, 123, 170, 160, 208, 341, 
    344, 281, 147, 89, 127, 163, 176, 132, 64, 27, 16, 27, 65, 94, 76, 48, 92, 164, 191, 200, 211, 215, 218, 181, 100, 67, 97, 127, 197, 332, 
    337, 286, 175, 94, 125, 198, 209, 159, 96, 41, 15, 6, 6, 26, 39, 23, 32, 130, 232, 268, 280, 265, 217, 156, 86, 48, 60, 97, 181, 321, 
    328, 321, 263, 185, 155, 187, 213, 179, 124, 73, 26, 1, 0, 0, 8, 13, 38, 142, 265, 315, 311, 306, 247, 120, 39, 31, 62, 108, 186, 316, 
    327, 340, 316, 251, 199, 202, 210, 175, 142, 103, 41, 3, 0, 2, 16, 36, 61, 122, 219, 279, 298, 300, 247, 121, 27, 21, 67, 121, 198, 317, 
    322, 318, 308, 280, 232, 206, 194, 162, 140, 116, 64, 18, 6, 13, 26, 51, 72, 93, 147, 205, 244, 263, 218, 103, 24, 20, 63, 120, 203, 318, 
    311, 304, 294, 277, 235, 185, 163, 145, 129, 113, 75, 35, 21, 26, 33, 44, 67, 94, 121, 152, 187, 220, 192, 92, 20, 21, 60, 114, 208, 321, 
    305, 300, 288, 276, 247, 180, 129, 122, 118, 102, 75, 51, 40, 45, 51, 56, 65, 82, 101, 123, 147, 175, 173, 101, 23, 24, 62, 124, 230, 330, 
    305, 309, 307, 298, 266, 191, 116, 96, 97, 90, 82, 74, 70, 74, 78, 79, 89, 106, 120, 130, 143, 155, 155, 116, 59, 51, 91, 173, 269, 342, 
    
    -- channel=148
    0, 0, 0, 0, 0, 15, 42, 31, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 19, 47, 44, 65, 76, 66, 83, 103, 98, 103, 96, 82, 73, 63, 59, 53, 33, 15, 7, 0, 0, 3, 9, 0, 0, 
    0, 0, 0, 0, 15, 91, 127, 109, 122, 129, 131, 151, 161, 183, 216, 210, 199, 190, 143, 104, 74, 29, 2, 15, 27, 33, 45, 26, 0, 0, 
    10, 9, 8, 11, 34, 94, 130, 110, 106, 80, 68, 83, 58, 66, 102, 123, 165, 194, 183, 140, 49, 0, 0, 12, 30, 52, 64, 51, 27, 11, 
    11, 10, 11, 29, 49, 57, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 57, 34, 0, 0, 6, 23, 61, 79, 61, 43, 25, 
    12, 9, 16, 53, 71, 67, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 64, 43, 33, 32, 22, 8, 0, 8, 30, 
    10, 7, 19, 46, 37, 53, 100, 24, 0, 0, 5, 0, 0, 27, 38, 14, 0, 0, 0, 0, 0, 43, 75, 56, 22, 0, 0, 6, 20, 30, 
    11, 9, 21, 40, 45, 92, 129, 32, 0, 76, 116, 122, 101, 48, 24, 16, 7, 8, 0, 0, 7, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    17, 11, 22, 79, 131, 163, 142, 26, 0, 32, 42, 83, 104, 47, 23, 25, 27, 42, 27, 8, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 16, 28, 72, 69, 63, 79, 64, 68, 85, 51, 62, 78, 54, 45, 56, 74, 88, 77, 58, 65, 56, 62, 86, 50, 8, 0, 0, 0, 0, 
    47, 38, 68, 87, 14, 0, 26, 57, 59, 63, 25, 5, 22, 46, 60, 69, 75, 56, 34, 52, 88, 89, 52, 12, 0, 0, 10, 8, 9, 10, 
    51, 79, 123, 137, 91, 67, 44, 0, 0, 0, 0, 0, 0, 1, 23, 13, 0, 0, 0, 0, 22, 43, 20, 0, 28, 79, 70, 28, 11, 9, 
    25, 82, 128, 122, 90, 83, 24, 0, 0, 0, 0, 30, 45, 28, 13, 8, 5, 13, 46, 75, 61, 52, 67, 89, 140, 184, 170, 102, 35, 9, 
    4, 83, 153, 128, 35, 0, 0, 0, 37, 79, 117, 134, 148, 121, 75, 66, 86, 124, 165, 179, 133, 89, 93, 121, 153, 172, 166, 126, 67, 18, 
    60, 124, 152, 107, 19, 0, 5, 58, 64, 40, 20, 1, 12, 32, 52, 89, 117, 128, 113, 86, 81, 102, 123, 130, 110, 83, 67, 33, 29, 24, 
    32, 73, 47, 0, 0, 68, 186, 141, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 34, 35, 0, 0, 112, 206, 107, 0, 0, 19, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 22, 33, 
    10, 61, 86, 25, 38, 113, 99, 7, 19, 68, 110, 146, 154, 112, 22, 0, 0, 9, 15, 25, 77, 45, 0, 0, 0, 26, 119, 124, 58, 13, 
    18, 46, 76, 58, 98, 122, 37, 0, 46, 85, 57, 39, 63, 89, 77, 61, 106, 107, 98, 119, 139, 130, 118, 101, 113, 145, 112, 52, 0, 0, 
    26, 46, 50, 15, 55, 90, 29, 6, 48, 65, 38, 0, 0, 0, 29, 116, 145, 74, 56, 86, 100, 71, 43, 57, 107, 112, 0, 0, 0, 0, 
    27, 68, 72, 0, 0, 9, 16, 3, 13, 30, 38, 0, 0, 0, 0, 49, 35, 0, 0, 0, 0, 0, 0, 0, 32, 29, 0, 0, 0, 0, 
    28, 90, 130, 56, 0, 0, 0, 0, 0, 0, 12, 29, 28, 40, 62, 16, 0, 0, 0, 0, 0, 0, 0, 0, 10, 15, 63, 99, 15, 0, 
    48, 105, 142, 85, 56, 0, 0, 0, 0, 0, 9, 45, 115, 172, 161, 38, 11, 94, 95, 9, 0, 0, 45, 180, 151, 38, 101, 136, 2, 0, 
    58, 71, 37, 0, 0, 0, 0, 3, 11, 0, 0, 13, 33, 65, 75, 33, 34, 32, 0, 0, 0, 0, 0, 110, 119, 26, 19, 0, 0, 0, 
    36, 3, 0, 0, 0, 0, 13, 56, 8, 0, 0, 2, 7, 4, 1, 1, 0, 0, 0, 0, 0, 0, 0, 37, 42, 28, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 13, 45, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 160, 160, 116, 132, 151, 61, 1, 0, 0, 0, 0, 
    0, 25, 61, 60, 30, 7, 46, 64, 19, 23, 21, 0, 0, 0, 0, 0, 0, 0, 69, 152, 130, 88, 114, 128, 44, 0, 0, 0, 0, 0, 
    23, 52, 55, 38, 23, 29, 77, 85, 25, 34, 27, 0, 0, 0, 0, 0, 19, 41, 49, 53, 51, 61, 95, 80, 14, 0, 0, 0, 0, 0, 
    48, 44, 24, 6, 11, 47, 68, 58, 22, 32, 25, 0, 0, 0, 0, 0, 0, 0, 1, 19, 41, 68, 96, 77, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 25, 38, 34, 37, 31, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 23, 0, 0, 0, 0, 0, 0, 
    
    -- channel=149
    0, 0, 0, 0, 0, 3, 24, 34, 23, 9, 4, 0, 0, 0, 0, 0, 0, 3, 9, 9, 16, 18, 15, 0, 0, 0, 8, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 35, 47, 33, 43, 45, 51, 57, 48, 44, 40, 30, 42, 38, 31, 28, 26, 11, 3, 6, 24, 17, 9, 2, 
    0, 0, 0, 0, 2, 13, 25, 48, 54, 53, 54, 56, 72, 84, 87, 94, 86, 77, 72, 66, 44, 29, 26, 21, 21, 24, 32, 38, 30, 10, 
    0, 0, 0, 1, 0, 6, 28, 39, 31, 28, 19, 10, 17, 20, 32, 54, 63, 80, 83, 72, 52, 24, 11, 15, 27, 30, 39, 57, 56, 27, 
    0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 43, 50, 34, 4, 6, 22, 30, 43, 58, 67, 47, 
    1, 0, 5, 12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 63, 40, 19, 11, 15, 13, 29, 52, 60, 
    0, 1, 2, 1, 8, 5, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 51, 63, 29, 7, 1, 4, 20, 45, 66, 
    1, 2, 0, 0, 14, 9, 0, 6, 18, 19, 35, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 30, 10, 0, 0, 0, 0, 6, 18, 
    5, 2, 1, 17, 29, 30, 9, 12, 5, 0, 15, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 19, 1, 0, 0, 0, 0, 0, 
    15, 6, 3, 0, 0, 3, 0, 41, 36, 19, 14, 11, 10, 4, 1, 8, 16, 13, 18, 13, 0, 13, 41, 49, 31, 5, 0, 0, 0, 0, 
    27, 19, 18, 0, 0, 0, 0, 31, 44, 28, 0, 0, 0, 9, 16, 19, 19, 10, 15, 27, 32, 31, 30, 34, 25, 5, 0, 0, 0, 0, 
    35, 40, 36, 39, 39, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 33, 36, 46, 52, 43, 26, 12, 2, 0, 
    30, 41, 36, 49, 51, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 10, 10, 13, 28, 41, 55, 72, 82, 88, 74, 46, 18, 0, 
    24, 41, 57, 56, 34, 0, 0, 0, 6, 30, 49, 67, 58, 42, 37, 41, 51, 63, 66, 61, 55, 55, 61, 74, 76, 76, 83, 69, 41, 6, 
    36, 45, 59, 67, 47, 18, 3, 4, 19, 8, 5, 15, 16, 26, 44, 62, 76, 80, 65, 58, 66, 73, 91, 84, 66, 44, 42, 50, 40, 14, 
    16, 11, 7, 38, 54, 73, 47, 35, 12, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 11, 8, 1, 0, 0, 17, 24, 20, 
    0, 0, 2, 28, 52, 65, 67, 52, 20, 26, 36, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 43, 36, 
    4, 3, 23, 54, 61, 29, 43, 59, 40, 44, 72, 81, 85, 47, 10, 1, 0, 8, 27, 27, 16, 14, 7, 0, 6, 17, 45, 64, 62, 42, 
    0, 0, 16, 71, 77, 31, 28, 56, 55, 40, 35, 43, 57, 63, 70, 46, 30, 36, 47, 46, 47, 50, 45, 55, 45, 30, 39, 46, 46, 34, 
    6, 0, 0, 45, 61, 42, 31, 45, 65, 60, 33, 15, 6, 24, 66, 74, 54, 37, 39, 44, 47, 36, 34, 55, 50, 22, 0, 7, 31, 35, 
    9, 0, 0, 6, 28, 25, 27, 28, 50, 66, 50, 23, 0, 0, 21, 55, 44, 19, 4, 8, 13, 0, 0, 6, 21, 23, 0, 0, 28, 42, 
    9, 8, 27, 35, 26, 0, 0, 3, 22, 46, 66, 67, 55, 32, 23, 45, 34, 0, 0, 0, 0, 0, 0, 0, 9, 66, 63, 41, 49, 44, 
    9, 4, 28, 76, 51, 5, 0, 0, 10, 37, 62, 83, 111, 90, 61, 68, 90, 70, 47, 27, 5, 26, 61, 36, 53, 78, 79, 65, 57, 37, 
    4, 0, 0, 8, 29, 19, 2, 0, 8, 27, 43, 57, 73, 71, 62, 68, 80, 49, 8, 0, 0, 0, 5, 21, 52, 56, 43, 35, 40, 30, 
    0, 0, 0, 0, 0, 15, 18, 0, 1, 10, 30, 47, 55, 54, 51, 49, 47, 34, 1, 0, 0, 0, 0, 0, 44, 55, 37, 23, 25, 21, 
    0, 0, 0, 0, 0, 14, 20, 2, 8, 7, 21, 42, 49, 48, 41, 22, 24, 59, 76, 74, 57, 45, 26, 26, 49, 52, 42, 26, 24, 18, 
    0, 6, 7, 0, 0, 23, 26, 21, 24, 17, 22, 33, 38, 38, 40, 39, 39, 60, 73, 73, 57, 35, 21, 24, 45, 48, 46, 32, 26, 17, 
    0, 4, 4, 0, 0, 29, 33, 40, 32, 25, 25, 32, 36, 38, 41, 49, 55, 59, 55, 52, 50, 39, 12, 18, 40, 51, 50, 34, 25, 10, 
    3, 0, 0, 0, 0, 18, 32, 44, 35, 33, 29, 30, 29, 31, 30, 32, 35, 38, 40, 46, 53, 56, 27, 20, 32, 48, 41, 17, 11, 0, 
    0, 0, 0, 0, 0, 0, 21, 49, 44, 35, 30, 20, 15, 13, 14, 14, 12, 8, 5, 7, 16, 24, 15, 1, 7, 18, 7, 0, 0, 0, 
    
    -- channel=150
    0, 0, 0, 0, 0, 3, 24, 29, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 16, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 17, 51, 69, 59, 75, 84, 92, 99, 97, 85, 78, 57, 54, 44, 43, 33, 24, 3, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 6, 40, 67, 98, 115, 103, 118, 124, 139, 172, 177, 176, 171, 146, 120, 91, 55, 30, 24, 21, 25, 26, 28, 21, 8, 0, 
    6, 5, 4, 9, 18, 39, 60, 84, 82, 62, 54, 44, 46, 58, 77, 112, 139, 154, 144, 106, 50, 6, 9, 19, 30, 37, 43, 54, 51, 19, 
    7, 7, 9, 23, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 48, 40, 20, 0, 6, 30, 39, 54, 61, 65, 41, 
    8, 5, 17, 39, 34, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 74, 55, 28, 19, 11, 0, 5, 39, 61, 
    6, 5, 15, 21, 15, 28, 8, 0, 2, 12, 0, 0, 0, 5, 7, 0, 0, 0, 0, 0, 18, 61, 80, 47, 0, 0, 0, 1, 47, 72, 
    7, 10, 9, 9, 31, 62, 35, 13, 44, 73, 87, 77, 39, 12, 2, 0, 0, 0, 0, 0, 0, 1, 25, 0, 0, 0, 0, 0, 0, 0, 
    14, 10, 11, 49, 90, 102, 46, 15, 20, 17, 45, 64, 45, 20, 9, 11, 16, 15, 13, 0, 0, 0, 12, 17, 0, 0, 0, 0, 0, 0, 
    34, 16, 17, 29, 19, 22, 16, 61, 76, 60, 46, 49, 43, 32, 30, 39, 56, 56, 55, 50, 30, 43, 78, 88, 50, 6, 0, 0, 0, 0, 
    51, 40, 47, 12, 0, 0, 0, 51, 70, 51, 12, 2, 9, 28, 45, 54, 53, 36, 32, 51, 63, 66, 56, 39, 22, 10, 6, 6, 7, 7, 
    66, 82, 90, 79, 62, 38, 0, 0, 0, 0, 0, 0, 0, 0, 9, 1, 0, 0, 0, 0, 24, 34, 26, 44, 76, 83, 57, 28, 9, 6, 
    53, 82, 83, 89, 84, 52, 0, 0, 0, 0, 9, 15, 11, 3, 4, 3, 7, 24, 41, 46, 52, 61, 88, 125, 153, 164, 135, 86, 36, 6, 
    32, 80, 107, 98, 44, 0, 0, 0, 37, 60, 97, 126, 110, 80, 62, 69, 93, 122, 130, 114, 93, 86, 99, 127, 146, 161, 159, 116, 67, 16, 
    71, 103, 109, 87, 30, 0, 24, 45, 44, 27, 6, 10, 8, 21, 47, 79, 110, 120, 97, 80, 78, 95, 131, 133, 118, 83, 75, 73, 57, 25, 
    30, 27, 2, 10, 39, 113, 116, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 35, 
    0, 3, 0, 1, 53, 126, 121, 69, 7, 7, 30, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 72, 59, 
    10, 23, 31, 49, 82, 66, 50, 42, 49, 82, 120, 128, 125, 84, 0, 0, 0, 12, 44, 56, 33, 15, 5, 0, 5, 46, 97, 120, 88, 55, 
    4, 4, 24, 84, 112, 50, 12, 46, 70, 66, 46, 52, 82, 83, 81, 97, 94, 78, 87, 99, 103, 100, 93, 89, 93, 90, 67, 52, 42, 37, 
    13, 0, 0, 42, 69, 45, 17, 42, 65, 62, 30, 0, 0, 10, 83, 116, 92, 59, 68, 78, 80, 57, 45, 83, 97, 48, 0, 0, 7, 35, 
    22, 17, 0, 0, 5, 7, 13, 10, 34, 61, 40, 0, 0, 0, 10, 68, 48, 5, 0, 0, 0, 0, 0, 0, 12, 6, 0, 0, 16, 47, 
    25, 42, 43, 22, 16, 0, 0, 0, 0, 24, 47, 60, 51, 46, 38, 28, 0, 0, 0, 0, 0, 0, 0, 0, 3, 60, 90, 82, 57, 47, 
    38, 43, 55, 81, 50, 0, 0, 0, 0, 6, 51, 96, 150, 139, 81, 57, 93, 109, 71, 20, 0, 18, 91, 96, 79, 96, 121, 90, 46, 41, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 39, 74, 73, 48, 61, 102, 56, 0, 0, 0, 0, 8, 26, 45, 52, 36, 14, 13, 37, 
    19, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 15, 29, 29, 27, 28, 13, 0, 0, 0, 0, 0, 0, 0, 32, 42, 12, 0, 2, 29, 
    2, 0, 0, 0, 0, 3, 24, 0, 0, 0, 0, 9, 18, 15, 4, 0, 0, 29, 112, 150, 120, 90, 66, 39, 38, 25, 12, 8, 9, 26, 
    4, 30, 35, 12, 1, 17, 41, 27, 18, 5, 0, 0, 0, 0, 0, 0, 14, 76, 127, 134, 102, 70, 54, 21, 20, 15, 22, 23, 15, 22, 
    25, 37, 26, 5, 0, 38, 55, 50, 30, 16, 2, 0, 0, 2, 12, 33, 50, 64, 66, 67, 72, 66, 38, 11, 7, 23, 35, 22, 8, 13, 
    28, 18, 2, 0, 0, 26, 40, 46, 30, 22, 9, 1, 0, 0, 0, 3, 11, 21, 31, 48, 69, 83, 40, 11, 0, 16, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 42, 42, 26, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 5, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=151
    69, 73, 69, 58, 56, 54, 61, 73, 67, 48, 52, 64, 70, 79, 77, 72, 68, 65, 73, 78, 76, 72, 72, 74, 81, 90, 95, 102, 101, 101, 
    58, 60, 62, 55, 51, 48, 44, 48, 46, 30, 28, 28, 33, 40, 37, 43, 50, 54, 77, 90, 82, 75, 71, 69, 72, 80, 91, 101, 101, 83, 
    46, 47, 48, 46, 48, 46, 26, 19, 15, 7, 5, 2, 6, 5, 9, 21, 26, 37, 67, 92, 92, 77, 67, 61, 64, 78, 99, 112, 107, 82, 
    40, 41, 41, 40, 39, 40, 25, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 43, 84, 95, 77, 60, 54, 66, 83, 101, 113, 108, 95, 
    40, 40, 40, 38, 38, 46, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 49, 86, 74, 54, 53, 59, 76, 96, 105, 111, 104, 
    40, 40, 39, 33, 33, 43, 24, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 44, 72, 60, 54, 55, 72, 97, 105, 106, 97, 
    40, 41, 39, 33, 33, 28, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 44, 68, 54, 62, 79, 89, 93, 85, 81, 
    40, 40, 40, 40, 30, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 22, 49, 56, 61, 63, 66, 76, 82, 73, 
    38, 39, 41, 34, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 33, 47, 43, 48, 58, 67, 71, 61, 
    34, 39, 40, 25, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 39, 47, 53, 57, 46, 41, 
    31, 35, 35, 38, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 27, 43, 41, 39, 39, 39, 39, 
    22, 25, 23, 31, 28, 9, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 29, 40, 40, 36, 37, 39, 39, 40, 40, 
    14, 20, 21, 29, 20, 21, 29, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 24, 24, 18, 19, 28, 33, 38, 41, 40, 
    23, 16, 19, 31, 27, 33, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 18, 17, 14, 12, 6, 1, 0, 20, 42, 40, 
    16, 13, 19, 41, 49, 40, 11, 0, 0, 0, 0, 7, 8, 17, 23, 22, 20, 20, 19, 25, 32, 30, 26, 15, 0, 0, 0, 0, 30, 42, 
    17, 35, 35, 45, 38, 24, 10, 4, 9, 24, 33, 30, 17, 21, 26, 32, 46, 52, 50, 54, 43, 42, 54, 45, 29, 6, 0, 0, 14, 38, 
    25, 32, 33, 40, 30, 19, 24, 33, 18, 25, 25, 18, 14, 17, 24, 51, 60, 54, 49, 49, 46, 52, 64, 52, 27, 7, 0, 0, 0, 36, 
    20, 27, 32, 38, 38, 36, 45, 41, 17, 7, 10, 20, 27, 18, 26, 39, 14, 12, 9, 1, 20, 30, 23, 17, 9, 0, 0, 0, 8, 36, 
    26, 34, 33, 32, 41, 53, 56, 35, 16, 20, 28, 25, 17, 25, 25, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 0, 10, 18, 12, 26, 
    25, 35, 33, 33, 43, 58, 53, 38, 37, 42, 36, 30, 26, 24, 9, 9, 19, 8, 0, 0, 5, 6, 12, 2, 0, 15, 19, 12, 9, 24, 
    19, 33, 43, 44, 42, 47, 48, 49, 52, 51, 47, 43, 29, 31, 23, 17, 25, 26, 17, 16, 22, 22, 28, 24, 17, 33, 30, 8, 0, 23, 
    9, 21, 35, 51, 49, 32, 45, 55, 60, 64, 59, 51, 35, 36, 31, 43, 55, 50, 33, 33, 35, 30, 41, 39, 21, 34, 25, 6, 6, 23, 
    0, 14, 31, 46, 56, 42, 36, 42, 53, 69, 61, 46, 36, 44, 63, 60, 41, 34, 37, 35, 27, 20, 17, 28, 44, 32, 24, 35, 26, 13, 
    0, 5, 35, 45, 46, 44, 25, 24, 51, 67, 70, 68, 58, 59, 76, 63, 29, 31, 56, 43, 37, 26, 17, 39, 68, 52, 47, 44, 18, 0, 
    0, 8, 35, 37, 27, 13, 18, 25, 47, 61, 72, 77, 78, 75, 71, 67, 62, 66, 66, 42, 29, 27, 37, 38, 53, 63, 57, 41, 6, 0, 
    0, 6, 14, 5, 2, 11, 26, 24, 39, 53, 64, 75, 81, 78, 75, 73, 65, 40, 21, 13, 15, 17, 32, 53, 66, 69, 56, 31, 0, 0, 
    0, 0, 0, 3, 11, 16, 27, 25, 31, 44, 64, 78, 82, 79, 74, 71, 58, 24, 4, 11, 14, 10, 27, 56, 77, 70, 49, 26, 2, 0, 
    0, 0, 0, 7, 17, 14, 23, 35, 33, 42, 62, 74, 77, 75, 67, 56, 48, 40, 29, 21, 9, 3, 23, 50, 73, 68, 48, 29, 7, 0, 
    0, 0, 0, 0, 10, 20, 27, 42, 39, 46, 59, 68, 68, 67, 63, 58, 52, 44, 35, 25, 14, 8, 31, 58, 66, 67, 51, 33, 10, 0, 
    0, 0, 0, 0, 3, 18, 33, 48, 46, 50, 60, 67, 61, 57, 54, 53, 51, 48, 39, 30, 27, 23, 33, 55, 65, 64, 53, 38, 8, 0, 
    
    -- channel=152
    0, 0, 0, 0, 9, 53, 32, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 12, 84, 77, 2, 15, 25, 9, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 119, 127, 42, 66, 65, 52, 84, 47, 25, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 36, 150, 192, 99, 109, 129, 115, 150, 128, 118, 125, 82, 68, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 36, 138, 237, 157, 122, 158, 161, 184, 173, 176, 195, 178, 162, 145, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 35, 31, 96, 243, 172, 80, 121, 144, 184, 189, 183, 197, 200, 198, 187, 155, 79, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 16, 55, 33, 97, 245, 157, 43, 87, 79, 142, 206, 184, 180, 176, 179, 188, 152, 140, 75, 0, 0, 0, 0, 0, 7, 16, 0, 0, 
    0, 0, 18, 64, 53, 123, 241, 145, 65, 124, 74, 107, 206, 194, 176, 169, 153, 180, 153, 131, 147, 21, 0, 0, 0, 0, 27, 31, 0, 0, 
    0, 0, 20, 92, 101, 135, 226, 136, 96, 177, 136, 122, 187, 188, 172, 167, 150, 170, 156, 124, 154, 79, 0, 0, 0, 0, 32, 36, 1, 0, 
    0, 0, 27, 125, 141, 166, 230, 147, 88, 149, 162, 154, 171, 177, 174, 168, 164, 164, 152, 124, 141, 118, 12, 0, 0, 0, 10, 14, 0, 0, 
    0, 0, 34, 103, 116, 176, 255, 179, 89, 109, 154, 174, 184, 178, 172, 167, 164, 154, 147, 140, 124, 110, 47, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 45, 68, 53, 141, 237, 184, 125, 124, 152, 175, 210, 205, 178, 164, 157, 145, 153, 171, 127, 78, 32, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 56, 57, 34, 87, 157, 163, 158, 160, 169, 164, 202, 210, 175, 151, 141, 131, 138, 158, 124, 68, 30, 0, 0, 0, 0, 0, 0, 0, 
    0, 59, 66, 24, 8, 28, 118, 175, 178, 181, 176, 145, 149, 166, 157, 142, 137, 140, 138, 140, 121, 91, 70, 43, 26, 30, 0, 0, 0, 0, 
    1, 95, 99, 0, 0, 0, 121, 196, 177, 169, 167, 156, 144, 141, 155, 142, 118, 121, 115, 115, 126, 111, 92, 74, 54, 72, 65, 0, 0, 0, 
    10, 116, 137, 0, 0, 8, 128, 162, 128, 117, 109, 140, 153, 140, 169, 143, 101, 114, 93, 92, 161, 143, 104, 89, 65, 92, 104, 0, 0, 0, 
    35, 124, 142, 0, 0, 97, 142, 81, 77, 93, 72, 90, 114, 129, 146, 101, 87, 107, 74, 62, 144, 142, 100, 94, 77, 107, 110, 36, 0, 0, 
    52, 140, 158, 0, 0, 152, 156, 41, 56, 102, 97, 70, 68, 80, 60, 45, 96, 90, 58, 51, 99, 104, 79, 58, 71, 147, 128, 47, 0, 0, 
    48, 154, 196, 24, 0, 133, 149, 70, 68, 100, 129, 111, 84, 68, 29, 25, 120, 124, 88, 97, 115, 105, 98, 59, 73, 173, 153, 60, 0, 0, 
    31, 147, 224, 94, 21, 94, 134, 109, 86, 77, 105, 114, 109, 110, 77, 40, 103, 129, 118, 117, 126, 108, 101, 107, 86, 129, 140, 88, 0, 0, 
    26, 137, 211, 113, 70, 91, 116, 129, 106, 70, 63, 70, 86, 133, 170, 76, 35, 101, 144, 124, 123, 92, 72, 161, 144, 54, 89, 128, 0, 0, 
    43, 153, 207, 70, 65, 101, 106, 145, 133, 85, 54, 35, 28, 99, 189, 77, 0, 43, 133, 99, 106, 71, 17, 177, 190, 18, 47, 120, 0, 0, 
    70, 178, 237, 62, 6, 62, 100, 170, 159, 103, 80, 53, 30, 59, 138, 74, 0, 0, 71, 61, 77, 68, 34, 151, 181, 55, 52, 86, 0, 0, 
    94, 182, 244, 121, 12, 19, 97, 181, 166, 124, 100, 81, 68, 64, 89, 82, 26, 0, 10, 62, 92, 105, 134, 192, 151, 76, 70, 62, 0, 0, 
    92, 135, 202, 164, 92, 30, 93, 177, 149, 140, 126, 92, 76, 74, 69, 81, 53, 0, 0, 33, 79, 84, 174, 242, 134, 64, 52, 50, 0, 0, 
    78, 91, 143, 172, 143, 60, 96, 169, 123, 142, 147, 103, 74, 72, 64, 65, 53, 0, 0, 12, 45, 64, 163, 240, 133, 53, 34, 49, 0, 0, 
    79, 93, 118, 151, 159, 82, 95, 155, 109, 133, 147, 109, 73, 70, 62, 48, 47, 22, 5, 36, 41, 62, 175, 229, 117, 50, 35, 51, 4, 0, 
    100, 113, 122, 129, 151, 123, 103, 128, 105, 123, 130, 106, 76, 69, 70, 63, 57, 59, 60, 59, 50, 58, 162, 219, 112, 49, 42, 49, 0, 0, 
    121, 127, 127, 122, 149, 175, 130, 96, 99, 118, 111, 98, 83, 75, 80, 83, 77, 73, 75, 71, 65, 64, 121, 194, 124, 52, 46, 34, 0, 10, 
    126, 126, 131, 132, 158, 207, 165, 84, 89, 102, 92, 90, 89, 85, 93, 94, 83, 78, 90, 91, 85, 85, 108, 159, 135, 73, 44, 15, 3, 49, 
    
    -- channel=153
    26, 25, 26, 22, 23, 32, 52, 57, 37, 18, 16, 16, 6, 0, 0, 0, 12, 26, 35, 41, 46, 48, 44, 32, 27, 32, 43, 54, 52, 39, 
    17, 18, 15, 12, 11, 22, 35, 49, 48, 34, 38, 40, 45, 48, 43, 47, 48, 49, 64, 69, 67, 59, 52, 40, 33, 39, 60, 66, 53, 36, 
    14, 15, 16, 17, 21, 29, 37, 48, 48, 39, 44, 47, 58, 69, 74, 78, 71, 69, 86, 90, 78, 59, 47, 44, 48, 59, 77, 83, 65, 45, 
    21, 21, 21, 21, 27, 45, 53, 53, 44, 29, 23, 25, 27, 32, 45, 56, 64, 76, 91, 96, 75, 48, 37, 41, 52, 66, 86, 95, 87, 63, 
    21, 21, 22, 24, 22, 23, 18, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 32, 63, 64, 40, 27, 31, 47, 64, 87, 99, 102, 80, 
    22, 22, 24, 28, 30, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 59, 47, 36, 40, 57, 66, 79, 92, 87, 
    22, 21, 23, 27, 31, 25, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 65, 70, 50, 40, 37, 37, 53, 73, 87, 
    22, 23, 23, 22, 21, 19, 8, 5, 9, 19, 30, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 41, 37, 24, 18, 31, 48, 54, 52, 
    25, 23, 24, 30, 34, 41, 20, 2, 0, 0, 3, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 17, 12, 12, 8, 2, 0, 0, 
    31, 24, 24, 29, 34, 33, 14, 23, 27, 19, 7, 11, 11, 0, 0, 0, 4, 8, 6, 0, 0, 2, 26, 42, 37, 23, 6, 0, 0, 0, 
    39, 31, 31, 23, 5, 0, 0, 36, 51, 37, 6, 0, 0, 4, 12, 18, 22, 21, 20, 26, 32, 37, 47, 53, 43, 26, 21, 21, 21, 21, 
    37, 41, 46, 50, 38, 17, 0, 10, 2, 0, 0, 0, 0, 0, 5, 7, 0, 0, 0, 4, 36, 51, 44, 36, 41, 44, 37, 28, 22, 21, 
    32, 45, 51, 59, 58, 52, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 29, 39, 47, 56, 71, 76, 63, 45, 29, 21, 
    24, 43, 58, 57, 42, 27, 13, 0, 0, 9, 34, 50, 48, 44, 37, 36, 45, 57, 67, 72, 64, 58, 61, 68, 71, 71, 68, 58, 42, 23, 
    29, 53, 73, 73, 45, 13, 8, 9, 15, 32, 44, 51, 47, 46, 51, 64, 78, 83, 79, 76, 73, 74, 84, 83, 72, 49, 35, 42, 45, 29, 
    31, 40, 38, 46, 45, 53, 54, 48, 17, 6, 0, 0, 0, 0, 15, 42, 55, 53, 34, 20, 23, 44, 68, 59, 29, 0, 0, 6, 27, 33, 
    3, 12, 15, 23, 38, 73, 92, 66, 22, 17, 17, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 28, 39, 
    13, 30, 40, 46, 53, 63, 77, 54, 32, 47, 70, 82, 74, 45, 14, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 35, 56, 53, 45, 
    16, 23, 37, 62, 75, 65, 53, 50, 51, 60, 56, 58, 70, 72, 51, 33, 39, 51, 53, 51, 57, 59, 57, 54, 44, 45, 54, 49, 35, 34, 
    17, 19, 26, 58, 76, 69, 49, 56, 68, 67, 48, 34, 25, 33, 55, 67, 51, 27, 27, 35, 41, 35, 31, 38, 48, 46, 22, 10, 14, 31, 
    17, 23, 18, 29, 46, 48, 47, 53, 69, 79, 67, 40, 5, 7, 37, 67, 68, 52, 42, 46, 47, 34, 24, 37, 50, 44, 8, 0, 15, 35, 
    7, 25, 41, 43, 39, 27, 27, 31, 48, 69, 73, 59, 37, 27, 40, 58, 39, 8, 0, 0, 0, 0, 0, 0, 19, 49, 41, 34, 39, 36, 
    4, 23, 52, 78, 64, 23, 0, 5, 37, 61, 77, 90, 107, 106, 92, 74, 64, 57, 44, 23, 12, 18, 38, 54, 69, 77, 91, 86, 51, 23, 
    2, 7, 24, 43, 49, 25, 3, 8, 38, 54, 70, 82, 93, 99, 92, 80, 85, 86, 62, 17, 4, 7, 40, 70, 82, 71, 67, 54, 25, 11, 
    4, 0, 0, 0, 0, 7, 26, 26, 31, 40, 57, 72, 78, 76, 74, 74, 68, 38, 0, 0, 0, 0, 0, 21, 64, 76, 58, 31, 8, 4, 
    0, 0, 0, 0, 0, 14, 31, 25, 27, 31, 50, 72, 80, 77, 69, 57, 47, 45, 53, 60, 52, 41, 44, 59, 77, 75, 55, 29, 9, 1, 
    0, 0, 7, 10, 15, 26, 37, 33, 34, 39, 53, 65, 68, 65, 60, 50, 40, 48, 71, 84, 67, 43, 48, 61, 74, 67, 52, 35, 17, 3, 
    0, 6, 10, 8, 8, 29, 49, 53, 43, 45, 54, 60, 62, 61, 61, 65, 68, 67, 60, 50, 40, 30, 34, 53, 66, 68, 59, 41, 19, 0, 
    2, 2, 0, 0, 5, 25, 48, 59, 49, 50, 56, 59, 56, 55, 53, 53, 53, 53, 51, 50, 51, 53, 49, 56, 60, 67, 58, 34, 8, 0, 
    0, 0, 0, 0, 0, 18, 42, 59, 58, 57, 57, 51, 43, 38, 36, 36, 35, 31, 27, 27, 32, 36, 38, 39, 43, 46, 33, 10, 0, 0, 
    
    -- channel=154
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 16, 20, 20, 16, 28, 29, 19, 13, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 18, 56, 61, 67, 74, 63, 76, 86, 87, 91, 77, 58, 32, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 79, 87, 71, 69, 63, 58, 60, 66, 79, 89, 91, 75, 44, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 30, 54, 22, 7, 9, 9, 4, 1, 7, 23, 34, 31, 24, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 21, 0, 0, 0, 0, 13, 19, 10, 8, 8, 3, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 43, 47, 32, 21, 18, 18, 47, 59, 45, 35, 29, 24, 17, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 41, 58, 58, 59, 67, 67, 57, 58, 58, 51, 41, 40, 36, 37, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 61, 67, 64, 61, 54, 61, 70, 76, 68, 61, 60, 53, 56, 53, 47, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 33, 46, 78, 98, 93, 75, 73, 81, 79, 74, 75, 79, 83, 84, 75, 68, 44, 27, 28, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 18, 64, 97, 97, 71, 54, 54, 71, 84, 84, 85, 80, 69, 65, 80, 76, 45, 16, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 22, 32, 34, 28, 25, 36, 46, 49, 30, 39, 64, 65, 52, 33, 14, 11, 38, 56, 42, 20, 8, 4, 0, 0, 0, 0, 
    0, 0, 4, 16, 20, 32, 32, 27, 17, 31, 49, 75, 73, 56, 61, 66, 67, 68, 67, 60, 58, 63, 65, 63, 62, 60, 51, 23, 0, 0, 
    0, 0, 25, 43, 16, 0, 0, 27, 70, 80, 96, 118, 129, 113, 94, 93, 102, 113, 124, 121, 106, 92, 88, 93, 97, 92, 79, 56, 11, 0, 
    0, 5, 32, 51, 25, 0, 0, 38, 81, 65, 52, 50, 57, 68, 68, 89, 115, 120, 119, 105, 91, 105, 119, 125, 123, 93, 66, 42, 13, 0, 
    0, 0, 0, 6, 5, 18, 63, 94, 59, 30, 4, 0, 0, 0, 0, 17, 26, 13, 3, 0, 0, 0, 25, 29, 37, 23, 4, 2, 0, 0, 
    0, 0, 0, 5, 2, 22, 79, 117, 55, 27, 48, 58, 38, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 33, 26, 4, 
    0, 0, 11, 34, 33, 28, 52, 83, 78, 60, 77, 101, 111, 94, 53, 10, 0, 22, 42, 38, 39, 37, 23, 17, 11, 15, 64, 91, 58, 11, 
    0, 0, 3, 48, 69, 57, 43, 55, 88, 89, 66, 64, 81, 87, 89, 79, 60, 61, 71, 77, 77, 79, 77, 70, 71, 64, 66, 72, 46, 2, 
    0, 0, 0, 26, 54, 66, 49, 49, 80, 96, 80, 57, 42, 40, 60, 102, 108, 75, 70, 83, 88, 80, 69, 65, 83, 88, 41, 15, 20, 5, 
    0, 0, 0, 19, 14, 34, 50, 40, 54, 76, 86, 70, 26, 0, 12, 71, 85, 40, 22, 40, 41, 28, 11, 0, 28, 77, 37, 3, 19, 16, 
    0, 0, 18, 54, 44, 12, 21, 13, 24, 53, 71, 87, 81, 65, 45, 58, 55, 12, 0, 0, 0, 0, 0, 0, 4, 72, 86, 76, 62, 22, 
    0, 4, 25, 66, 82, 41, 0, 0, 15, 46, 64, 84, 113, 123, 106, 76, 77, 90, 67, 41, 24, 17, 38, 66, 77, 75, 93, 103, 75, 24, 
    16, 6, 0, 1, 21, 35, 18, 8, 26, 34, 51, 66, 79, 87, 90, 78, 84, 82, 28, 0, 0, 0, 0, 23, 77, 72, 68, 64, 47, 26, 
    19, 0, 0, 0, 0, 7, 33, 30, 33, 20, 31, 56, 69, 69, 68, 65, 60, 47, 4, 0, 0, 0, 0, 0, 51, 77, 69, 50, 35, 26, 
    10, 0, 0, 0, 0, 14, 30, 31, 41, 27, 27, 48, 62, 62, 58, 47, 30, 33, 61, 76, 69, 50, 33, 43, 63, 68, 68, 54, 43, 32, 
    1, 9, 22, 28, 21, 22, 42, 47, 52, 43, 37, 41, 49, 50, 49, 51, 52, 57, 76, 93, 80, 56, 33, 38, 62, 60, 63, 62, 53, 34, 
    16, 25, 25, 21, 19, 26, 52, 69, 57, 51, 45, 41, 45, 49, 51, 57, 66, 73, 74, 74, 70, 64, 49, 31, 48, 65, 66, 65, 55, 28, 
    32, 34, 25, 16, 10, 21, 49, 73, 57, 53, 52, 46, 41, 44, 44, 45, 49, 53, 55, 60, 66, 71, 64, 44, 37, 59, 62, 52, 35, 11, 
    21, 12, 5, 4, 5, 7, 29, 66, 67, 60, 47, 39, 33, 30, 30, 32, 31, 26, 21, 23, 29, 35, 38, 32, 20, 26, 31, 19, 0, 0, 
    
    -- channel=155
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=156
    247, 239, 245, 248, 241, 210, 203, 210, 202, 191, 193, 203, 199, 207, 221, 241, 266, 276, 276, 265, 266, 268, 269, 243, 219, 223, 238, 218, 198, 202, 
    264, 262, 260, 266, 249, 203, 185, 212, 224, 218, 233, 240, 257, 280, 285, 295, 297, 292, 297, 283, 267, 268, 279, 268, 258, 250, 251, 231, 229, 230, 
    282, 282, 282, 286, 271, 213, 178, 200, 208, 213, 224, 217, 237, 261, 267, 292, 295, 292, 295, 283, 262, 265, 277, 275, 274, 263, 247, 249, 259, 247, 
    294, 294, 294, 292, 268, 192, 147, 164, 165, 176, 178, 161, 170, 175, 183, 215, 228, 245, 266, 270, 262, 265, 265, 263, 270, 255, 236, 254, 276, 264, 
    294, 294, 296, 291, 259, 168, 98, 110, 133, 138, 136, 125, 131, 127, 121, 130, 137, 151, 187, 235, 271, 279, 262, 254, 255, 237, 221, 233, 268, 281, 
    294, 293, 295, 280, 262, 192, 103, 111, 153, 158, 150, 145, 154, 167, 161, 150, 143, 137, 142, 192, 261, 301, 286, 264, 237, 218, 197, 198, 235, 280, 
    293, 295, 287, 255, 251, 211, 121, 151, 213, 234, 235, 217, 190, 201, 209, 201, 193, 185, 184, 192, 215, 270, 298, 268, 236, 224, 202, 188, 203, 258, 
    293, 296, 280, 247, 250, 204, 126, 164, 215, 228, 260, 247, 198, 196, 202, 208, 206, 200, 215, 213, 193, 229, 266, 255, 251, 242, 214, 179, 176, 217, 
    294, 294, 279, 249, 234, 191, 134, 166, 189, 180, 214, 215, 192, 190, 194, 203, 211, 201, 214, 226, 202, 225, 264, 277, 276, 263, 218, 183, 185, 207, 
    294, 294, 276, 212, 177, 153, 118, 168, 186, 177, 183, 182, 181, 181, 187, 197, 204, 197, 214, 230, 219, 233, 270, 299, 306, 293, 262, 251, 251, 258, 
    291, 296, 272, 199, 172, 125, 89, 124, 151, 164, 153, 150, 159, 163, 169, 171, 169, 168, 185, 206, 214, 212, 226, 267, 303, 299, 293, 294, 294, 294, 
    276, 287, 253, 215, 207, 149, 74, 63, 101, 139, 145, 140, 132, 134, 139, 135, 133, 143, 153, 157, 171, 182, 208, 264, 304, 307, 303, 299, 295, 294, 
    249, 251, 212, 191, 188, 148, 97, 84, 107, 139, 159, 166, 145, 123, 122, 133, 152, 175, 174, 147, 143, 164, 205, 254, 287, 304, 316, 319, 307, 294, 
    227, 206, 181, 165, 155, 128, 128, 118, 149, 162, 161, 172, 160, 138, 130, 141, 158, 175, 171, 147, 136, 141, 164, 197, 219, 234, 271, 317, 324, 298, 
    216, 164, 138, 154, 173, 169, 135, 109, 137, 117, 95, 98, 100, 109, 111, 113, 117, 116, 104, 100, 106, 113, 131, 141, 155, 167, 199, 273, 317, 305, 
    186, 123, 81, 129, 190, 203, 134, 112, 113, 97, 73, 58, 53, 67, 48, 36, 43, 37, 36, 46, 32, 31, 51, 61, 103, 128, 147, 232, 295, 308, 
    183, 121, 84, 132, 178, 144, 99, 117, 127, 139, 154, 140, 127, 107, 49, 42, 40, 29, 65, 86, 40, 21, 24, 46, 101, 133, 159, 219, 286, 317, 
    204, 136, 107, 156, 170, 70, 54, 115, 138, 133, 151, 163, 185, 151, 133, 156, 147, 150, 188, 199, 171, 161, 150, 161, 181, 167, 172, 201, 275, 318, 
    208, 130, 90, 149, 156, 59, 45, 97, 116, 101, 88, 95, 121, 135, 190, 199, 167, 169, 192, 194, 185, 183, 178, 209, 205, 145, 126, 157, 246, 308, 
    218, 135, 63, 102, 118, 76, 57, 66, 86, 94, 75, 60, 65, 92, 148, 170, 153, 137, 142, 143, 141, 135, 138, 168, 157, 111, 92, 124, 226, 304, 
    226, 152, 71, 66, 80, 69, 58, 41, 54, 75, 80, 82, 79, 74, 76, 109, 130, 119, 98, 99, 102, 106, 116, 105, 97, 118, 121, 119, 209, 303, 
    229, 158, 99, 95, 86, 58, 55, 36, 28, 40, 77, 113, 142, 111, 47, 70, 125, 119, 77, 84, 86, 113, 146, 83, 58, 143, 168, 131, 206, 300, 
    227, 146, 82, 112, 110, 89, 81, 45, 26, 30, 58, 91, 147, 121, 59, 79, 161, 171, 145, 147, 134, 166, 206, 112, 75, 122, 132, 117, 206, 293, 
    220, 127, 41, 60, 102, 140, 128, 63, 39, 29, 30, 39, 64, 60, 49, 66, 110, 133, 144, 137, 129, 141, 137, 74, 67, 71, 64, 83, 192, 282, 
    207, 136, 61, 46, 92, 151, 142, 82, 55, 31, 21, 22, 26, 29, 35, 34, 55, 131, 184, 180, 167, 163, 108, 39, 41, 53, 58, 88, 185, 267, 
    210, 191, 150, 116, 112, 152, 135, 89, 79, 49, 20, 17, 21, 24, 30, 23, 53, 167, 246, 259, 241, 232, 146, 51, 31, 44, 74, 106, 184, 259, 
    213, 217, 199, 161, 130, 155, 133, 101, 100, 67, 29, 15, 18, 24, 37, 53, 78, 139, 182, 201, 209, 202, 124, 39, 25, 43, 82, 111, 185, 255, 
    209, 202, 188, 167, 135, 145, 119, 109, 101, 74, 41, 26, 28, 35, 46, 66, 85, 108, 122, 143, 169, 177, 100, 28, 23, 48, 82, 108, 186, 251, 
    202, 193, 180, 167, 137, 119, 96, 103, 94, 75, 50, 36, 35, 41, 46, 52, 63, 78, 94, 118, 143, 161, 101, 37, 19, 47, 72, 101, 191, 244, 
    190, 186, 179, 172, 138, 91, 75, 96, 89, 71, 57, 46, 42, 46, 50, 51, 58, 67, 74, 86, 103, 119, 93, 41, 20, 40, 64, 116, 201, 233, 
    
    -- channel=157
    236, 230, 228, 233, 243, 232, 187, 162, 176, 186, 187, 191, 194, 198, 216, 231, 246, 255, 252, 243, 237, 230, 234, 231, 220, 200, 193, 177, 163, 160, 
    264, 263, 262, 267, 267, 254, 202, 168, 185, 191, 204, 214, 213, 228, 244, 247, 255, 251, 239, 229, 218, 216, 228, 242, 245, 232, 208, 180, 177, 198, 
    291, 288, 288, 289, 291, 275, 214, 171, 179, 185, 190, 198, 190, 197, 207, 213, 230, 228, 203, 193, 188, 199, 227, 245, 242, 228, 197, 170, 177, 207, 
    297, 296, 296, 297, 286, 249, 185, 133, 141, 161, 165, 167, 160, 155, 161, 165, 172, 176, 162, 147, 159, 196, 232, 246, 235, 214, 184, 155, 159, 193, 
    298, 296, 298, 302, 285, 238, 182, 122, 127, 166, 180, 189, 188, 187, 185, 178, 169, 161, 153, 150, 158, 204, 242, 254, 238, 205, 165, 136, 133, 174, 
    297, 295, 300, 298, 272, 249, 215, 152, 149, 207, 227, 242, 252, 251, 250, 237, 227, 219, 195, 191, 196, 202, 232, 256, 232, 193, 153, 132, 129, 157, 
    295, 296, 296, 282, 255, 256, 225, 175, 196, 264, 274, 279, 275, 255, 250, 250, 246, 248, 244, 232, 215, 190, 200, 232, 224, 211, 200, 165, 135, 139, 
    295, 296, 294, 284, 269, 257, 212, 163, 182, 231, 243, 256, 256, 238, 237, 242, 244, 247, 247, 247, 235, 206, 188, 218, 240, 241, 224, 173, 132, 138, 
    292, 293, 295, 295, 257, 224, 187, 165, 182, 217, 223, 231, 231, 226, 230, 234, 242, 244, 242, 250, 251, 238, 229, 246, 268, 273, 253, 220, 205, 212, 
    280, 291, 294, 264, 211, 191, 175, 156, 156, 182, 193, 197, 198, 203, 211, 218, 222, 219, 221, 240, 247, 248, 243, 235, 259, 285, 293, 287, 285, 286, 
    263, 287, 295, 259, 213, 203, 171, 117, 92, 124, 160, 177, 186, 182, 179, 179, 172, 165, 175, 196, 199, 191, 184, 192, 241, 284, 298, 297, 297, 298, 
    249, 272, 268, 236, 205, 198, 148, 95, 89, 130, 173, 188, 196, 178, 149, 140, 143, 157, 174, 175, 147, 130, 150, 186, 239, 272, 280, 288, 296, 297, 
    236, 247, 225, 187, 163, 147, 133, 142, 163, 185, 200, 206, 208, 189, 157, 155, 176, 203, 209, 183, 137, 115, 132, 160, 196, 227, 243, 257, 286, 297, 
    236, 237, 195, 142, 121, 123, 156, 175, 180, 190, 167, 151, 140, 134, 123, 122, 130, 140, 135, 117, 94, 88, 104, 125, 150, 171, 195, 216, 261, 295, 
    227, 198, 135, 89, 110, 163, 191, 170, 131, 120, 80, 64, 62, 68, 75, 65, 49, 45, 33, 32, 48, 46, 50, 56, 76, 117, 158, 185, 237, 288, 
    201, 169, 110, 71, 114, 179, 164, 114, 97, 107, 95, 104, 102, 91, 68, 15, 0, 0, 0, 0, 26, 0, 0, 0, 37, 107, 158, 188, 229, 275, 
    231, 200, 141, 89, 122, 138, 88, 45, 90, 134, 140, 147, 150, 142, 103, 65, 74, 84, 106, 129, 132, 96, 65, 80, 121, 176, 202, 201, 214, 254, 
    239, 203, 142, 94, 114, 96, 35, 22, 81, 113, 94, 89, 113, 115, 122, 159, 203, 193, 189, 206, 213, 195, 184, 181, 197, 213, 174, 143, 165, 229, 
    239, 205, 139, 82, 79, 66, 27, 25, 47, 63, 56, 43, 44, 65, 110, 148, 171, 150, 148, 159, 160, 147, 139, 161, 176, 164, 114, 94, 134, 216, 
    241, 211, 133, 59, 42, 41, 30, 18, 14, 24, 37, 36, 42, 55, 84, 104, 127, 140, 139, 133, 128, 116, 120, 142, 135, 107, 95, 107, 136, 206, 
    242, 225, 149, 56, 45, 41, 26, 10, 0, 0, 0, 23, 57, 80, 81, 36, 32, 77, 89, 71, 68, 70, 74, 112, 92, 60, 110, 147, 143, 193, 
    254, 228, 158, 63, 46, 53, 38, 31, 1, 0, 0, 25, 82, 102, 72, 10, 22, 95, 119, 98, 104, 120, 142, 157, 101, 63, 113, 129, 115, 180, 
    263, 224, 131, 44, 27, 61, 91, 83, 30, 0, 0, 0, 15, 28, 10, 0, 40, 93, 121, 124, 132, 155, 175, 143, 65, 21, 37, 48, 76, 182, 
    259, 208, 116, 26, 27, 85, 137, 119, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 112, 141, 147, 142, 100, 21, 0, 0, 13, 76, 191, 
    241, 212, 166, 120, 101, 116, 140, 123, 58, 16, 0, 0, 0, 0, 0, 0, 0, 11, 119, 218, 230, 223, 190, 112, 8, 0, 0, 26, 99, 198, 
    229, 241, 237, 208, 164, 134, 135, 120, 75, 48, 1, 0, 0, 0, 0, 0, 0, 46, 139, 206, 211, 212, 186, 93, 0, 0, 0, 45, 116, 202, 
    239, 247, 235, 205, 169, 146, 129, 110, 79, 58, 13, 0, 0, 0, 0, 0, 13, 50, 88, 121, 146, 169, 156, 72, 0, 0, 0, 47, 113, 199, 
    245, 237, 220, 198, 168, 145, 108, 81, 69, 54, 17, 0, 0, 0, 0, 0, 4, 28, 56, 87, 123, 155, 133, 64, 0, 0, 0, 37, 105, 203, 
    233, 225, 214, 201, 180, 144, 86, 50, 54, 45, 14, 0, 0, 0, 0, 0, 0, 14, 36, 60, 85, 111, 98, 52, 0, 0, 0, 27, 112, 220, 
    221, 219, 221, 218, 197, 150, 81, 33, 36, 24, 8, 0, 0, 1, 10, 12, 13, 23, 42, 56, 69, 82, 79, 44, 0, 0, 0, 54, 155, 246, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    117, 124, 122, 123, 113, 107, 95, 91, 96, 104, 108, 105, 118, 128, 132, 128, 111, 105, 102, 110, 107, 104, 106, 120, 134, 136, 134, 125, 128, 136, 
    112, 114, 117, 117, 115, 101, 78, 52, 37, 36, 27, 24, 21, 19, 20, 31, 40, 58, 70, 86, 91, 97, 101, 110, 116, 123, 117, 126, 128, 130, 
    98, 98, 100, 96, 93, 67, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 51, 79, 93, 101, 104, 101, 106, 111, 123, 124, 123, 
    84, 85, 85, 84, 78, 58, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 70, 105, 109, 110, 106, 105, 110, 107, 107, 114, 
    83, 83, 82, 75, 80, 79, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 93, 117, 114, 108, 106, 101, 100, 97, 106, 
    83, 84, 78, 65, 66, 67, 40, 7, 0, 18, 37, 22, 0, 0, 0, 0, 0, 0, 0, 0, 19, 41, 82, 102, 111, 124, 134, 128, 109, 96, 
    84, 85, 78, 74, 72, 42, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 52, 83, 113, 133, 147, 131, 110, 95, 
    85, 84, 82, 77, 55, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 65, 102, 120, 129, 129, 134, 137, 131, 
    83, 84, 83, 51, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 79, 97, 113, 135, 165, 181, 171, 
    76, 83, 80, 55, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 49, 84, 116, 130, 137, 130, 
    70, 72, 68, 77, 67, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 54, 78, 84, 84, 85, 84, 
    70, 56, 50, 53, 44, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 34, 46, 58, 73, 83, 85, 
    83, 62, 59, 55, 51, 35, 35, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 65, 84, 
    106, 80, 54, 54, 81, 105, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 78, 
    98, 70, 41, 51, 92, 117, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 68, 
    118, 100, 86, 83, 86, 53, 8, 0, 0, 10, 58, 67, 62, 40, 25, 21, 26, 34, 53, 62, 54, 41, 17, 17, 6, 0, 2, 8, 34, 60, 
    130, 105, 89, 86, 78, 31, 0, 0, 0, 1, 3, 0, 10, 19, 62, 106, 142, 147, 139, 132, 134, 146, 152, 139, 100, 49, 8, 0, 9, 41, 
    98, 73, 49, 51, 51, 47, 16, 0, 0, 0, 0, 0, 0, 0, 17, 47, 48, 27, 0, 0, 4, 14, 30, 34, 18, 0, 0, 0, 0, 32, 
    96, 80, 45, 18, 18, 41, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 
    91, 81, 59, 24, 21, 26, 23, 2, 0, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 13, 37, 
    79, 69, 65, 53, 53, 39, 22, 22, 7, 0, 0, 4, 30, 34, 2, 0, 0, 0, 0, 0, 0, 8, 27, 17, 0, 0, 14, 17, 14, 30, 
    60, 43, 30, 37, 41, 57, 46, 46, 39, 23, 6, 0, 0, 0, 5, 13, 36, 57, 72, 64, 58, 66, 79, 60, 36, 0, 0, 0, 0, 24, 
    28, 23, 7, 4, 19, 47, 63, 54, 43, 34, 5, 0, 0, 0, 0, 0, 0, 0, 5, 21, 29, 20, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 19, 43, 41, 46, 38, 27, 34, 31, 36, 27, 14, 0, 0, 0, 0, 0, 0, 35, 77, 83, 59, 22, 15, 0, 0, 6, 7, 3, 1, 
    0, 42, 82, 101, 70, 33, 6, 14, 24, 41, 41, 32, 26, 23, 22, 18, 24, 52, 78, 100, 92, 82, 61, 42, 17, 10, 21, 19, 2, 0, 
    8, 31, 45, 43, 31, 21, 12, 14, 16, 31, 40, 37, 32, 31, 34, 47, 49, 18, 0, 0, 0, 0, 0, 10, 17, 24, 19, 5, 0, 0, 
    8, 0, 0, 0, 3, 8, 2, 1, 0, 12, 32, 45, 47, 44, 42, 44, 32, 0, 0, 0, 0, 0, 0, 15, 27, 33, 14, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 6, 26, 43, 46, 41, 32, 17, 4, 0, 0, 0, 0, 0, 0, 23, 36, 27, 8, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 6, 23, 36, 42, 38, 33, 28, 20, 11, 1, 0, 0, 0, 0, 18, 40, 30, 15, 11, 0, 0, 
    0, 0, 0, 0, 6, 7, 6, 0, 0, 6, 27, 41, 46, 43, 39, 35, 36, 38, 34, 24, 13, 3, 13, 30, 50, 48, 44, 42, 18, 0, 
    
    
    others => 0);
end gold_package;
