-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(36-1 downto 0);
        ADDR : in std_logic_vector(9-1 downto 0);
        DO   : out std_logic_vector(36-1 downto 0)
    );
    attribute dont_touch : string;
    attribute dont_touch of bram_single : entity is "true";
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(8-1 downto 0);
    signal bram_addr     : std_logic_vector(9-1 downto 0);
    signal bram_di     : std_logic_vector(44-1 downto 0);
    signal bram_do     : std_logic_vector(44-1 downto 0);
    constant bram_par     : std_logic_vector(8-1 downto 0) := "00000000";

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(9-1 downto 0);
    bram_di <= bram_par & DI;
    DO <= bram_do(36-1 downto 0);


    MEM_IWGHT_LAYER0_INSTANCE0 : if BRAM_NAME = "iwght_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000089400000000fffffa57ffffffff000004fe00000000fffff05bffffffff",
            INIT_01 => X"00001869000000000000112a00000000000008a4000000000000001d00000000",
            INIT_02 => X"000013d200000000fffffebaffffffffffffdeecfffffffffffffcf0ffffffff",
            INIT_03 => X"00001da300000000ffffcfa0ffffffff00000a4b000000000000188d00000000",
            INIT_04 => X"fffffff7ffffffff0000000a0000000000000022000000000000001f00000000",
            INIT_05 => X"00000004000000000000000000000000ffffffe5ffffffffffffffcaffffffff",
            INIT_06 => X"ffffffd3ffffffff0000002e000000000000002c000000000000000300000000",
            INIT_07 => X"0000001800000000ffffffddffffffffffffffffffffffff0000003800000000",
            INIT_08 => X"0000001800000000000000200000000000000021000000000000003500000000",
            INIT_09 => X"ffffffedffffffffffffffc3ffffffffffffffccffffffffffffffc9ffffffff",
            INIT_0A => X"ffffffe6ffffffff0000000b00000000ffffffdaffffffffffffffc6ffffffff",
            INIT_0B => X"ffffffc0ffffffffffffffd3ffffffff0000001f000000000000001b00000000",
            INIT_0C => X"fffffff5ffffffff0000001000000000ffffffe2ffffffffffffffc6ffffffff",
            INIT_0D => X"0000000f00000000000000250000000000000018000000000000001700000000",
            INIT_0E => X"ffffffd3fffffffffffffff6ffffffffffffffd8ffffffffffffffd8ffffffff",
            INIT_0F => X"fffffff3ffffffff000000320000000000000007000000000000000700000000",
            INIT_10 => X"ffffffd8ffffffff00000033000000000000001d000000000000002600000000",
            INIT_11 => X"0000001300000000ffffffcfffffffff0000000c000000000000000600000000",
            INIT_12 => X"000000240000000000000005000000000000002000000000fffffff3ffffffff",
            INIT_13 => X"ffffffebffffffff0000000b00000000fffffffbffffffffffffffffffffffff",
            INIT_14 => X"ffffffdcffffffffffffffc1fffffffffffffffaffffffffffffffdfffffffff",
            INIT_15 => X"ffffffdbffffffff0000000e00000000ffffffecfffffffffffffff4ffffffff",
            INIT_16 => X"ffffffe1ffffffff000000270000000000000009000000000000003200000000",
            INIT_17 => X"00000018000000000000002d0000000000000037000000000000000600000000",
            INIT_18 => X"ffffffe6ffffffff000000020000000000000012000000000000002400000000",
            INIT_19 => X"0000001600000000ffffffeeffffffff0000002d000000000000002100000000",
            INIT_1A => X"fffffffbfffffffffffffff8ffffffffffffffc6ffffffffffffffe7ffffffff",
            INIT_1B => X"ffffffd2fffffffffffffffcffffffff0000003700000000ffffffc2ffffffff",
            INIT_1C => X"0000004000000000ffffffc2ffffffff0000001e00000000ffffffe6ffffffff",
            INIT_1D => X"0000001000000000000000340000000000000000000000000000001f00000000",
            INIT_1E => X"ffffffccffffffff0000001e000000000000005200000000fffffff5ffffffff",
            INIT_1F => X"fffffff6ffffffffffffffe6ffffffffffffffc6ffffffffffffffe5ffffffff",
            INIT_20 => X"0000002b000000000000004d00000000ffffffebffffffff0000002b00000000",
            INIT_21 => X"fffffffcffffffffffffffafffffffffffffffbefffffffffffffffaffffffff",
            INIT_22 => X"00000022000000000000002b00000000fffffffdffffffffffffffcdffffffff",
            INIT_23 => X"ffffffc2ffffffffffffffe1ffffffff00000039000000000000004400000000",
            INIT_24 => X"0000000b0000000000000039000000000000000100000000ffffffe1ffffffff",
            INIT_25 => X"0000002c00000000fffffff9fffffffffffffffaffffffff0000003300000000",
            INIT_26 => X"0000002f000000000000001f0000000000000026000000000000002800000000",
            INIT_27 => X"fffffffaffffffff0000002f0000000000000045000000000000003b00000000",
            INIT_28 => X"ffffffe6fffffffffffffff0ffffffffffffffefffffffff0000001b00000000",
            INIT_29 => X"fffffff8ffffffff0000002100000000ffffffe4ffffffff0000001800000000",
            INIT_2A => X"0000000400000000ffffffd2ffffffffffffffd6ffffffffffffffd5ffffffff",
            INIT_2B => X"fffffff4ffffffffffffffc6ffffffffffffffcaffffffffffffffe5ffffffff",
            INIT_2C => X"00000000000000000000001900000000ffffffd6ffffffffffffffe9ffffffff",
            INIT_2D => X"0000003300000000000000300000000000000004000000000000001c00000000",
            INIT_2E => X"ffffffbeffffffff00000044000000000000000d00000000ffffffd6ffffffff",
            INIT_2F => X"ffffffc1ffffffffffffffb3ffffffff0000000500000000fffffffcffffffff",
            INIT_30 => X"fffffff5ffffffffffffffd0fffffffffffffff0ffffffff0000002200000000",
            INIT_31 => X"ffffffbcffffffff0000001c00000000ffffffe4ffffffff0000000900000000",
            INIT_32 => X"00000000000000000000000f0000000000000025000000000000001000000000",
            INIT_33 => X"0000001100000000000000400000000000000026000000000000000e00000000",
            INIT_34 => X"0000001f00000000ffffffeaffffffff0000002d000000000000003300000000",
            INIT_35 => X"ffffffcdfffffffffffffff0ffffffff00000000000000000000003400000000",
            INIT_36 => X"ffffffc9ffffffff0000000900000000fffffff5fffffffffffffff6ffffffff",
            INIT_37 => X"0000002100000000ffffffd3ffffffffffffffbbffffffffffffffc4ffffffff",
            INIT_38 => X"ffffffbaffffffffffffffc7ffffffff0000000a000000000000001c00000000",
            INIT_39 => X"0000002800000000ffffffc6fffffffffffffff2ffffffff0000000000000000",
            INIT_3A => X"0000003400000000ffffffffffffffff0000002d000000000000001500000000",
            INIT_3B => X"ffffffcbfffffffffffffff7ffffffff00000033000000000000003c00000000",
            INIT_3C => X"ffffffdeffffffff00000003000000000000002f00000000ffffffc7ffffffff",
            INIT_3D => X"ffffffd1ffffffff0000001700000000fffffff7fffffffffffffff8ffffffff",
            INIT_3E => X"0000000a00000000fffffff8ffffffffffffffc5ffffffffffffffc9ffffffff",
            INIT_3F => X"0000001c0000000000000039000000000000000b00000000fffffffcffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000300000000fffffff9ffffffffffffffd5fffffffffffffff7ffffffff",
            INIT_41 => X"fffffff8fffffffffffffffafffffffffffffffbffffffff0000000200000000",
            INIT_42 => X"fffffff0ffffffffffffffc5ffffffffffffffc1ffffffff0000001600000000",
            INIT_43 => X"0000001d00000000ffffffdfffffffff0000001e000000000000002b00000000",
            INIT_44 => X"0000002d00000000000000310000000000000017000000000000001b00000000",
            INIT_45 => X"00000028000000000000003b000000000000002000000000fffffff3ffffffff",
            INIT_46 => X"fffffff7ffffffff00000006000000000000002900000000ffffffe9ffffffff",
            INIT_47 => X"0000003d00000000000000140000000000000027000000000000002c00000000",
            INIT_48 => X"ffffffd2fffffffffffffff5ffffffff00000025000000000000002500000000",
            INIT_49 => X"0000001d00000000ffffffc8ffffffffffffffd8fffffffffffffff1ffffffff",
            INIT_4A => X"ffffffe4ffffffff0000001e0000000000000031000000000000001000000000",
            INIT_4B => X"ffffffaeffffffffffffffbfffffffff00000021000000000000001200000000",
            INIT_4C => X"fffffff3ffffffff00000045000000000000001d00000000ffffffe6ffffffff",
            INIT_4D => X"00000010000000000000003500000000ffffffdaffffffffffffffdcffffffff",
            INIT_4E => X"0000001c00000000ffffffddffffffffffffffedffffffffffffffcbffffffff",
            INIT_4F => X"ffffffd5ffffffffffffffe6fffffffffffffff7ffffffffffffffd0ffffffff",
            INIT_50 => X"fffffffdffffffffffffffd9ffffffffffffffe0ffffffffffffffecffffffff",
            INIT_51 => X"fffffff9ffffffffffffffe2ffffffffffffffe3ffffffff0000002600000000",
            INIT_52 => X"0000002f000000000000001f0000000000000001000000000000001500000000",
            INIT_53 => X"0000002c00000000ffffffeaffffffff00000033000000000000001600000000",
            INIT_54 => X"0000003300000000fffffffbffffffffffffffe5ffffffff0000003300000000",
            INIT_55 => X"ffffffe0ffffffff0000003e00000000ffffffdbffffffffffffffc5ffffffff",
            INIT_56 => X"0000002800000000ffffffd7ffffffff0000001b00000000fffffff9ffffffff",
            INIT_57 => X"00000026000000000000000500000000ffffffd7fffffffffffffff8ffffffff",
            INIT_58 => X"fffffff3ffffffff0000004b000000000000000a000000000000000300000000",
            INIT_59 => X"fffffffeffffffffffffffd8ffffffff00000030000000000000003a00000000",
            INIT_5A => X"ffffffffffffffff0000002900000000ffffffc7fffffffffffffff9ffffffff",
            INIT_5B => X"ffffffddfffffffffffffffaffffffffffffffebffffffffffffffd7ffffffff",
            INIT_5C => X"ffffffe4ffffffffffffffdfffffffffffffffd9ffffffffffffffc9ffffffff",
            INIT_5D => X"fffffffeffffffff0000004d00000000fffffff9ffffffff0000003400000000",
            INIT_5E => X"ffffffecffffffffffffffbfffffffffffffffffffffffffffffffd6ffffffff",
            INIT_5F => X"00000003000000000000003d0000000000000013000000000000001900000000",
            INIT_60 => X"ffffffbcfffffffffffffff2ffffffffffffffdbffffffff0000001b00000000",
            INIT_61 => X"0000003600000000ffffffffffffffff0000000700000000ffffffe9ffffffff",
            INIT_62 => X"0000003800000000fffffffbffffffff0000003e00000000ffffffe8ffffffff",
            INIT_63 => X"0000000a00000000000000120000000000000024000000000000000f00000000",
            INIT_64 => X"ffffffe4ffffffff0000000a000000000000002d000000000000002300000000",
            INIT_65 => X"00000029000000000000001500000000fffffffaffffffff0000001000000000",
            INIT_66 => X"ffffffd1fffffffffffffffdfffffffffffffff7ffffffffffffffd1ffffffff",
            INIT_67 => X"00000019000000000000000900000000ffffffe0ffffffffffffffdfffffffff",
            INIT_68 => X"0000001a00000000fffffff7ffffffff0000001000000000ffffffdaffffffff",
            INIT_69 => X"ffffffddffffffff0000000d00000000fffffff5ffffffffffffffebffffffff",
            INIT_6A => X"0000001300000000ffffffefffffffffffffffe1ffffffff0000001800000000",
            INIT_6B => X"00000031000000000000000200000000ffffffd2ffffffffffffffe4ffffffff",
            INIT_6C => X"fffffff0ffffffff000000260000000000000046000000000000001400000000",
            INIT_6D => X"ffffffdbfffffffffffffff5ffffffff0000002b000000000000004200000000",
            INIT_6E => X"ffffffe4fffffffffffffff7fffffffffffffff8ffffffffffffffcfffffffff",
            INIT_6F => X"ffffffccfffffffffffffff2ffffffff0000002300000000ffffffdaffffffff",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE0 : if BRAM_NAME = "iwght_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffff170fffffffffffffe76fffffffffffff509fffffffffffff8e0ffffffff",
            INIT_01 => X"00002a0c00000000ffffb7b0ffffffff00003001000000000000007300000000",
            INIT_02 => X"ffffe731ffffffffffffe7efffffffff000006a4000000000000052100000000",
            INIT_03 => X"000016b30000000000000b7a00000000000015ce0000000000000dc200000000",
            INIT_04 => X"0000234200000000fffff083fffffffffffffd10fffffffffffff645ffffffff",
            INIT_05 => X"00000a6300000000fffff8a1ffffffff000023230000000000000bd500000000",
            INIT_06 => X"ffffddffffffffff000017c200000000000002700000000000000f0a00000000",
            INIT_07 => X"00002a4900000000000018e600000000ffffee1effffffff000007d600000000",
            INIT_08 => X"0000000000000000fffffff2fffffffffffffff5ffffffff0000000600000000",
            INIT_09 => X"fffffff7ffffffffffffffedfffffffffffffffaffffffffffffffedffffffff",
            INIT_0A => X"ffffffd7ffffffffffffffefffffffff0000000500000000fffffff2ffffffff",
            INIT_0B => X"ffffffddffffffff0000001700000000fffffffdffffffffffffffcfffffffff",
            INIT_0C => X"ffffffe4fffffffffffffffdffffffffffffffe9ffffffff0000001000000000",
            INIT_0D => X"ffffffdcffffffffffffffebffffffffffffffebffffffff0000000500000000",
            INIT_0E => X"ffffffe2ffffffffffffffdcffffffff0000000200000000fffffff5ffffffff",
            INIT_0F => X"fffffff5ffffffff00000004000000000000000800000000ffffffd1ffffffff",
            INIT_10 => X"ffffffdcffffffffffffffdfffffffffffffffd3fffffffffffffffeffffffff",
            INIT_11 => X"0000000c00000000fffffff7ffffffffffffffdeffffffffffffffeaffffffff",
            INIT_12 => X"ffffffe8ffffffff0000000000000000fffffffbffffffffffffffffffffffff",
            INIT_13 => X"0000001300000000000000090000000000000014000000000000001c00000000",
            INIT_14 => X"0000000400000000fffffff6ffffffffffffffeaffffffff0000000000000000",
            INIT_15 => X"fffffff5fffffffffffffffcffffffff0000001500000000fffffff9ffffffff",
            INIT_16 => X"00000013000000000000001600000000fffffffaffffffffffffffe4ffffffff",
            INIT_17 => X"ffffffeafffffffffffffffafffffffffffffffcffffffffffffffecffffffff",
            INIT_18 => X"ffffffe4ffffffffffffffeaffffffff0000000900000000fffffff9ffffffff",
            INIT_19 => X"00000004000000000000001a00000000fffffff2ffffffff0000001c00000000",
            INIT_1A => X"fffffff4fffffffffffffff3ffffffff0000000700000000ffffffedffffffff",
            INIT_1B => X"0000001500000000fffffff5ffffffffffffffe2ffffffffffffffe4ffffffff",
            INIT_1C => X"0000000f00000000fffffff0ffffffff0000000000000000fffffff8ffffffff",
            INIT_1D => X"ffffffd9ffffffffffffffe2fffffffffffffff1ffffffffffffffdbffffffff",
            INIT_1E => X"fffffff5fffffffffffffff4ffffffffffffffd7ffffffffffffffd4ffffffff",
            INIT_1F => X"ffffffdaffffffffffffffefffffffffffffffdaffffffffffffffe2ffffffff",
            INIT_20 => X"ffffffe4ffffffffffffffd0ffffffffffffffe3fffffffffffffff8ffffffff",
            INIT_21 => X"0000000c00000000ffffffe8ffffffff00000016000000000000000000000000",
            INIT_22 => X"ffffffddffffffffffffffd0ffffffffffffffe6fffffffffffffff9ffffffff",
            INIT_23 => X"00000003000000000000000e00000000fffffff2ffffffff0000000500000000",
            INIT_24 => X"ffffffdbffffffffffffffe3ffffffffffffffedfffffffffffffff3ffffffff",
            INIT_25 => X"0000000d000000000000001700000000fffffffaffffffffffffffe0ffffffff",
            INIT_26 => X"ffffffe7ffffffff0000000000000000ffffffefffffffff0000000600000000",
            INIT_27 => X"ffffffdefffffffffffffffbffffffffffffffe5ffffffff0000001300000000",
            INIT_28 => X"ffffffeaffffffffffffffeaffffffffffffffe6ffffffff0000000400000000",
            INIT_29 => X"0000000d000000000000000a0000000000000005000000000000001200000000",
            INIT_2A => X"0000000000000000fffffffcfffffffffffffffafffffffffffffff9ffffffff",
            INIT_2B => X"fffffff5ffffffffffffffe0ffffffffffffffdaffffffffffffffdcffffffff",
            INIT_2C => X"00000009000000000000002c0000000000000015000000000000001400000000",
            INIT_2D => X"ffffffeefffffffffffffff5ffffffff0000001e000000000000000a00000000",
            INIT_2E => X"ffffffffffffffff000000160000000000000016000000000000000e00000000",
            INIT_2F => X"ffffffedffffffff0000001300000000fffffffeffffffff0000000a00000000",
            INIT_30 => X"0000000b00000000000000080000000000000014000000000000001400000000",
            INIT_31 => X"ffffffe8ffffffff0000000000000000ffffffeafffffffffffffffdffffffff",
            INIT_32 => X"00000030000000000000000000000000fffffff6ffffffffffffffeeffffffff",
            INIT_33 => X"0000000f000000000000000d0000000000000015000000000000002600000000",
            INIT_34 => X"ffffffe2ffffffffffffffcbffffffffffffffd2fffffffffffffff1ffffffff",
            INIT_35 => X"0000002900000000000000120000000000000036000000000000002700000000",
            INIT_36 => X"0000003c0000000000000004000000000000004f000000000000005700000000",
            INIT_37 => X"0000000c0000000000000036000000000000000a000000000000002e00000000",
            INIT_38 => X"ffffffdfffffffffffffffecfffffffffffffff4ffffffff0000000900000000",
            INIT_39 => X"0000001a000000000000001100000000ffffffd9ffffffffffffffd4ffffffff",
            INIT_3A => X"000000070000000000000000000000000000000a00000000ffffffedffffffff",
            INIT_3B => X"0000000400000000ffffffe6ffffffffffffffc1ffffffffffffffafffffffff",
            INIT_3C => X"fffffffafffffffffffffff8ffffffff00000031000000000000001d00000000",
            INIT_3D => X"ffffffd7ffffffffffffffc3ffffffffffffffe0fffffffffffffff0ffffffff",
            INIT_3E => X"0000003d00000000000000110000000000000058000000000000001400000000",
            INIT_3F => X"0000000f00000000fffffff0ffffffff00000030000000000000006800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000030000000000000000a000000000000000f00000000ffffffdeffffffff",
            INIT_41 => X"ffffffd4fffffffffffffff7ffffffff0000001200000000ffffffe8ffffffff",
            INIT_42 => X"0000003f000000000000003a00000000ffffffddffffffff0000000100000000",
            INIT_43 => X"0000006200000000000000600000000000000059000000000000004e00000000",
            INIT_44 => X"0000001700000000000000370000000000000049000000000000002900000000",
            INIT_45 => X"ffffffe6fffffffffffffff6ffffffff0000000b000000000000001200000000",
            INIT_46 => X"ffffffeaffffffff0000000300000000ffffffe6ffffffff0000000600000000",
            INIT_47 => X"0000001700000000fffffff8ffffffff00000011000000000000001000000000",
            INIT_48 => X"fffffffbfffffffffffffffaffffffff0000000500000000fffffffbffffffff",
            INIT_49 => X"ffffffbfffffffffffffffc7ffffffffffffffecffffffff0000001a00000000",
            INIT_4A => X"0000001e0000000000000021000000000000002b00000000ffffffeeffffffff",
            INIT_4B => X"0000003d00000000000000210000000000000004000000000000001200000000",
            INIT_4C => X"fffffff8ffffffff00000009000000000000000d000000000000003500000000",
            INIT_4D => X"0000000b00000000ffffffe3ffffffffffffffe9ffffffffffffffd2ffffffff",
            INIT_4E => X"0000000200000000000000060000000000000022000000000000001c00000000",
            INIT_4F => X"ffffffcaffffffffffffffc8ffffffffffffffdaffffffffffffffdeffffffff",
            INIT_50 => X"0000001e00000000ffffffefffffffffffffffc5ffffffff0000000900000000",
            INIT_51 => X"ffffffe4ffffffff00000032000000000000000600000000ffffffbfffffffff",
            INIT_52 => X"00000002000000000000001700000000ffffffd2ffffffff0000000900000000",
            INIT_53 => X"ffffffcefffffffffffffff6ffffffff0000000400000000ffffffe2ffffffff",
            INIT_54 => X"0000001f0000000000000011000000000000002c00000000fffffff6ffffffff",
            INIT_55 => X"fffffff4ffffffff0000001b00000000ffffffcafffffffffffffff2ffffffff",
            INIT_56 => X"0000003b0000000000000007000000000000000800000000fffffff8ffffffff",
            INIT_57 => X"ffffffb2ffffffff0000005f000000000000001900000000ffffffaeffffffff",
            INIT_58 => X"fffffffeffffffffffffffd7ffffffff0000005e000000000000001300000000",
            INIT_59 => X"0000000100000000ffffffd9ffffffffffffffd0ffffffff0000001200000000",
            INIT_5A => X"fffffffbffffffffffffffeaffffffffffffffe4fffffffffffffff3ffffffff",
            INIT_5B => X"0000001a00000000ffffffeeffffffff0000001e00000000fffffffcffffffff",
            INIT_5C => X"0000001f000000000000000000000000ffffffcffffffffffffffff7ffffffff",
            INIT_5D => X"0000005600000000ffffffa4ffffffff00000005000000000000000300000000",
            INIT_5E => X"0000000b000000000000008b00000000ffffff63ffffffff0000001700000000",
            INIT_5F => X"0000001f000000000000001d000000000000004600000000ffffff8affffffff",
            INIT_60 => X"ffffffeaffffffff0000001400000000ffffffddffffffff0000000b00000000",
            INIT_61 => X"ffffffffffffffffffffffd4ffffffff0000001600000000fffffff3ffffffff",
            INIT_62 => X"0000001b00000000ffffffe6fffffffffffffff0ffffffff0000001400000000",
            INIT_63 => X"ffffffdcfffffffffffffff4fffffffffffffff7ffffffffffffffeaffffffff",
            INIT_64 => X"0000001700000000fffffff7ffffffffffffffe2fffffffffffffff7ffffffff",
            INIT_65 => X"00000022000000000000001400000000ffffffe1fffffffffffffff6ffffffff",
            INIT_66 => X"ffffffe5ffffffff0000003300000000ffffffeffffffffffffffff5ffffffff",
            INIT_67 => X"ffffffedffffffff00000002000000000000006200000000fffffff0ffffffff",
            INIT_68 => X"ffffffdbfffffffffffffffeffffffff00000023000000000000000f00000000",
            INIT_69 => X"0000005000000000ffffff92ffffffff00000013000000000000004500000000",
            INIT_6A => X"0000001c000000000000001a00000000ffffffbbffffffff0000000500000000",
            INIT_6B => X"ffffff49ffffffff0000000c000000000000004700000000ffffff73ffffffff",
            INIT_6C => X"0000005400000000ffffff68ffffffff0000001b000000000000005700000000",
            INIT_6D => X"fffffffaffffffffffffffd2ffffffff00000012000000000000000e00000000",
            INIT_6E => X"0000001900000000ffffffe9ffffffffffffffd6fffffffffffffff2ffffffff",
            INIT_6F => X"00000003000000000000000800000000fffffff6fffffffffffffffdffffffff",
            INIT_70 => X"fffffffdfffffffffffffff8ffffffff00000022000000000000001200000000",
            INIT_71 => X"00000042000000000000000100000000ffffffd5ffffffff0000000400000000",
            INIT_72 => X"ffffffc9ffffffff00000045000000000000000100000000ffffffaaffffffff",
            INIT_73 => X"ffffffd8fffffffffffffffbfffffffffffffffaffffffff0000000d00000000",
            INIT_74 => X"0000003000000000fffffff4ffffffff0000001c000000000000001b00000000",
            INIT_75 => X"0000000000000000ffffffddfffffffffffffff4ffffffffffffffe3ffffffff",
            INIT_76 => X"0000001e00000000fffffff8ffffffff0000001600000000fffffffbffffffff",
            INIT_77 => X"ffffffdcffffffff0000001100000000ffffffebfffffffffffffff3ffffffff",
            INIT_78 => X"ffffffe6ffffffffffffffaeffffffff00000036000000000000001600000000",
            INIT_79 => X"0000003b000000000000000b00000000ffffffeeffffffff0000001e00000000",
            INIT_7A => X"ffffffb5ffffffff0000002d00000000fffffff3ffffffff0000000600000000",
            INIT_7B => X"ffffffc4ffffffffffffff83ffffffffffffffe3ffffffffffffffdeffffffff",
            INIT_7C => X"0000004000000000ffffffefffffffffffffffa7ffffffff0000000a00000000",
            INIT_7D => X"fffffff5ffffffff00000024000000000000000000000000ffffffc5ffffffff",
            INIT_7E => X"0000001a00000000000000160000000000000014000000000000004200000000",
            INIT_7F => X"ffffffeeffffffff0000000e000000000000000a00000000ffffffe3ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE0;


    MEM_IWGHT_LAYER1_INSTANCE1 : if BRAM_NAME = "iwght_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffd9ffffffff0000000900000000ffffffe3ffffffffffffffe6ffffffff",
            INIT_01 => X"0000002a000000000000001600000000fffffffbfffffffffffffff0ffffffff",
            INIT_02 => X"0000001c000000000000001c000000000000004c000000000000004700000000",
            INIT_03 => X"00000029000000000000000400000000fffffffeffffffff0000004700000000",
            INIT_04 => X"ffffffc8ffffffff0000001100000000ffffffe8ffffffffffffffdfffffffff",
            INIT_05 => X"fffffff0fffffffffffffff9ffffffffffffffe1ffffffffffffffdbffffffff",
            INIT_06 => X"ffffffcdffffffffffffffe6ffffffffffffffe2ffffffff0000001f00000000",
            INIT_07 => X"0000000000000000ffffffacffffffff0000000800000000ffffffc1ffffffff",
            INIT_08 => X"0000002d00000000ffffffefffffffffffffffdefffffffffffffff9ffffffff",
            INIT_09 => X"ffffffd7ffffffff00000016000000000000001100000000ffffffefffffffff",
            INIT_0A => X"ffffffceffffffff000000000000000000000030000000000000000f00000000",
            INIT_0B => X"0000000d00000000ffffffcaffffffffffffffceffffffffffffffcdffffffff",
            INIT_0C => X"ffffffd9ffffffff0000000200000000ffffffc8ffffffffffffff94ffffffff",
            INIT_0D => X"0000000e00000000ffffffedffffffff0000000b00000000fffffff9ffffffff",
            INIT_0E => X"0000002800000000000000170000000000000001000000000000003f00000000",
            INIT_0F => X"00000050000000000000004d0000000000000042000000000000001600000000",
            INIT_10 => X"0000002a0000000000000049000000000000003c000000000000004f00000000",
            INIT_11 => X"00000039000000000000003100000000ffffffcafffffffffffffff2ffffffff",
            INIT_12 => X"0000003a00000000ffffffeaffffffff00000032000000000000000f00000000",
            INIT_13 => X"0000001200000000ffffffe2ffffffff00000021000000000000002a00000000",
            INIT_14 => X"00000019000000000000001b00000000ffffffc4ffffffff0000000c00000000",
            INIT_15 => X"ffffffe9ffffffff00000006000000000000002900000000ffffffdbffffffff",
            INIT_16 => X"ffffff9fffffffffffffffc0ffffffffffffff8cffffffffffffffaeffffffff",
            INIT_17 => X"ffffffecffffffffffffffd2ffffffffffffffaaffffffffffffffdcffffffff",
            INIT_18 => X"fffffff6fffffffffffffff0ffffffff00000015000000000000000f00000000",
            INIT_19 => X"0000003400000000ffffffecffffffffffffffd5ffffffff0000000a00000000",
            INIT_1A => X"0000000600000000ffffffe7ffffffff0000001800000000ffffffd5ffffffff",
            INIT_1B => X"fffffffeffffffff0000000b00000000ffffffe0ffffffff0000000500000000",
            INIT_1C => X"fffffff4fffffffffffffff8fffffffffffffffcfffffffffffffff2ffffffff",
            INIT_1D => X"0000002500000000ffffffccffffffff0000002c000000000000000500000000",
            INIT_1E => X"0000000c000000000000002700000000ffffffc0ffffffff0000002f00000000",
            INIT_1F => X"0000006100000000ffffffdaffffffffffffffd2ffffffff0000004400000000",
            INIT_20 => X"ffffffc8ffffffff0000004a00000000ffffffe5ffffffffffffffacffffffff",
            INIT_21 => X"ffffffcaffffffffffffffe5fffffffffffffff0ffffffff0000000300000000",
            INIT_22 => X"ffffffc4ffffffff0000001d00000000ffffffd5ffffffffffffffccffffffff",
            INIT_23 => X"ffffffeeffffffff0000000c00000000fffffffdffffffff0000000e00000000",
            INIT_24 => X"fffffff1ffffffffffffffd8ffffffff0000002e000000000000000c00000000",
            INIT_25 => X"ffffffbbffffffff0000001b00000000ffffffc5ffffffff0000001900000000",
            INIT_26 => X"0000006800000000ffffff38ffffffff00000039000000000000001900000000",
            INIT_27 => X"0000002b000000000000005f00000000ffffff6affffffff0000003100000000",
            INIT_28 => X"0000003300000000ffffffe6ffffffff00000019000000000000000500000000",
            INIT_29 => X"ffffffc7ffffffff00000039000000000000000f000000000000000500000000",
            INIT_2A => X"fffffffbfffffffffffffff3ffffffff00000003000000000000000000000000",
            INIT_2B => X"0000000700000000ffffffccffffffffffffffddfffffffffffffffbffffffff",
            INIT_2C => X"ffffffeefffffffffffffff7ffffffff0000000f00000000ffffffc4ffffffff",
            INIT_2D => X"0000002900000000fffffff1ffffffff0000000000000000fffffff8ffffffff",
            INIT_2E => X"0000002c00000000ffffffd1ffffffffffffffebfffffffffffffffcffffffff",
            INIT_2F => X"ffffffe1ffffffff0000003e00000000ffffffcbffffffffffffffe9ffffffff",
            INIT_30 => X"0000001d00000000ffffffd3ffffffff0000003900000000ffffffbfffffffff",
            INIT_31 => X"ffffffa5ffffffff0000001e000000000000002300000000ffffffdaffffffff",
            INIT_32 => X"0000005b00000000ffffff78ffffffff0000002a000000000000002a00000000",
            INIT_33 => X"00000054000000000000001200000000ffffffd0ffffffff0000001c00000000",
            INIT_34 => X"ffffff67ffffffff00000059000000000000004e00000000ffffff86ffffffff",
            INIT_35 => X"fffffff3ffffffff000000040000000000000020000000000000007f00000000",
            INIT_36 => X"0000000f000000000000001700000000ffffffe2ffffffff0000001e00000000",
            INIT_37 => X"00000016000000000000000d00000000fffffffaffffffff0000000300000000",
            INIT_38 => X"ffffffc4ffffffff0000001c00000000fffffffeffffffffffffffe8ffffffff",
            INIT_39 => X"ffffffdeffffffffffffffe7ffffffff00000000000000000000003100000000",
            INIT_3A => X"0000006000000000ffffffd3ffffffffffffffc9ffffffff0000003300000000",
            INIT_3B => X"ffffffacffffffff0000004c000000000000000900000000ffffff81ffffffff",
            INIT_3C => X"fffffff0fffffffffffffff1ffffffffffffffefffffffff0000001300000000",
            INIT_3D => X"00000004000000000000000700000000ffffffecfffffffffffffff1ffffffff",
            INIT_3E => X"0000001900000000fffffff4ffffffff0000001000000000fffffff9ffffffff",
            INIT_3F => X"ffffffdbffffffffffffffe0ffffffffffffffffffffffffffffffc6ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffaffffffff0000001100000000ffffffc5ffffffffffffffbeffffffff",
            INIT_41 => X"00000011000000000000001000000000ffffffe9ffffffff0000002300000000",
            INIT_42 => X"0000002f00000000000000210000000000000001000000000000000f00000000",
            INIT_43 => X"00000008000000000000000a000000000000000c000000000000000500000000",
            INIT_44 => X"ffffffedfffffffffffffffdffffffff0000003a000000000000001100000000",
            INIT_45 => X"ffffff69ffffffffffffff88ffffffffffffff90ffffffffffffff91ffffffff",
            INIT_46 => X"ffffff7dffffffffffffff7dffffffffffffff8bffffffffffffff23ffffffff",
            INIT_47 => X"fffffff9ffffffff0000000c000000000000002200000000ffffff94ffffffff",
            INIT_48 => X"0000003800000000ffffffe6fffffffffffffffaffffffff0000001a00000000",
            INIT_49 => X"00000027000000000000000e00000000ffffffe1ffffffff0000001700000000",
            INIT_4A => X"00000009000000000000002300000000fffffffdffffffff0000001200000000",
            INIT_4B => X"0000000d00000000ffffffe8ffffffff0000000f00000000fffffffdffffffff",
            INIT_4C => X"ffffffecffffffffffffffefffffffff00000015000000000000001600000000",
            INIT_4D => X"000000090000000000000012000000000000000f000000000000001f00000000",
            INIT_4E => X"ffffffc5ffffffffffffffebffffffffffffffd6ffffffff0000000600000000",
            INIT_4F => X"ffffffa5ffffffffffffffaeffffffffffffffa8ffffffffffffffb1ffffffff",
            INIT_50 => X"ffffffe3ffffffff0000000a00000000ffffffdeffffffffffffff9bffffffff",
            INIT_51 => X"fffffffeffffffffffffffdbfffffffffffffff6ffffffff0000001700000000",
            INIT_52 => X"ffffffb7ffffffffffffffe7ffffffff0000001500000000fffffff0ffffffff",
            INIT_53 => X"ffffff84ffffffffffffff87ffffffffffffffc3fffffffffffffff7ffffffff",
            INIT_54 => X"0000000f00000000ffffff8effffffffffffff94ffffffffffffffbcffffffff",
            INIT_55 => X"fffffffffffffffffffffffeffffffff0000001f00000000ffffffedffffffff",
            INIT_56 => X"0000000b000000000000000100000000ffffffe7ffffffff0000002000000000",
            INIT_57 => X"000000100000000000000007000000000000002300000000ffffffe3ffffffff",
            INIT_58 => X"0000002f00000000000000140000000000000007000000000000002800000000",
            INIT_59 => X"ffffffa9ffffffffffffff7effffffffffffff8fffffffff0000000200000000",
            INIT_5A => X"ffffffadffffffffffffffb0ffffffffffffff70ffffffffffffff71ffffffff",
            INIT_5B => X"0000000200000000fffffff7ffffffffffffffe3ffffffffffffffc8ffffffff",
            INIT_5C => X"ffffffcdffffffffffffffe5ffffffff0000001200000000ffffffe2ffffffff",
            INIT_5D => X"fffffff8ffffffff00000001000000000000000c000000000000001c00000000",
            INIT_5E => X"0000001e000000000000000000000000ffffffeeffffffff0000000d00000000",
            INIT_5F => X"0000002200000000000000190000000000000013000000000000000a00000000",
            INIT_60 => X"fffffff7fffffffffffffffcffffffff00000028000000000000001600000000",
            INIT_61 => X"0000003b000000000000002600000000fffffff0ffffffff0000001d00000000",
            INIT_62 => X"ffffffddffffffff0000002f000000000000001b000000000000001700000000",
            INIT_63 => X"ffffffd5ffffffff0000000d00000000fffffff3fffffffffffffffdffffffff",
            INIT_64 => X"00000010000000000000003200000000ffffffd3ffffffffffffffd9ffffffff",
            INIT_65 => X"000000080000000000000004000000000000002a000000000000002800000000",
            INIT_66 => X"0000002c000000000000000c0000000000000003000000000000001400000000",
            INIT_67 => X"fffffff7ffffffff0000001d00000000ffffffeaffffffff0000002f00000000",
            INIT_68 => X"fffffff0ffffffff0000001800000000fffffffdffffffff0000000d00000000",
            INIT_69 => X"0000003000000000ffffffd7ffffffff0000004200000000fffffffdffffffff",
            INIT_6A => X"0000000a000000000000001b0000000000000021000000000000003000000000",
            INIT_6B => X"fffffff2ffffffffffffffe3ffffffffffffffc3ffffffff0000000d00000000",
            INIT_6C => X"0000004400000000fffffffffffffffffffffffbffffffffffffffefffffffff",
            INIT_6D => X"0000000600000000ffffffeaffffffff0000000b000000000000003f00000000",
            INIT_6E => X"0000002f00000000000000190000000000000021000000000000000300000000",
            INIT_6F => X"ffffffacffffffff0000000f0000000000000035000000000000001900000000",
            INIT_70 => X"fffffffcfffffffffffffffcffffffffffffffaeffffffffffffff9bffffffff",
            INIT_71 => X"000000130000000000000027000000000000001d000000000000000100000000",
            INIT_72 => X"fffffff7ffffffffffffffddffffffffffffffdbffffffffffffffecffffffff",
            INIT_73 => X"0000003c00000000fffffff1ffffffffffffffe6ffffffff0000000200000000",
            INIT_74 => X"0000000f0000000000000008000000000000002b000000000000001600000000",
            INIT_75 => X"00000019000000000000000000000000fffffff3fffffffffffffffbffffffff",
            INIT_76 => X"000000250000000000000033000000000000000d00000000ffffffdfffffffff",
            INIT_77 => X"ffffffe7ffffffff0000001600000000fffffffaffffffff0000002800000000",
            INIT_78 => X"0000003700000000ffffffcfffffffff0000000d00000000fffffffdffffffff",
            INIT_79 => X"0000000f00000000000000050000000000000006000000000000001000000000",
            INIT_7A => X"0000000e00000000ffffffcdffffffffffffffcdffffffff0000000e00000000",
            INIT_7B => X"0000002700000000000000360000000000000026000000000000001800000000",
            INIT_7C => X"ffffffbeffffffffffffffe9ffffffff0000000600000000fffffff9ffffffff",
            INIT_7D => X"ffffffeaffffffff0000000a000000000000001600000000ffffffe2ffffffff",
            INIT_7E => X"0000000200000000ffffffd8ffffffffffffffe5ffffffff0000000f00000000",
            INIT_7F => X"0000000900000000ffffffc5ffffffffffffffdfffffffffffffffd6ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE1;


    MEM_IWGHT_LAYER1_INSTANCE2 : if BRAM_NAME = "iwght_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001f000000000000001c000000000000002000000000fffffff0ffffffff",
            INIT_01 => X"ffffffd6ffffffff000000290000000000000018000000000000002d00000000",
            INIT_02 => X"ffffffd5ffffffffffffffcdffffffff00000009000000000000000600000000",
            INIT_03 => X"ffffffc4ffffffffffffffdeffffffffffffffedffffffff0000002600000000",
            INIT_04 => X"fffffff6ffffffffffffffc7ffffffffffffffdeffffffffffffffddffffffff",
            INIT_05 => X"0000001f000000000000000200000000ffffffe9ffffffffffffffdeffffffff",
            INIT_06 => X"0000000000000000ffffffd7ffffffffffffffeeffffffff0000001600000000",
            INIT_07 => X"ffffffedffffffffffffffecffffffffffffffd8ffffffffffffffd6ffffffff",
            INIT_08 => X"0000000100000000fffffff1ffffffff0000000200000000ffffffd3ffffffff",
            INIT_09 => X"fffffff5fffffffffffffffefffffffffffffff9ffffffff0000001c00000000",
            INIT_0A => X"00000002000000000000000a000000000000000000000000fffffff7ffffffff",
            INIT_0B => X"fffffff8fffffffffffffff4fffffffffffffffbffffffffffffffffffffffff",
            INIT_0C => X"0000000600000000ffffffefffffffffffffffdcffffffff0000000000000000",
            INIT_0D => X"0000003c00000000fffffff6ffffffff0000002a000000000000002600000000",
            INIT_0E => X"0000004800000000000000440000000000000013000000000000003b00000000",
            INIT_0F => X"fffffff7ffffffff0000000a00000000fffffff5ffffffff0000002700000000",
            INIT_10 => X"00000024000000000000001200000000fffffffffffffffffffffff5ffffffff",
            INIT_11 => X"0000002600000000000000000000000000000007000000000000002600000000",
            INIT_12 => X"0000002e00000000000000030000000000000018000000000000003000000000",
            INIT_13 => X"ffffffcdffffffff0000000c00000000fffffff3ffffffff0000001600000000",
            INIT_14 => X"ffffffaeffffffffffffffc1ffffffffffffffaaffffffffffffff92ffffffff",
            INIT_15 => X"ffffff6bffffffffffffffa0ffffffffffffff9dffffffffffffff82ffffffff",
            INIT_16 => X"0000000400000000fffffff4ffffffffffffffdaffffffff0000002300000000",
            INIT_17 => X"0000000600000000ffffffcfffffffffffffffe1ffffffff0000001e00000000",
            INIT_18 => X"0000000b00000000ffffffdfffffffff0000000000000000ffffffefffffffff",
            INIT_19 => X"0000001500000000ffffffdffffffffffffffff1fffffffffffffff8ffffffff",
            INIT_1A => X"00000020000000000000002b00000000ffffffdeffffffff0000001b00000000",
            INIT_1B => X"0000000c000000000000003d0000000000000021000000000000000100000000",
            INIT_1C => X"000000220000000000000021000000000000001e000000000000000200000000",
            INIT_1D => X"fffffffffffffffffffffff9ffffffff00000020000000000000000000000000",
            INIT_1E => X"ffffffecffffffff0000000000000000ffffffffffffffff0000000200000000",
            INIT_1F => X"0000000800000000fffffff1ffffffff0000001500000000fffffffbffffffff",
            INIT_20 => X"fffffff5ffffffff00000002000000000000002000000000ffffffe2ffffffff",
            INIT_21 => X"ffffffe0ffffffffffffffd0fffffffffffffff2ffffffff0000000e00000000",
            INIT_22 => X"ffffffc8ffffffffffffffd1ffffffffffffffdfffffffff0000001300000000",
            INIT_23 => X"fffffff0ffffffffffffffd0ffffffffffffffd8ffffffffffffffd8ffffffff",
            INIT_24 => X"0000000b00000000ffffffe2fffffffffffffff4ffffffffffffffe1ffffffff",
            INIT_25 => X"00000000000000000000000d00000000fffffff8ffffffff0000000800000000",
            INIT_26 => X"fffffff8fffffffffffffffbffffffffffffffd4fffffffffffffff2ffffffff",
            INIT_27 => X"fffffffcffffffffffffffeaffffffffffffffecffffffffffffffd0ffffffff",
            INIT_28 => X"fffffff1ffffffff00000015000000000000000d000000000000001900000000",
            INIT_29 => X"ffffffcaffffffff0000000000000000fffffff5fffffffffffffffbffffffff",
            INIT_2A => X"0000002b000000000000001b00000000ffffffe8ffffffffffffffb6ffffffff",
            INIT_2B => X"0000001c00000000fffffff9ffffffff0000000c00000000fffffff8ffffffff",
            INIT_2C => X"000000010000000000000009000000000000002500000000fffffff0ffffffff",
            INIT_2D => X"0000002000000000fffffff1fffffffffffffff6ffffffffffffffe4ffffffff",
            INIT_2E => X"fffffffcffffffff0000001500000000ffffffe7ffffffffffffffe5ffffffff",
            INIT_2F => X"0000002000000000000000270000000000000010000000000000001200000000",
            INIT_30 => X"000000140000000000000012000000000000000f000000000000001200000000",
            INIT_31 => X"ffffff8dffffffffffffffd6ffffffffffffffc6ffffffff0000001500000000",
            INIT_32 => X"0000000f00000000ffffffd2ffffffff0000002100000000ffffffb7ffffffff",
            INIT_33 => X"0000002200000000000000020000000000000023000000000000000400000000",
            INIT_34 => X"fffffff9ffffffff0000001200000000fffffffeffffffff0000000600000000",
            INIT_35 => X"fffffff9ffffffff0000001a00000000ffffffe5ffffffffffffffecffffffff",
            INIT_36 => X"0000001d000000000000001a00000000ffffffefffffffff0000001400000000",
            INIT_37 => X"0000001d0000000000000011000000000000001600000000fffffff3ffffffff",
            INIT_38 => X"000000160000000000000026000000000000000c000000000000000c00000000",
            INIT_39 => X"0000000f000000000000000e0000000000000015000000000000002000000000",
            INIT_3A => X"00000005000000000000000c0000000000000026000000000000002700000000",
            INIT_3B => X"0000002e000000000000000a00000000fffffff9ffffffff0000000e00000000",
            INIT_3C => X"ffffffffffffffff0000001a000000000000002c000000000000000000000000",
            INIT_3D => X"0000000300000000ffffffebffffffffffffffd7ffffffff0000000a00000000",
            INIT_3E => X"0000003f00000000fffffffeffffffffffffffd0ffffffffffffffe0ffffffff",
            INIT_3F => X"00000021000000000000003d0000000000000049000000000000001800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffc4ffffffff000000290000000000000039000000000000003f00000000",
            INIT_41 => X"fffffff8ffffffffffffffd3fffffffffffffff6ffffffffffffffd7ffffffff",
            INIT_42 => X"fffffffdffffffff0000001000000000fffffff3fffffffffffffff3ffffffff",
            INIT_43 => X"ffffffeaffffffffffffffebffffffffffffffdeffffffff0000003100000000",
            INIT_44 => X"ffffffe5fffffffffffffff0ffffffffffffffd8ffffffffffffffaaffffffff",
            INIT_45 => X"ffffffc4ffffffffffffffd3ffffffff0000000d000000000000001a00000000",
            INIT_46 => X"ffffffe4fffffffffffffff8fffffffffffffff6ffffffffffffffd2ffffffff",
            INIT_47 => X"0000001300000000000000230000000000000028000000000000002900000000",
            INIT_48 => X"fffffff1ffffffffffffffe6fffffffffffffff4fffffffffffffff3ffffffff",
            INIT_49 => X"0000001800000000ffffffdeffffffffffffffbdffffffffffffffd1ffffffff",
            INIT_4A => X"fffffff1fffffffffffffffdfffffffffffffff1ffffffff0000001e00000000",
            INIT_4B => X"fffffff8ffffffffffffffcbffffffffffffffe4ffffffffffffffceffffffff",
            INIT_4C => X"ffffffedffffffffffffffc5ffffffffffffffe8ffffffff0000002e00000000",
            INIT_4D => X"0000002400000000fffffff7ffffffffffffffe8fffffffffffffffbffffffff",
            INIT_4E => X"fffffff5ffffffff0000000400000000fffffff7ffffffff0000000400000000",
            INIT_4F => X"00000038000000000000000a000000000000001d000000000000002a00000000",
            INIT_50 => X"00000013000000000000001c00000000fffffffdfffffffffffffff2ffffffff",
            INIT_51 => X"fffffffdffffffffffffffebfffffffffffffff1ffffffff0000001400000000",
            INIT_52 => X"00000034000000000000000400000000ffffffedffffffff0000000200000000",
            INIT_53 => X"00000025000000000000002600000000fffffff7ffffffff0000000f00000000",
            INIT_54 => X"00000007000000000000001c000000000000001c00000000fffffffbffffffff",
            INIT_55 => X"0000006500000000000000020000000000000006000000000000000c00000000",
            INIT_56 => X"000000170000000000000035000000000000002a000000000000003800000000",
            INIT_57 => X"ffffffddfffffffffffffff7ffffffffffffffe0ffffffff0000000600000000",
            INIT_58 => X"ffffffe5ffffffffffffffc3ffffffffffffffddffffffffffffffe8ffffffff",
            INIT_59 => X"ffffffcbffffffffffffffddffffffffffffffcafffffffffffffff9ffffffff",
            INIT_5A => X"ffffff62ffffffffffffff78ffffffffffffffa7ffffffffffffffbcffffffff",
            INIT_5B => X"0000003500000000ffffff9cffffffffffffff96fffffffffffffff5ffffffff",
            INIT_5C => X"ffffffbdffffffffffffffc7ffffffff00000005000000000000003b00000000",
            INIT_5D => X"ffffffd7ffffffffffffffbfffffffffffffffdcffffffffffffffe9ffffffff",
            INIT_5E => X"00000004000000000000001000000000ffffffc7ffffffff0000002e00000000",
            INIT_5F => X"0000002300000000fffffff7ffffffffffffffdcffffffff0000001d00000000",
            INIT_60 => X"000000000000000000000008000000000000000a00000000fffffff5ffffffff",
            INIT_61 => X"fffffffaffffffffffffffe9ffffffffffffffe2ffffffff0000001900000000",
            INIT_62 => X"0000001e00000000000000000000000000000003000000000000001100000000",
            INIT_63 => X"0000001e0000000000000012000000000000001900000000fffffff7ffffffff",
            INIT_64 => X"fffffff6ffffffff00000023000000000000001b000000000000001c00000000",
            INIT_65 => X"fffffff8fffffffffffffffaffffffff0000001a000000000000000e00000000",
            INIT_66 => X"0000000f000000000000001b000000000000002b00000000fffffff2ffffffff",
            INIT_67 => X"fffffff2ffffffffffffffc1ffffffffffffffa1ffffffffffffffb1ffffffff",
            INIT_68 => X"ffffffccfffffffffffffffaffffffffffffffa5ffffffffffffffc1ffffffff",
            INIT_69 => X"ffffffeaffffffff0000000e000000000000000500000000ffffffb4ffffffff",
            INIT_6A => X"0000000a000000000000003e000000000000003c000000000000004000000000",
            INIT_6B => X"0000000800000000ffffffe5ffffffff00000030000000000000003700000000",
            INIT_6C => X"fffffff7ffffffffffffffe9fffffffffffffff1ffffffff0000001600000000",
            INIT_6D => X"ffffffe7ffffffffffffffedffffffff0000001400000000ffffffebffffffff",
            INIT_6E => X"00000005000000000000002c000000000000000100000000fffffff8ffffffff",
            INIT_6F => X"000000280000000000000029000000000000002b000000000000000800000000",
            INIT_70 => X"0000000100000000ffffffebffffffff0000000500000000ffffffe8ffffffff",
            INIT_71 => X"0000001800000000fffffffbfffffffffffffffeffffffff0000000000000000",
            INIT_72 => X"fffffff4ffffffffffffffe4ffffffff0000002100000000fffffffbffffffff",
            INIT_73 => X"ffffffe7ffffffff0000004b0000000000000033000000000000001100000000",
            INIT_74 => X"000000110000000000000029000000000000002200000000fffffff5ffffffff",
            INIT_75 => X"0000001c000000000000000a0000000000000024000000000000001d00000000",
            INIT_76 => X"fffffff9fffffffffffffff3ffffffffffffffe7ffffffffffffffe6ffffffff",
            INIT_77 => X"0000001e0000000000000005000000000000003400000000ffffffedffffffff",
            INIT_78 => X"ffffffe1ffffffffffffffe6fffffffffffffff1ffffffffffffffedffffffff",
            INIT_79 => X"000000120000000000000018000000000000001d00000000fffffffbffffffff",
            INIT_7A => X"0000001b0000000000000023000000000000001e000000000000001300000000",
            INIT_7B => X"ffffffe1ffffffff0000000d0000000000000013000000000000001200000000",
            INIT_7C => X"0000001300000000fffffffeffffffff00000024000000000000001400000000",
            INIT_7D => X"00000001000000000000003c00000000ffffffceffffffff0000000d00000000",
            INIT_7E => X"00000004000000000000003c000000000000001d00000000ffffffe7ffffffff",
            INIT_7F => X"0000001600000000000000320000000000000035000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE2;


    MEM_IWGHT_LAYER1_INSTANCE3 : if BRAM_NAME = "iwght_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000032000000000000004200000000ffffffedffffffff0000000000000000",
            INIT_01 => X"00000025000000000000001b000000000000001b000000000000003e00000000",
            INIT_02 => X"000000410000000000000015000000000000002000000000fffffffcffffffff",
            INIT_03 => X"0000003a000000000000002b000000000000002a000000000000006200000000",
            INIT_04 => X"0000000900000000fffffffdffffffff00000018000000000000004400000000",
            INIT_05 => X"ffffffe8ffffffff0000001700000000fffffffaffffffff0000000d00000000",
            INIT_06 => X"00000019000000000000000700000000ffffffcaffffffffffffffccffffffff",
            INIT_07 => X"0000004e00000000000000520000000000000036000000000000000000000000",
            INIT_08 => X"ffffffefffffffff000000410000000000000038000000000000001400000000",
            INIT_09 => X"000000230000000000000000000000000000000200000000fffffffbffffffff",
            INIT_0A => X"fffffff9ffffffff0000001100000000fffffffdffffffff0000002a00000000",
            INIT_0B => X"000000020000000000000014000000000000001e000000000000001b00000000",
            INIT_0C => X"ffffffe2fffffffffffffff8ffffffffffffffefffffffff0000000400000000",
            INIT_0D => X"fffffff2fffffffffffffff0ffffffff0000000a000000000000000900000000",
            INIT_0E => X"0000001900000000ffffffd4ffffffffffffffdeffffffff0000001000000000",
            INIT_0F => X"0000001300000000fffffff4ffffffffffffffc9fffffffffffffff2ffffffff",
            INIT_10 => X"fffffffaffffffff0000000a00000000fffffff9fffffffffffffffcffffffff",
            INIT_11 => X"fffffffafffffffffffffffdffffffffffffffd3ffffffffffffffd9ffffffff",
            INIT_12 => X"0000001e00000000fffffffbffffffff00000023000000000000000900000000",
            INIT_13 => X"fffffff8ffffffff0000000900000000fffffff7ffffffff0000000000000000",
            INIT_14 => X"000000040000000000000021000000000000000000000000ffffffeaffffffff",
            INIT_15 => X"0000001300000000fffffff7ffffffff0000002b000000000000000800000000",
            INIT_16 => X"0000001700000000fffffffdffffffff0000001f000000000000000300000000",
            INIT_17 => X"fffffffbffffffff0000001e000000000000001400000000ffffffe4ffffffff",
            INIT_18 => X"0000000700000000000000050000000000000035000000000000002d00000000",
            INIT_19 => X"ffffffeaffffffff0000001000000000ffffffdcffffffff0000001600000000",
            INIT_1A => X"fffffff6fffffffffffffffcffffffff0000001300000000ffffffe1ffffffff",
            INIT_1B => X"ffffffdcffffffffffffffd5ffffffff0000002a000000000000001a00000000",
            INIT_1C => X"0000001500000000ffffffbbffffffffffffffcefffffffffffffff0ffffffff",
            INIT_1D => X"ffffff4affffffffffffffe5ffffffffffffffd8ffffffffffffffaeffffffff",
            INIT_1E => X"ffffff73ffffffffffffff74ffffffffffffff63ffffffffffffff45ffffffff",
            INIT_1F => X"ffffffe4ffffffff0000000f000000000000000000000000ffffff65ffffffff",
            INIT_20 => X"fffffff6ffffffff000000000000000000000004000000000000000e00000000",
            INIT_21 => X"00000013000000000000003100000000ffffffe9ffffffff0000001a00000000",
            INIT_22 => X"ffffffe7ffffffff00000022000000000000005b00000000ffffffc9ffffffff",
            INIT_23 => X"fffffff7ffffffffffffffdaffffffff00000018000000000000003700000000",
            INIT_24 => X"00000003000000000000002800000000ffffffcbfffffffffffffffaffffffff",
            INIT_25 => X"000000060000000000000020000000000000005100000000ffffffd8ffffffff",
            INIT_26 => X"0000000200000000ffffffc5ffffffffffffffd7ffffffffffffffe2ffffffff",
            INIT_27 => X"0000002d000000000000004b00000000fffffffaffffffff0000001100000000",
            INIT_28 => X"00000037000000000000002b00000000ffffffeeffffffff0000001d00000000",
            INIT_29 => X"ffffffcbffffffff00000032000000000000001e00000000ffffffdbffffffff",
            INIT_2A => X"ffffff7effffffffffffffc1ffffffff0000000e000000000000000100000000",
            INIT_2B => X"ffffffd3ffffffffffffffc9ffffffffffffffc9ffffffffffffffccffffffff",
            INIT_2C => X"0000001600000000ffffffebffffffffffffffc6ffffffffffffffcbffffffff",
            INIT_2D => X"00000020000000000000000b0000000000000006000000000000000100000000",
            INIT_2E => X"00000019000000000000002d00000000fffffff5ffffffff0000001300000000",
            INIT_2F => X"0000003f000000000000000c0000000000000005000000000000003200000000",
            INIT_30 => X"000000370000000000000033000000000000001b000000000000002600000000",
            INIT_31 => X"00000022000000000000000c00000000fffffffaffffffff0000001500000000",
            INIT_32 => X"ffffffcbffffffffffffffd1ffffffffffffff99ffffffffffffff82ffffffff",
            INIT_33 => X"00000025000000000000001800000000fffffff3ffffffffffffffc3ffffffff",
            INIT_34 => X"0000001900000000fffffffbffffffff0000001800000000fffffff8ffffffff",
            INIT_35 => X"0000000200000000ffffffcdffffffffffffffe9ffffffff0000000100000000",
            INIT_36 => X"0000001500000000fffffff8ffffffff0000002700000000ffffffd9ffffffff",
            INIT_37 => X"0000001a00000000000000190000000000000018000000000000001900000000",
            INIT_38 => X"ffffffe6fffffffffffffffaffffffffffffffe0ffffffffffffffecffffffff",
            INIT_39 => X"fffffffeffffffff0000001200000000ffffffeeffffffffffffffddffffffff",
            INIT_3A => X"ffffffdfffffffff0000001100000000fffffff0ffffffff0000001800000000",
            INIT_3B => X"fffffff8ffffffffffffffd9ffffffff0000000c000000000000000c00000000",
            INIT_3C => X"fffffff4ffffffff0000000500000000ffffffdcfffffffffffffffbffffffff",
            INIT_3D => X"00000011000000000000000500000000fffffffcffffffff0000001200000000",
            INIT_3E => X"ffffffffffffffff0000001600000000ffffffe1ffffffffffffffeeffffffff",
            INIT_3F => X"00000000000000000000000000000000fffffff9ffffffff0000001100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffecffffffffffffffe2fffffffffffffff6ffffffff0000000e00000000",
            INIT_41 => X"ffffffcdffffffffffffffa3ffffffffffffff9fffffffffffffffceffffffff",
            INIT_42 => X"ffffffecffffffff0000001200000000ffffffbfffffffffffffffc8ffffffff",
            INIT_43 => X"0000001f000000000000000f000000000000000c00000000ffffffffffffffff",
            INIT_44 => X"0000001300000000000000070000000000000014000000000000000a00000000",
            INIT_45 => X"fffffffeffffffffffffffeeffffffff0000001800000000fffffff9ffffffff",
            INIT_46 => X"ffffffefffffffffffffffdbffffffffffffffdefffffffffffffffcffffffff",
            INIT_47 => X"ffffffafffffffff0000001200000000fffffff1ffffffffffffffcfffffffff",
            INIT_48 => X"ffffffb0ffffffffffffffafffffffffffffffd2ffffffffffffffd0ffffffff",
            INIT_49 => X"ffffffd6ffffffffffffffcaffffffffffffffeeffffffffffffffddffffffff",
            INIT_4A => X"ffffffefffffffffffffff97ffffffffffffffa8ffffffffffffff96ffffffff",
            INIT_4B => X"0000001300000000fffffff4ffffffffffffffe9ffffffffffffffbdffffffff",
            INIT_4C => X"0000000100000000fffffffdffffffff0000000600000000fffffff0ffffffff",
            INIT_4D => X"0000001f0000000000000023000000000000001700000000fffffffeffffffff",
            INIT_4E => X"ffffff63ffffffffffffffadffffffff00000006000000000000002300000000",
            INIT_4F => X"ffffffc5ffffffffffffffb5ffffffffffffffc2ffffffffffffff95ffffffff",
            INIT_50 => X"0000001700000000ffffffdeffffffffffffffe2ffffffffffffffc4ffffffff",
            INIT_51 => X"0000000800000000ffffffe1fffffffffffffff8ffffffff0000001400000000",
            INIT_52 => X"fffffff0ffffffff00000009000000000000000a00000000fffffffbffffffff",
            INIT_53 => X"000000120000000000000003000000000000001e000000000000000b00000000",
            INIT_54 => X"0000000e000000000000001700000000fffffff0fffffffffffffff7ffffffff",
            INIT_55 => X"ffffffb1ffffffff0000000000000000fffffff1ffffffff0000001100000000",
            INIT_56 => X"0000001f00000000ffffffefffffffffffffffcfffffffffffffffe8ffffffff",
            INIT_57 => X"fffffffbffffffffffffffecffffffff00000014000000000000002800000000",
            INIT_58 => X"00000008000000000000000f000000000000000d00000000fffffff3ffffffff",
            INIT_59 => X"fffffff3ffffffffffffffdefffffffffffffffbffffffffffffffe3ffffffff",
            INIT_5A => X"0000000b00000000ffffffefffffffffffffffd0ffffffffffffffd7ffffffff",
            INIT_5B => X"fffffff7ffffffff0000002800000000fffffffdffffffffffffffcdffffffff",
            INIT_5C => X"ffffffd9ffffffff00000001000000000000000d00000000ffffffcdffffffff",
            INIT_5D => X"000000230000000000000001000000000000001c00000000fffffffeffffffff",
            INIT_5E => X"fffffff9ffffffffffffffefffffffff00000010000000000000002a00000000",
            INIT_5F => X"0000000a00000000ffffffecffffffffffffffe0ffffffff0000000e00000000",
            INIT_60 => X"fffffff2ffffffff0000000300000000ffffffddfffffffffffffffbffffffff",
            INIT_61 => X"fffffff5ffffffffffffffdfffffffffffffffffffffffff0000001100000000",
            INIT_62 => X"000000030000000000000010000000000000000a000000000000001b00000000",
            INIT_63 => X"fffffff2ffffffffffffffedffffffff00000016000000000000000300000000",
            INIT_64 => X"fffffff1fffffffffffffff1fffffffffffffffdffffffff0000000300000000",
            INIT_65 => X"0000006a000000000000002c0000000000000014000000000000003d00000000",
            INIT_66 => X"0000004d0000000000000069000000000000005c000000000000005f00000000",
            INIT_67 => X"ffffffb6ffffffffffffffc6ffffffffffffffbbffffffff0000007500000000",
            INIT_68 => X"0000002000000000fffffffbfffffffffffffff8ffffffffffffffaeffffffff",
            INIT_69 => X"ffffffd2ffffffffffffffc0ffffffff00000029000000000000001e00000000",
            INIT_6A => X"ffffffc6ffffffffffffff95ffffffffffffffa9ffffffffffffffc3ffffffff",
            INIT_6B => X"ffffff9bffffffffffffffe9ffffffffffffffcbffffffffffffffd3ffffffff",
            INIT_6C => X"ffffffb5ffffffffffffffbdffffffffffffffbdffffffffffffffa7ffffffff",
            INIT_6D => X"000000130000000000000027000000000000001b00000000ffffffb5ffffffff",
            INIT_6E => X"0000002c00000000ffffffe2ffffffff00000007000000000000002b00000000",
            INIT_6F => X"0000001e00000000ffffffe9ffffffff00000014000000000000004400000000",
            INIT_70 => X"00000011000000000000001e00000000fffffff1ffffffff0000000200000000",
            INIT_71 => X"00000000000000000000000100000000fffffff1ffffffff0000000000000000",
            INIT_72 => X"00000019000000000000001c000000000000000f00000000ffffffeeffffffff",
            INIT_73 => X"0000000900000000000000070000000000000002000000000000000500000000",
            INIT_74 => X"0000002900000000ffffffd1fffffffffffffff9ffffffff0000001000000000",
            INIT_75 => X"ffffffecffffffff000000070000000000000019000000000000000300000000",
            INIT_76 => X"fffffffeffffffffffffffd8fffffffffffffffdffffffff0000000b00000000",
            INIT_77 => X"fffffff5ffffffff00000002000000000000001e000000000000000c00000000",
            INIT_78 => X"ffffffe2ffffffff0000000c0000000000000015000000000000000e00000000",
            INIT_79 => X"fffffffdfffffffffffffff7fffffffffffffffcffffffff0000000700000000",
            INIT_7A => X"000000600000000000000028000000000000003a000000000000004f00000000",
            INIT_7B => X"fffffff2ffffffffffffffcfffffffff00000032000000000000003b00000000",
            INIT_7C => X"ffffffedffffffff0000001800000000fffffffbfffffffffffffff4ffffffff",
            INIT_7D => X"fffffffaffffffff0000003800000000fffffffffffffffffffffffbffffffff",
            INIT_7E => X"ffffffe6fffffffffffffff8fffffffffffffff6ffffffffffffffe3ffffffff",
            INIT_7F => X"00000008000000000000001600000000fffffff6fffffffffffffffbffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE3;


    MEM_IWGHT_LAYER1_INSTANCE4 : if BRAM_NAME = "iwght_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001800000000fffffffdfffffffffffffff0ffffffff0000000600000000",
            INIT_01 => X"fffffff0fffffffffffffffefffffffffffffffaffffffff0000000700000000",
            INIT_02 => X"0000002e000000000000000000000000ffffffdffffffffffffffff0ffffffff",
            INIT_03 => X"ffffffb6ffffffff0000000600000000fffffffaffffffffffffffe1ffffffff",
            INIT_04 => X"fffffffefffffffffffffffdfffffffffffffff2ffffffffffffffdbffffffff",
            INIT_05 => X"ffffffecffffffffffffffe1ffffffffffffffdfffffffff0000001f00000000",
            INIT_06 => X"0000001900000000000000010000000000000009000000000000000000000000",
            INIT_07 => X"00000008000000000000001e000000000000001f000000000000000600000000",
            INIT_08 => X"ffffffebffffffff0000000500000000fffffffeffffffff0000000500000000",
            INIT_09 => X"fffffef2ffffffffffffffe3ffffffffffffff56ffffffffffffff63ffffffff",
            INIT_0A => X"ffffff1effffffffffffff33ffffffffffffff1bfffffffffffffeb6ffffffff",
            INIT_0B => X"ffffffedffffffff0000002b000000000000003c00000000ffffff2fffffffff",
            INIT_0C => X"0000003b00000000fffffff3ffffffff00000019000000000000002900000000",
            INIT_0D => X"fffffffdffffffff000000190000000000000000000000000000002700000000",
            INIT_0E => X"fffffff2ffffffff00000003000000000000003900000000fffffff8ffffffff",
            INIT_0F => X"0000001e00000000ffffffeaffffffff0000000c000000000000001100000000",
            INIT_10 => X"00000004000000000000000f000000000000000000000000fffffff6ffffffff",
            INIT_11 => X"0000002a0000000000000019000000000000005100000000fffffffbffffffff",
            INIT_12 => X"0000002d000000000000001000000000ffffffd7ffffffff0000000000000000",
            INIT_13 => X"fffffff5ffffffff00000013000000000000002c00000000ffffffefffffffff",
            INIT_14 => X"0000000b000000000000000d000000000000002400000000fffffff3ffffffff",
            INIT_15 => X"fffffffdffffffff0000001f00000000fffffff5ffffffffffffffebffffffff",
            INIT_16 => X"ffffffd3fffffffffffffff0ffffffffffffffffffffffff0000000f00000000",
            INIT_17 => X"ffffffdeffffffffffffffe3ffffffffffffffddffffffffffffffeaffffffff",
            INIT_18 => X"fffffffefffffffffffffffaffffffffffffffc7ffffffffffffffe6ffffffff",
            INIT_19 => X"fffffffbffffffffffffffdeffffffff0000000100000000fffffffdffffffff",
            INIT_1A => X"ffffffe4ffffffffffffffd7fffffffffffffff2ffffffff0000001c00000000",
            INIT_1B => X"0000001700000000ffffffeaffffffff0000001e000000000000002400000000",
            INIT_1C => X"fffffffcffffffff0000000600000000ffffffdcfffffffffffffff7ffffffff",
            INIT_1D => X"0000000e00000000ffffff7cffffffffffffff88fffffffffffffff8ffffffff",
            INIT_1E => X"ffffff6bffffffffffffff5dffffffffffffff3affffffffffffff12ffffffff",
            INIT_1F => X"00000003000000000000001f00000000ffffff84ffffffffffffff38ffffffff",
            INIT_20 => X"000000010000000000000021000000000000001100000000fffffff8ffffffff",
            INIT_21 => X"ffffffcdffffffffffffffecfffffffffffffffeffffffffffffffedffffffff",
            INIT_22 => X"ffffffe5ffffffffffffffd1fffffffffffffff0fffffffffffffff5ffffffff",
            INIT_23 => X"0000001300000000ffffffeaffffffff0000000000000000fffffff9ffffffff",
            INIT_24 => X"ffffffe7fffffffffffffff6ffffffff0000002e000000000000003300000000",
            INIT_25 => X"000000330000000000000030000000000000001d000000000000001600000000",
            INIT_26 => X"0000001a00000000fffffff4ffffffff0000002f000000000000000b00000000",
            INIT_27 => X"0000001600000000ffffffdfffffffff00000001000000000000002900000000",
            INIT_28 => X"0000000f00000000fffffffafffffffffffffff4fffffffffffffff4ffffffff",
            INIT_29 => X"ffffffe9ffffffffffffffd0fffffffffffffffbffffffff0000001500000000",
            INIT_2A => X"ffffffffffffffffffffffd0ffffffffffffffc8fffffffffffffff9ffffffff",
            INIT_2B => X"0000000300000000fffffff9fffffffffffffffdffffffffffffffecffffffff",
            INIT_2C => X"0000000900000000ffffffdcffffffffffffffe5ffffffffffffffedffffffff",
            INIT_2D => X"fffffff6fffffffffffffff3ffffffffffffffecffffffffffffffdaffffffff",
            INIT_2E => X"ffffffebffffffffffffffd1ffffffff0000000700000000ffffffb0ffffffff",
            INIT_2F => X"ffffffe0ffffffffffffffe3ffffffffffffffe6ffffffff0000000100000000",
            INIT_30 => X"ffffffe5fffffffffffffff2fffffffffffffffeffffffffffffffeeffffffff",
            INIT_31 => X"ffffffb3ffffffffffffffceffffffff0000000100000000ffffffe7ffffffff",
            INIT_32 => X"ffffffc3ffffffffffffffaeffffffffffffffc4ffffffffffffffabffffffff",
            INIT_33 => X"ffffff52ffffffffffffffbeffffffffffffff8dffffffffffffff92ffffffff",
            INIT_34 => X"ffffff75ffffffffffffff83ffffffffffffffd6ffffffffffffffa2ffffffff",
            INIT_35 => X"ffffff90ffffffffffffff75ffffffffffffff94ffffffffffffffb4ffffffff",
            INIT_36 => X"ffffffcaffffffffffffffdfffffffffffffffd9ffffffffffffffd3ffffffff",
            INIT_37 => X"ffffffc7ffffffffffffffc2ffffffffffffffd6ffffffffffffffe5ffffffff",
            INIT_38 => X"000000010000000000000025000000000000002b00000000ffffffc4ffffffff",
            INIT_39 => X"00000014000000000000001f000000000000001f000000000000002700000000",
            INIT_3A => X"ffffffeeffffffff000000210000000000000001000000000000001700000000",
            INIT_3B => X"ffffffeafffffffffffffff9ffffffffffffffebffffffff0000001000000000",
            INIT_3C => X"0000000b000000000000000700000000ffffffe4fffffffffffffff1ffffffff",
            INIT_3D => X"0000000000000000000000070000000000000027000000000000001400000000",
            INIT_3E => X"ffffffffffffffff00000023000000000000001c000000000000000a00000000",
            INIT_3F => X"00000016000000000000000e000000000000003f00000000fffffffdffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003600000000000000280000000000000028000000000000004a00000000",
            INIT_41 => X"ffffffc0ffffffff0000001c00000000ffffffe9ffffffff0000003f00000000",
            INIT_42 => X"00000019000000000000000100000000ffffffecffffffffffffffcbffffffff",
            INIT_43 => X"0000000800000000ffffffdbffffffff0000000f000000000000000c00000000",
            INIT_44 => X"fffffffeffffffffffffffddffffffff00000000000000000000001000000000",
            INIT_45 => X"0000002600000000ffffffe5ffffffffffffffebffffffffffffffceffffffff",
            INIT_46 => X"000000650000000000000038000000000000000d000000000000001d00000000",
            INIT_47 => X"00000073000000000000007e000000000000004d000000000000006900000000",
            INIT_48 => X"fffffffcffffffff00000007000000000000002b000000000000002800000000",
            INIT_49 => X"ffffffe3ffffffffffffffeafffffffffffffffeffffffff0000001200000000",
            INIT_4A => X"ffffffb9ffffffffffffff8dffffffffffffffbeffffffffffffffd5ffffffff",
            INIT_4B => X"0000003600000000000000240000000000000020000000000000001900000000",
            INIT_4C => X"0000001900000000000000110000000000000046000000000000002d00000000",
            INIT_4D => X"fffffff1fffffffffffffff4ffffffff00000016000000000000000700000000",
            INIT_4E => X"ffffffc8fffffffffffffff0fffffffffffffff4ffffffffffffffdcffffffff",
            INIT_4F => X"0000001e000000000000000800000000ffffffe8ffffffffffffffbbffffffff",
            INIT_50 => X"000000250000000000000020000000000000001a00000000ffffffe6ffffffff",
            INIT_51 => X"0000000e0000000000000022000000000000001d000000000000004100000000",
            INIT_52 => X"fffffff0ffffffff0000002a000000000000001b000000000000001700000000",
            INIT_53 => X"000000200000000000000050000000000000003600000000ffffffcfffffffff",
            INIT_54 => X"ffffffd8fffffffffffffff8ffffffffffffffedffffffff0000001200000000",
            INIT_55 => X"00000048000000000000004f00000000ffffffd7ffffffffffffffaaffffffff",
            INIT_56 => X"0000000400000000ffffffe9ffffffffffffffecffffffff0000002300000000",
            INIT_57 => X"0000006200000000ffffffd9ffffffffffffffa2ffffffffffffffd0ffffffff",
            INIT_58 => X"0000001d0000000000000004000000000000004d000000000000007d00000000",
            INIT_59 => X"ffffffabffffffffffffff8effffffffffffffb7fffffffffffffffaffffffff",
            INIT_5A => X"0000001d00000000000000260000000000000032000000000000004200000000",
            INIT_5B => X"ffffffdaffffffffffffffbfffffffff0000001a000000000000001700000000",
            INIT_5C => X"fffffff6ffffffffffffffdaffffffffffffffe0ffffffffffffffeaffffffff",
            INIT_5D => X"0000000f00000000000000150000000000000016000000000000001300000000",
            INIT_5E => X"ffffffb7ffffffffffffffc0ffffffff00000024000000000000000400000000",
            INIT_5F => X"ffffffffffffffff00000010000000000000000e00000000ffffffc1ffffffff",
            INIT_60 => X"ffffffdbffffffff000000210000000000000029000000000000002a00000000",
            INIT_61 => X"0000000b00000000fffffff1ffffffffffffffb5ffffffffffffffa6ffffffff",
            INIT_62 => X"0000003100000000000000460000000000000041000000000000000700000000",
            INIT_63 => X"ffffffe8ffffffff0000001100000000fffffff7fffffffffffffffeffffffff",
            INIT_64 => X"ffffffd8fffffffffffffff9ffffffffffffffe1fffffffffffffff5ffffffff",
            INIT_65 => X"fffffff3ffffffff0000000b000000000000002500000000ffffffe5ffffffff",
            INIT_66 => X"0000002b00000000000000110000000000000015000000000000001600000000",
            INIT_67 => X"0000000400000000fffffffdfffffffffffffffeffffffff0000000000000000",
            INIT_68 => X"00000019000000000000001000000000fffffffaffffffff0000003300000000",
            INIT_69 => X"0000001900000000ffffffc3ffffffffffffffddffffffffffffffe2ffffffff",
            INIT_6A => X"0000000d00000000000000100000000000000028000000000000002f00000000",
            INIT_6B => X"ffffffc0ffffffffffffffcbffffffffffffffddffffffff0000000400000000",
            INIT_6C => X"fffffff8ffffffffffffffefffffffffffffffe9fffffffffffffffbffffffff",
            INIT_6D => X"ffffffe7ffffffffffffffcafffffffffffffffeffffffff0000000000000000",
            INIT_6E => X"ffffffdffffffffffffffff3ffffffff0000000a00000000ffffffdcffffffff",
            INIT_6F => X"0000002400000000000000060000000000000037000000000000001400000000",
            INIT_70 => X"0000002300000000fffffff2ffffffff00000025000000000000000300000000",
            INIT_71 => X"0000002e00000000fffffff3ffffffff00000001000000000000003600000000",
            INIT_72 => X"0000002300000000fffffff9ffffffff0000000200000000fffffff2ffffffff",
            INIT_73 => X"000000100000000000000000000000000000001a000000000000002a00000000",
            INIT_74 => X"0000000c00000000fffffffaffffffff00000014000000000000001600000000",
            INIT_75 => X"0000003600000000fffffffeffffffff00000013000000000000002e00000000",
            INIT_76 => X"0000002000000000000000060000000000000008000000000000000100000000",
            INIT_77 => X"ffffffe6ffffffffffffffe3ffffffffffffffdcfffffffffffffff5ffffffff",
            INIT_78 => X"fffffff1ffffffff0000000300000000ffffffefffffffffffffffecffffffff",
            INIT_79 => X"0000000f00000000fffffffbfffffffffffffff8fffffffffffffff7ffffffff",
            INIT_7A => X"00000013000000000000000a0000000000000001000000000000001000000000",
            INIT_7B => X"0000000b00000000000000380000000000000012000000000000002700000000",
            INIT_7C => X"0000005a000000000000006000000000ffffffe8ffffffff0000001f00000000",
            INIT_7D => X"00000049000000000000003a0000000000000042000000000000001f00000000",
            INIT_7E => X"0000002200000000fffffff4ffffffff00000017000000000000002100000000",
            INIT_7F => X"000000160000000000000026000000000000002c000000000000003d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE4;


    MEM_IWGHT_LAYER1_INSTANCE5 : if BRAM_NAME = "iwght_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000028000000000000000000000000ffffffe9ffffffff0000001a00000000",
            INIT_01 => X"ffffffe3ffffffff00000024000000000000000c00000000fffffff5ffffffff",
            INIT_02 => X"fffffff7ffffffff000000150000000000000004000000000000000e00000000",
            INIT_03 => X"ffffffc7ffffffff00000026000000000000001b00000000ffffffe9ffffffff",
            INIT_04 => X"0000001e00000000ffffffd8ffffffffffffffdbfffffffffffffff7ffffffff",
            INIT_05 => X"0000002b000000000000001f000000000000001c00000000fffffffdffffffff",
            INIT_06 => X"000000300000000000000013000000000000001d000000000000002800000000",
            INIT_07 => X"fffffff2ffffffff0000002300000000fffffffbffffffffffffffd1ffffffff",
            INIT_08 => X"ffffffd7ffffffffffffffdaffffffffffffffdcffffffffffffffe8ffffffff",
            INIT_09 => X"ffffffe5ffffffff0000001000000000fffffff1ffffffffffffffe3ffffffff",
            INIT_0A => X"0000002100000000000000080000000000000005000000000000002800000000",
            INIT_0B => X"0000001d00000000fffffff8fffffffffffffffcffffffff0000001100000000",
            INIT_0C => X"fffffff3ffffffffffffffefffffffff0000001a00000000ffffffeaffffffff",
            INIT_0D => X"ffffffc6ffffffffffffffe7fffffffffffffff0ffffffffffffffeaffffffff",
            INIT_0E => X"ffffffd3ffffffffffffffb5ffffffffffffffb8ffffffffffffffbeffffffff",
            INIT_0F => X"ffffffa8ffffffffffffffcaffffffffffffffd3ffffffffffffffcdffffffff",
            INIT_10 => X"0000003d0000000000000011000000000000002d000000000000003100000000",
            INIT_11 => X"0000003300000000000000190000000000000020000000000000003600000000",
            INIT_12 => X"00000052000000000000002d0000000000000045000000000000002100000000",
            INIT_13 => X"000000630000000000000000000000000000000f000000000000004300000000",
            INIT_14 => X"0000001100000000000000360000000000000015000000000000002500000000",
            INIT_15 => X"0000005700000000fffffff6ffffffff00000002000000000000001500000000",
            INIT_16 => X"ffffffe4ffffffff00000037000000000000002a000000000000000e00000000",
            INIT_17 => X"ffffff8bffffffffffffffa7ffffffffffffff96fffffffffffffff2ffffffff",
            INIT_18 => X"0000001800000000ffffffa8ffffffffffffffbfffffffffffffffa6ffffffff",
            INIT_19 => X"ffffffbbffffffff0000001200000000ffffffe3ffffffffffffffcbffffffff",
            INIT_1A => X"ffffffffffffffffffffffe6ffffffff0000002900000000ffffffe0ffffffff",
            INIT_1B => X"ffffffd7ffffffff0000000d00000000ffffffe7ffffffff0000001200000000",
            INIT_1C => X"ffffffcfffffffffffffffeaffffffff0000000400000000ffffffe1ffffffff",
            INIT_1D => X"ffffffbfffffffffffffffb7ffffffff0000000b00000000fffffffbffffffff",
            INIT_1E => X"0000000e00000000ffffffcaffffffffffffffe3ffffffffffffffb1ffffffff",
            INIT_1F => X"ffffffe2ffffffff000000030000000000000003000000000000000a00000000",
            INIT_20 => X"0000000a00000000fffffff4ffffffffffffffe7fffffffffffffffeffffffff",
            INIT_21 => X"00000021000000000000002900000000ffffffe9ffffffff0000002000000000",
            INIT_22 => X"fffffff1ffffffffffffffe6fffffffffffffff4ffffffffffffffe5ffffffff",
            INIT_23 => X"0000000a00000000ffffffdfffffffff0000000c000000000000001100000000",
            INIT_24 => X"ffffffcdffffffff0000000100000000fffffff0ffffffff0000003000000000",
            INIT_25 => X"ffffffbeffffffffffffffd2ffffffffffffffc8ffffffffffffffdbffffffff",
            INIT_26 => X"0000003d00000000ffffffcefffffffffffffffeffffffffffffffe1ffffffff",
            INIT_27 => X"0000001000000000fffffffaffffffff0000000f000000000000000600000000",
            INIT_28 => X"00000023000000000000003200000000fffffff5fffffffffffffffdffffffff",
            INIT_29 => X"ffffffd2ffffffff0000000f0000000000000027000000000000001b00000000",
            INIT_2A => X"fffffffaffffffffffffffefffffffff00000019000000000000000e00000000",
            INIT_2B => X"0000000400000000000000010000000000000008000000000000003c00000000",
            INIT_2C => X"0000003e00000000000000040000000000000020000000000000002c00000000",
            INIT_2D => X"0000002b00000000ffffffebffffffffffffffffffffffff0000001a00000000",
            INIT_2E => X"fffffff5ffffffff0000004900000000fffffffaffffffffffffffd9ffffffff",
            INIT_2F => X"0000002300000000000000090000000000000022000000000000003100000000",
            INIT_30 => X"000000220000000000000024000000000000000f00000000fffffff0ffffffff",
            INIT_31 => X"00000040000000000000002e00000000fffffff8ffffffffffffffe1ffffffff",
            INIT_32 => X"00000044000000000000004d000000000000003f000000000000005600000000",
            INIT_33 => X"000000300000000000000020000000000000002c000000000000004e00000000",
            INIT_34 => X"0000000f00000000ffffffe7fffffffffffffffaffffffff0000001c00000000",
            INIT_35 => X"00000020000000000000000b00000000fffffffcffffffff0000001500000000",
            INIT_36 => X"ffffffc9ffffffffffffffc4fffffffffffffff9ffffffffffffffedffffffff",
            INIT_37 => X"ffffffcbffffffffffffffdcffffffffffffffbaffffffffffffffa8ffffffff",
            INIT_38 => X"ffffffe4fffffffffffffff2ffffffffffffffcdffffffffffffffbdffffffff",
            INIT_39 => X"000000020000000000000000000000000000001b000000000000000e00000000",
            INIT_3A => X"fffffff5ffffffff000000090000000000000000000000000000000b00000000",
            INIT_3B => X"0000001f0000000000000016000000000000000300000000ffffffebffffffff",
            INIT_3C => X"fffffff5ffffffff000000080000000000000025000000000000000000000000",
            INIT_3D => X"ffffffe8fffffffffffffffbfffffffffffffffbffffffffffffffedffffffff",
            INIT_3E => X"0000001b00000000ffffffddffffffffffffffdeffffffffffffffebffffffff",
            INIT_3F => X"fffffffffffffffffffffffdffffffff00000019000000000000003500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001800000000000000090000000000000003000000000000001c00000000",
            INIT_41 => X"0000000f00000000fffffff9ffffffff00000026000000000000002900000000",
            INIT_42 => X"ffffffe7fffffffffffffff3ffffffff0000000b00000000ffffffe7ffffffff",
            INIT_43 => X"ffffffdeffffffffffffffeaffffffff00000015000000000000001900000000",
            INIT_44 => X"fffffff4ffffffffffffffd9ffffffffffffffc9fffffffffffffff5ffffffff",
            INIT_45 => X"ffffffccffffffffffffffb6ffffffffffffffd6ffffffffffffffe8ffffffff",
            INIT_46 => X"ffffffdeffffffffffffffffffffffff0000000a00000000fffffff8ffffffff",
            INIT_47 => X"ffffffe7fffffffffffffffdffffffff0000000700000000ffffffdbffffffff",
            INIT_48 => X"0000001200000000fffffff7ffffffff0000001900000000fffffff7ffffffff",
            INIT_49 => X"0000001000000000ffffffefffffffff00000011000000000000001300000000",
            INIT_4A => X"ffffffe4fffffffffffffffbffffffff00000017000000000000000700000000",
            INIT_4B => X"0000000900000000fffffffdffffffff0000000f00000000fffffffdffffffff",
            INIT_4C => X"ffffffddffffffff0000000700000000ffffffeeffffffff0000000400000000",
            INIT_4D => X"ffffffcefffffffffffffffaffffffffffffffe0ffffffffffffffd7ffffffff",
            INIT_4E => X"fffffff7fffffffffffffff9ffffffffffffffe4ffffffffffffffecffffffff",
            INIT_4F => X"0000001000000000fffffff0ffffffff0000001a00000000fffffffaffffffff",
            INIT_50 => X"0000002400000000ffffffe1ffffffffffffffe8ffffffff0000000a00000000",
            INIT_51 => X"ffffffc7ffffffffffffffc9ffffffffffffffc1ffffffff0000001700000000",
            INIT_52 => X"ffffffc6ffffffff0000000900000000ffffffb9ffffffffffffffcfffffffff",
            INIT_53 => X"00000016000000000000001c00000000ffffffcfffffffffffffffbcffffffff",
            INIT_54 => X"ffffffefffffffff00000019000000000000001e000000000000000f00000000",
            INIT_55 => X"ffffffe6ffffffff000000020000000000000001000000000000001e00000000",
            INIT_56 => X"00000004000000000000000a00000000ffffffe0ffffffff0000000600000000",
            INIT_57 => X"ffffffffffffffffffffffdffffffffffffffff2ffffffffffffffefffffffff",
            INIT_58 => X"0000001900000000000000190000000000000014000000000000000500000000",
            INIT_59 => X"0000003500000000fffffff2ffffffff00000012000000000000000200000000",
            INIT_5A => X"00000003000000000000000000000000ffffffecffffffff0000002200000000",
            INIT_5B => X"fffffff5ffffffff0000000a00000000ffffffd7ffffffffffffffd3ffffffff",
            INIT_5C => X"ffffffc2ffffffffffffffc0ffffffff0000000300000000ffffffebffffffff",
            INIT_5D => X"ffffffd1ffffffffffffffdfffffffffffffffd2fffffffffffffff7ffffffff",
            INIT_5E => X"ffffffdaffffffffffffffe6fffffffffffffff6ffffffff0000000500000000",
            INIT_5F => X"ffffffe4ffffffffffffffe3ffffffffffffffd2ffffffffffffffefffffffff",
            INIT_60 => X"fffffff4ffffffffffffffe9ffffffffffffffe6ffffffffffffffecffffffff",
            INIT_61 => X"fffffff8fffffffffffffff8ffffffff00000015000000000000002500000000",
            INIT_62 => X"fffffffafffffffffffffff6ffffffff0000002300000000fffffff9ffffffff",
            INIT_63 => X"000000140000000000000021000000000000000d000000000000000200000000",
            INIT_64 => X"0000002100000000fffffff1ffffffff0000000b00000000fffffffcffffffff",
            INIT_65 => X"ffffffe3ffffffffffffffedffffffff00000010000000000000000800000000",
            INIT_66 => X"ffffffe9ffffffffffffffcaffffffffffffffc5ffffffffffffffdfffffffff",
            INIT_67 => X"ffffffe9ffffffffffffffddfffffffffffffff3ffffffff0000001200000000",
            INIT_68 => X"ffffffe0ffffffffffffffe3ffffffffffffffd2fffffffffffffff7ffffffff",
            INIT_69 => X"ffffffe3ffffffffffffffdeffffffffffffffedffffffffffffffe6ffffffff",
            INIT_6A => X"0000000400000000fffffffbffffffff0000000f000000000000000f00000000",
            INIT_6B => X"fffffffbffffffff0000001b00000000fffffff1fffffffffffffff5ffffffff",
            INIT_6C => X"ffffffeeffffffff00000003000000000000001300000000ffffffe0ffffffff",
            INIT_6D => X"fffffff7ffffffff000000050000000000000006000000000000000600000000",
            INIT_6E => X"0000002300000000000000080000000000000002000000000000001500000000",
            INIT_6F => X"0000001a0000000000000019000000000000000e000000000000000100000000",
            INIT_70 => X"000000070000000000000031000000000000000c00000000fffffffeffffffff",
            INIT_71 => X"ffffffe3fffffffffffffff3ffffffff0000000800000000fffffffaffffffff",
            INIT_72 => X"ffffffdbffffffffffffffdafffffffffffffffdffffffffffffffd5ffffffff",
            INIT_73 => X"00000006000000000000003e000000000000002c000000000000000400000000",
            INIT_74 => X"000000350000000000000008000000000000003f000000000000000f00000000",
            INIT_75 => X"00000005000000000000000a00000000fffffff4ffffffff0000001600000000",
            INIT_76 => X"ffffffd0ffffffff0000000000000000ffffffdbfffffffffffffff5ffffffff",
            INIT_77 => X"ffffffddffffffffffffffe6ffffffff0000000b00000000ffffffefffffffff",
            INIT_78 => X"0000000800000000fffffff5ffffffff0000000b000000000000000e00000000",
            INIT_79 => X"0000000e00000000fffffff8ffffffffffffffe7ffffffff0000001d00000000",
            INIT_7A => X"0000001e0000000000000010000000000000002d000000000000003600000000",
            INIT_7B => X"0000001b000000000000002b0000000000000010000000000000003700000000",
            INIT_7C => X"000000170000000000000007000000000000000b00000000ffffffe4ffffffff",
            INIT_7D => X"fffffff0ffffffffffffffffffffffff00000019000000000000000800000000",
            INIT_7E => X"ffffffebffffffff000000000000000000000011000000000000000c00000000",
            INIT_7F => X"fffffffeffffffffffffffc5ffffffffffffffc5ffffffffffffffc3ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE5;


    MEM_IWGHT_LAYER1_INSTANCE6 : if BRAM_NAME = "iwght_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe7ffffffff0000000e00000000ffffffdbffffffffffffffd1ffffffff",
            INIT_01 => X"ffffffebfffffffffffffff5ffffffffffffffd7fffffffffffffff7ffffffff",
            INIT_02 => X"0000001b00000000fffffff0ffffffffffffffd7ffffffffffffffd3ffffffff",
            INIT_03 => X"ffffffdbffffffff000000080000000000000001000000000000001400000000",
            INIT_04 => X"0000000b000000000000000c00000000fffffff9ffffffffffffffe8ffffffff",
            INIT_05 => X"ffffffdaffffffffffffffefffffffffffffffd0ffffffffffffffedffffffff",
            INIT_06 => X"ffffffc1ffffffffffffffd8ffffffffffffffe5fffffffffffffff8ffffffff",
            INIT_07 => X"0000001c00000000ffffffeafffffffffffffff2ffffffff0000000b00000000",
            INIT_08 => X"0000002200000000000000280000000000000017000000000000001500000000",
            INIT_09 => X"0000000000000000ffffffe7ffffffff00000025000000000000000d00000000",
            INIT_0A => X"ffffffffffffffff0000001400000000ffffffe2ffffffff0000000400000000",
            INIT_0B => X"fffffff4ffffffff0000000a00000000fffffff4ffffffff0000000600000000",
            INIT_0C => X"fffffff0ffffffff0000000600000000ffffffe6ffffffffffffffd4ffffffff",
            INIT_0D => X"fffffff5ffffffffffffffe7ffffffffffffffe2ffffffffffffffe8ffffffff",
            INIT_0E => X"fffffff7ffffffff0000000100000000fffffffcffffffff0000003500000000",
            INIT_0F => X"ffffffceffffffff00000014000000000000000b00000000ffffffecffffffff",
            INIT_10 => X"000000060000000000000011000000000000001c00000000fffffffcffffffff",
            INIT_11 => X"fffffff3ffffffff00000009000000000000001800000000ffffffefffffffff",
            INIT_12 => X"00000009000000000000000e00000000ffffffecffffffff0000000800000000",
            INIT_13 => X"fffffff4fffffffffffffff6ffffffff00000028000000000000001b00000000",
            INIT_14 => X"fffffffbffffffffffffffffffffffffffffffedffffffff0000000d00000000",
            INIT_15 => X"00000000000000000000000000000000fffffff2fffffffffffffff8ffffffff",
            INIT_16 => X"ffffffcbffffffffffffffc4fffffffffffffff8ffffffffffffffbeffffffff",
            INIT_17 => X"fffffff6ffffffff0000001000000000fffffff0ffffffff0000000000000000",
            INIT_18 => X"000000280000000000000018000000000000000600000000fffffff7ffffffff",
            INIT_19 => X"ffffffcfffffffffffffffdcffffffffffffffd5ffffffff0000000700000000",
            INIT_1A => X"ffffffcbffffffffffffffd0fffffffffffffff0ffffffffffffffc2ffffffff",
            INIT_1B => X"0000000700000000fffffff1ffffffffffffffceffffffffffffffc9ffffffff",
            INIT_1C => X"fffffff9ffffffffffffffdcffffffffffffffe5ffffffff0000000800000000",
            INIT_1D => X"ffffffdcffffffffffffffd9fffffffffffffff8fffffffffffffffcffffffff",
            INIT_1E => X"fffffffeffffffffffffffedffffffff00000002000000000000000800000000",
            INIT_1F => X"0000000d000000000000001b000000000000000e000000000000002c00000000",
            INIT_20 => X"ffffffdeffffffffffffffdfffffffffffffffe1fffffffffffffff9ffffffff",
            INIT_21 => X"fffffff5ffffffff0000000400000000ffffffffffffffff0000001700000000",
            INIT_22 => X"ffffffe4ffffffff0000000600000000fffffff8ffffffff0000001700000000",
            INIT_23 => X"ffffffeaffffffffffffffeeffffffff0000001d00000000fffffff1ffffffff",
            INIT_24 => X"0000001f000000000000003700000000ffffffefffffffffffffffe9ffffffff",
            INIT_25 => X"fffffff3ffffffff0000000c000000000000000900000000ffffffe2ffffffff",
            INIT_26 => X"00000039000000000000000c0000000000000010000000000000000000000000",
            INIT_27 => X"0000001f000000000000000c0000000000000020000000000000001a00000000",
            INIT_28 => X"fffffffaffffffff0000001c000000000000002600000000fffffffbffffffff",
            INIT_29 => X"ffffffeffffffffffffffff3ffffffff0000000b000000000000001b00000000",
            INIT_2A => X"0000000a000000000000001400000000fffffff4fffffffffffffff2ffffffff",
            INIT_2B => X"ffffffdbfffffffffffffff1ffffffffffffffeefffffffffffffff7ffffffff",
            INIT_2C => X"ffffffe9ffffffffffffffd5ffffffffffffffc4ffffffffffffffdfffffffff",
            INIT_2D => X"ffffffccffffffff000000200000000000000005000000000000000100000000",
            INIT_2E => X"ffffffc0ffffffffffffffe1ffffffff0000000000000000ffffffd1ffffffff",
            INIT_2F => X"ffffffceffffffffffffffb7ffffffff0000001f000000000000000000000000",
            INIT_30 => X"ffffffa5ffffffffffffffd4ffffffffffffffbeffffffffffffffb9ffffffff",
            INIT_31 => X"0000003c0000000000000036000000000000003b000000000000000300000000",
            INIT_32 => X"0000000100000000fffffff1fffffffffffffff7ffffffffffffffe3ffffffff",
            INIT_33 => X"fffffffefffffffffffffff3fffffffffffffff1fffffffffffffff1ffffffff",
            INIT_34 => X"000000090000000000000030000000000000001a000000000000001c00000000",
            INIT_35 => X"ffffffedffffffff000000000000000000000027000000000000000b00000000",
            INIT_36 => X"00000010000000000000000a00000000fffffff2ffffffff0000000e00000000",
            INIT_37 => X"fffffff9ffffffff000000240000000000000035000000000000002600000000",
            INIT_38 => X"0000000a00000000fffffff8ffffffff0000001900000000ffffffe7ffffffff",
            INIT_39 => X"00000005000000000000000900000000ffffffe0ffffffffffffffecffffffff",
            INIT_3A => X"ffffffe6fffffffffffffff8fffffffffffffff2ffffffffffffffe4ffffffff",
            INIT_3B => X"0000000100000000ffffffdeffffffff0000000100000000fffffffaffffffff",
            INIT_3C => X"00000017000000000000000b00000000ffffffa7ffffffffffffffdbffffffff",
            INIT_3D => X"ffffffe8ffffffff00000003000000000000001500000000ffffffe0ffffffff",
            INIT_3E => X"0000001000000000fffffffdffffffff00000014000000000000001900000000",
            INIT_3F => X"fffffff2ffffffff0000001700000000fffffff2ffffffffffffffe7ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe3fffffffffffffff1fffffffffffffffdffffffff0000000100000000",
            INIT_41 => X"ffffff9dffffffff0000000e00000000fffffff0ffffffff0000001f00000000",
            INIT_42 => X"0000000600000000ffffffccffffffffffffffefffffffff0000000000000000",
            INIT_43 => X"fffffffdffffffff0000000600000000ffffffebfffffffffffffff0ffffffff",
            INIT_44 => X"fffffff4ffffffffffffffdfffffffff0000000700000000ffffffe2ffffffff",
            INIT_45 => X"00000017000000000000000b000000000000000b000000000000001300000000",
            INIT_46 => X"0000000400000000000000180000000000000030000000000000000d00000000",
            INIT_47 => X"0000000e000000000000000200000000ffffffdcfffffffffffffff4ffffffff",
            INIT_48 => X"0000000b000000000000002200000000ffffff8bfffffffffffffffaffffffff",
            INIT_49 => X"00000001000000000000002a000000000000005000000000fffffffeffffffff",
            INIT_4A => X"fffffff5ffffffff000000070000000000000039000000000000003b00000000",
            INIT_4B => X"ffffffeaffffffff0000001a00000000fffffff5ffffffffffffffeaffffffff",
            INIT_4C => X"000000190000000000000020000000000000002e00000000fffffffcffffffff",
            INIT_4D => X"fffffff0ffffffffffffffe4ffffffff0000001500000000ffffffddffffffff",
            INIT_4E => X"0000000d000000000000000500000000fffffffbffffffffffffffe0ffffffff",
            INIT_4F => X"0000002900000000000000130000000000000014000000000000000700000000",
            INIT_50 => X"fffffff6ffffffff00000056000000000000003c000000000000000800000000",
            INIT_51 => X"0000002d0000000000000042000000000000003e000000000000000700000000",
            INIT_52 => X"000000370000000000000060000000000000004c000000000000003300000000",
            INIT_53 => X"000000140000000000000057000000000000003e000000000000003d00000000",
            INIT_54 => X"0000004100000000000000450000000000000015000000000000004700000000",
            INIT_55 => X"0000001b000000000000002b0000000000000011000000000000006b00000000",
            INIT_56 => X"0000001500000000000000390000000000000024000000000000001f00000000",
            INIT_57 => X"fffffff9ffffffff0000001c0000000000000024000000000000000700000000",
            INIT_58 => X"fffffffffffffffffffffff1ffffffff00000018000000000000001500000000",
            INIT_59 => X"0000000600000000fffffffdffffffffffffffe2ffffffff0000000b00000000",
            INIT_5A => X"ffffffe3ffffffffffffffdfffffffff0000000500000000ffffffe7ffffffff",
            INIT_5B => X"0000000100000000ffffffb7ffffffffffffffc7fffffffffffffffdffffffff",
            INIT_5C => X"0000000a00000000fffffff4ffffffffffffffbfffffffffffffffe5ffffffff",
            INIT_5D => X"ffffffdfffffffff0000001000000000ffffffe6ffffffffffffffd2ffffffff",
            INIT_5E => X"ffffffc9ffffffff0000000e000000000000003a00000000ffffffa8ffffffff",
            INIT_5F => X"fffffffeffffffffffffffe5ffffffffffffffd9ffffffffffffffefffffffff",
            INIT_60 => X"ffffffe6ffffffffffffffdcffffffffffffffabffffffffffffffcaffffffff",
            INIT_61 => X"ffffffdcffffffffffffffdafffffffffffffff6ffffffffffffffccffffffff",
            INIT_62 => X"0000001f00000000ffffffe7ffffffff0000000300000000ffffffffffffffff",
            INIT_63 => X"00000005000000000000000900000000fffffffaffffffff0000001700000000",
            INIT_64 => X"00000023000000000000002000000000ffffffe0ffffffff0000001800000000",
            INIT_65 => X"ffffffbfffffffff00000008000000000000000d000000000000000100000000",
            INIT_66 => X"ffffffcafffffffffffffff9ffffffffffffffd8ffffffffffffffe3ffffffff",
            INIT_67 => X"ffffffdfffffffffffffffccffffffffffffffe3ffffffffffffffbeffffffff",
            INIT_68 => X"0000000300000000fffffffcfffffffffffffff7ffffffffffffffebffffffff",
            INIT_69 => X"fffffff9ffffffff0000001300000000fffffff9ffffffffffffffffffffffff",
            INIT_6A => X"0000001600000000fffffff2ffffffff00000034000000000000000000000000",
            INIT_6B => X"0000003600000000ffffffcafffffffffffffff1ffffffff0000002a00000000",
            INIT_6C => X"ffffffcaffffffff0000000600000000ffffffaaffffffff0000000300000000",
            INIT_6D => X"ffffffedffffffffffffffd5ffffffff0000002700000000ffffffb4ffffffff",
            INIT_6E => X"0000003300000000ffffffeeffffffffffffffefffffffff0000002e00000000",
            INIT_6F => X"0000002f000000000000006300000000ffffffc0ffffffff0000001a00000000",
            INIT_70 => X"00000002000000000000004e000000000000004000000000fffffff8ffffffff",
            INIT_71 => X"0000001900000000ffffffc9ffffffff0000001b000000000000003400000000",
            INIT_72 => X"0000002400000000ffffffbbffffffff00000004000000000000000600000000",
            INIT_73 => X"ffffffebffffffff00000023000000000000001d000000000000002e00000000",
            INIT_74 => X"000000090000000000000015000000000000000300000000ffffffefffffffff",
            INIT_75 => X"ffffffc5ffffffffffffffdfffffffff00000021000000000000000000000000",
            INIT_76 => X"0000000900000000ffffffa4ffffffffffffffeaffffffff0000004800000000",
            INIT_77 => X"ffffffedffffffffffffffe3ffffffffffffffb3ffffffff0000001100000000",
            INIT_78 => X"0000000200000000fffffff2ffffffff0000001e000000000000000a00000000",
            INIT_79 => X"0000000b000000000000001800000000fffffff3ffffffff0000001d00000000",
            INIT_7A => X"fffffff5ffffffff0000001900000000ffffffe2ffffffffffffffeaffffffff",
            INIT_7B => X"ffffffedffffffffffffffe6ffffffffffffffe7ffffffffffffffdbffffffff",
            INIT_7C => X"ffffffcaffffffffffffffe0ffffffff0000000200000000ffffffe7ffffffff",
            INIT_7D => X"0000003100000000ffffffb1ffffffffffffffe8ffffffff0000004300000000",
            INIT_7E => X"00000026000000000000000900000000ffffffc5ffffffff0000001f00000000",
            INIT_7F => X"0000003000000000000000130000000000000010000000000000002100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE6;


    MEM_IWGHT_LAYER1_INSTANCE7 : if BRAM_NAME = "iwght_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffffffffffff0000001800000000fffffffaffffffffffffffffffffffff",
            INIT_01 => X"ffffff9fffffffff0000003800000000fffffffdffffffffffffffe2ffffffff",
            INIT_02 => X"ffffffbefffffffffffffff4ffffffff0000005600000000fffffffeffffffff",
            INIT_03 => X"ffffffb3ffffffff0000000c00000000ffffffe3ffffffffffffffb9ffffffff",
            INIT_04 => X"ffffff85fffffffffffffff4fffffffffffffffcffffffffffffff5dffffffff",
            INIT_05 => X"ffffffc5ffffffffffffffe1ffffffff0000000200000000fffffff8ffffffff",
            INIT_06 => X"ffffffe6ffffffffffffffd1ffffffffffffffd3fffffffffffffff7ffffffff",
            INIT_07 => X"ffffffe4ffffffff0000001000000000ffffffecffffffff0000000e00000000",
            INIT_08 => X"ffffffdeffffffff00000016000000000000000900000000ffffffd6ffffffff",
            INIT_09 => X"0000001b00000000ffffffe6ffffffff0000001a000000000000001400000000",
            INIT_0A => X"0000002a00000000ffffffebffffffff00000013000000000000002f00000000",
            INIT_0B => X"00000059000000000000001f00000000ffffffcaffffffff0000005900000000",
            INIT_0C => X"0000000b000000000000001d00000000fffffff2ffffffffffffffe1ffffffff",
            INIT_0D => X"fffffffeffffffff0000002c0000000000000009000000000000001500000000",
            INIT_0E => X"ffffffc2ffffffffffffffeaffffffffffffffc8fffffffffffffff4ffffffff",
            INIT_0F => X"0000000600000000fffffff2fffffffffffffff4ffffffff0000001300000000",
            INIT_10 => X"ffffffecffffffff0000000c00000000ffffffd4ffffffffffffffdfffffffff",
            INIT_11 => X"0000000000000000ffffffe8ffffffff00000013000000000000001200000000",
            INIT_12 => X"00000007000000000000000700000000ffffffeeffffffff0000000100000000",
            INIT_13 => X"00000000000000000000000e0000000000000007000000000000000300000000",
            INIT_14 => X"0000001900000000000000180000000000000000000000000000001600000000",
            INIT_15 => X"0000007400000000000000290000000000000037000000000000005700000000",
            INIT_16 => X"0000005600000000000000360000000000000072000000000000008300000000",
            INIT_17 => X"fffffff6ffffffff0000000900000000fffffffaffffffff0000002f00000000",
            INIT_18 => X"fffffff3fffffffffffffff7fffffffffffffff2ffffffffffffffeeffffffff",
            INIT_19 => X"0000001300000000fffffff0fffffffffffffffdffffffff0000000600000000",
            INIT_1A => X"ffffffeeffffffff0000003300000000ffffffecffffffff0000000d00000000",
            INIT_1B => X"0000000f000000000000001b000000000000000a000000000000000c00000000",
            INIT_1C => X"0000001700000000ffffffeeffffffff0000001b000000000000001400000000",
            INIT_1D => X"ffffffdffffffffffffffff9ffffffffffffffd1ffffffffffffffe9ffffffff",
            INIT_1E => X"000000080000000000000038000000000000002e00000000fffffff8ffffffff",
            INIT_1F => X"fffffff4ffffffffffffffecffffffffffffffe5ffffffff0000002600000000",
            INIT_20 => X"ffffffddffffffff0000000800000000ffffffe5ffffffffffffffd6ffffffff",
            INIT_21 => X"0000000000000000fffffff4ffffffff0000000100000000ffffffe8ffffffff",
            INIT_22 => X"0000000f0000000000000022000000000000001f00000000fffffffaffffffff",
            INIT_23 => X"0000003a00000000000000390000000000000058000000000000002f00000000",
            INIT_24 => X"0000000f0000000000000020000000000000001a000000000000003600000000",
            INIT_25 => X"0000002700000000ffffffdffffffffffffffffbffffffff0000000e00000000",
            INIT_26 => X"ffffffd6fffffffffffffffdffffffffffffffe7ffffffffffffffd3ffffffff",
            INIT_27 => X"00000003000000000000000c00000000fffffff8ffffffff0000000000000000",
            INIT_28 => X"0000002b00000000000000010000000000000030000000000000000400000000",
            INIT_29 => X"000000310000000000000034000000000000001e000000000000002600000000",
            INIT_2A => X"0000003c0000000000000030000000000000002a000000000000002900000000",
            INIT_2B => X"ffffffe5ffffffff0000001e000000000000003f000000000000002f00000000",
            INIT_2C => X"ffffffefffffffffffffffedffffffff0000000400000000fffffff4ffffffff",
            INIT_2D => X"00000007000000000000001400000000fffffff9ffffffffffffffe8ffffffff",
            INIT_2E => X"ffffffd1ffffffff00000012000000000000001200000000ffffffd7ffffffff",
            INIT_2F => X"ffffffd3ffffffffffffffefffffffff0000000b000000000000000000000000",
            INIT_30 => X"ffffffcbffffffff000000060000000000000000000000000000000700000000",
            INIT_31 => X"ffffffc5ffffffffffffffd7ffffffffffffffdbffffffffffffffe5ffffffff",
            INIT_32 => X"00000004000000000000000600000000fffffff4fffffffffffffff1ffffffff",
            INIT_33 => X"0000004d00000000fffffffcffffffff0000001a000000000000001c00000000",
            INIT_34 => X"0000000d00000000ffffffe9ffffffff0000001e000000000000003500000000",
            INIT_35 => X"ffffffe3ffffffffffffffe0ffffffff0000001100000000fffffffcffffffff",
            INIT_36 => X"0000001f00000000000000030000000000000001000000000000001b00000000",
            INIT_37 => X"ffffffffffffffff0000001400000000ffffffddffffffffffffffe5ffffffff",
            INIT_38 => X"000000190000000000000013000000000000000c000000000000001600000000",
            INIT_39 => X"fffffff7ffffffff0000001c000000000000002a000000000000000c00000000",
            INIT_3A => X"fffffffcffffffff000000210000000000000008000000000000003100000000",
            INIT_3B => X"00000003000000000000000000000000ffffffc9ffffffff0000002200000000",
            INIT_3C => X"ffffffafffffffffffffffd0ffffffffffffffaeffffffffffffffc3ffffffff",
            INIT_3D => X"0000000000000000fffffff9ffffffffffffffa5ffffffffffffffd1ffffffff",
            INIT_3E => X"ffffffe9ffffffffffffffbbffffffffffffffdcfffffffffffffff9ffffffff",
            INIT_3F => X"fffffff1ffffffffffffffc0ffffffffffffffe2fffffffffffffff3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffff9bffffffffffffff96ffffffff0000005d000000000000002300000000",
            INIT_41 => X"ffffffb1ffffffffffffffd2ffffffffffffffaafffffffffffffff8ffffffff",
            INIT_42 => X"ffffffd8ffffffff0000000a00000000fffffffeffffffffffffffe9ffffffff",
            INIT_43 => X"0000000700000000ffffffcdffffffff0000002400000000ffffffe0ffffffff",
            INIT_44 => X"fffffffbffffffff0000000f000000000000000a00000000ffffffdcffffffff",
            INIT_45 => X"000000140000000000000016000000000000000200000000fffffffcffffffff",
            INIT_46 => X"0000000a000000000000001c00000000ffffffe9fffffffffffffff4ffffffff",
            INIT_47 => X"0000003a00000000000000040000000000000005000000000000000800000000",
            INIT_48 => X"fffffffdffffffff0000000c00000000ffffffdffffffffffffffffeffffffff",
            INIT_49 => X"ffffffffffffffff0000001c0000000000000028000000000000000b00000000",
            INIT_4A => X"0000003600000000000000250000000000000045000000000000004000000000",
            INIT_4B => X"fffffffbffffffffffffffedfffffffffffffff9fffffffffffffff5ffffffff",
            INIT_4C => X"ffffffd6ffffffffffffffefffffffffffffffeffffffffffffffff8ffffffff",
            INIT_4D => X"0000000300000000ffffffffffffffff0000001d000000000000000100000000",
            INIT_4E => X"0000000400000000000000190000000000000033000000000000000400000000",
            INIT_4F => X"ffffffe9fffffffffffffff6ffffffff0000002b000000000000001c00000000",
            INIT_50 => X"ffffffd5ffffffffffffffd9ffffffffffffffcdffffffff0000001b00000000",
            INIT_51 => X"ffffffecffffffffffffffc4fffffffffffffff4ffffffffffffffe8ffffffff",
            INIT_52 => X"0000001500000000fffffff5ffffffff00000019000000000000001500000000",
            INIT_53 => X"0000000000000000fffffffafffffffffffffff4ffffffff0000003300000000",
            INIT_54 => X"0000001b00000000ffffffe8fffffffffffffff6fffffffffffffff8ffffffff",
            INIT_55 => X"00000022000000000000002b00000000fffffffcfffffffffffffff8ffffffff",
            INIT_56 => X"ffffffecffffffff000000030000000000000006000000000000003700000000",
            INIT_57 => X"0000001000000000ffffffe8fffffffffffffff5ffffffff0000000d00000000",
            INIT_58 => X"0000000900000000000000040000000000000017000000000000000e00000000",
            INIT_59 => X"fffffff1ffffffffffffffe6fffffffffffffffafffffffffffffffdffffffff",
            INIT_5A => X"00000026000000000000000f00000000ffffffefffffffff0000000a00000000",
            INIT_5B => X"000000080000000000000012000000000000001400000000fffffffeffffffff",
            INIT_5C => X"fffffff6ffffffff0000001d000000000000000d000000000000001200000000",
            INIT_5D => X"fffffff7ffffffff0000002300000000ffffffecffffffff0000000000000000",
            INIT_5E => X"00000032000000000000002f0000000000000019000000000000000900000000",
            INIT_5F => X"ffffffe0fffffffffffffff0ffffffff00000017000000000000004500000000",
            INIT_60 => X"000000370000000000000007000000000000003f000000000000003e00000000",
            INIT_61 => X"fffffff0fffffffffffffff4ffffffff00000030000000000000003800000000",
            INIT_62 => X"0000001500000000ffffffc5ffffffffffffffe5fffffffffffffff7ffffffff",
            INIT_63 => X"0000000d000000000000002d00000000ffffffc6ffffffffffffffd0ffffffff",
            INIT_64 => X"ffffffcfffffffffffffffe8ffffffffffffffbcffffffff0000000100000000",
            INIT_65 => X"fffffff1ffffffffffffffc4ffffffffffffffc3ffffffffffffffd7ffffffff",
            INIT_66 => X"fffffff1fffffffffffffff2fffffffffffffff3ffffffff0000002f00000000",
            INIT_67 => X"ffffffebffffffffffffffc2ffffffffffffffe9ffffffff0000003200000000",
            INIT_68 => X"00000009000000000000000e00000000ffffffecffffffffffffffe6ffffffff",
            INIT_69 => X"0000002c000000000000000100000000fffffff3ffffffff0000003100000000",
            INIT_6A => X"ffffffdbffffffffffffffe4ffffffff0000002300000000fffffff6ffffffff",
            INIT_6B => X"ffffffcfffffffff0000000000000000ffffffccffffffff0000002100000000",
            INIT_6C => X"fffffff3fffffffffffffff9ffffffffffffffe3ffffffffffffffc8ffffffff",
            INIT_6D => X"ffffffdaffffffff000000030000000000000000000000000000000f00000000",
            INIT_6E => X"0000001000000000ffffffe0fffffffffffffffbffffffff0000000a00000000",
            INIT_6F => X"ffffffcdffffffffffffffeaffffffffffffffb0ffffffffffffffa8ffffffff",
            INIT_70 => X"ffffffe8ffffffffffffffc2ffffffff0000000f00000000ffffffc3ffffffff",
            INIT_71 => X"0000002d000000000000001800000000fffffff9ffffffff0000000500000000",
            INIT_72 => X"0000002400000000fffffff9ffffffffffffffe6ffffffffffffffedffffffff",
            INIT_73 => X"fffffffbffffffff0000001a0000000000000037000000000000001600000000",
            INIT_74 => X"0000000700000000000000040000000000000021000000000000001000000000",
            INIT_75 => X"ffffffd0ffffffff0000000a0000000000000003000000000000001c00000000",
            INIT_76 => X"ffffffe4ffffffffffffffbdffffffffffffffeeffffffffffffffe4ffffffff",
            INIT_77 => X"ffffffe3ffffffff0000003400000000fffffff0ffffffffffffffbcffffffff",
            INIT_78 => X"0000001200000000ffffffddffffffff00000009000000000000000c00000000",
            INIT_79 => X"ffffffe2ffffffff0000000700000000ffffffe8ffffffffffffffeaffffffff",
            INIT_7A => X"000000430000000000000003000000000000001400000000ffffffe4ffffffff",
            INIT_7B => X"00000000000000000000003c0000000000000001000000000000002000000000",
            INIT_7C => X"ffffffedffffffff00000000000000000000003900000000fffffffbffffffff",
            INIT_7D => X"00000026000000000000000300000000ffffffd5ffffffff0000001f00000000",
            INIT_7E => X"0000002a000000000000001e000000000000002100000000fffffffbffffffff",
            INIT_7F => X"ffffffb1ffffffff0000000e00000000ffffffd4ffffffffffffffe8ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE7;


    MEM_IWGHT_LAYER1_INSTANCE8 : if BRAM_NAME = "iwght_layer1_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001c00000000ffffffe2fffffffffffffffdffffffff0000001d00000000",
            INIT_01 => X"ffffffbaffffffff0000000900000000ffffffdbffffffffffffff9affffffff",
            INIT_02 => X"fffffffbfffffffffffffff6ffffffffffffffe7fffffffffffffff4ffffffff",
            INIT_03 => X"fffffffbffffffff0000001e00000000fffffffdffffffffffffffe2ffffffff",
            INIT_04 => X"ffffffe7ffffffffffffffe6ffffffff0000000000000000fffffff1ffffffff",
            INIT_05 => X"0000002300000000ffffffddfffffffffffffff5fffffffffffffffbffffffff",
            INIT_06 => X"00000053000000000000003200000000ffffffe6ffffffff0000004600000000",
            INIT_07 => X"000000160000000000000034000000000000001f000000000000001600000000",
            INIT_08 => X"ffffffd5ffffffff0000002900000000fffffff1ffffffff0000001800000000",
            INIT_09 => X"0000000000000000ffffffecffffffff0000001600000000ffffffd1ffffffff",
            INIT_0A => X"0000002000000000ffffffb6fffffffffffffff9ffffffff0000001d00000000",
            INIT_0B => X"ffffffaaffffffffffffffe0ffffffffffffffb7ffffffffffffffa8ffffffff",
            INIT_0C => X"0000000100000000ffffffdfffffffffffffffe7ffffffffffffffa4ffffffff",
            INIT_0D => X"ffffffd6ffffffff0000001800000000ffffffe0ffffffffffffffdbffffffff",
            INIT_0E => X"00000007000000000000002f000000000000003b00000000ffffffe4ffffffff",
            INIT_0F => X"ffffff8effffffffffffffb9ffffffff0000005d00000000ffffffa7ffffffff",
            INIT_10 => X"ffffffdeffffffffffffffc2ffffffffffffff85ffffffff0000002100000000",
            INIT_11 => X"0000001900000000fffffff9ffffffff00000037000000000000001600000000",
            INIT_12 => X"0000002a00000000000000310000000000000005000000000000002800000000",
            INIT_13 => X"ffffffddffffffff0000001e000000000000002100000000ffffffd7ffffffff",
            INIT_14 => X"0000004300000000fffffff8ffffffff0000005a000000000000003c00000000",
            INIT_15 => X"0000003f000000000000002400000000fffffff3ffffffff0000005400000000",
            INIT_16 => X"ffffffe4ffffffff00000030000000000000001c00000000ffffffeeffffffff",
            INIT_17 => X"ffffffffffffffff0000001100000000fffffff9ffffffff0000001d00000000",
            INIT_18 => X"fffffff7ffffffffffffffe0fffffffffffffffeffffffff0000000800000000",
            INIT_19 => X"000000130000000000000017000000000000000800000000ffffffebffffffff",
            INIT_1A => X"ffffffd7ffffffff0000002300000000ffffffb5ffffffff0000000a00000000",
            INIT_1B => X"ffffffb8ffffffffffffffc0fffffffffffffffaffffffffffffffd0ffffffff",
            INIT_1C => X"0000000200000000fffffff1ffffffffffffffd2ffffffff0000000f00000000",
            INIT_1D => X"0000001900000000ffffffe8ffffffff0000000000000000ffffffe9ffffffff",
            INIT_1E => X"fffffff4ffffffffffffffecffffffffffffffecffffffff0000000a00000000",
            INIT_1F => X"0000001200000000fffffff3fffffffffffffffcffffffff0000002700000000",
            INIT_20 => X"fffffff5ffffffffffffffe8ffffffff0000000400000000fffffffdffffffff",
            INIT_21 => X"0000001e00000000fffffff2ffffffff0000001b000000000000000d00000000",
            INIT_22 => X"0000001d00000000000000240000000000000017000000000000003700000000",
            INIT_23 => X"00000012000000000000001000000000ffffffd8fffffffffffffffcffffffff",
            INIT_24 => X"0000000a00000000000000390000000000000017000000000000001800000000",
            INIT_25 => X"fffffffdffffffff0000001b0000000000000031000000000000003900000000",
            INIT_26 => X"000000520000000000000023000000000000003c000000000000004000000000",
            INIT_27 => X"ffffffecffffffff0000001d0000000000000007000000000000004700000000",
            INIT_28 => X"0000000400000000000000190000000000000001000000000000001e00000000",
            INIT_29 => X"ffffffe2ffffffffffffffe4ffffffff00000022000000000000002300000000",
            INIT_2A => X"ffffffeeffffffffffffffd6ffffffff00000015000000000000001000000000",
            INIT_2B => X"0000002700000000ffffffb3fffffffffffffff2fffffffffffffff8ffffffff",
            INIT_2C => X"0000000a000000000000002a0000000000000047000000000000001a00000000",
            INIT_2D => X"0000001a00000000fffffffbfffffffffffffff4ffffffff0000004800000000",
            INIT_2E => X"ffffffc3ffffffff0000000d00000000ffffffe8ffffffffffffffd6ffffffff",
            INIT_2F => X"ffffff9cffffffffffffffb1ffffffffffffffb3ffffffffffffffbeffffffff",
            INIT_30 => X"ffffffe1ffffffffffffffe8fffffffffffffffeffffffffffffffe0ffffffff",
            INIT_31 => X"0000002a00000000fffffff6fffffffffffffffcffffffff0000002100000000",
            INIT_32 => X"ffffffe6ffffffffffffffc0ffffffff00000012000000000000003100000000",
            INIT_33 => X"ffffff84ffffffffffffff6bffffffffffffff82ffffffffffffffc6ffffffff",
            INIT_34 => X"ffffffe5ffffffffffffff6affffffffffffff53ffffffffffffff67ffffffff",
            INIT_35 => X"00000002000000000000000100000000ffffffecffffffffffffffe1ffffffff",
            INIT_36 => X"000000320000000000000015000000000000001a00000000ffffffebffffffff",
            INIT_37 => X"ffffffc6ffffffff0000000000000000ffffffddffffffffffffffd8ffffffff",
            INIT_38 => X"ffffff9dffffffffffffffefffffffffffffff8dffffffffffffffa4ffffffff",
            INIT_39 => X"fffffffeffffffff00000001000000000000000e00000000ffffffabffffffff",
            INIT_3A => X"000000180000000000000023000000000000003d000000000000000500000000",
            INIT_3B => X"ffffffeeffffffff0000000e0000000000000035000000000000002f00000000",
            INIT_3C => X"fffffff2ffffffff000000100000000000000022000000000000000600000000",
            INIT_3D => X"0000000b000000000000000c0000000000000022000000000000000000000000",
            INIT_3E => X"0000002b00000000ffffffccfffffffffffffff1ffffffff0000003400000000",
            INIT_3F => X"ffffffeeffffffffffffffe0ffffffffffffffcdffffffff0000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff1ffffffff0000000f000000000000000000000000ffffffeeffffffff",
            INIT_41 => X"00000020000000000000000000000000ffffffe8fffffffffffffffeffffffff",
            INIT_42 => X"ffffffa8ffffffffffffffdfffffffffffffffd2ffffffff0000001a00000000",
            INIT_43 => X"ffffffe3fffffffffffffff2fffffffffffffff0ffffffffffffffd1ffffffff",
            INIT_44 => X"ffffffdbffffffffffffffd4ffffffffffffffeffffffffffffffff2ffffffff",
            INIT_45 => X"ffffffddffffffffffffffeeffffffffffffffdbffffffffffffffd0ffffffff",
            INIT_46 => X"ffffffedffffffff0000000000000000ffffffedfffffffffffffff3ffffffff",
            INIT_47 => X"ffffffe9ffffffffffffffdeffffffffffffffddffffffffffffffc0ffffffff",
            INIT_48 => X"fffffffdffffffffffffffeeffffffffffffffd8fffffffffffffff1ffffffff",
            INIT_49 => X"00000016000000000000000c000000000000000900000000ffffffffffffffff",
            INIT_4A => X"0000000d000000000000000b0000000000000004000000000000000000000000",
            INIT_4B => X"0000001a000000000000000900000000fffffff4ffffffff0000002200000000",
            INIT_4C => X"00000007000000000000000d00000000ffffffffffffffff0000001200000000",
            INIT_4D => X"ffffffe2ffffffff00000011000000000000001d000000000000002100000000",
            INIT_4E => X"fffffffbffffffff0000000c00000000fffffff5ffffffffffffffeeffffffff",
            INIT_4F => X"fffffff8ffffffff000000070000000000000015000000000000001a00000000",
            INIT_50 => X"fffffff7ffffffff00000006000000000000001900000000ffffffe2ffffffff",
            INIT_51 => X"ffffffddffffffffffffffefffffffffffffffdfffffffffffffffeaffffffff",
            INIT_52 => X"fffffff3ffffffffffffffe9ffffffff0000000d00000000fffffff5ffffffff",
            INIT_53 => X"fffffff8ffffffffffffffe7fffffffffffffff8ffffffffffffffeeffffffff",
            INIT_54 => X"ffffffe8ffffffffffffffecffffffffffffffeeffffffffffffffecffffffff",
            INIT_55 => X"fffffff6ffffffff000000200000000000000006000000000000000700000000",
            INIT_56 => X"fffffffeffffffffffffffe0ffffffff00000013000000000000002200000000",
            INIT_57 => X"ffffffe7ffffffff0000000e00000000ffffffe1ffffffffffffffe6ffffffff",
            INIT_58 => X"ffffffd6fffffffffffffffdffffffffffffffe7fffffffffffffff8ffffffff",
            INIT_59 => X"ffffffebffffffffffffffe6ffffffffffffffbdffffffffffffffc2ffffffff",
            INIT_5A => X"0000000e000000000000000200000000ffffffc7ffffffffffffffffffffffff",
            INIT_5B => X"0000002c000000000000000e0000000000000037000000000000001400000000",
            INIT_5C => X"0000000600000000000000340000000000000019000000000000002800000000",
            INIT_5D => X"fffffff2fffffffffffffff9fffffffffffffffeffffffff0000000d00000000",
            INIT_5E => X"ffffffd7fffffffffffffff9ffffffffffffffecffffffffffffffebffffffff",
            INIT_5F => X"00000004000000000000000500000000fffffff8ffffffff0000000900000000",
            INIT_60 => X"ffffffffffffffffffffffe9ffffffff0000000d00000000fffffff7ffffffff",
            INIT_61 => X"00000028000000000000000b000000000000000e000000000000001c00000000",
            INIT_62 => X"0000001d00000000000000260000000000000017000000000000001900000000",
            INIT_63 => X"fffffff0fffffffffffffffcffffffff0000002200000000fffffff5ffffffff",
            INIT_64 => X"fffffffbffffffffffffffe3ffffffffffffffecfffffffffffffff9ffffffff",
            INIT_65 => X"ffffffb2ffffffffffffffcfffffffffffffffefffffffffffffffe2ffffffff",
            INIT_66 => X"fffffff6ffffffffffffffeefffffffffffffff4ffffffffffffffc3ffffffff",
            INIT_67 => X"0000003d000000000000001400000000fffffff4ffffffff0000000100000000",
            INIT_68 => X"ffffffdfffffffff0000000f00000000ffffffefffffffff0000001200000000",
            INIT_69 => X"0000001600000000ffffffddffffffffffffffdcffffffff0000001700000000",
            INIT_6A => X"00000015000000000000001b000000000000000600000000ffffffe5ffffffff",
            INIT_6B => X"ffffffebfffffffffffffffcffffffff00000011000000000000000f00000000",
            INIT_6C => X"0000002800000000000000060000000000000017000000000000000e00000000",
            INIT_6D => X"ffffffc3ffffffffffffffadffffffffffffffeffffffffffffffff3ffffffff",
            INIT_6E => X"0000000500000000ffffffe0ffffffffffffffd2ffffffffffffffeeffffffff",
            INIT_6F => X"0000000200000000fffffff9fffffffffffffff3ffffffffffffffe8ffffffff",
            INIT_70 => X"ffffff88fffffffffffffffeffffffffffffffe9ffffffffffffffbdffffffff",
            INIT_71 => X"fffffffcffffffffffffffd4ffffffffffffffbaffffffffffffffd2ffffffff",
            INIT_72 => X"0000000000000000ffffffcdffffffffffffffd2ffffffff0000000200000000",
            INIT_73 => X"ffffffe2fffffffffffffffcffffffffffffffccfffffffffffffff1ffffffff",
            INIT_74 => X"ffffffbdffffffffffffffb1ffffffff00000039000000000000002900000000",
            INIT_75 => X"ffffffe1ffffffffffffffc9ffffffffffffffc0ffffffffffffffdbffffffff",
            INIT_76 => X"ffffffc5fffffffffffffffaffffffffffffffe1ffffffffffffffdeffffffff",
            INIT_77 => X"ffffffbdffffffffffffffccffffffffffffffe2ffffffffffffffcdffffffff",
            INIT_78 => X"00000020000000000000002000000000ffffffeeffffffffffffffedffffffff",
            INIT_79 => X"00000000000000000000001300000000ffffffedffffffff0000001a00000000",
            INIT_7A => X"0000000600000000fffffff9ffffffff0000000200000000fffffff1ffffffff",
            INIT_7B => X"fffffffbffffffffffffffedffffffffffffffe4ffffffff0000001300000000",
            INIT_7C => X"0000001f000000000000000b000000000000000000000000fffffff2ffffffff",
            INIT_7D => X"000000010000000000000017000000000000002900000000ffffffe1ffffffff",
            INIT_7E => X"0000001500000000000000160000000000000013000000000000002c00000000",
            INIT_7F => X"00000009000000000000001600000000fffffff3ffffffff0000000d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE8;


    MEM_IWGHT_LAYER1_INSTANCE9 : if BRAM_NAME = "iwght_layer1_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000017000000000000000f0000000000000001000000000000001a00000000",
            INIT_01 => X"ffffffadffffffffffffffedffffffff00000005000000000000002700000000",
            INIT_02 => X"0000001100000000fffffff2ffffffff0000000d00000000fffffffdffffffff",
            INIT_03 => X"0000001600000000000000190000000000000019000000000000001a00000000",
            INIT_04 => X"fffffff8ffffffff0000000c00000000ffffffd7ffffffff0000002400000000",
            INIT_05 => X"0000002300000000fffffff0fffffffffffffff8ffffffffffffffbeffffffff",
            INIT_06 => X"00000017000000000000002d00000000ffffffd3ffffffff0000000f00000000",
            INIT_07 => X"000000130000000000000003000000000000002c000000000000003b00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER1_INSTANCE9;


    MEM_IWGHT_LAYER2_INSTANCE0 : if BRAM_NAME = "iwght_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffb98fffffffffffff23efffffffffffff546ffffffffffffd97fffffffff",
            INIT_01 => X"fffffa16ffffffff000010170000000000004a5700000000fffff88dffffffff",
            INIT_02 => X"0000417100000000000021850000000000000a320000000000000ea500000000",
            INIT_03 => X"00001a1000000000fffff2beffffffffffffda53ffffffff0000027700000000",
            INIT_04 => X"00000d1f00000000fffff3efffffffff000044f200000000000041b400000000",
            INIT_05 => X"ffffed1bffffffff00000aed0000000000002f1d000000000000130500000000",
            INIT_06 => X"fffff844ffffffffffffd00fffffffff00002f0600000000fffffb1bffffffff",
            INIT_07 => X"00002a6e00000000fffff25effffffff00001b8c00000000fffffa92ffffffff",
            INIT_08 => X"0000172900000000000026570000000000004eda0000000000001aee00000000",
            INIT_09 => X"000005d900000000ffffd5f5ffffffff00001e3d00000000000022b700000000",
            INIT_0A => X"0000091d00000000ffffe848ffffffff0000136100000000ffffed40ffffffff",
            INIT_0B => X"fffff0afffffffff00001eef00000000fffff538ffffffffffffd2aaffffffff",
            INIT_0C => X"fffffaefffffffff0000227f0000000000002c7a0000000000000be800000000",
            INIT_0D => X"fffff967fffffffffffffec7ffffffff00002c6e000000000000175600000000",
            INIT_0E => X"000025710000000000002da400000000000018cc0000000000000ac300000000",
            INIT_0F => X"00002be40000000000001e3c00000000ffffe100ffffffff0000380e00000000",
            INIT_10 => X"0000000600000000fffffff4ffffffff0000000a00000000ffffffedffffffff",
            INIT_11 => X"ffffffffffffffff00000019000000000000000000000000ffffffebffffffff",
            INIT_12 => X"0000001f00000000fffffff0fffffffffffffff3ffffffff0000001000000000",
            INIT_13 => X"ffffffe6ffffffff0000001d000000000000000b00000000fffffffbffffffff",
            INIT_14 => X"0000002a000000000000002700000000ffffffe0fffffffffffffffaffffffff",
            INIT_15 => X"00000034000000000000008f0000000000000028000000000000002d00000000",
            INIT_16 => X"0000001400000000000000230000000000000064000000000000002800000000",
            INIT_17 => X"0000000b00000000fffffff6fffffffffffffffeffffffff0000003800000000",
            INIT_18 => X"ffffffd6ffffffffffffffd6ffffffff0000000600000000fffffff9ffffffff",
            INIT_19 => X"000000540000000000000043000000000000003f000000000000001100000000",
            INIT_1A => X"00000060000000000000003a0000000000000045000000000000008d00000000",
            INIT_1B => X"ffffffe6ffffffff0000001a0000000000000000000000000000000700000000",
            INIT_1C => X"000000240000000000000000000000000000000f000000000000001900000000",
            INIT_1D => X"0000000000000000fffffffeffffffff00000011000000000000001f00000000",
            INIT_1E => X"0000002100000000fffffffcffffffffffffffd3ffffffff0000001b00000000",
            INIT_1F => X"0000000000000000fffffffeffffffffffffffecffffffffffffffd8ffffffff",
            INIT_20 => X"fffffff0ffffffffffffffddffffffffffffffecfffffffffffffffeffffffff",
            INIT_21 => X"fffffff2ffffffffffffffdffffffffffffffff7ffffffffffffffd8ffffffff",
            INIT_22 => X"fffffffdffffffff000000180000000000000003000000000000002000000000",
            INIT_23 => X"ffffffeeffffffff00000002000000000000003b000000000000001200000000",
            INIT_24 => X"00000009000000000000001a00000000fffffff4fffffffffffffff4ffffffff",
            INIT_25 => X"fffffff8ffffffff0000000400000000fffffffefffffffffffffffcffffffff",
            INIT_26 => X"0000002600000000ffffffe5ffffffff0000000500000000fffffffaffffffff",
            INIT_27 => X"fffffffcffffffff0000000d00000000fffffffcffffffff0000001100000000",
            INIT_28 => X"0000000800000000ffffffeaffffffffffffffd8ffffffffffffffe8ffffffff",
            INIT_29 => X"fffffffaffffffff0000000700000000ffffffdcfffffffffffffffbffffffff",
            INIT_2A => X"00000003000000000000000900000000ffffffc8ffffffffffffffdcffffffff",
            INIT_2B => X"0000000700000000000000020000000000000011000000000000000f00000000",
            INIT_2C => X"0000000e000000000000000b00000000fffffffdffffffffffffffefffffffff",
            INIT_2D => X"00000025000000000000000f0000000000000010000000000000002200000000",
            INIT_2E => X"00000000000000000000001500000000fffffff7ffffffffffffffe3ffffffff",
            INIT_2F => X"fffffff8ffffffff00000000000000000000000400000000fffffffaffffffff",
            INIT_30 => X"000000100000000000000015000000000000001000000000ffffffcbffffffff",
            INIT_31 => X"00000010000000000000000a0000000000000024000000000000000200000000",
            INIT_32 => X"ffffffcffffffffffffffff7ffffffffffffffd9ffffffff0000000300000000",
            INIT_33 => X"fffffff1ffffffffffffffe9ffffffff0000000100000000fffffff0ffffffff",
            INIT_34 => X"fffffff5ffffffff0000000e0000000000000009000000000000001100000000",
            INIT_35 => X"fffffff0ffffffff000000010000000000000037000000000000001100000000",
            INIT_36 => X"000000130000000000000020000000000000000700000000ffffffdfffffffff",
            INIT_37 => X"ffffffe5ffffffff0000000c00000000fffffff3fffffffffffffffdffffffff",
            INIT_38 => X"ffffffd2ffffffffffffffbdffffffff0000000000000000ffffffe7ffffffff",
            INIT_39 => X"ffffffd7ffffffffffffffb7ffffffffffffffffffffffffffffffc6ffffffff",
            INIT_3A => X"ffffffeeffffffffffffffdfffffffffffffff91ffffffffffffffd4ffffffff",
            INIT_3B => X"0000000100000000fffffff4fffffffffffffff9ffffffff0000000800000000",
            INIT_3C => X"000000120000000000000000000000000000002200000000fffffffaffffffff",
            INIT_3D => X"fffffff4ffffffffffffffd8fffffffffffffff7ffffffffffffffe5ffffffff",
            INIT_3E => X"fffffff0ffffffff0000000200000000fffffff2ffffffffffffffdeffffffff",
            INIT_3F => X"ffffffe4fffffffffffffff6ffffffff0000000900000000fffffffcffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001000000000fffffff6ffffffffffffffffffffffff0000001100000000",
            INIT_41 => X"0000000500000000fffffff8ffffffff00000018000000000000000100000000",
            INIT_42 => X"0000000200000000fffffff0fffffffffffffff0fffffffffffffff5ffffffff",
            INIT_43 => X"0000000100000000ffffffefffffffffffffffebffffffff0000000200000000",
            INIT_44 => X"00000007000000000000000c000000000000000200000000fffffff7ffffffff",
            INIT_45 => X"0000001a00000000ffffffe3fffffffffffffff8ffffffff0000002c00000000",
            INIT_46 => X"0000000d00000000ffffffedffffffff00000010000000000000000700000000",
            INIT_47 => X"ffffffe6ffffffff0000001300000000ffffffc7ffffffff0000000600000000",
            INIT_48 => X"00000030000000000000000e000000000000000d00000000ffffff98ffffffff",
            INIT_49 => X"fffffff6ffffffff00000011000000000000001200000000fffffffbffffffff",
            INIT_4A => X"ffffffeeffffffff000000030000000000000004000000000000000800000000",
            INIT_4B => X"0000001a00000000fffffffeffffffff0000001d000000000000002200000000",
            INIT_4C => X"0000000a00000000ffffffdcffffffffffffffe3ffffffffffffffffffffffff",
            INIT_4D => X"0000000000000000ffffffe8ffffffff0000001600000000fffffffcffffffff",
            INIT_4E => X"0000002100000000ffffffeeffffffff00000008000000000000001b00000000",
            INIT_4F => X"0000001000000000000000020000000000000019000000000000001900000000",
            INIT_50 => X"ffffffedffffffffffffffd5ffffffff00000012000000000000001500000000",
            INIT_51 => X"0000001400000000ffffffe0ffffffff0000001c00000000ffffffdbffffffff",
            INIT_52 => X"ffffffe7fffffffffffffffafffffffffffffffcfffffffffffffff5ffffffff",
            INIT_53 => X"0000000400000000ffffffebfffffffffffffffbffffffff0000000e00000000",
            INIT_54 => X"00000016000000000000000300000000ffffffe9ffffffff0000000200000000",
            INIT_55 => X"ffffffffffffffff00000019000000000000001400000000ffffffffffffffff",
            INIT_56 => X"0000001d0000000000000006000000000000001000000000ffffffebffffffff",
            INIT_57 => X"ffffffe8ffffffffffffffccfffffffffffffffdffffffff0000000400000000",
            INIT_58 => X"0000001e00000000000000120000000000000001000000000000000000000000",
            INIT_59 => X"000000000000000000000023000000000000000200000000fffffff0ffffffff",
            INIT_5A => X"ffffffdeffffffffffffffc6ffffffffffffffddfffffffffffffffdffffffff",
            INIT_5B => X"000000250000000000000005000000000000000000000000ffffffd7ffffffff",
            INIT_5C => X"ffffffe2ffffffff00000011000000000000002c000000000000006e00000000",
            INIT_5D => X"ffffffebffffffff00000026000000000000002400000000ffffffceffffffff",
            INIT_5E => X"fffffff6ffffffff00000043000000000000002a000000000000006900000000",
            INIT_5F => X"ffffff9bffffffff0000000900000000ffffffaffffffffffffffff6ffffffff",
            INIT_60 => X"0000003b000000000000001c00000000fffffff3ffffffff0000000000000000",
            INIT_61 => X"00000014000000000000000700000000fffffff1fffffffffffffff7ffffffff",
            INIT_62 => X"00000046000000000000003f000000000000003e000000000000003900000000",
            INIT_63 => X"ffffffe5ffffffff0000000700000000fffffff1ffffffff0000002200000000",
            INIT_64 => X"ffffffbbfffffffffffffffeffffffff0000005100000000fffffff5ffffffff",
            INIT_65 => X"00000021000000000000000200000000ffffffedffffffffffffffbeffffffff",
            INIT_66 => X"ffffffddfffffffffffffffdffffffffffffffeaffffffff0000003300000000",
            INIT_67 => X"0000001000000000ffffffeaffffffffffffffb4ffffffffffffffb2ffffffff",
            INIT_68 => X"ffffffc6ffffffffffffffd0ffffffff00000003000000000000000200000000",
            INIT_69 => X"00000011000000000000000c000000000000001900000000ffffffbfffffffff",
            INIT_6A => X"fffffff8fffffffffffffff2fffffffffffffffeffffffffffffffecffffffff",
            INIT_6B => X"0000002000000000000000000000000000000014000000000000001200000000",
            INIT_6C => X"0000000400000000000000220000000000000034000000000000001400000000",
            INIT_6D => X"0000001800000000000000080000000000000022000000000000001300000000",
            INIT_6E => X"0000000900000000ffffffedffffffffffffffd7fffffffffffffff5ffffffff",
            INIT_6F => X"000000200000000000000029000000000000001200000000fffffff2ffffffff",
            INIT_70 => X"ffffffffffffffffffffffdcffffffff00000021000000000000001f00000000",
            INIT_71 => X"00000036000000000000005400000000ffffffe2ffffffff0000000300000000",
            INIT_72 => X"fffffffaffffffffffffffe1ffffffff0000002300000000ffffffdaffffffff",
            INIT_73 => X"0000000600000000ffffffdafffffffffffffffcffffffff0000001100000000",
            INIT_74 => X"ffffffcfffffffffffffffbaffffffffffffffd0ffffffff0000000300000000",
            INIT_75 => X"0000000e0000000000000043000000000000003900000000ffffffc1ffffffff",
            INIT_76 => X"0000001200000000ffffffe4ffffffffffffffddffffffffffffffd9ffffffff",
            INIT_77 => X"ffffffefffffffffffffffdcffffffff00000038000000000000002500000000",
            INIT_78 => X"00000018000000000000003e000000000000002500000000ffffffd5ffffffff",
            INIT_79 => X"0000001900000000ffffffc6ffffffffffffffcdffffffffffffffccffffffff",
            INIT_7A => X"0000000400000000000000050000000000000018000000000000001f00000000",
            INIT_7B => X"ffffff8effffffffffffff97ffffffffffffffd9fffffffffffffffeffffffff",
            INIT_7C => X"ffffffefffffffff000000420000000000000031000000000000003400000000",
            INIT_7D => X"0000002a000000000000000500000000fffffff4ffffffff0000000c00000000",
            INIT_7E => X"0000000d00000000000000330000000000000030000000000000001700000000",
            INIT_7F => X"ffffffe2ffffffff00000005000000000000001e000000000000002300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE0;


    MEM_IWGHT_LAYER2_INSTANCE1 : if BRAM_NAME = "iwght_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000230000000000000004000000000000000500000000fffffffdffffffff",
            INIT_01 => X"00000010000000000000004d000000000000000700000000ffffffe7ffffffff",
            INIT_02 => X"0000000500000000fffffff7ffffffff0000001d00000000fffffffaffffffff",
            INIT_03 => X"0000002200000000fffffff9fffffffffffffffcffffffff0000000400000000",
            INIT_04 => X"ffffffe5ffffffffffffffe0fffffffffffffff2fffffffffffffffdffffffff",
            INIT_05 => X"0000001d0000000000000003000000000000001a00000000fffffffeffffffff",
            INIT_06 => X"fffffff7ffffffff00000000000000000000000d000000000000000800000000",
            INIT_07 => X"000000100000000000000004000000000000001b00000000ffffffe0ffffffff",
            INIT_08 => X"ffffffe6ffffffff00000000000000000000001f000000000000000900000000",
            INIT_09 => X"fffffffeffffffff0000000700000000ffffffe3ffffffffffffffd2ffffffff",
            INIT_0A => X"00000007000000000000000d00000000fffffff7fffffffffffffff0ffffffff",
            INIT_0B => X"ffffffdaffffffffffffffddfffffffffffffff0ffffffffffffffd4ffffffff",
            INIT_0C => X"000000490000000000000031000000000000000000000000fffffffeffffffff",
            INIT_0D => X"ffffffd8ffffffffffffffdcffffffffffffffe7ffffffff0000002300000000",
            INIT_0E => X"0000002800000000fffffff1ffffffffffffffb6ffffffffffffffdeffffffff",
            INIT_0F => X"ffffffd3ffffffff0000004d00000000ffffffc7ffffffffffffffadffffffff",
            INIT_10 => X"fffffff6ffffffffffffffdeffffffffffffffeaffffffffffffffccffffffff",
            INIT_11 => X"0000001400000000ffffffefffffffffffffffceffffffffffffffe0ffffffff",
            INIT_12 => X"0000003800000000000000300000000000000031000000000000002400000000",
            INIT_13 => X"00000020000000000000002a0000000000000013000000000000001600000000",
            INIT_14 => X"ffffffeeffffffffffffffc3fffffffffffffff3ffffffff0000001100000000",
            INIT_15 => X"0000002400000000ffffffcefffffffffffffff6ffffffff0000001500000000",
            INIT_16 => X"ffffffeeffffffffffffffbbffffffff00000000000000000000001400000000",
            INIT_17 => X"fffffff1ffffffffffffffbbffffffff0000000400000000fffffffbffffffff",
            INIT_18 => X"00000026000000000000000e000000000000000100000000ffffffedffffffff",
            INIT_19 => X"00000005000000000000000000000000ffffffffffffffff0000003b00000000",
            INIT_1A => X"fffffffaffffffffffffffc2ffffffff0000001a00000000ffffffb7ffffffff",
            INIT_1B => X"fffffff3ffffffff0000000300000000ffffffd9ffffffffffffffdaffffffff",
            INIT_1C => X"ffffffeeffffffffffffffe4ffffffff0000000800000000ffffffe4ffffffff",
            INIT_1D => X"00000032000000000000001800000000ffffffe9ffffffffffffffe1ffffffff",
            INIT_1E => X"0000001300000000ffffffeffffffffffffffff7ffffffff0000001300000000",
            INIT_1F => X"ffffffddffffffffffffffe6ffffffffffffffe6fffffffffffffffbffffffff",
            INIT_20 => X"fffffff2ffffffff000000140000000000000022000000000000001100000000",
            INIT_21 => X"0000000000000000fffffff9ffffffff0000000700000000ffffffeeffffffff",
            INIT_22 => X"0000000800000000fffffff6ffffffff0000000200000000fffffff8ffffffff",
            INIT_23 => X"0000001c00000000ffffffb3ffffffffffffffdffffffffffffffff5ffffffff",
            INIT_24 => X"ffffffeeffffffffffffffe9ffffffffffffffe5ffffffff0000001900000000",
            INIT_25 => X"ffffffefffffffffffffffd9ffffffffffffffc7fffffffffffffffdffffffff",
            INIT_26 => X"0000000d000000000000000b000000000000000f00000000fffffffcffffffff",
            INIT_27 => X"0000001f0000000000000059000000000000001d000000000000001f00000000",
            INIT_28 => X"000000190000000000000035000000000000000e000000000000003c00000000",
            INIT_29 => X"ffffffeeffffffffffffffd9ffffffffffffffd3ffffffffffffffc5ffffffff",
            INIT_2A => X"fffffff3ffffffff00000006000000000000000100000000ffffffc4ffffffff",
            INIT_2B => X"0000000d000000000000000a00000000fffffffcffffffff0000002500000000",
            INIT_2C => X"fffffff4ffffffff0000000a0000000000000026000000000000000600000000",
            INIT_2D => X"fffffffffffffffffffffffdffffffff0000001e000000000000000c00000000",
            INIT_2E => X"00000004000000000000000600000000ffffffd9fffffffffffffff5ffffffff",
            INIT_2F => X"0000003500000000ffffffeaffffffffffffffdcffffffffffffffddffffffff",
            INIT_30 => X"ffffffe4ffffffff000000000000000000000018000000000000001a00000000",
            INIT_31 => X"ffffffeffffffffffffffff1ffffffff0000000f00000000ffffffcaffffffff",
            INIT_32 => X"0000000d00000000ffffffd2ffffffff0000002200000000ffffffe7ffffffff",
            INIT_33 => X"00000010000000000000003700000000fffffffbffffffff0000000000000000",
            INIT_34 => X"00000038000000000000003100000000ffffffffffffffffffffffe0ffffffff",
            INIT_35 => X"ffffffcfffffffff0000002e000000000000001900000000ffffffd6ffffffff",
            INIT_36 => X"fffffffcffffffff0000001c000000000000002800000000ffffffe2ffffffff",
            INIT_37 => X"ffffffe3ffffffff0000001e000000000000001f00000000fffffffbffffffff",
            INIT_38 => X"0000001900000000ffffffe3fffffffffffffffcfffffffffffffffdffffffff",
            INIT_39 => X"0000002600000000fffffffcffffffff0000000f00000000fffffff8ffffffff",
            INIT_3A => X"0000002c000000000000002400000000ffffffe9ffffffff0000001100000000",
            INIT_3B => X"ffffffeaffffffff0000001300000000ffffffe8fffffffffffffff3ffffffff",
            INIT_3C => X"0000000c00000000ffffffe7ffffffff0000000f000000000000000200000000",
            INIT_3D => X"000000380000000000000007000000000000001d000000000000001600000000",
            INIT_3E => X"0000001b00000000ffffffd8ffffffffffffffd8ffffffffffffffd6ffffffff",
            INIT_3F => X"fffffffdffffffff0000000f000000000000000200000000fffffffcffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffeafffffffffffffffeffffffff0000000800000000ffffffd4ffffffff",
            INIT_41 => X"ffffffd2ffffffff0000000500000000fffffff4ffffffffffffffceffffffff",
            INIT_42 => X"0000000400000000ffffffcfffffffff0000003600000000ffffffecffffffff",
            INIT_43 => X"0000002c00000000ffffffceffffffffffffffc8ffffffff0000003800000000",
            INIT_44 => X"0000002300000000fffffff6fffffffffffffff0ffffffff0000002d00000000",
            INIT_45 => X"00000007000000000000003100000000ffffffcfffffffffffffffd4ffffffff",
            INIT_46 => X"0000003c0000000000000001000000000000000a00000000fffffff0ffffffff",
            INIT_47 => X"ffffffc6ffffffff00000028000000000000000800000000ffffffe5ffffffff",
            INIT_48 => X"ffffffc9ffffffff00000006000000000000002400000000ffffffe5ffffffff",
            INIT_49 => X"0000001f0000000000000000000000000000001f00000000ffffffddffffffff",
            INIT_4A => X"0000000100000000fffffff8ffffffffffffffe6fffffffffffffff4ffffffff",
            INIT_4B => X"00000011000000000000001800000000ffffffe6ffffffffffffffffffffffff",
            INIT_4C => X"0000000900000000fffffffbfffffffffffffff6ffffffff0000000000000000",
            INIT_4D => X"0000000f00000000ffffffe9ffffffffffffffe6ffffffff0000001f00000000",
            INIT_4E => X"00000004000000000000000b000000000000000d000000000000001000000000",
            INIT_4F => X"ffffffe8fffffffffffffffeffffffff0000002400000000fffffffaffffffff",
            INIT_50 => X"fffffff2ffffffff0000000700000000fffffff6ffffffff0000002300000000",
            INIT_51 => X"0000001d00000000fffffff3ffffffff00000002000000000000000000000000",
            INIT_52 => X"0000002200000000fffffffaffffffffffffffd8ffffffff0000003100000000",
            INIT_53 => X"00000000000000000000001f00000000ffffffccffffffffffffffc9ffffffff",
            INIT_54 => X"00000014000000000000001600000000ffffffb7fffffffffffffff3ffffffff",
            INIT_55 => X"ffffffcbffffffff0000000300000000fffffff8ffffffffffffffeeffffffff",
            INIT_56 => X"0000001b000000000000000d000000000000003200000000ffffffebffffffff",
            INIT_57 => X"0000003600000000000000260000000000000022000000000000002700000000",
            INIT_58 => X"ffffffe0ffffffffffffffebffffffff00000003000000000000003000000000",
            INIT_59 => X"0000003700000000ffffffb7ffffffffffffffe8fffffffffffffffdffffffff",
            INIT_5A => X"ffffffffffffffffffffffdcffffffffffffffe3ffffffff0000001d00000000",
            INIT_5B => X"0000002300000000ffffffd9ffffffffffffffc3ffffffff0000002300000000",
            INIT_5C => X"ffffffe4ffffffff0000002000000000ffffffedffffffffffffffbeffffffff",
            INIT_5D => X"fffffffcffffffffffffffe9ffffffff0000002d000000000000002e00000000",
            INIT_5E => X"0000002c00000000ffffffe8ffffffffffffffe5ffffffff0000003000000000",
            INIT_5F => X"0000000f000000000000001f0000000000000017000000000000000200000000",
            INIT_60 => X"0000004400000000000000250000000000000049000000000000003e00000000",
            INIT_61 => X"0000001c000000000000001300000000fffffff8ffffffff0000002c00000000",
            INIT_62 => X"ffffffd8ffffffff00000035000000000000000f00000000ffffffdcffffffff",
            INIT_63 => X"fffffffcffffffff0000000500000000fffffffcffffffffffffffe3ffffffff",
            INIT_64 => X"0000001a0000000000000013000000000000003000000000ffffffcaffffffff",
            INIT_65 => X"ffffffebffffffff00000006000000000000001b000000000000001200000000",
            INIT_66 => X"ffffffffffffffffffffffbfffffffff0000002900000000fffffff4ffffffff",
            INIT_67 => X"0000003e000000000000000300000000ffffffc0ffffffff0000000e00000000",
            INIT_68 => X"000000030000000000000000000000000000000000000000fffffffdffffffff",
            INIT_69 => X"ffffffeeffffffff0000000c00000000fffffffbfffffffffffffffdffffffff",
            INIT_6A => X"0000000a00000000ffffffe4fffffffffffffff0ffffffff0000000800000000",
            INIT_6B => X"fffffff6fffffffffffffff3fffffffffffffff8ffffffffffffffeaffffffff",
            INIT_6C => X"ffffffedffffffff0000000600000000fffffff3ffffffffffffffeaffffffff",
            INIT_6D => X"fffffff6fffffffffffffff4ffffffffffffffe7ffffffff0000000b00000000",
            INIT_6E => X"fffffff0ffffffff00000000000000000000000e00000000fffffff6ffffffff",
            INIT_6F => X"ffffffe8fffffffffffffff0fffffffffffffff5ffffffff0000000800000000",
            INIT_70 => X"fffffffdffffffff0000000500000000ffffffebffffffff0000000d00000000",
            INIT_71 => X"000000000000000000000005000000000000000000000000ffffffecffffffff",
            INIT_72 => X"ffffffeeffffffff0000000300000000fffffff6fffffffffffffffaffffffff",
            INIT_73 => X"fffffff4ffffffff0000000700000000fffffff1ffffffffffffffedffffffff",
            INIT_74 => X"00000011000000000000000200000000fffffffbffffffff0000000000000000",
            INIT_75 => X"fffffff4fffffffffffffffbfffffffffffffff6ffffffff0000000600000000",
            INIT_76 => X"fffffff3fffffffffffffff7fffffffffffffff0fffffffffffffff3ffffffff",
            INIT_77 => X"0000000d00000000fffffffdfffffffffffffffdffffffff0000000600000000",
            INIT_78 => X"ffffffeeffffffff000000070000000000000005000000000000000a00000000",
            INIT_79 => X"0000000000000000ffffffddffffffffffffffebffffffff0000000000000000",
            INIT_7A => X"00000009000000000000000200000000ffffffe7ffffffff0000000c00000000",
            INIT_7B => X"ffffffecfffffffffffffff9ffffffff00000007000000000000000400000000",
            INIT_7C => X"ffffffffffffffff0000000800000000ffffffedfffffffffffffffcffffffff",
            INIT_7D => X"fffffff9fffffffffffffff7ffffffff00000002000000000000000200000000",
            INIT_7E => X"0000000f00000000ffffffebfffffffffffffffffffffffffffffffcffffffff",
            INIT_7F => X"000000100000000000000000000000000000000300000000fffffff2ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE1;


    MEM_IWGHT_LAYER2_INSTANCE2 : if BRAM_NAME = "iwght_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffebffffffffffffffdffffffffffffffffaffffffffffffffeaffffffff",
            INIT_01 => X"0000000700000000fffffff8ffffffff0000001100000000fffffff8ffffffff",
            INIT_02 => X"0000000800000000fffffffcfffffffffffffff2ffffffff0000000400000000",
            INIT_03 => X"fffffff4ffffffff0000000500000000fffffff8ffffffff0000000500000000",
            INIT_04 => X"fffffff4ffffffff0000000200000000ffffffebffffffff0000000000000000",
            INIT_05 => X"ffffffe2fffffffffffffffdffffffffffffffe1fffffffffffffffcffffffff",
            INIT_06 => X"0000000000000000fffffff2ffffffff0000000b000000000000000a00000000",
            INIT_07 => X"ffffffeeffffffff00000001000000000000000000000000fffffffdffffffff",
            INIT_08 => X"00000012000000000000000800000000ffffffeefffffffffffffff9ffffffff",
            INIT_09 => X"fffffff8fffffffffffffff5ffffffff0000000b000000000000000700000000",
            INIT_0A => X"00000005000000000000000300000000fffffff1ffffffffffffffecffffffff",
            INIT_0B => X"fffffff5fffffffffffffffbfffffffffffffffbfffffffffffffff2ffffffff",
            INIT_0C => X"fffffff7ffffffff0000000000000000fffffff0ffffffff0000000b00000000",
            INIT_0D => X"0000000000000000fffffffbffffffffffffffffffffffffffffffe8ffffffff",
            INIT_0E => X"ffffffecffffffff0000000600000000ffffffffffffffffffffffedffffffff",
            INIT_0F => X"ffffffe7ffffffffffffffe9ffffffffffffffefffffffffffffffebffffffff",
            INIT_10 => X"0000000000000000fffffff4fffffffffffffffafffffffffffffffdffffffff",
            INIT_11 => X"fffffff2ffffffff0000000a00000000fffffff6fffffffffffffffeffffffff",
            INIT_12 => X"ffffffeafffffffffffffff8fffffffffffffff4fffffffffffffff5ffffffff",
            INIT_13 => X"0000000000000000fffffff1fffffffffffffffeffffffff0000000c00000000",
            INIT_14 => X"ffffffebfffffffffffffff4ffffffffffffffe7fffffffffffffff0ffffffff",
            INIT_15 => X"fffffff9ffffffffffffffedffffffff0000000f00000000ffffffecffffffff",
            INIT_16 => X"fffffff3fffffffffffffffbffffffffffffffebfffffffffffffffbffffffff",
            INIT_17 => X"00000004000000000000000300000000fffffff4ffffffffffffffedffffffff",
            INIT_18 => X"ffffffeeffffffff0000000700000000fffffffaffffffff0000000100000000",
            INIT_19 => X"0000000c00000000fffffffefffffffffffffff2ffffffff0000000b00000000",
            INIT_1A => X"ffffffebffffffff0000000000000000ffffffe9ffffffff0000000500000000",
            INIT_1B => X"0000000400000000fffffffcffffffffffffffe7fffffffffffffff8ffffffff",
            INIT_1C => X"0000000000000000ffffffeafffffffffffffffcffffffff0000000300000000",
            INIT_1D => X"ffffffedfffffffffffffff2ffffffff0000000300000000fffffff8ffffffff",
            INIT_1E => X"ffffffeaffffffffffffffffffffffff0000000500000000ffffffeaffffffff",
            INIT_1F => X"0000000000000000fffffffcffffffff0000000500000000ffffffe8ffffffff",
            INIT_20 => X"0000000100000000fffffff0ffffffffffffffeeffffffffffffffe0ffffffff",
            INIT_21 => X"fffffff0fffffffffffffff6ffffffff0000000900000000fffffff3ffffffff",
            INIT_22 => X"0000000200000000fffffffbffffffffffffffedffffffff0000000900000000",
            INIT_23 => X"0000000100000000000000000000000000000011000000000000000400000000",
            INIT_24 => X"0000000b00000000ffffffecffffffff00000005000000000000000000000000",
            INIT_25 => X"00000008000000000000001000000000ffffffeaffffffff0000000b00000000",
            INIT_26 => X"ffffffe8fffffffffffffff6ffffffff0000000200000000ffffffecffffffff",
            INIT_27 => X"fffffff0fffffffffffffffefffffffffffffff2ffffffffffffffeaffffffff",
            INIT_28 => X"fffffff5fffffffffffffff1fffffffffffffff1fffffffffffffff9ffffffff",
            INIT_29 => X"00000007000000000000000700000000fffffff6ffffffff0000000900000000",
            INIT_2A => X"00000001000000000000000b000000000000000b00000000ffffffedffffffff",
            INIT_2B => X"fffffff6ffffffff0000000900000000fffffff1fffffffffffffffaffffffff",
            INIT_2C => X"0000000d000000000000000800000000fffffffaffffffff0000000600000000",
            INIT_2D => X"fffffff3fffffffffffffff4fffffffffffffffbffffffff0000000900000000",
            INIT_2E => X"00000012000000000000000400000000ffffffe3ffffffffffffffefffffffff",
            INIT_2F => X"fffffff0ffffffff0000000800000000fffffff7fffffffffffffff3ffffffff",
            INIT_30 => X"fffffffbffffffff00000017000000000000001b000000000000000900000000",
            INIT_31 => X"00000001000000000000000c000000000000000100000000fffffff6ffffffff",
            INIT_32 => X"ffffffe3ffffffffffffffd5ffffffffffffffe3fffffffffffffffcffffffff",
            INIT_33 => X"ffffffe6fffffffffffffffaffffffff0000003e000000000000001200000000",
            INIT_34 => X"ffffffd6ffffffffffffffb6fffffffffffffff3ffffffffffffffeeffffffff",
            INIT_35 => X"ffffffd9fffffffffffffff7ffffffff0000000c00000000ffffffeaffffffff",
            INIT_36 => X"ffffffe6ffffffff00000007000000000000001e000000000000001100000000",
            INIT_37 => X"ffffffbeffffffffffffffe4ffffffff0000003200000000ffffffceffffffff",
            INIT_38 => X"ffffffc2ffffffffffffffe4ffffffffffffffdfffffffffffffffd5ffffffff",
            INIT_39 => X"0000000a00000000ffffffcdffffffffffffffceffffffffffffffd0ffffffff",
            INIT_3A => X"ffffffd6fffffffffffffff8ffffffffffffffd0ffffffffffffffd1ffffffff",
            INIT_3B => X"ffffffd3ffffffffffffffc3ffffffffffffffc3ffffffffffffffe5ffffffff",
            INIT_3C => X"fffffffeffffffffffffffe9ffffffffffffffeaffffffffffffffbfffffffff",
            INIT_3D => X"0000002500000000000000230000000000000016000000000000001600000000",
            INIT_3E => X"fffffffbffffffff0000000f000000000000001b000000000000003100000000",
            INIT_3F => X"ffffffffffffffff00000036000000000000001c000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff7ffffffffffffffe1ffffffff00000018000000000000001600000000",
            INIT_41 => X"fffffff2ffffffff0000001f000000000000000e00000000ffffffedffffffff",
            INIT_42 => X"0000002b00000000fffffff6ffffffff00000008000000000000000700000000",
            INIT_43 => X"0000000e000000000000000300000000fffffff1ffffffff0000001100000000",
            INIT_44 => X"fffffff0ffffffffffffffc3fffffffffffffff9ffffffff0000002400000000",
            INIT_45 => X"ffffffd7ffffffffffffffabffffffffffffffcfffffffffffffffb6ffffffff",
            INIT_46 => X"000000030000000000000009000000000000000f00000000ffffffdeffffffff",
            INIT_47 => X"0000000e000000000000003a0000000000000028000000000000000000000000",
            INIT_48 => X"ffffffe9ffffffff0000001d000000000000000f00000000fffffffaffffffff",
            INIT_49 => X"0000002400000000fffffff4ffffffff00000001000000000000001400000000",
            INIT_4A => X"ffffffdcffffffffffffffeefffffffffffffffdfffffffffffffff0ffffffff",
            INIT_4B => X"fffffff4fffffffffffffff7ffffffff0000001a000000000000001600000000",
            INIT_4C => X"ffffffe0fffffffffffffff5ffffffff0000000000000000ffffffdeffffffff",
            INIT_4D => X"0000001c000000000000003800000000fffffff3ffffffffffffffdfffffffff",
            INIT_4E => X"ffffffb2ffffffffffffffaaffffffffffffffcfffffffffffffffb5ffffffff",
            INIT_4F => X"0000000000000000ffffffeaffffffffffffffe2ffffffffffffffebffffffff",
            INIT_50 => X"fffffff2fffffffffffffffaffffffffffffffffffffffff0000000000000000",
            INIT_51 => X"0000000f000000000000000c0000000000000003000000000000001600000000",
            INIT_52 => X"ffffffe0ffffffffffffffefffffffff0000000000000000fffffffaffffffff",
            INIT_53 => X"ffffffc8ffffffffffffffe5fffffffffffffffcffffffff0000000000000000",
            INIT_54 => X"0000002a00000000ffffffe8ffffffff0000000d000000000000002700000000",
            INIT_55 => X"0000003500000000000000120000000000000060000000000000004100000000",
            INIT_56 => X"00000017000000000000001a000000000000000f000000000000001d00000000",
            INIT_57 => X"fffffff9ffffffff00000022000000000000003f00000000ffffffedffffffff",
            INIT_58 => X"0000000000000000000000060000000000000037000000000000004600000000",
            INIT_59 => X"0000000c000000000000002c000000000000000600000000fffffff8ffffffff",
            INIT_5A => X"0000001600000000ffffffd4ffffffff0000000000000000ffffffe4ffffffff",
            INIT_5B => X"00000001000000000000000d000000000000000a00000000fffffffdffffffff",
            INIT_5C => X"0000000200000000fffffffeffffffff00000004000000000000000200000000",
            INIT_5D => X"0000000d000000000000001f0000000000000018000000000000002b00000000",
            INIT_5E => X"fffffffbffffffff000000130000000000000016000000000000001300000000",
            INIT_5F => X"0000000e00000000ffffffe6ffffffff00000002000000000000000400000000",
            INIT_60 => X"00000014000000000000001500000000ffffffdfffffffff0000001000000000",
            INIT_61 => X"0000001b00000000ffffffdaffffffff0000000d00000000fffffffaffffffff",
            INIT_62 => X"ffffffe3ffffffffffffffeeffffffffffffffcefffffffffffffff0ffffffff",
            INIT_63 => X"fffffff5ffffffff0000000200000000ffffffecfffffffffffffff7ffffffff",
            INIT_64 => X"0000003f000000000000002200000000fffffffffffffffffffffff2ffffffff",
            INIT_65 => X"000000110000000000000012000000000000001a000000000000003200000000",
            INIT_66 => X"0000002e00000000ffffffe7ffffffffffffffceffffffff0000001700000000",
            INIT_67 => X"ffffffecffffffff0000002300000000ffffffd6fffffffffffffff5ffffffff",
            INIT_68 => X"ffffffdaffffffffffffffdaffffffffffffffedffffffffffffffbeffffffff",
            INIT_69 => X"fffffff1ffffffffffffffd6ffffffff0000002e00000000ffffffe7ffffffff",
            INIT_6A => X"ffffffe0ffffffffffffffccffffffff00000008000000000000000500000000",
            INIT_6B => X"ffffffeeffffffffffffffe9ffffffffffffffd4ffffffffffffffe5ffffffff",
            INIT_6C => X"0000000b00000000000000280000000000000006000000000000000800000000",
            INIT_6D => X"ffffffe9ffffffff0000000600000000ffffffd5fffffffffffffff8ffffffff",
            INIT_6E => X"fffffffdfffffffffffffff7ffffffff0000001c00000000ffffffe9ffffffff",
            INIT_6F => X"ffffffd9ffffffff0000001500000000ffffffb6ffffffffffffffa7ffffffff",
            INIT_70 => X"ffffffd7ffffffffffffffbcffffffffffffffd1ffffffffffffffc7ffffffff",
            INIT_71 => X"ffffffd9fffffffffffffffcffffffff0000000d00000000fffffff3ffffffff",
            INIT_72 => X"0000001400000000fffffff1ffffffff00000003000000000000002400000000",
            INIT_73 => X"0000000500000000000000290000000000000011000000000000000600000000",
            INIT_74 => X"ffffffe9fffffffffffffff7ffffffff0000000c000000000000001400000000",
            INIT_75 => X"fffffff6fffffffffffffff0ffffffff0000000f000000000000001100000000",
            INIT_76 => X"0000000a00000000ffffffe5ffffffffffffffecffffffffffffffebffffffff",
            INIT_77 => X"fffffff6ffffffffffffffecffffffffffffffdbffffffffffffffe9ffffffff",
            INIT_78 => X"fffffffffffffffffffffffdffffffffffffffecffffffff0000000f00000000",
            INIT_79 => X"fffffff5fffffffffffffff8ffffffff0000001c00000000fffffff0ffffffff",
            INIT_7A => X"000000050000000000000026000000000000003800000000fffffff9ffffffff",
            INIT_7B => X"fffffff3ffffffffffffffe9fffffffffffffff1ffffffff0000000c00000000",
            INIT_7C => X"ffffffadfffffffffffffffaffffffff0000002c000000000000000e00000000",
            INIT_7D => X"ffffffadffffffffffffff9fffffffffffffffcbffffffffffffff92ffffffff",
            INIT_7E => X"fffffffbffffffffffffffd5ffffffffffffffe7ffffffff0000003600000000",
            INIT_7F => X"ffffffe5ffffffffffffffd0ffffffffffffffc4ffffffffffffff8dffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE2;


    MEM_IWGHT_LAYER2_INSTANCE3 : if BRAM_NAME = "iwght_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffeffffffffffffffdbffffffff0000000400000000ffffffcbffffffff",
            INIT_01 => X"fffffff0ffffffffffffffecffffffffffffffb7fffffffffffffff2ffffffff",
            INIT_02 => X"fffffff7ffffffffffffffd1ffffffffffffffc6ffffffffffffff9effffffff",
            INIT_03 => X"000000220000000000000035000000000000002300000000ffffffebffffffff",
            INIT_04 => X"000000000000000000000031000000000000001a000000000000001200000000",
            INIT_05 => X"ffffffd8ffffffffffffffe0ffffffffffffffedfffffffffffffffdffffffff",
            INIT_06 => X"ffffffd8fffffffffffffffdfffffffffffffff3ffffffffffffffdeffffffff",
            INIT_07 => X"0000001b00000000fffffffcfffffffffffffff2ffffffff0000000800000000",
            INIT_08 => X"ffffffefffffffff000000070000000000000012000000000000000a00000000",
            INIT_09 => X"0000001900000000ffffffeeffffffffffffffe3ffffffff0000001c00000000",
            INIT_0A => X"ffffffbafffffffffffffff4ffffffffffffffd4fffffffffffffffeffffffff",
            INIT_0B => X"fffffff1ffffffffffffffd3ffffffffffffffe0ffffffffffffffb7ffffffff",
            INIT_0C => X"0000000d000000000000002400000000fffffffaffffffff0000000c00000000",
            INIT_0D => X"0000001500000000fffffff1ffffffff00000018000000000000002d00000000",
            INIT_0E => X"ffffffd7fffffffffffffffaffffffff00000000000000000000001800000000",
            INIT_0F => X"ffffffe0ffffffffffffffe4ffffffffffffffefffffffffffffffdfffffffff",
            INIT_10 => X"ffffffe8ffffffff000000580000000000000016000000000000000e00000000",
            INIT_11 => X"00000000000000000000000700000000ffffffe0ffffffffffffffdcffffffff",
            INIT_12 => X"ffffffbeffffffffffffffe2ffffffff0000001000000000ffffffbdffffffff",
            INIT_13 => X"000000000000000000000010000000000000000d00000000fffffffcffffffff",
            INIT_14 => X"ffffffeeffffffff00000001000000000000000700000000fffffffdffffffff",
            INIT_15 => X"0000000000000000000000140000000000000010000000000000000600000000",
            INIT_16 => X"0000001a00000000000000160000000000000012000000000000001900000000",
            INIT_17 => X"0000000800000000000000190000000000000010000000000000000b00000000",
            INIT_18 => X"ffffffeffffffffffffffffeffffffffffffffe4ffffffff0000001a00000000",
            INIT_19 => X"0000000400000000fffffff9ffffffffffffffeeffffffffffffffe3ffffffff",
            INIT_1A => X"00000011000000000000000f0000000000000012000000000000002000000000",
            INIT_1B => X"ffffffd5ffffffff00000000000000000000000e00000000fffffff8ffffffff",
            INIT_1C => X"ffffffe9ffffffffffffffddffffffffffffffd1ffffffffffffffe5ffffffff",
            INIT_1D => X"ffffffedffffffffffffffd7ffffffff0000000100000000ffffffbcffffffff",
            INIT_1E => X"00000016000000000000000300000000fffffffdffffffff0000000200000000",
            INIT_1F => X"0000001400000000fffffff8ffffffff0000000f000000000000003e00000000",
            INIT_20 => X"0000000700000000fffffff9ffffffffffffffd3fffffffffffffffdffffffff",
            INIT_21 => X"fffffffaffffffff0000000a00000000fffffffeffffffffffffffc4ffffffff",
            INIT_22 => X"0000000000000000ffffffe2ffffffff00000022000000000000001500000000",
            INIT_23 => X"0000000d00000000000000020000000000000011000000000000001200000000",
            INIT_24 => X"0000000a000000000000000700000000ffffffdbffffffff0000002300000000",
            INIT_25 => X"0000002300000000000000210000000000000025000000000000001400000000",
            INIT_26 => X"0000000500000000ffffffe7ffffffff00000034000000000000001c00000000",
            INIT_27 => X"0000002f0000000000000005000000000000000c000000000000000d00000000",
            INIT_28 => X"fffffffdffffffff0000003c0000000000000027000000000000000900000000",
            INIT_29 => X"0000000b00000000fffffff4ffffffffffffffffffffffff0000000500000000",
            INIT_2A => X"ffffffe9ffffffff00000016000000000000000500000000ffffffe5ffffffff",
            INIT_2B => X"ffffffedffffffffffffffc8ffffffff0000000600000000ffffffedffffffff",
            INIT_2C => X"fffffffaffffffffffffffd2fffffffffffffff8ffffffffffffffe5ffffffff",
            INIT_2D => X"0000002b0000000000000013000000000000000f000000000000000a00000000",
            INIT_2E => X"fffffffbffffffffffffffdeffffffffffffffb3ffffffff0000001c00000000",
            INIT_2F => X"fffffff9ffffffff0000003300000000fffffff1fffffffffffffff8ffffffff",
            INIT_30 => X"ffffffeefffffffffffffff2ffffffff0000001b00000000ffffffe2ffffffff",
            INIT_31 => X"000000150000000000000005000000000000000e000000000000000700000000",
            INIT_32 => X"0000002100000000000000220000000000000031000000000000001a00000000",
            INIT_33 => X"ffffffd2ffffffff0000000a000000000000002e00000000fffffff7ffffffff",
            INIT_34 => X"fffffff7ffffffffffffffecffffffff00000004000000000000004400000000",
            INIT_35 => X"0000000700000000ffffffc3fffffffffffffff9fffffffffffffff1ffffffff",
            INIT_36 => X"00000002000000000000000000000000ffffffffffffffff0000000500000000",
            INIT_37 => X"ffffffd4ffffffffffffffbdffffffffffffff78ffffffffffffffbeffffffff",
            INIT_38 => X"ffffffd5fffffffffffffff0ffffffffffffffcdffffffffffffffb8ffffffff",
            INIT_39 => X"00000015000000000000000b000000000000000f00000000ffffffd3ffffffff",
            INIT_3A => X"0000001e0000000000000030000000000000002100000000fffffffcffffffff",
            INIT_3B => X"0000001d000000000000000b00000000fffffff8ffffffffffffffeaffffffff",
            INIT_3C => X"0000001a00000000000000190000000000000004000000000000001000000000",
            INIT_3D => X"00000017000000000000002f00000000fffffffbfffffffffffffffcffffffff",
            INIT_3E => X"000000170000000000000037000000000000001e000000000000001900000000",
            INIT_3F => X"ffffffc6ffffffff0000000c000000000000002500000000fffffff8ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff1fffffffffffffff1ffffffffffffffe5ffffffffffffffd8ffffffff",
            INIT_41 => X"fffffff2fffffffffffffff9fffffffffffffffbffffffffffffffeaffffffff",
            INIT_42 => X"00000029000000000000002a000000000000002600000000ffffffebffffffff",
            INIT_43 => X"fffffff7ffffffff000000150000000000000025000000000000003200000000",
            INIT_44 => X"0000000e000000000000000000000000ffffffb8ffffffffffffffbbffffffff",
            INIT_45 => X"0000002600000000ffffffeaffffffffffffffe2fffffffffffffffdffffffff",
            INIT_46 => X"fffffff6ffffffff0000001a00000000fffffff5ffffffffffffffe5ffffffff",
            INIT_47 => X"ffffffdaffffffffffffffd6ffffffff00000031000000000000001200000000",
            INIT_48 => X"0000002300000000ffffffedffffffffffffffe8ffffffff0000000d00000000",
            INIT_49 => X"0000002e00000000ffffffeaffffffff0000001c00000000ffffffdaffffffff",
            INIT_4A => X"0000001a00000000fffffff0ffffffff00000016000000000000003500000000",
            INIT_4B => X"0000000500000000000000080000000000000004000000000000000700000000",
            INIT_4C => X"00000027000000000000001c0000000000000036000000000000001500000000",
            INIT_4D => X"0000000200000000000000380000000000000033000000000000003100000000",
            INIT_4E => X"ffffffedfffffffffffffff9ffffffff00000019000000000000002400000000",
            INIT_4F => X"fffffff2ffffffffffffffd3ffffffffffffffcdfffffffffffffff2ffffffff",
            INIT_50 => X"ffffffa1ffffffffffffffb5fffffffffffffff1fffffffffffffff1ffffffff",
            INIT_51 => X"ffffffcbffffffffffffffceffffffffffffffdfffffffffffffffabffffffff",
            INIT_52 => X"0000005300000000000000220000000000000026000000000000002800000000",
            INIT_53 => X"00000003000000000000000e0000000000000037000000000000003f00000000",
            INIT_54 => X"fffffff6fffffffffffffff2fffffffffffffffbfffffffffffffff0ffffffff",
            INIT_55 => X"00000014000000000000000b0000000000000001000000000000000a00000000",
            INIT_56 => X"fffffffeffffffff00000005000000000000000c00000000fffffff0ffffffff",
            INIT_57 => X"0000000b000000000000000a000000000000001b000000000000001700000000",
            INIT_58 => X"0000000b00000000ffffffddfffffffffffffff1ffffffffffffffdeffffffff",
            INIT_59 => X"000000000000000000000002000000000000002100000000ffffffefffffffff",
            INIT_5A => X"0000003000000000fffffffdfffffffffffffffcffffffff0000004000000000",
            INIT_5B => X"ffffffe5ffffffff000000200000000000000021000000000000002100000000",
            INIT_5C => X"fffffff5ffffffffffffffe8ffffffff00000013000000000000001900000000",
            INIT_5D => X"ffffffe7ffffffffffffffc4ffffffffffffffdefffffffffffffff2ffffffff",
            INIT_5E => X"ffffffeeffffffffffffffcaffffffffffffffc1ffffffffffffffccffffffff",
            INIT_5F => X"00000025000000000000000a00000000ffffffd2ffffffffffffffddffffffff",
            INIT_60 => X"00000023000000000000003a0000000000000022000000000000002c00000000",
            INIT_61 => X"00000018000000000000001300000000fffffff3ffffffff0000000600000000",
            INIT_62 => X"fffffffefffffffffffffffffffffffffffffff7fffffffffffffff0ffffffff",
            INIT_63 => X"0000002c000000000000001a00000000ffffffe4ffffffff0000000e00000000",
            INIT_64 => X"ffffffabfffffffffffffff5ffffffff00000002000000000000001100000000",
            INIT_65 => X"ffffff95ffffffffffffffaeffffffffffffffedffffffffffffffb3ffffffff",
            INIT_66 => X"000000130000000000000005000000000000001a00000000ffffffa3ffffffff",
            INIT_67 => X"fffffff5ffffffff0000002f0000000000000016000000000000002200000000",
            INIT_68 => X"0000000c00000000ffffffd3ffffffff00000006000000000000000800000000",
            INIT_69 => X"0000003100000000fffffffaffffffffffffffd5ffffffff0000001600000000",
            INIT_6A => X"000000340000000000000011000000000000003400000000ffffffecffffffff",
            INIT_6B => X"0000001600000000fffffff6ffffffff0000001d000000000000003200000000",
            INIT_6C => X"fffffff1fffffffffffffff5fffffffffffffff0ffffffffffffffefffffffff",
            INIT_6D => X"ffffffceffffffff0000000400000000ffffffeeffffffff0000000400000000",
            INIT_6E => X"0000000400000000fffffffcffffffffffffffe9fffffffffffffffdffffffff",
            INIT_6F => X"0000001a00000000000000270000000000000025000000000000001500000000",
            INIT_70 => X"0000001f00000000fffffffbffffffff00000016000000000000000e00000000",
            INIT_71 => X"0000002d00000000000000290000000000000011000000000000001500000000",
            INIT_72 => X"0000000f00000000000000020000000000000017000000000000001f00000000",
            INIT_73 => X"0000000b00000000ffffffe3ffffffffffffffd0ffffffffffffffe5ffffffff",
            INIT_74 => X"0000000a00000000ffffffe9ffffffffffffffffffffffff0000001200000000",
            INIT_75 => X"fffffffbffffffffffffffebffffffffffffffe5fffffffffffffffeffffffff",
            INIT_76 => X"ffffffe8ffffffffffffffcefffffffffffffffaffffffff0000002b00000000",
            INIT_77 => X"ffffffefffffffffffffffbbffffffffffffffacffffffffffffffdcffffffff",
            INIT_78 => X"000000130000000000000002000000000000000700000000ffffffcdffffffff",
            INIT_79 => X"ffffffc6ffffffffffffffb6ffffffffffffffacffffffffffffffb0ffffffff",
            INIT_7A => X"00000011000000000000001900000000ffffffabffffffffffffffb6ffffffff",
            INIT_7B => X"0000002400000000fffffffeffffffffffffffecffffffff0000000300000000",
            INIT_7C => X"0000001a000000000000000300000000ffffffffffffffffffffffe0ffffffff",
            INIT_7D => X"fffffff8ffffffff0000000b00000000ffffffecffffffff0000000a00000000",
            INIT_7E => X"ffffffb7ffffffffffffffbaffffffffffffffb6ffffffffffffffbaffffffff",
            INIT_7F => X"ffffffcdfffffffffffffffefffffffffffffff8fffffffffffffffcffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE3;


    MEM_IWGHT_LAYER2_INSTANCE4 : if BRAM_NAME = "iwght_layer2_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004e00000000fffffff4ffffffff0000002f000000000000001000000000",
            INIT_01 => X"ffffffdeffffffffffffffe2ffffffff00000009000000000000002e00000000",
            INIT_02 => X"ffffffe4ffffffffffffffb3ffffffffffffffd3fffffffffffffff0ffffffff",
            INIT_03 => X"0000000500000000fffffff6ffffffffffffffc3ffffffffffffffc3ffffffff",
            INIT_04 => X"0000000000000000ffffffefffffffffffffffd3ffffffff0000000600000000",
            INIT_05 => X"fffffff9fffffffffffffffefffffffffffffff8ffffffff0000001000000000",
            INIT_06 => X"ffffffefffffffff00000013000000000000001f00000000fffffff5ffffffff",
            INIT_07 => X"0000001e000000000000001000000000fffffffeffffffff0000001600000000",
            INIT_08 => X"fffffff5ffffffff0000000c000000000000000f00000000fffffffdffffffff",
            INIT_09 => X"00000012000000000000000c000000000000000e000000000000000b00000000",
            INIT_0A => X"ffffffecfffffffffffffffefffffffffffffff2fffffffffffffffbffffffff",
            INIT_0B => X"ffffffe5fffffffffffffff4fffffffffffffffbffffffff0000000c00000000",
            INIT_0C => X"00000001000000000000000900000000ffffffe7fffffffffffffffaffffffff",
            INIT_0D => X"0000000000000000fffffff3ffffffff0000000100000000fffffffcffffffff",
            INIT_0E => X"ffffffe6fffffffffffffffaffffffff0000000200000000fffffff8ffffffff",
            INIT_0F => X"0000000000000000fffffff5ffffffffffffffeaffffffff0000000100000000",
            INIT_10 => X"0000000000000000fffffff6ffffffffffffffffffffffff0000000500000000",
            INIT_11 => X"ffffffe5ffffffff0000000300000000ffffffeefffffffffffffff4ffffffff",
            INIT_12 => X"ffffffebffffffffffffffeefffffffffffffffafffffffffffffff6ffffffff",
            INIT_13 => X"ffffffe9ffffffffffffffecffffffff00000001000000000000000600000000",
            INIT_14 => X"fffffff4ffffffff000000000000000000000009000000000000000a00000000",
            INIT_15 => X"fffffffeffffffff00000005000000000000000100000000fffffff4ffffffff",
            INIT_16 => X"ffffffebffffffff0000001100000000fffffffffffffffffffffffbffffffff",
            INIT_17 => X"ffffffeffffffffffffffff9ffffffffffffffedfffffffffffffff5ffffffff",
            INIT_18 => X"ffffffe8ffffffff00000004000000000000000600000000fffffff6ffffffff",
            INIT_19 => X"0000000400000000fffffff5ffffffff00000007000000000000000500000000",
            INIT_1A => X"fffffffbfffffffffffffff6fffffffffffffff1ffffffffffffffe0ffffffff",
            INIT_1B => X"ffffffe3ffffffffffffffffffffffff00000005000000000000000500000000",
            INIT_1C => X"0000000600000000fffffff0ffffffff00000000000000000000000500000000",
            INIT_1D => X"0000001400000000ffffffefffffffff0000000b00000000fffffffcffffffff",
            INIT_1E => X"fffffff1ffffffffffffffe3ffffffff0000000600000000ffffffedffffffff",
            INIT_1F => X"0000000000000000ffffffe3ffffffffffffffe5fffffffffffffffcffffffff",
            INIT_20 => X"0000000300000000ffffffe7ffffffff0000000000000000ffffffe5ffffffff",
            INIT_21 => X"fffffffdffffffff0000000d00000000fffffff4fffffffffffffffcffffffff",
            INIT_22 => X"0000000c00000000fffffffafffffffffffffff2ffffffff0000000800000000",
            INIT_23 => X"0000000700000000000000130000000000000013000000000000000600000000",
            INIT_24 => X"fffffff8ffffffff0000000d00000000ffffffebffffffffffffffeeffffffff",
            INIT_25 => X"fffffff9fffffffffffffff3fffffffffffffffaffffffff0000001300000000",
            INIT_26 => X"fffffff2ffffffff00000000000000000000000400000000fffffff8ffffffff",
            INIT_27 => X"0000000000000000000000030000000000000000000000000000000700000000",
            INIT_28 => X"0000000e00000000fffffff7ffffffffffffffeafffffffffffffffdffffffff",
            INIT_29 => X"ffffffe4ffffffffffffffffffffffff0000000d00000000fffffff8ffffffff",
            INIT_2A => X"ffffffedffffffff00000008000000000000000400000000fffffff8ffffffff",
            INIT_2B => X"fffffffdfffffffffffffff0fffffffffffffff2ffffffff0000000b00000000",
            INIT_2C => X"00000000000000000000000100000000ffffffeafffffffffffffff0ffffffff",
            INIT_2D => X"fffffffdffffffff0000000c00000000fffffffefffffffffffffff7ffffffff",
            INIT_2E => X"fffffff7fffffffffffffffbfffffffffffffff8fffffffffffffff0ffffffff",
            INIT_2F => X"0000000500000000fffffff2ffffffffffffffecfffffffffffffffdffffffff",
            INIT_30 => X"0000000300000000ffffffe7ffffffff0000000400000000fffffff0ffffffff",
            INIT_31 => X"ffffffedffffffffffffffeefffffffffffffffefffffffffffffffbffffffff",
            INIT_32 => X"fffffff8fffffffffffffff4ffffffff00000009000000000000000700000000",
            INIT_33 => X"0000000900000000ffffffe7ffffffffffffffe9ffffffff0000000000000000",
            INIT_34 => X"ffffffe9fffffffffffffff3ffffffff00000001000000000000000600000000",
            INIT_35 => X"ffffffeafffffffffffffffffffffffffffffff2fffffffffffffff5ffffffff",
            INIT_36 => X"ffffffeffffffffffffffff9fffffffffffffff1ffffffffffffffe3ffffffff",
            INIT_37 => X"fffffff8ffffffffffffffeffffffffffffffffcffffffff0000000800000000",
            INIT_38 => X"fffffffcffffffff0000000200000000ffffffe7ffffffff0000000a00000000",
            INIT_39 => X"0000000900000000fffffff9ffffffff0000000500000000fffffff1ffffffff",
            INIT_3A => X"fffffff1ffffffff00000011000000000000000e00000000fffffffcffffffff",
            INIT_3B => X"fffffff8fffffffffffffff5ffffffff0000000e00000000ffffffeeffffffff",
            INIT_3C => X"ffffffe6fffffffffffffff6fffffffffffffff9fffffffffffffffbffffffff",
            INIT_3D => X"ffffffeafffffffffffffffafffffffffffffff0fffffffffffffff9ffffffff",
            INIT_3E => X"fffffff7ffffffff0000000b000000000000000100000000fffffff5ffffffff",
            INIT_3F => X"ffffffecffffffff0000000400000000ffffffe1fffffffffffffffdffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000300000000ffffffe6fffffffffffffffcffffffffffffffeaffffffff",
            INIT_41 => X"ffffffdafffffffffffffff1fffffffffffffff1fffffffffffffff1ffffffff",
            INIT_42 => X"fffffff5ffffffff0000001000000000ffffffecffffffff0000000000000000",
            INIT_43 => X"000000070000000000000002000000000000001100000000fffffff3ffffffff",
            INIT_44 => X"0000000f00000000ffffffefffffffff00000007000000000000001400000000",
            INIT_45 => X"ffffffedffffffff00000003000000000000000a00000000fffffffaffffffff",
            INIT_46 => X"ffffffedfffffffffffffffeffffffff00000001000000000000000400000000",
            INIT_47 => X"fffffff7ffffffff0000000d00000000ffffffffffffffffffffffe8ffffffff",
            INIT_48 => X"0000000a000000000000000000000000fffffff2fffffffffffffff1ffffffff",
            INIT_49 => X"00000002000000000000000100000000fffffffcffffffff0000000000000000",
            INIT_4A => X"0000000100000000fffffff8fffffffffffffffffffffffffffffffdffffffff",
            INIT_4B => X"000000060000000000000004000000000000000500000000fffffff5ffffffff",
            INIT_4C => X"00000006000000000000000500000000fffffffeffffffff0000000100000000",
            INIT_4D => X"fffffffcfffffffffffffffcffffffff0000000800000000fffffff6ffffffff",
            INIT_4E => X"0000000000000000fffffff0ffffffff0000000300000000ffffffe9ffffffff",
            INIT_4F => X"00000000000000000000000b00000000ffffffebffffffffffffffecffffffff",
            INIT_50 => X"ffffffebffffffff0000000f00000000fffffff9ffffffff0000000000000000",
            INIT_51 => X"fffffffdfffffffffffffff7fffffffffffffffdffffffff0000000300000000",
            INIT_52 => X"fffffffcffffffff0000000400000000fffffff1ffffffff0000000a00000000",
            INIT_53 => X"ffffffdcffffffffffffffdbffffffff00000015000000000000000200000000",
            INIT_54 => X"ffffffeeffffffff0000002200000000ffffffd9ffffffffffffffb8ffffffff",
            INIT_55 => X"000000210000000000000010000000000000001900000000fffffff7ffffffff",
            INIT_56 => X"0000001c00000000000000050000000000000005000000000000002e00000000",
            INIT_57 => X"0000003000000000fffffff4ffffffff0000000a000000000000002f00000000",
            INIT_58 => X"0000002200000000000000480000000000000002000000000000002e00000000",
            INIT_59 => X"fffffff6ffffffff0000002800000000ffffffedffffffffffffffe6ffffffff",
            INIT_5A => X"000000420000000000000036000000000000001e000000000000001400000000",
            INIT_5B => X"00000011000000000000001d00000000fffffff7ffffffff0000001900000000",
            INIT_5C => X"0000002700000000ffffffedffffffff00000048000000000000002b00000000",
            INIT_5D => X"0000000f00000000ffffffddffffffff00000034000000000000003b00000000",
            INIT_5E => X"fffffffeffffffffffffffc9ffffffffffffffdcffffffff0000000a00000000",
            INIT_5F => X"00000024000000000000002900000000fffffff4ffffffffffffffd5ffffffff",
            INIT_60 => X"ffffffdafffffffffffffffffffffffffffffff1ffffffff0000000d00000000",
            INIT_61 => X"00000016000000000000000c00000000ffffffe6fffffffffffffffdffffffff",
            INIT_62 => X"ffffffe3ffffffff0000000300000000fffffffeffffffffffffffe8ffffffff",
            INIT_63 => X"ffffffeaffffffff0000001c000000000000001a00000000ffffffeeffffffff",
            INIT_64 => X"0000002f000000000000001000000000ffffffdcffffffff0000001000000000",
            INIT_65 => X"00000006000000000000000000000000ffffffd1ffffffffffffffedffffffff",
            INIT_66 => X"ffffffebffffffffffffffecffffffff0000000100000000fffffff0ffffffff",
            INIT_67 => X"ffffffffffffffffffffffdfffffffffffffffbeffffffff0000000200000000",
            INIT_68 => X"fffffffaffffffffffffffe2ffffffffffffffc7ffffffffffffffb9ffffffff",
            INIT_69 => X"fffffffaffffffffffffffefffffffff0000000600000000fffffffcffffffff",
            INIT_6A => X"0000001500000000fffffff4ffffffffffffffe8ffffffff0000000f00000000",
            INIT_6B => X"fffffffbffffffffffffffdeffffffffffffffebfffffffffffffff5ffffffff",
            INIT_6C => X"ffffffefffffffffffffffd9ffffffff0000001700000000fffffffcffffffff",
            INIT_6D => X"ffffffceffffffff0000000a00000000fffffff0fffffffffffffff3ffffffff",
            INIT_6E => X"ffffffbfffffffff0000000300000000ffffffeeffffffff0000000000000000",
            INIT_6F => X"fffffff7ffffffffffffffebfffffffffffffff8ffffffffffffffd9ffffffff",
            INIT_70 => X"0000000f000000000000000d00000000fffffff0ffffffff0000001300000000",
            INIT_71 => X"fffffffdffffffff00000000000000000000000200000000fffffff9ffffffff",
            INIT_72 => X"ffffffeaffffffff0000000600000000ffffffe7ffffffffffffffd1ffffffff",
            INIT_73 => X"ffffffdeffffffffffffffc9ffffffffffffffdfffffffffffffffe0ffffffff",
            INIT_74 => X"ffffffbdffffffff0000001500000000fffffff9ffffffff0000001800000000",
            INIT_75 => X"ffffffdeffffffffffffffaaffffffffffffffd6ffffffff0000002400000000",
            INIT_76 => X"0000002e000000000000001300000000ffffffefffffffff0000000a00000000",
            INIT_77 => X"ffffffc0ffffffff0000000000000000ffffffd9ffffffffffffffc1ffffffff",
            INIT_78 => X"fffffff4ffffffff0000001200000000fffffff0ffffffffffffffefffffffff",
            INIT_79 => X"0000002e00000000000000310000000000000011000000000000000700000000",
            INIT_7A => X"ffffffeafffffffffffffffbffffffff0000002e000000000000000e00000000",
            INIT_7B => X"0000000400000000fffffffcffffffff0000000000000000ffffffe7ffffffff",
            INIT_7C => X"ffffffefffffffff00000005000000000000000200000000fffffffaffffffff",
            INIT_7D => X"fffffff0ffffffff000000220000000000000004000000000000000100000000",
            INIT_7E => X"fffffffafffffffffffffffeffffffff0000000200000000fffffff5ffffffff",
            INIT_7F => X"fffffffaffffffff0000000900000000ffffffdffffffffffffffff1ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE4;


    MEM_IWGHT_LAYER2_INSTANCE5 : if BRAM_NAME = "iwght_layer2_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffcffffffff0000000400000000fffffffbffffffff0000000f00000000",
            INIT_01 => X"fffffff2ffffffffffffffb3fffffffffffffff0ffffffffffffffeaffffffff",
            INIT_02 => X"0000000500000000fffffff7ffffffffffffffdaffffffff0000002300000000",
            INIT_03 => X"ffffffcbfffffffffffffffbffffffffffffffdcfffffffffffffff4ffffffff",
            INIT_04 => X"ffffffe6ffffffffffffffb1ffffffff0000001800000000fffffffaffffffff",
            INIT_05 => X"0000001600000000ffffffe0ffffffffffffffa2ffffffff0000000f00000000",
            INIT_06 => X"0000001e000000000000004d00000000ffffffd5ffffffffffffffc4ffffffff",
            INIT_07 => X"ffffffe5ffffffff000000080000000000000024000000000000000200000000",
            INIT_08 => X"ffffffd9ffffffffffffffecfffffffffffffffffffffffffffffff0ffffffff",
            INIT_09 => X"ffffffbcffffffffffffffe3ffffffffffffffeeffffffffffffffd1ffffffff",
            INIT_0A => X"0000000900000000ffffffe8ffffffff0000001200000000fffffffcffffffff",
            INIT_0B => X"0000002400000000ffffffe2ffffffff0000000c000000000000000c00000000",
            INIT_0C => X"ffffffebffffffff0000000a00000000ffffffcffffffffffffffff8ffffffff",
            INIT_0D => X"0000000800000000ffffffdeffffffff0000001a00000000fffffff8ffffffff",
            INIT_0E => X"ffffffe4ffffffffffffffcdffffffffffffffdfffffffff0000000500000000",
            INIT_0F => X"0000002a000000000000001d000000000000002a000000000000001400000000",
            INIT_10 => X"000000690000000000000056000000000000002a000000000000001600000000",
            INIT_11 => X"00000004000000000000002500000000ffffffe9ffffffff0000003800000000",
            INIT_12 => X"ffffffd6fffffffffffffff5fffffffffffffffbffffffffffffffcbffffffff",
            INIT_13 => X"00000003000000000000001a00000000fffffff6ffffffffffffff9bffffffff",
            INIT_14 => X"fffffffefffffffffffffff6ffffffffffffffe9ffffffff0000001500000000",
            INIT_15 => X"0000000a0000000000000028000000000000000500000000ffffffd6ffffffff",
            INIT_16 => X"0000000600000000fffffffcffffffff0000000700000000fffffffdffffffff",
            INIT_17 => X"0000000e0000000000000018000000000000001f000000000000001700000000",
            INIT_18 => X"fffffff7ffffffffffffffe9ffffffffffffffebffffffff0000000500000000",
            INIT_19 => X"0000000f00000000000000010000000000000002000000000000001e00000000",
            INIT_1A => X"fffffff0fffffffffffffffeffffffff0000001e00000000fffffff0ffffffff",
            INIT_1B => X"000000190000000000000022000000000000002f000000000000002c00000000",
            INIT_1C => X"ffffffd4ffffffffffffffe4ffffffff00000000000000000000001600000000",
            INIT_1D => X"00000012000000000000001100000000fffffff9ffffffffffffffe5ffffffff",
            INIT_1E => X"000000270000000000000010000000000000001a00000000fffffff8ffffffff",
            INIT_1F => X"00000037000000000000000500000000ffffffe5fffffffffffffff3ffffffff",
            INIT_20 => X"0000000600000000000000350000000000000025000000000000000600000000",
            INIT_21 => X"0000001000000000ffffffecffffffffffffffd0ffffffffffffffefffffffff",
            INIT_22 => X"00000046000000000000000000000000ffffffdaffffffff0000000000000000",
            INIT_23 => X"0000002200000000fffffffdfffffffffffffff4ffffffffffffffeaffffffff",
            INIT_24 => X"00000006000000000000000800000000fffffff9ffffffff0000002600000000",
            INIT_25 => X"fffffff5fffffffffffffffcffffffff0000001a000000000000000000000000",
            INIT_26 => X"00000005000000000000000d000000000000001d00000000ffffffdfffffffff",
            INIT_27 => X"0000002000000000000000180000000000000008000000000000002600000000",
            INIT_28 => X"00000013000000000000002800000000fffffff3ffffffff0000000000000000",
            INIT_29 => X"fffffff3ffffffff0000000900000000fffffffbffffffffffffffebffffffff",
            INIT_2A => X"0000001100000000ffffffd0ffffffffffffffe7ffffffffffffffefffffffff",
            INIT_2B => X"fffffff1ffffffffffffffecfffffffffffffff2ffffffff0000001100000000",
            INIT_2C => X"00000022000000000000000800000000ffffffd9ffffffffffffffd0ffffffff",
            INIT_2D => X"ffffffe8ffffffff0000001800000000ffffffebffffffffffffffc1ffffffff",
            INIT_2E => X"00000014000000000000002d000000000000002000000000ffffffd1ffffffff",
            INIT_2F => X"00000014000000000000000d000000000000003100000000fffffff7ffffffff",
            INIT_30 => X"ffffffd7ffffffffffffffeafffffffffffffffdffffffff0000001300000000",
            INIT_31 => X"ffffffe4ffffffffffffffc8ffffffff0000000800000000ffffffe1ffffffff",
            INIT_32 => X"fffffffbffffffffffffffdfffffffffffffffcfffffffff0000000d00000000",
            INIT_33 => X"fffffffdffffffff00000011000000000000001a00000000fffffff8ffffffff",
            INIT_34 => X"00000000000000000000000d000000000000000e00000000fffffffcffffffff",
            INIT_35 => X"fffffffbffffffff0000001f000000000000000d000000000000000400000000",
            INIT_36 => X"ffffffc9ffffffff0000000000000000fffffff7fffffffffffffff0ffffffff",
            INIT_37 => X"fffffff6ffffffffffffffffffffffffffffffeffffffffffffffff1ffffffff",
            INIT_38 => X"ffffffcfffffffffffffffd2fffffffffffffffcffffffff0000001600000000",
            INIT_39 => X"ffffffc0ffffffffffffffcffffffffffffffff9ffffffff0000001900000000",
            INIT_3A => X"ffffffe4ffffffffffffffe9ffffffff0000001200000000fffffffdffffffff",
            INIT_3B => X"00000049000000000000000200000000ffffffd9ffffffff0000004700000000",
            INIT_3C => X"00000018000000000000000d00000000fffffffcffffffff0000000200000000",
            INIT_3D => X"ffffffefffffffff000000140000000000000013000000000000000800000000",
            INIT_3E => X"ffffffe5ffffffffffffffd2ffffffffffffffe6ffffffff0000000400000000",
            INIT_3F => X"ffffffd9ffffffff0000003000000000ffffffe3ffffffffffffffc0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000600000000ffffffd3ffffffff0000001000000000fffffff0ffffffff",
            INIT_41 => X"0000003500000000fffffffdffffffffffffffdffffffffffffffff4ffffffff",
            INIT_42 => X"0000000c000000000000000f00000000ffffffedfffffffffffffffbffffffff",
            INIT_43 => X"00000011000000000000001c0000000000000013000000000000001700000000",
            INIT_44 => X"000000160000000000000002000000000000002e00000000ffffffffffffffff",
            INIT_45 => X"0000001600000000fffffffcffffffff00000012000000000000001b00000000",
            INIT_46 => X"ffffffdaffffffff00000004000000000000000a00000000ffffffe2ffffffff",
            INIT_47 => X"00000012000000000000000200000000fffffff2fffffffffffffff3ffffffff",
            INIT_48 => X"ffffffe9ffffffff0000000b00000000fffffff3ffffffff0000001900000000",
            INIT_49 => X"0000001b00000000fffffff1ffffffff0000000200000000fffffff7ffffffff",
            INIT_4A => X"0000002d00000000fffffff4ffffffffffffffe9ffffffff0000000000000000",
            INIT_4B => X"ffffffebffffffff0000000800000000ffffffeeffffffff0000000a00000000",
            INIT_4C => X"0000000a000000000000003000000000ffffffefffffffffffffffe9ffffffff",
            INIT_4D => X"ffffffd6fffffffffffffff4ffffffff0000002300000000ffffffccffffffff",
            INIT_4E => X"0000001300000000ffffffedffffffff0000001d000000000000002100000000",
            INIT_4F => X"0000005300000000000000250000000000000046000000000000004800000000",
            INIT_50 => X"ffffffe9ffffffff000000100000000000000038000000000000004f00000000",
            INIT_51 => X"00000020000000000000000a000000000000003b000000000000002100000000",
            INIT_52 => X"ffffffeaffffffffffffffd5ffffffffffffffe1ffffffff0000001800000000",
            INIT_53 => X"0000002d00000000ffffffcbffffffffffffff98ffffffff0000002100000000",
            INIT_54 => X"00000002000000000000001e00000000fffffffbffffffffffffffdeffffffff",
            INIT_55 => X"fffffffdffffffff0000002c000000000000001400000000ffffffe1ffffffff",
            INIT_56 => X"fffffff8ffffffff0000001a000000000000003c00000000ffffffe0ffffffff",
            INIT_57 => X"fffffff2ffffffffffffffeaffffffffffffffdefffffffffffffffcffffffff",
            INIT_58 => X"0000004e000000000000004500000000fffffff3ffffffff0000002b00000000",
            INIT_59 => X"0000002d00000000fffffff9ffffffffffffffdaffffffff0000002100000000",
            INIT_5A => X"0000000900000000fffffff8ffffffffffffffe1ffffffff0000000000000000",
            INIT_5B => X"00000034000000000000001700000000ffffffd8ffffffffffffffd0ffffffff",
            INIT_5C => X"ffffffddffffffff000000010000000000000029000000000000000c00000000",
            INIT_5D => X"ffffffaeffffffffffffffd9ffffffffffffffd6ffffffff0000000a00000000",
            INIT_5E => X"ffffffd0ffffffffffffff9bffffffff0000002400000000ffffffe5ffffffff",
            INIT_5F => X"0000004f000000000000001100000000ffffffd9ffffffff0000001700000000",
            INIT_60 => X"fffffffefffffffffffffff9fffffffffffffffefffffffffffffffcffffffff",
            INIT_61 => X"0000000a00000000000000080000000000000000000000000000000300000000",
            INIT_62 => X"ffffffaeffffffffffffffb7ffffffff0000000200000000ffffffffffffffff",
            INIT_63 => X"0000001700000000ffffffafffffffffffffffb0ffffffff0000001300000000",
            INIT_64 => X"0000002800000000ffffffddfffffffffffffff1ffffffffffffffffffffffff",
            INIT_65 => X"00000050000000000000002a00000000ffffffdcffffffff0000004300000000",
            INIT_66 => X"ffffffe6ffffffff0000001d00000000fffffffbffffffff0000000600000000",
            INIT_67 => X"0000001400000000fffffff5fffffffffffffffbffffffff0000000100000000",
            INIT_68 => X"00000030000000000000002d00000000ffffffe5ffffffff0000002a00000000",
            INIT_69 => X"0000000d00000000fffffffaffffffff0000002c00000000ffffffe9ffffffff",
            INIT_6A => X"fffffff9ffffffffffffffe3ffffffff00000045000000000000006e00000000",
            INIT_6B => X"0000001800000000ffffffedffffffffffffffe9ffffffff0000001600000000",
            INIT_6C => X"ffffffe6ffffffff0000002c000000000000000900000000ffffffe5ffffffff",
            INIT_6D => X"ffffffe0ffffffff00000000000000000000000500000000fffffffcffffffff",
            INIT_6E => X"fffffff8ffffffff0000000600000000fffffff1ffffffffffffffd4ffffffff",
            INIT_6F => X"000000060000000000000003000000000000001e000000000000002700000000",
            INIT_70 => X"ffffffe9ffffffff0000000500000000ffffffdbfffffffffffffffbffffffff",
            INIT_71 => X"ffffffe0ffffffffffffffe2ffffffff00000005000000000000000200000000",
            INIT_72 => X"fffffff9ffffffff0000002700000000ffffffdbfffffffffffffffaffffffff",
            INIT_73 => X"ffffffe8ffffffff00000017000000000000000400000000fffffff2ffffffff",
            INIT_74 => X"ffffffa5ffffffffffffffe3fffffffffffffff2ffffffff0000000b00000000",
            INIT_75 => X"0000000400000000ffffffbbffffffffffffffd0ffffffff0000002100000000",
            INIT_76 => X"ffffffd2ffffffffffffffe9ffffffffffffffc8ffffffffffffffd2ffffffff",
            INIT_77 => X"0000000a00000000ffffffd6ffffffff00000007000000000000001600000000",
            INIT_78 => X"fffffff3fffffffffffffffbffffffff00000009000000000000000a00000000",
            INIT_79 => X"ffffffeeffffffffffffffdeffffffff00000016000000000000000d00000000",
            INIT_7A => X"ffffffddfffffffffffffffbffffffffffffffe1ffffffff0000000800000000",
            INIT_7B => X"00000009000000000000001e000000000000001e00000000ffffffe2ffffffff",
            INIT_7C => X"0000002b0000000000000016000000000000000d000000000000000700000000",
            INIT_7D => X"ffffffbbffffffffffffffd7ffffffff00000012000000000000001200000000",
            INIT_7E => X"0000003300000000ffffffc3ffffffff00000000000000000000006400000000",
            INIT_7F => X"ffffffe6ffffffffffffffd0ffffffffffffffbdffffffffffffffe8ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE5;


    MEM_IWGHT_LAYER2_INSTANCE6 : if BRAM_NAME = "iwght_layer2_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000003000000000000000c00000000ffffffe6ffffffff0000002900000000",
            INIT_01 => X"fffffff2ffffffffffffffdfffffffffffffffd9ffffffffffffffdfffffffff",
            INIT_02 => X"00000036000000000000000f000000000000000a000000000000000700000000",
            INIT_03 => X"0000000a00000000000000030000000000000013000000000000002600000000",
            INIT_04 => X"fffffffaffffffffffffff7cffffffffffffffcdffffffff0000002a00000000",
            INIT_05 => X"ffffffb9fffffffffffffff4ffffffffffffffa2ffffffffffffff9affffffff",
            INIT_06 => X"ffffffe4fffffffffffffff2ffffffff0000001800000000ffffffcfffffffff",
            INIT_07 => X"0000002700000000ffffffd7fffffffffffffff1ffffffff0000004000000000",
            INIT_08 => X"0000000b00000000fffffff0ffffffffffffffddfffffffffffffff0ffffffff",
            INIT_09 => X"ffffffeeffffffff0000001900000000ffffffeaffffffff0000000d00000000",
            INIT_0A => X"fffffff3ffffffff00000000000000000000001b00000000fffffff8ffffffff",
            INIT_0B => X"fffffffeffffffff000000010000000000000034000000000000002b00000000",
            INIT_0C => X"0000000e00000000000000140000000000000005000000000000001d00000000",
            INIT_0D => X"000000110000000000000004000000000000001e000000000000001c00000000",
            INIT_0E => X"0000001f00000000fffffffaffffffffffffffeeffffffff0000000900000000",
            INIT_0F => X"000000100000000000000000000000000000001300000000ffffffeaffffffff",
            INIT_10 => X"0000000000000000000000260000000000000012000000000000000700000000",
            INIT_11 => X"fffffff7ffffffffffffffeeffffffff0000000000000000fffffffcffffffff",
            INIT_12 => X"ffffffe8ffffffff0000000f00000000fffffff3fffffffffffffffcffffffff",
            INIT_13 => X"000000070000000000000018000000000000001c000000000000000000000000",
            INIT_14 => X"0000000300000000ffffffeaffffffff00000027000000000000001100000000",
            INIT_15 => X"fffffff5ffffffff0000000e00000000ffffffefffffffff0000002a00000000",
            INIT_16 => X"ffffffcbffffffff00000058000000000000002a00000000ffffffc9ffffffff",
            INIT_17 => X"ffffffe3fffffffffffffff3ffffffff00000053000000000000001400000000",
            INIT_18 => X"ffffffdaffffffffffffffd7ffffffff00000006000000000000002800000000",
            INIT_19 => X"0000000b00000000fffffff1fffffffffffffffcffffffff0000001500000000",
            INIT_1A => X"00000007000000000000000f00000000fffffff2fffffffffffffffdffffffff",
            INIT_1B => X"fffffffbfffffffffffffff9ffffffff0000003300000000ffffffd6ffffffff",
            INIT_1C => X"0000000000000000ffffffc3ffffffffffffffe6ffffffff0000000900000000",
            INIT_1D => X"0000000100000000ffffffeeffffffffffffffecffffffffffffffe1ffffffff",
            INIT_1E => X"0000001a00000000fffffff8fffffffffffffff9fffffffffffffffcffffffff",
            INIT_1F => X"fffffff9ffffffff000000170000000000000026000000000000001800000000",
            INIT_20 => X"fffffff8ffffffffffffffd8fffffffffffffffaffffffff0000000700000000",
            INIT_21 => X"fffffff8ffffffff0000001300000000fffffff3ffffffff0000000900000000",
            INIT_22 => X"ffffffe6ffffffff0000000a00000000ffffffecffffffff0000001800000000",
            INIT_23 => X"0000001f00000000fffffff4ffffffffffffffe7ffffffffffffffe7ffffffff",
            INIT_24 => X"ffffffecfffffffffffffffeffffffff0000000d000000000000000a00000000",
            INIT_25 => X"fffffff7ffffffffffffffedffffffff00000016000000000000000900000000",
            INIT_26 => X"000000080000000000000026000000000000000300000000fffffff9ffffffff",
            INIT_27 => X"ffffffe9ffffffff000000070000000000000020000000000000000f00000000",
            INIT_28 => X"fffffff4ffffffff000000070000000000000010000000000000000400000000",
            INIT_29 => X"ffffffdafffffffffffffffffffffffffffffff6ffffffff0000000900000000",
            INIT_2A => X"ffffffa8ffffffffffffffbeffffffffffffff99fffffffffffffff8ffffffff",
            INIT_2B => X"ffffffa4ffffffffffffffa9ffffffffffffff74ffffffffffffff8affffffff",
            INIT_2C => X"00000021000000000000001200000000ffffffccffffffffffffffa0ffffffff",
            INIT_2D => X"0000001500000000000000370000000000000010000000000000002200000000",
            INIT_2E => X"00000024000000000000001a00000000fffffffbffffffff0000002b00000000",
            INIT_2F => X"00000000000000000000002200000000fffffffeffffffffffffffe3ffffffff",
            INIT_30 => X"ffffffe4fffffffffffffffcfffffffffffffff6ffffffffffffffe4ffffffff",
            INIT_31 => X"0000005f000000000000002c0000000000000029000000000000004600000000",
            INIT_32 => X"0000002900000000000000510000000000000004000000000000001500000000",
            INIT_33 => X"fffffff8ffffffff00000004000000000000000d00000000fffffff1ffffffff",
            INIT_34 => X"000000020000000000000006000000000000001d000000000000000000000000",
            INIT_35 => X"ffffffffffffffffffffffe2ffffffffffffffeeffffffffffffffe6ffffffff",
            INIT_36 => X"0000000b00000000fffffff3fffffffffffffffcffffffffffffffebffffffff",
            INIT_37 => X"fffffff1fffffffffffffff6fffffffffffffffdffffffff0000001900000000",
            INIT_38 => X"0000000a0000000000000017000000000000001f000000000000002400000000",
            INIT_39 => X"fffffff7ffffffff0000003c0000000000000028000000000000000b00000000",
            INIT_3A => X"ffffffcfffffffff0000000300000000fffffffdfffffffffffffffdffffffff",
            INIT_3B => X"ffffffc8ffffffffffffffc3ffffffffffffffd7ffffffffffffffa1ffffffff",
            INIT_3C => X"ffffffffffffffffffffffe9fffffffffffffff5ffffffff0000001600000000",
            INIT_3D => X"fffffff9ffffffffffffffedfffffffffffffff0ffffffffffffffedffffffff",
            INIT_3E => X"ffffffe2ffffffffffffffd2ffffffff0000002500000000fffffff7ffffffff",
            INIT_3F => X"ffffffcfffffffffffffffa0ffffffffffffffd2ffffffffffffffe5ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdcfffffffffffffff9ffffffffffffffc9fffffffffffffff0ffffffff",
            INIT_41 => X"00000004000000000000001800000000ffffffdfffffffffffffffd8ffffffff",
            INIT_42 => X"ffffffebffffffffffffffeaffffffff0000000900000000ffffffe5ffffffff",
            INIT_43 => X"0000000c00000000ffffffefffffffffffffffe5ffffffffffffffe8ffffffff",
            INIT_44 => X"0000001d000000000000001b00000000ffffffeaffffffff0000000900000000",
            INIT_45 => X"00000002000000000000001b000000000000000d000000000000001000000000",
            INIT_46 => X"00000015000000000000001300000000fffffff5fffffffffffffffaffffffff",
            INIT_47 => X"fffffffffffffffffffffffefffffffffffffffcffffffff0000000e00000000",
            INIT_48 => X"00000002000000000000000700000000ffffffe8ffffffffffffffe4ffffffff",
            INIT_49 => X"ffffffe8fffffffffffffff2ffffffffffffffe1fffffffffffffff8ffffffff",
            INIT_4A => X"ffffffe8ffffffff0000001400000000ffffffd9fffffffffffffff5ffffffff",
            INIT_4B => X"0000000c0000000000000018000000000000002b00000000ffffffe8ffffffff",
            INIT_4C => X"ffffffb1ffffffffffffffefffffffffffffffd3ffffffffffffffb0ffffffff",
            INIT_4D => X"ffffffeeffffffffffffffe0fffffffffffffff0ffffffffffffffd7ffffffff",
            INIT_4E => X"ffffffd6ffffffffffffffd9fffffffffffffff9ffffffff0000000f00000000",
            INIT_4F => X"0000000d000000000000000300000000ffffffecfffffffffffffff8ffffffff",
            INIT_50 => X"0000002900000000fffffff0ffffffff0000000600000000fffffffeffffffff",
            INIT_51 => X"fffffff6ffffffff0000000b00000000fffffff6ffffffff0000001900000000",
            INIT_52 => X"0000000500000000ffffffe4ffffffffffffffebfffffffffffffff4ffffffff",
            INIT_53 => X"00000017000000000000000500000000fffffffeffffffff0000000a00000000",
            INIT_54 => X"00000005000000000000001e000000000000000f00000000fffffffaffffffff",
            INIT_55 => X"00000014000000000000000700000000fffffffcfffffffffffffff8ffffffff",
            INIT_56 => X"fffffffdffffffff0000001c00000000ffffffedffffffff0000000600000000",
            INIT_57 => X"fffffffcfffffffffffffff2ffffffffffffffe9ffffffffffffffdeffffffff",
            INIT_58 => X"0000001200000000ffffffecfffffffffffffff6ffffffffffffffe9ffffffff",
            INIT_59 => X"ffffffe5ffffffffffffffefffffffff0000000a00000000fffffffbffffffff",
            INIT_5A => X"0000000800000000fffffff9ffffffffffffffe4fffffffffffffff4ffffffff",
            INIT_5B => X"00000027000000000000001400000000fffffff6fffffffffffffff3ffffffff",
            INIT_5C => X"fffffff6ffffffffffffffebffffffff00000012000000000000000500000000",
            INIT_5D => X"00000004000000000000000800000000fffffff0ffffffff0000001200000000",
            INIT_5E => X"00000000000000000000000f00000000fffffffffffffffffffffffeffffffff",
            INIT_5F => X"0000001000000000ffffffd0ffffffff0000002a00000000fffffff1ffffffff",
            INIT_60 => X"000000200000000000000014000000000000001d000000000000003100000000",
            INIT_61 => X"000000080000000000000009000000000000001b000000000000000800000000",
            INIT_62 => X"fffffffefffffffffffffff7fffffffffffffff1ffffffffffffffedffffffff",
            INIT_63 => X"000000060000000000000006000000000000001e000000000000001400000000",
            INIT_64 => X"fffffffdffffffff0000003a0000000000000001000000000000000000000000",
            INIT_65 => X"ffffffe7ffffffff00000003000000000000000500000000ffffffeaffffffff",
            INIT_66 => X"0000000000000000fffffffcffffffff00000014000000000000001f00000000",
            INIT_67 => X"0000000300000000000000110000000000000029000000000000003400000000",
            INIT_68 => X"0000002100000000000000090000000000000003000000000000003100000000",
            INIT_69 => X"00000015000000000000000900000000ffffffdbffffffff0000000c00000000",
            INIT_6A => X"fffffff5ffffffff0000002e000000000000000200000000ffffffe1ffffffff",
            INIT_6B => X"0000001100000000000000030000000000000000000000000000000c00000000",
            INIT_6C => X"fffffff7ffffffff0000000d000000000000000d000000000000000f00000000",
            INIT_6D => X"0000001700000000ffffffddfffffffffffffff6ffffffff0000000200000000",
            INIT_6E => X"00000017000000000000001a0000000000000015000000000000000000000000",
            INIT_6F => X"0000000a0000000000000018000000000000002d000000000000001e00000000",
            INIT_70 => X"fffffff7ffffffffffffffdfffffffff00000001000000000000000800000000",
            INIT_71 => X"fffffff8ffffffff00000007000000000000000a00000000ffffffebffffffff",
            INIT_72 => X"fffffff3ffffffff0000000a0000000000000004000000000000000000000000",
            INIT_73 => X"0000000500000000ffffffedffffffff0000002d000000000000002300000000",
            INIT_74 => X"0000002e000000000000000b00000000ffffffaeffffffffffffffceffffffff",
            INIT_75 => X"fffffff3ffffffff00000006000000000000001e000000000000005600000000",
            INIT_76 => X"0000000400000000ffffffefffffffffffffffe4ffffffffffffffedffffffff",
            INIT_77 => X"0000000c00000000ffffffc6ffffffff00000000000000000000001500000000",
            INIT_78 => X"0000001300000000fffffff2ffffffffffffffbaffffffff0000002a00000000",
            INIT_79 => X"fffffff3ffffffff00000022000000000000001b000000000000003700000000",
            INIT_7A => X"ffffffd7fffffffffffffff1ffffffffffffffd8ffffffff0000000600000000",
            INIT_7B => X"ffffffe1ffffffffffffffb3ffffffffffffffd9ffffffffffffffd0ffffffff",
            INIT_7C => X"00000029000000000000000f00000000ffffffb1ffffffff0000000c00000000",
            INIT_7D => X"fffffff3ffffffff000000190000000000000044000000000000002900000000",
            INIT_7E => X"0000001700000000ffffffeaffffffffffffffdfffffffff0000001200000000",
            INIT_7F => X"0000000b00000000ffffffe1ffffffffffffffe3fffffffffffffff4ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE6;


    MEM_IWGHT_LAYER2_INSTANCE7 : if BRAM_NAME = "iwght_layer2_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001f00000000fffffff1ffffffff00000013000000000000000500000000",
            INIT_01 => X"ffffffeaffffffffffffffefffffffff0000000200000000ffffffffffffffff",
            INIT_02 => X"00000028000000000000001a000000000000001100000000ffffffedffffffff",
            INIT_03 => X"ffffffd5ffffffffffffffe2ffffffff0000002100000000fffffffeffffffff",
            INIT_04 => X"fffffff0ffffffffffffffe8ffffffffffffffd5ffffffffffffffe5ffffffff",
            INIT_05 => X"fffffff5ffffffffffffffd7ffffffffffffffe3ffffffffffffffeeffffffff",
            INIT_06 => X"00000000000000000000001100000000fffffffbffffffffffffffe0ffffffff",
            INIT_07 => X"ffffffedfffffffffffffffeffffffff0000003300000000ffffffe4ffffffff",
            INIT_08 => X"0000001700000000ffffffddffffffffffffffeffffffffffffffff9ffffffff",
            INIT_09 => X"ffffffdefffffffffffffff7fffffffffffffff2fffffffffffffff2ffffffff",
            INIT_0A => X"fffffff8ffffffffffffffe8fffffffffffffffbffffffffffffffe9ffffffff",
            INIT_0B => X"0000001200000000ffffffd6ffffffffffffffd8fffffffffffffffaffffffff",
            INIT_0C => X"0000001e00000000000000080000000000000008000000000000000400000000",
            INIT_0D => X"0000003100000000000000050000000000000005000000000000003100000000",
            INIT_0E => X"ffffffe7ffffffff000000090000000000000015000000000000001e00000000",
            INIT_0F => X"ffffffadffffffff0000000300000000ffffffeaffffffff0000000300000000",
            INIT_10 => X"0000000900000000ffffffccffffffff0000004400000000ffffffaeffffffff",
            INIT_11 => X"00000000000000000000003d000000000000001d000000000000003600000000",
            INIT_12 => X"00000011000000000000000c0000000000000019000000000000000c00000000",
            INIT_13 => X"0000001800000000ffffffe5ffffffff00000003000000000000001500000000",
            INIT_14 => X"0000000300000000ffffffdbffffffffffffffe9ffffffff0000000d00000000",
            INIT_15 => X"ffffffdcffffffff0000001e00000000ffffffbfffffffff0000000c00000000",
            INIT_16 => X"0000000200000000fffffff6ffffffffffffffd7ffffffffffffffd6ffffffff",
            INIT_17 => X"ffffffe2fffffffffffffff9fffffffffffffff6ffffffffffffffc5ffffffff",
            INIT_18 => X"0000003400000000fffffffcffffffff0000002600000000ffffffdaffffffff",
            INIT_19 => X"0000004d000000000000004d0000000000000010000000000000002500000000",
            INIT_1A => X"0000000100000000ffffffedffffffffffffffffffffffff0000001c00000000",
            INIT_1B => X"ffffffd8ffffffff0000001000000000ffffffebffffffffffffffdfffffffff",
            INIT_1C => X"0000001800000000ffffffffffffffff00000026000000000000002500000000",
            INIT_1D => X"ffffffecffffffff0000000b00000000ffffffeeffffffff0000002400000000",
            INIT_1E => X"ffffffecffffffff00000000000000000000000000000000ffffffdcffffffff",
            INIT_1F => X"0000001600000000ffffffe8ffffffffffffffedfffffffffffffffdffffffff",
            INIT_20 => X"0000000c000000000000002000000000ffffffe2fffffffffffffff1ffffffff",
            INIT_21 => X"fffffffeffffffffffffffcaffffffff0000001f000000000000000700000000",
            INIT_22 => X"0000000000000000fffffffaffffffffffffffdffffffffffffffff4ffffffff",
            INIT_23 => X"fffffff4ffffffff0000000c00000000fffffff5ffffffffffffffecffffffff",
            INIT_24 => X"00000010000000000000000c00000000ffffffebffffffffffffffbcffffffff",
            INIT_25 => X"000000280000000000000011000000000000002b000000000000001b00000000",
            INIT_26 => X"000000260000000000000031000000000000006d000000000000001000000000",
            INIT_27 => X"ffffffe5ffffffffffffffdcfffffffffffffff9ffffffff0000003b00000000",
            INIT_28 => X"00000028000000000000001300000000fffffff8ffffffffffffffe5ffffffff",
            INIT_29 => X"fffffff0fffffffffffffff1ffffffff0000000400000000fffffffbffffffff",
            INIT_2A => X"fffffffffffffffffffffff6ffffffffffffffbfffffffffffffffecffffffff",
            INIT_2B => X"0000001a00000000fffffff2ffffffff00000017000000000000000900000000",
            INIT_2C => X"0000000b000000000000000600000000fffffff9ffffffffffffffedffffffff",
            INIT_2D => X"0000000e000000000000000500000000ffffffe0ffffffffffffffdbffffffff",
            INIT_2E => X"fffffff7ffffffff00000006000000000000001000000000fffffff3ffffffff",
            INIT_2F => X"fffffffdffffffff000000350000000000000013000000000000001800000000",
            INIT_30 => X"fffffff9fffffffffffffff1ffffffff0000000a000000000000000f00000000",
            INIT_31 => X"ffffffdeffffffffffffffdaffffffff0000000200000000ffffffffffffffff",
            INIT_32 => X"ffffffecffffffffffffffe2ffffffff00000019000000000000000800000000",
            INIT_33 => X"ffffffdeffffffff0000000600000000fffffff7fffffffffffffff7ffffffff",
            INIT_34 => X"0000000000000000ffffffe5ffffffff0000000600000000fffffffaffffffff",
            INIT_35 => X"fffffffaffffffff000000110000000000000005000000000000000200000000",
            INIT_36 => X"0000001b00000000fffffffeffffffff0000000b000000000000000100000000",
            INIT_37 => X"000000280000000000000018000000000000001f000000000000001d00000000",
            INIT_38 => X"fffffff7ffffffff0000000100000000fffffffbffffffff0000000800000000",
            INIT_39 => X"fffffff9ffffffff000000140000000000000000000000000000001d00000000",
            INIT_3A => X"fffffff8ffffffff0000001000000000fffffff1fffffffffffffffeffffffff",
            INIT_3B => X"ffffffeefffffffffffffff8fffffffffffffff7fffffffffffffffaffffffff",
            INIT_3C => X"fffffff8ffffffffffffffe0ffffffff0000002300000000fffffff5ffffffff",
            INIT_3D => X"00000017000000000000002a00000000fffffff7ffffffffffffffcaffffffff",
            INIT_3E => X"0000001c00000000000000590000000000000060000000000000005100000000",
            INIT_3F => X"ffffffe6ffffffffffffffdbffffffff00000008000000000000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdbfffffffffffffff2ffffffff0000001900000000fffffff5ffffffff",
            INIT_41 => X"0000002500000000ffffffb1ffffffffffffffd9fffffffffffffff8ffffffff",
            INIT_42 => X"00000027000000000000004f00000000ffffffd4ffffffff0000000d00000000",
            INIT_43 => X"0000001300000000000000150000000000000007000000000000001400000000",
            INIT_44 => X"0000000a000000000000000300000000ffffffddffffffffffffffecffffffff",
            INIT_45 => X"0000000a00000000ffffffeeffffffff0000000100000000ffffffe6ffffffff",
            INIT_46 => X"0000000800000000ffffffe1ffffffffffffffe3ffffffff0000001900000000",
            INIT_47 => X"fffffff9fffffffffffffff4fffffffffffffff2ffffffff0000000b00000000",
            INIT_48 => X"0000000200000000ffffffedffffffff0000001f00000000ffffffd8ffffffff",
            INIT_49 => X"0000001e0000000000000016000000000000000c000000000000000000000000",
            INIT_4A => X"0000001400000000ffffffbbffffffffffffffd8ffffffff0000000400000000",
            INIT_4B => X"ffffffedffffffff0000001c00000000ffffffd9ffffffff0000001600000000",
            INIT_4C => X"fffffffefffffffffffffffaffffffffffffffecffffffff0000000000000000",
            INIT_4D => X"0000000f00000000fffffff3ffffffff0000002f000000000000002700000000",
            INIT_4E => X"fffffff2ffffffffffffffe2ffffffffffffffdbffffffff0000000b00000000",
            INIT_4F => X"fffffff8ffffffff00000007000000000000000600000000ffffffc4ffffffff",
            INIT_50 => X"ffffffeffffffffffffffffefffffffffffffff0ffffffffffffffdaffffffff",
            INIT_51 => X"fffffffeffffffffffffffeeffffffff0000001d00000000fffffff1ffffffff",
            INIT_52 => X"fffffffeffffffff0000002c0000000000000001000000000000003200000000",
            INIT_53 => X"fffffffaffffffff00000002000000000000000e00000000ffffffefffffffff",
            INIT_54 => X"ffffffdcffffffffffffffd1ffffffff0000001400000000fffffff5ffffffff",
            INIT_55 => X"0000002d0000000000000008000000000000000a00000000fffffff9ffffffff",
            INIT_56 => X"0000000c00000000ffffffdfffffffff00000018000000000000000b00000000",
            INIT_57 => X"0000000e00000000000000150000000000000006000000000000001300000000",
            INIT_58 => X"0000000000000000000000020000000000000001000000000000001000000000",
            INIT_59 => X"ffffffe4ffffffff0000001000000000ffffffe2ffffffff0000001200000000",
            INIT_5A => X"fffffffdffffffffffffffedffffffff0000000a00000000ffffffd5ffffffff",
            INIT_5B => X"ffffffd3ffffffff00000000000000000000001200000000fffffff6ffffffff",
            INIT_5C => X"00000071000000000000002d000000000000002f000000000000002500000000",
            INIT_5D => X"fffffffcffffffff000000230000000000000060000000000000004a00000000",
            INIT_5E => X"00000005000000000000000d00000000ffffffe5ffffffff0000001f00000000",
            INIT_5F => X"00000012000000000000000c0000000000000015000000000000000500000000",
            INIT_60 => X"0000000100000000ffffffffffffffffffffffedffffffff0000000700000000",
            INIT_61 => X"fffffff3ffffffffffffffd6ffffffff0000000200000000fffffff2ffffffff",
            INIT_62 => X"fffffff7fffffffffffffff0ffffffffffffffdbffffffffffffffdbffffffff",
            INIT_63 => X"ffffffc7fffffffffffffff9ffffffff0000002400000000ffffffe2ffffffff",
            INIT_64 => X"fffffffbfffffffffffffff1fffffffffffffff7ffffffffffffffd0ffffffff",
            INIT_65 => X"fffffff2ffffffff0000002a0000000000000013000000000000000600000000",
            INIT_66 => X"00000004000000000000000100000000ffffffe1ffffffffffffffcaffffffff",
            INIT_67 => X"0000001f00000000fffffffdfffffffffffffff4ffffffff0000000400000000",
            INIT_68 => X"0000001700000000ffffffe3fffffffffffffff9ffffffffffffffcdffffffff",
            INIT_69 => X"fffffff8fffffffffffffff3fffffffffffffffefffffffffffffffbffffffff",
            INIT_6A => X"fffffff3ffffffff0000000c000000000000002400000000fffffff0ffffffff",
            INIT_6B => X"0000000000000000ffffffefffffffff00000003000000000000001500000000",
            INIT_6C => X"fffffff7ffffffff00000003000000000000001c00000000ffffffebffffffff",
            INIT_6D => X"fffffff0ffffffffffffffc1ffffffffffffffeaffffffff0000002400000000",
            INIT_6E => X"fffffff5ffffffffffffffe3ffffffff00000010000000000000000900000000",
            INIT_6F => X"00000002000000000000001400000000ffffffddffffffffffffffeeffffffff",
            INIT_70 => X"00000000000000000000000000000000ffffffffffffffff0000000000000000",
            INIT_71 => X"00000013000000000000000300000000ffffffebffffffff0000000800000000",
            INIT_72 => X"0000000f00000000fffffffcffffffff00000015000000000000002600000000",
            INIT_73 => X"fffffff7ffffffff0000002a000000000000000e00000000ffffffe1ffffffff",
            INIT_74 => X"ffffffd8ffffffffffffffd3ffffffffffffffecffffffff0000000300000000",
            INIT_75 => X"ffffffeefffffffffffffff3ffffffff0000000700000000ffffffe7ffffffff",
            INIT_76 => X"00000027000000000000001d000000000000001400000000fffffff2ffffffff",
            INIT_77 => X"fffffff9fffffffffffffffcfffffffffffffff5ffffffffffffffc2ffffffff",
            INIT_78 => X"fffffff3ffffffff0000002300000000fffffffbfffffffffffffff6ffffffff",
            INIT_79 => X"0000002d000000000000003200000000fffffffeffffffffffffffe5ffffffff",
            INIT_7A => X"ffffffe9ffffffff0000004200000000fffffff3fffffffffffffffaffffffff",
            INIT_7B => X"000000000000000000000032000000000000001400000000fffffffbffffffff",
            INIT_7C => X"fffffff2ffffffffffffffd7fffffffffffffffaffffffff0000002700000000",
            INIT_7D => X"ffffffeffffffffffffffff6fffffffffffffff3fffffffffffffff9ffffffff",
            INIT_7E => X"0000001d00000000fffffff8fffffffffffffff9ffffffff0000001900000000",
            INIT_7F => X"fffffff0fffffffffffffffdffffffff0000000a000000000000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE7;


    MEM_IWGHT_LAYER2_INSTANCE8 : if BRAM_NAME = "iwght_layer2_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000009000000000000001e00000000ffffffecffffffffffffffefffffffff",
            INIT_01 => X"0000001c000000000000002a000000000000000b000000000000001400000000",
            INIT_02 => X"fffffffdffffffff000000130000000000000027000000000000001c00000000",
            INIT_03 => X"ffffffd6ffffffff0000000c0000000000000006000000000000002c00000000",
            INIT_04 => X"fffffffeffffffff0000000e000000000000000d00000000ffffffd4ffffffff",
            INIT_05 => X"0000003400000000000000520000000000000014000000000000001100000000",
            INIT_06 => X"0000002c00000000000000270000000000000021000000000000004100000000",
            INIT_07 => X"0000003d000000000000002b000000000000001f000000000000003800000000",
            INIT_08 => X"ffffffdefffffffffffffffcffffffff00000002000000000000000e00000000",
            INIT_09 => X"0000003400000000ffffffe0fffffffffffffffcffffffff0000002d00000000",
            INIT_0A => X"fffffff7ffffffff0000000500000000ffffffe3ffffffff0000005000000000",
            INIT_0B => X"00000032000000000000000c00000000fffffff3ffffffffffffffe7ffffffff",
            INIT_0C => X"0000002f000000000000000f00000000fffffff7ffffffffffffffffffffffff",
            INIT_0D => X"ffffffddffffffff00000002000000000000001d000000000000000f00000000",
            INIT_0E => X"ffffffbaffffffffffffffd6ffffffffffffffd6fffffffffffffff9ffffffff",
            INIT_0F => X"fffffffcfffffffffffffff4ffffffff0000000f000000000000000600000000",
            INIT_10 => X"00000026000000000000000b000000000000000200000000ffffffe7ffffffff",
            INIT_11 => X"00000003000000000000001e000000000000001c000000000000000a00000000",
            INIT_12 => X"fffffffefffffffffffffff0ffffffff00000024000000000000002c00000000",
            INIT_13 => X"ffffffe0ffffffffffffffe4fffffffffffffff4ffffffff0000000200000000",
            INIT_14 => X"00000023000000000000001e0000000000000008000000000000000400000000",
            INIT_15 => X"00000000000000000000000000000000ffffffdfffffffffffffffdaffffffff",
            INIT_16 => X"fffffff3ffffffff0000002500000000fffffffdfffffffffffffff3ffffffff",
            INIT_17 => X"ffffffe5fffffffffffffff0ffffffff0000000200000000ffffffe6ffffffff",
            INIT_18 => X"0000000f00000000ffffffe9ffffffffffffffd6fffffffffffffff8ffffffff",
            INIT_19 => X"0000000900000000ffffffddffffffff0000000200000000ffffffdfffffffff",
            INIT_1A => X"ffffffeaffffffffffffffdcffffffff0000001800000000fffffff3ffffffff",
            INIT_1B => X"ffffffc8ffffffff00000007000000000000000500000000ffffffd2ffffffff",
            INIT_1C => X"0000000700000000ffffffe6fffffffffffffff7ffffffffffffffe3ffffffff",
            INIT_1D => X"fffffff2ffffffffffffffcefffffffffffffff6ffffffff0000000400000000",
            INIT_1E => X"0000001c00000000000000050000000000000001000000000000002900000000",
            INIT_1F => X"0000001b00000000fffffffdffffffff0000001e000000000000001500000000",
            INIT_20 => X"00000017000000000000000100000000ffffffe0ffffffff0000000100000000",
            INIT_21 => X"ffffffc5ffffffff0000001a000000000000003d000000000000004200000000",
            INIT_22 => X"ffffffc8ffffffffffffffa3ffffffff0000000a00000000fffffff3ffffffff",
            INIT_23 => X"ffffffefffffffff0000000d00000000ffffffe1ffffffff0000001000000000",
            INIT_24 => X"0000000a00000000fffffff6ffffffffffffffd1ffffffff0000004300000000",
            INIT_25 => X"ffffffffffffffffffffffebffffffffffffffc2ffffffffffffffebffffffff",
            INIT_26 => X"0000001c00000000fffffff9ffffffffffffffe2ffffffff0000002600000000",
            INIT_27 => X"00000022000000000000000100000000fffffff7ffffffff0000000900000000",
            INIT_28 => X"ffffffe1ffffffffffffffd3ffffffff00000002000000000000000c00000000",
            INIT_29 => X"ffffffdfffffffffffffffe3ffffffffffffffbeffffffff0000001e00000000",
            INIT_2A => X"fffffff5ffffffff0000000400000000fffffff9ffffffff0000002000000000",
            INIT_2B => X"fffffff3ffffffffffffffddfffffffffffffff3ffffffff0000000500000000",
            INIT_2C => X"fffffff1ffffffffffffffe8ffffffff0000001c000000000000001100000000",
            INIT_2D => X"ffffffd7ffffffff0000001f00000000fffffff1ffffffff0000002300000000",
            INIT_2E => X"fffffff5ffffffffffffffeaffffffff0000001800000000ffffffe0ffffffff",
            INIT_2F => X"00000023000000000000002a0000000000000001000000000000001000000000",
            INIT_30 => X"0000000b000000000000001600000000fffffffdffffffffffffffe3ffffffff",
            INIT_31 => X"fffffff7fffffffffffffff8ffffffff00000006000000000000001100000000",
            INIT_32 => X"0000001e00000000fffffff4ffffffffffffffccffffffff0000000a00000000",
            INIT_33 => X"0000003a0000000000000024000000000000003400000000fffffff0ffffffff",
            INIT_34 => X"ffffffd6ffffffff0000000100000000fffffff8fffffffffffffff8ffffffff",
            INIT_35 => X"ffffffddffffffffffffffe7ffffffff0000000100000000ffffffc5ffffffff",
            INIT_36 => X"00000025000000000000004b000000000000002900000000fffffff2ffffffff",
            INIT_37 => X"fffffff5ffffffffffffffedffffffff00000020000000000000003200000000",
            INIT_38 => X"ffffffe0ffffffffffffffe5fffffffffffffffcfffffffffffffffbffffffff",
            INIT_39 => X"ffffffeeffffffffffffffeaffffffff00000012000000000000001e00000000",
            INIT_3A => X"ffffffecfffffffffffffffeffffffff0000000000000000fffffff5ffffffff",
            INIT_3B => X"0000002800000000ffffffedfffffffffffffffcffffffff0000003200000000",
            INIT_3C => X"ffffffdfffffffff00000005000000000000001d000000000000001400000000",
            INIT_3D => X"0000000400000000ffffffe6ffffffff0000000c00000000fffffff6ffffffff",
            INIT_3E => X"0000001100000000ffffffeaffffffff0000000c000000000000001700000000",
            INIT_3F => X"0000001500000000000000030000000000000058000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001c000000000000001900000000ffffffe7ffffffff0000005c00000000",
            INIT_41 => X"0000000d00000000ffffff99ffffffffffffffc0ffffffffffffffd0ffffffff",
            INIT_42 => X"fffffffefffffffffffffff6ffffffffffffffe3ffffffffffffffe7ffffffff",
            INIT_43 => X"fffffff8ffffffff0000000500000000fffffff6ffffffff0000001500000000",
            INIT_44 => X"00000002000000000000000000000000fffffff4ffffffff0000000d00000000",
            INIT_45 => X"0000000000000000000000290000000000000006000000000000000a00000000",
            INIT_46 => X"fffffffafffffffffffffff2ffffffff00000013000000000000000f00000000",
            INIT_47 => X"fffffffefffffffffffffffeffffffff00000004000000000000002000000000",
            INIT_48 => X"000000020000000000000009000000000000000900000000fffffff4ffffffff",
            INIT_49 => X"0000000b000000000000000c0000000000000017000000000000001300000000",
            INIT_4A => X"00000036000000000000001b000000000000002a000000000000000d00000000",
            INIT_4B => X"0000000e0000000000000010000000000000000000000000fffffff4ffffffff",
            INIT_4C => X"0000000a0000000000000039000000000000001d000000000000002100000000",
            INIT_4D => X"ffffffffffffffff000000190000000000000042000000000000002500000000",
            INIT_4E => X"ffffffdcffffffff000000170000000000000018000000000000001500000000",
            INIT_4F => X"ffffffcdffffffffffffffd0ffffffff0000001300000000ffffffe1ffffffff",
            INIT_50 => X"ffffffc5ffffffffffffffb9ffffffffffffffbfffffffffffffffe1ffffffff",
            INIT_51 => X"00000010000000000000002c0000000000000021000000000000001b00000000",
            INIT_52 => X"fffffffaffffffffffffffe8ffffffff00000040000000000000004300000000",
            INIT_53 => X"0000000f000000000000000c00000000fffffff6ffffffff0000000500000000",
            INIT_54 => X"0000001e0000000000000000000000000000001500000000ffffffdbffffffff",
            INIT_55 => X"0000001800000000fffffffdfffffffffffffffafffffffffffffff6ffffffff",
            INIT_56 => X"fffffffbffffffff000000180000000000000002000000000000003200000000",
            INIT_57 => X"0000000000000000ffffffeaffffffffffffffe6fffffffffffffffeffffffff",
            INIT_58 => X"00000007000000000000001300000000ffffffeaffffffffffffffffffffffff",
            INIT_59 => X"00000018000000000000000a00000000ffffffe8ffffffff0000000000000000",
            INIT_5A => X"0000001e00000000fffffff5ffffffffffffffd0ffffffff0000000d00000000",
            INIT_5B => X"fffffffbffffffff0000002800000000fffffff0ffffffff0000000a00000000",
            INIT_5C => X"00000000000000000000001a0000000000000005000000000000000000000000",
            INIT_5D => X"ffffffefffffffffffffffebffffffff0000000300000000fffffffcffffffff",
            INIT_5E => X"fffffff0ffffffff00000015000000000000000c00000000fffffff0ffffffff",
            INIT_5F => X"0000001b000000000000001500000000fffffffaffffffff0000000c00000000",
            INIT_60 => X"0000001f000000000000001a0000000000000017000000000000001b00000000",
            INIT_61 => X"0000000d00000000ffffffc7ffffffff00000027000000000000001300000000",
            INIT_62 => X"ffffffe6ffffffff0000002d000000000000000300000000fffffff2ffffffff",
            INIT_63 => X"00000000000000000000002c000000000000000e00000000ffffffffffffffff",
            INIT_64 => X"ffffffe1ffffffffffffffe1ffffffff0000000c00000000ffffffe7ffffffff",
            INIT_65 => X"00000006000000000000000d00000000fffffff7ffffffffffffffd1ffffffff",
            INIT_66 => X"ffffffddffffffff000000090000000000000019000000000000000f00000000",
            INIT_67 => X"0000001500000000000000170000000000000011000000000000001500000000",
            INIT_68 => X"fffffff3ffffffffffffffeaffffffffffffffcaffffffff0000003400000000",
            INIT_69 => X"0000000c00000000fffffff9ffffffff0000001100000000ffffffffffffffff",
            INIT_6A => X"0000000d00000000000000050000000000000033000000000000002200000000",
            INIT_6B => X"ffffffe9ffffffff0000000000000000fffffff4ffffffff0000000900000000",
            INIT_6C => X"fffffff4ffffffffffffffe5ffffffff00000034000000000000000200000000",
            INIT_6D => X"0000002200000000ffffffffffffffff0000002f000000000000000600000000",
            INIT_6E => X"0000001c000000000000001b0000000000000025000000000000001200000000",
            INIT_6F => X"ffffffd6fffffffffffffff6ffffffff0000001a00000000fffffff1ffffffff",
            INIT_70 => X"ffffffccffffffffffffff9bffffffffffffffeaffffffff0000000100000000",
            INIT_71 => X"ffffffccfffffffffffffff0ffffffffffffffc7ffffffffffffffccffffffff",
            INIT_72 => X"0000000000000000ffffffd6ffffffff0000001500000000ffffffd3ffffffff",
            INIT_73 => X"fffffffbfffffffffffffff8ffffffff0000000e00000000fffffffbffffffff",
            INIT_74 => X"fffffff2ffffffff00000008000000000000000b000000000000000600000000",
            INIT_75 => X"ffffffdaffffffffffffffdaffffffff0000000000000000ffffffeeffffffff",
            INIT_76 => X"0000000c00000000ffffffecfffffffffffffff1ffffffffffffffd6ffffffff",
            INIT_77 => X"fffffff8ffffffff0000001b0000000000000016000000000000000800000000",
            INIT_78 => X"0000001d00000000ffffffe5ffffffffffffffedffffffffffffffe5ffffffff",
            INIT_79 => X"00000024000000000000001b000000000000000e00000000fffffff9ffffffff",
            INIT_7A => X"0000001f00000000ffffffebfffffffffffffffdffffffff0000003500000000",
            INIT_7B => X"ffffffdbffffffffffffffebffffffffffffffdeffffffff0000000500000000",
            INIT_7C => X"0000000d00000000ffffffdcffffffff0000000e000000000000001200000000",
            INIT_7D => X"ffffffe1ffffffff00000020000000000000001000000000ffffffe7ffffffff",
            INIT_7E => X"0000000700000000ffffffd5ffffffffffffffc2fffffffffffffff3ffffffff",
            INIT_7F => X"fffffff0ffffffff0000001d00000000ffffffcdffffffffffffffe9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE8;


    MEM_IWGHT_LAYER2_INSTANCE9 : if BRAM_NAME = "iwght_layer2_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffcbffffffffffffffeefffffffffffffff8ffffffff0000001900000000",
            INIT_01 => X"ffffffebfffffffffffffffdffffffff0000000d000000000000001b00000000",
            INIT_02 => X"00000025000000000000001900000000fffffff6ffffffff0000000e00000000",
            INIT_03 => X"ffffffe7fffffffffffffff4ffffffff0000001900000000fffffff9ffffffff",
            INIT_04 => X"fffffff5ffffffffffffffe0ffffffff0000000a00000000fffffff1ffffffff",
            INIT_05 => X"ffffffe1fffffffffffffffafffffffffffffffefffffffffffffff2ffffffff",
            INIT_06 => X"ffffffd5ffffffffffffffdaffffffff0000000200000000fffffff2ffffffff",
            INIT_07 => X"ffffffc0ffffffff0000001000000000ffffffdbffffffffffffffdaffffffff",
            INIT_08 => X"ffffffd4ffffffffffffffddffffffffffffffeaffffffffffffffbbffffffff",
            INIT_09 => X"fffffff3ffffffffffffffe7ffffffffffffffe6ffffffffffffffc4ffffffff",
            INIT_0A => X"0000000300000000ffffffddfffffffffffffff2fffffffffffffff1ffffffff",
            INIT_0B => X"ffffffe5ffffffffffffffe9ffffffffffffffebffffffff0000000100000000",
            INIT_0C => X"ffffffd1ffffffffffffffdbffffffffffffffd9ffffffffffffffc5ffffffff",
            INIT_0D => X"0000002500000000ffffffeeffffffff0000000f00000000fffffff1ffffffff",
            INIT_0E => X"00000000000000000000000e0000000000000043000000000000003900000000",
            INIT_0F => X"ffffffd4ffffffffffffffdcffffffffffffffecffffffff0000000000000000",
            INIT_10 => X"fffffff1ffffffff00000016000000000000000d00000000fffffff0ffffffff",
            INIT_11 => X"ffffffffffffffff00000005000000000000001500000000fffffff9ffffffff",
            INIT_12 => X"ffffffe9ffffffffffffffe2ffffffffffffffdffffffffffffffffbffffffff",
            INIT_13 => X"0000001f0000000000000027000000000000000100000000fffffffaffffffff",
            INIT_14 => X"ffffffc7ffffffff0000000e0000000000000014000000000000000500000000",
            INIT_15 => X"ffffffa6ffffffffffffffb3ffffffffffffffc6ffffffffffffffe1ffffffff",
            INIT_16 => X"0000001b00000000ffffffa9ffffffffffffffa9ffffffffffffffe4ffffffff",
            INIT_17 => X"ffffffc5fffffffffffffff2ffffffffffffffb3ffffffffffffffb6ffffffff",
            INIT_18 => X"ffffff94ffffffff0000001e000000000000001900000000ffffffa7ffffffff",
            INIT_19 => X"ffffffa0ffffffffffffffc6ffffffffffffffa8ffffffffffffffdaffffffff",
            INIT_1A => X"fffffff4ffffffffffffffc4ffffffffffffff9bffffffffffffffc5ffffffff",
            INIT_1B => X"ffffffeaffffffffffffffd4ffffffffffffffc1ffffffffffffffa8ffffffff",
            INIT_1C => X"fffffffbffffffff0000001500000000fffffff0ffffffffffffffdaffffffff",
            INIT_1D => X"fffffff2fffffffffffffff4ffffffff00000010000000000000000b00000000",
            INIT_1E => X"ffffffe1ffffffff0000000b00000000fffffff3ffffffffffffffdbffffffff",
            INIT_1F => X"0000002900000000ffffffcaffffffff00000000000000000000000a00000000",
            INIT_20 => X"00000026000000000000003100000000fffffff1ffffffff0000001d00000000",
            INIT_21 => X"ffffffdbffffffff0000000a0000000000000027000000000000000c00000000",
            INIT_22 => X"ffffffe6ffffffff000000220000000000000000000000000000000100000000",
            INIT_23 => X"0000001700000000fffffffcffffffff00000015000000000000001700000000",
            INIT_24 => X"0000003600000000ffffffecffffffffffffffe9ffffffff0000000a00000000",
            INIT_25 => X"fffffff0ffffffff0000002700000000ffffffd4fffffffffffffffeffffffff",
            INIT_26 => X"0000000800000000fffffff6ffffffff00000047000000000000002100000000",
            INIT_27 => X"ffffffffffffffff0000000700000000fffffff2ffffffff0000001600000000",
            INIT_28 => X"ffffff86ffffffff0000000100000000fffffff8fffffffffffffffdffffffff",
            INIT_29 => X"ffffff7affffffffffffffd1ffffffffffffffbdffffffffffffff9cffffffff",
            INIT_2A => X"ffffffe8fffffffffffffff5ffffffff0000001500000000ffffffbeffffffff",
            INIT_2B => X"0000000300000000ffffffd1fffffffffffffff2ffffffffffffffe2ffffffff",
            INIT_2C => X"fffffffefffffffffffffff2fffffffffffffff4ffffffff0000000000000000",
            INIT_2D => X"ffffffe8ffffffff00000000000000000000000700000000fffffff5ffffffff",
            INIT_2E => X"0000001700000000ffffffecfffffffffffffff2fffffffffffffffeffffffff",
            INIT_2F => X"ffffffccffffffffffffffadffffffff0000000000000000ffffffe4ffffffff",
            INIT_30 => X"ffffffdfffffffffffffffaeffffffffffffffd4ffffffffffffffe3ffffffff",
            INIT_31 => X"ffffffd9ffffffffffffffd6ffffffffffffffe3ffffffffffffffd0ffffffff",
            INIT_32 => X"00000016000000000000001100000000fffffff5ffffffffffffffebffffffff",
            INIT_33 => X"0000001700000000000000130000000000000008000000000000002f00000000",
            INIT_34 => X"0000001200000000000000100000000000000026000000000000003300000000",
            INIT_35 => X"0000000c0000000000000002000000000000000c000000000000000200000000",
            INIT_36 => X"ffffffd8ffffffffffffffeefffffffffffffff1ffffffffffffffdeffffffff",
            INIT_37 => X"fffffffafffffffffffffff6ffffffffffffffe4fffffffffffffff4ffffffff",
            INIT_38 => X"0000001c000000000000001100000000fffffffbffffffffffffffe9ffffffff",
            INIT_39 => X"ffffffdaffffffffffffffd8ffffffffffffffeeffffffff0000001000000000",
            INIT_3A => X"fffffffbffffffffffffffc0ffffffffffffffbaffffffffffffffb0ffffffff",
            INIT_3B => X"00000024000000000000002e000000000000001a000000000000003400000000",
            INIT_3C => X"fffffffaffffffff0000002d000000000000001d000000000000001e00000000",
            INIT_3D => X"fffffff9fffffffffffffff0ffffffffffffffebffffffffffffffe7ffffffff",
            INIT_3E => X"fffffffaffffffff0000000000000000ffffffefffffffff0000001500000000",
            INIT_3F => X"00000005000000000000000000000000fffffff0fffffffffffffffcffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000001700000000fffffff8fffffffffffffffcffffffff",
            INIT_41 => X"0000000000000000000000060000000000000000000000000000002800000000",
            INIT_42 => X"0000002a000000000000000c000000000000001300000000ffffffeeffffffff",
            INIT_43 => X"00000005000000000000001a0000000000000004000000000000000b00000000",
            INIT_44 => X"fffffffbffffffff0000001100000000fffffff4ffffffff0000002900000000",
            INIT_45 => X"fffffff5ffffffff0000001e00000000fffffff7ffffffff0000000300000000",
            INIT_46 => X"0000004f0000000000000033000000000000001a000000000000000600000000",
            INIT_47 => X"00000054000000000000007a000000000000002f000000000000006d00000000",
            INIT_48 => X"fffffffbffffffff00000013000000000000002a000000000000006400000000",
            INIT_49 => X"0000000d00000000fffffff4ffffffff00000003000000000000003200000000",
            INIT_4A => X"fffffff7fffffffffffffff8ffffffffffffffd5ffffffff0000001000000000",
            INIT_4B => X"0000001e00000000fffffff9ffffffffffffffedffffffff0000002300000000",
            INIT_4C => X"fffffff8ffffffff0000003a00000000ffffffffffffffff0000000300000000",
            INIT_4D => X"0000000d000000000000001b000000000000001300000000fffffff2ffffffff",
            INIT_4E => X"fffffff3ffffffff0000000b00000000fffffffdfffffffffffffff1ffffffff",
            INIT_4F => X"ffffffb1fffffffffffffff6ffffffffffffffbbfffffffffffffff8ffffffff",
            INIT_50 => X"ffffffd2ffffffffffffffeaffffffffffffffb9ffffffffffffffa3ffffffff",
            INIT_51 => X"000000060000000000000015000000000000001800000000ffffffafffffffff",
            INIT_52 => X"00000015000000000000000000000000ffffffe8ffffffffffffffddffffffff",
            INIT_53 => X"00000020000000000000002700000000fffffffffffffffffffffff8ffffffff",
            INIT_54 => X"000000010000000000000021000000000000001200000000fffffffcffffffff",
            INIT_55 => X"ffffffdfffffffffffffffd3fffffffffffffff6fffffffffffffff5ffffffff",
            INIT_56 => X"ffffffeefffffffffffffff5ffffffff0000000600000000fffffff1ffffffff",
            INIT_57 => X"0000003700000000000000150000000000000014000000000000001a00000000",
            INIT_58 => X"fffffffefffffffffffffff9fffffffffffffff9ffffffff0000000000000000",
            INIT_59 => X"fffffff0ffffffff0000000a000000000000000f00000000fffffffaffffffff",
            INIT_5A => X"ffffff99ffffffffffffff8bffffffffffffffb6ffffffff0000000600000000",
            INIT_5B => X"fffffff6ffffffffffffffcfffffffffffffff86ffffffffffffffacffffffff",
            INIT_5C => X"0000004700000000ffffffdcffffffffffffffd6ffffffffffffffcaffffffff",
            INIT_5D => X"0000001400000000000000070000000000000002000000000000004200000000",
            INIT_5E => X"fffffffbffffffffffffffd7ffffffffffffffe8ffffffffffffffe8ffffffff",
            INIT_5F => X"0000000900000000fffffff1ffffffff00000044000000000000001600000000",
            INIT_60 => X"ffffffcfffffffffffffffe0ffffffff0000000100000000ffffffe3ffffffff",
            INIT_61 => X"0000001c00000000000000210000000000000030000000000000003000000000",
            INIT_62 => X"fffffffeffffffff00000011000000000000004d000000000000000600000000",
            INIT_63 => X"0000001e000000000000003e0000000000000019000000000000000f00000000",
            INIT_64 => X"00000007000000000000001f000000000000001f000000000000001f00000000",
            INIT_65 => X"ffffffd7ffffffffffffffdcffffffff00000013000000000000001800000000",
            INIT_66 => X"ffffffe5ffffffffffffffd7fffffffffffffff0ffffffffffffffc2ffffffff",
            INIT_67 => X"fffffffaffffffff0000000300000000ffffffebffffffffffffffd1ffffffff",
            INIT_68 => X"0000001e00000000000000160000000000000010000000000000001900000000",
            INIT_69 => X"0000000900000000000000190000000000000024000000000000000500000000",
            INIT_6A => X"ffffffddfffffffffffffff8ffffffffffffffe4fffffffffffffffaffffffff",
            INIT_6B => X"ffffffd1ffffffffffffffd9ffffffffffffffefffffffffffffffcbffffffff",
            INIT_6C => X"ffffffefffffffffffffffe4ffffffffffffffa2ffffffff0000000000000000",
            INIT_6D => X"ffffffe5ffffffff0000000400000000fffffffbffffffffffffffc1ffffffff",
            INIT_6E => X"ffffffbcffffffffffffffe7ffffffffffffffdfffffffff0000000900000000",
            INIT_6F => X"ffffffddffffffffffffffcdfffffffffffffffbffffffffffffffcbffffffff",
            INIT_70 => X"ffffffc9ffffffffffffffe6ffffffffffffffdfffffffff0000000d00000000",
            INIT_71 => X"ffffffe3ffffffffffffffebffffffff0000001300000000ffffffd0ffffffff",
            INIT_72 => X"ffffffddffffffffffffffd6ffffffff0000001200000000ffffffe1ffffffff",
            INIT_73 => X"fffffff5ffffffff0000001100000000fffffff4ffffffff0000000000000000",
            INIT_74 => X"0000001100000000fffffff9ffffffff0000000f000000000000000100000000",
            INIT_75 => X"ffffffd4ffffffffffffffd3ffffffffffffffcfffffffff0000001800000000",
            INIT_76 => X"ffffffc9ffffffffffffffe1ffffffffffffffd2fffffffffffffff4ffffffff",
            INIT_77 => X"ffffffebfffffffffffffffbffffffff0000000600000000ffffffeeffffffff",
            INIT_78 => X"ffffffebfffffffffffffffefffffffffffffff3ffffffff0000001200000000",
            INIT_79 => X"ffffffc3ffffffffffffffd6ffffffff0000000000000000fffffff3ffffffff",
            INIT_7A => X"0000000a00000000ffffffd6fffffffffffffff6ffffffffffffffe7ffffffff",
            INIT_7B => X"00000024000000000000003900000000fffffff4ffffffff0000000600000000",
            INIT_7C => X"ffffffa6ffffffffffffffa7ffffffffffffffeaffffffffffffffd5ffffffff",
            INIT_7D => X"ffffffbfffffffffffffffc7ffffffffffffffbeffffffffffffffc5ffffffff",
            INIT_7E => X"ffffffdcffffffffffffffbfffffffffffffffdeffffffffffffffb7ffffffff",
            INIT_7F => X"0000001c00000000ffffffe3ffffffffffffffefffffffff0000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE9;


    MEM_IWGHT_LAYER2_INSTANCE10 : if BRAM_NAME = "iwght_layer2_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000e000000000000001e00000000ffffffe6ffffffff0000000000000000",
            INIT_01 => X"0000000700000000ffffffe9ffffffffffffffe8ffffffff0000002700000000",
            INIT_02 => X"0000000800000000ffffffefffffffff0000000000000000ffffffaaffffffff",
            INIT_03 => X"00000027000000000000000f000000000000000600000000fffffffeffffffff",
            INIT_04 => X"0000002f000000000000001700000000fffffff9ffffffff0000002200000000",
            INIT_05 => X"ffffffefffffffff00000020000000000000000f00000000ffffffebffffffff",
            INIT_06 => X"0000001600000000fffffff9ffffffff00000003000000000000001000000000",
            INIT_07 => X"fffffffffffffffffffffffcfffffffffffffff8ffffffff0000001900000000",
            INIT_08 => X"00000001000000000000000c0000000000000008000000000000000a00000000",
            INIT_09 => X"ffffffdaffffffffffffffc2ffffffff00000016000000000000001a00000000",
            INIT_0A => X"ffffffe4fffffffffffffff5ffffffffffffffccffffffffffffffc5ffffffff",
            INIT_0B => X"0000001800000000fffffffdffffffffffffffebffffffff0000000c00000000",
            INIT_0C => X"0000001500000000000000190000000000000011000000000000000a00000000",
            INIT_0D => X"fffffffaffffffff0000000c00000000fffffff6ffffffffffffffefffffffff",
            INIT_0E => X"ffffffb7ffffffffffffffffffffffff0000002b00000000ffffffedffffffff",
            INIT_0F => X"ffffffdeffffffffffffffa4ffffffff0000000500000000fffffff2ffffffff",
            INIT_10 => X"00000025000000000000002a0000000000000010000000000000000600000000",
            INIT_11 => X"fffffff5ffffffff0000000500000000fffffff2ffffffffffffffffffffffff",
            INIT_12 => X"fffffffbffffffffffffffe7ffffffff0000000500000000ffffffe6ffffffff",
            INIT_13 => X"fffffffafffffffffffffff3fffffffffffffff0ffffffff0000000f00000000",
            INIT_14 => X"ffffffebfffffffffffffff8ffffffff0000000900000000fffffff3ffffffff",
            INIT_15 => X"0000000800000000ffffffe5ffffffffffffffe0ffffffffffffffc8ffffffff",
            INIT_16 => X"00000004000000000000000000000000ffffffbefffffffffffffff6ffffffff",
            INIT_17 => X"0000000800000000000000370000000000000013000000000000001c00000000",
            INIT_18 => X"ffffffadffffffffffffffe3fffffffffffffff2ffffffff0000000000000000",
            INIT_19 => X"ffffffd9ffffffff0000000500000000fffffffaffffffff0000001200000000",
            INIT_1A => X"ffffffe1ffffffffffffffdffffffffffffffff2ffffffffffffffd6ffffffff",
            INIT_1B => X"00000032000000000000001900000000ffffffcbffffffff0000000200000000",
            INIT_1C => X"00000011000000000000001f00000000fffffff8ffffffff0000000c00000000",
            INIT_1D => X"000000000000000000000017000000000000001a00000000fffffff8ffffffff",
            INIT_1E => X"000000160000000000000012000000000000000000000000ffffffebffffffff",
            INIT_1F => X"0000000400000000fffffffdffffffff0000002a00000000fffffffdffffffff",
            INIT_20 => X"0000000d000000000000001400000000ffffffeeffffffffffffffeeffffffff",
            INIT_21 => X"ffffffe9ffffffff00000000000000000000000a000000000000000300000000",
            INIT_22 => X"0000003e000000000000000f0000000000000016000000000000001700000000",
            INIT_23 => X"fffffff5ffffffff0000000a000000000000001c000000000000000500000000",
            INIT_24 => X"0000000000000000ffffffe9ffffffff00000003000000000000000000000000",
            INIT_25 => X"0000000e000000000000001b00000000fffffffcffffffff0000000100000000",
            INIT_26 => X"ffffffceffffffff0000001c000000000000000a00000000fffffff4ffffffff",
            INIT_27 => X"000000060000000000000032000000000000000f00000000ffffffe3ffffffff",
            INIT_28 => X"00000000000000000000000b000000000000002f00000000ffffffe7ffffffff",
            INIT_29 => X"0000000b000000000000000200000000fffffffcffffffffffffffeeffffffff",
            INIT_2A => X"fffffffcffffffff00000022000000000000000800000000fffffffbffffffff",
            INIT_2B => X"00000003000000000000001800000000fffffff7ffffffff0000000700000000",
            INIT_2C => X"ffffffefffffffff0000000900000000ffffffeeffffffffffffffedffffffff",
            INIT_2D => X"0000001b00000000000000000000000000000022000000000000000400000000",
            INIT_2E => X"0000001800000000000000010000000000000003000000000000000f00000000",
            INIT_2F => X"ffffffeaffffffff0000000f00000000ffffffffffffffffffffffeeffffffff",
            INIT_30 => X"0000001700000000ffffffe5ffffffff00000025000000000000000000000000",
            INIT_31 => X"0000005000000000000000180000000000000048000000000000003100000000",
            INIT_32 => X"0000001b00000000ffffffc7ffffffffffffffddffffffff0000001e00000000",
            INIT_33 => X"00000001000000000000002800000000ffffffdcffffffff0000003400000000",
            INIT_34 => X"fffffff2ffffffff00000022000000000000001100000000fffffff7ffffffff",
            INIT_35 => X"ffffffa9ffffffffffffffd8fffffffffffffffeffffffffffffffedffffffff",
            INIT_36 => X"00000000000000000000001b00000000ffffffd0ffffffffffffffe2ffffffff",
            INIT_37 => X"ffffffe5ffffffff0000000d00000000fffffff9ffffffff0000001100000000",
            INIT_38 => X"0000000d00000000fffffff2ffffffff0000000900000000ffffffe6ffffffff",
            INIT_39 => X"ffffffcaffffffffffffffd3ffffffff0000002c00000000fffffff0ffffffff",
            INIT_3A => X"ffffffebffffffffffffffd4ffffffffffffffc4ffffffffffffffc8ffffffff",
            INIT_3B => X"ffffffe7ffffffff000000240000000000000026000000000000002300000000",
            INIT_3C => X"fffffff9fffffffffffffff9ffffffff0000000800000000ffffffe1ffffffff",
            INIT_3D => X"00000020000000000000002b0000000000000014000000000000001300000000",
            INIT_3E => X"000000110000000000000019000000000000001b00000000fffffff7ffffffff",
            INIT_3F => X"ffffffddfffffffffffffff2ffffffff0000004300000000fffffff7ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdfffffffffffffffe5ffffffffffffffecffffffffffffffdeffffffff",
            INIT_41 => X"0000004a000000000000003e000000000000003d000000000000002c00000000",
            INIT_42 => X"fffffff8ffffffffffffffe4ffffffff00000021000000000000004600000000",
            INIT_43 => X"ffffffc6ffffffffffffffc2ffffffffffffffbeffffffff0000000000000000",
            INIT_44 => X"ffffffecffffffffffffffb4ffffffffffffffd1ffffffffffffffc7ffffffff",
            INIT_45 => X"ffffffefffffffffffffffd1ffffffff0000000c000000000000001c00000000",
            INIT_46 => X"0000000f0000000000000025000000000000002100000000ffffffdfffffffff",
            INIT_47 => X"ffffffb6fffffffffffffff6fffffffffffffffeffffffffffffffe2ffffffff",
            INIT_48 => X"ffffffdeffffffffffffffe1ffffffff0000000300000000fffffffaffffffff",
            INIT_49 => X"fffffff8ffffffff00000031000000000000000200000000ffffffd3ffffffff",
            INIT_4A => X"0000000d00000000ffffffcdffffffffffffffe9ffffffffffffffbaffffffff",
            INIT_4B => X"fffffffaffffffffffffffe9fffffffffffffff5ffffffffffffffffffffffff",
            INIT_4C => X"0000001e00000000ffffffe5fffffffffffffff0ffffffffffffffeaffffffff",
            INIT_4D => X"00000013000000000000000e000000000000000a000000000000000000000000",
            INIT_4E => X"ffffffedfffffffffffffffbffffffff0000002e000000000000001100000000",
            INIT_4F => X"00000016000000000000001e0000000000000021000000000000000400000000",
            INIT_50 => X"0000000e000000000000001300000000fffffff1fffffffffffffff5ffffffff",
            INIT_51 => X"0000002d0000000000000052000000000000000300000000ffffffdcffffffff",
            INIT_52 => X"ffffffceffffffff000000000000000000000000000000000000001a00000000",
            INIT_53 => X"ffffffccfffffffffffffff6fffffffffffffff1fffffffffffffff6ffffffff",
            INIT_54 => X"ffffffe2ffffffffffffffe9ffffffffffffffd0ffffffffffffffacffffffff",
            INIT_55 => X"00000012000000000000001200000000ffffffeafffffffffffffff8ffffffff",
            INIT_56 => X"fffffff4ffffffffffffffafffffffffffffffa5ffffffffffffffd8ffffffff",
            INIT_57 => X"ffffffd4fffffffffffffff5ffffffffffffffe1ffffffffffffffefffffffff",
            INIT_58 => X"fffffff7ffffffffffffffd7ffffffffffffffb2ffffffffffffffbcffffffff",
            INIT_59 => X"0000002a000000000000000c0000000000000034000000000000000e00000000",
            INIT_5A => X"0000000e00000000fffffffefffffffffffffffdfffffffffffffff7ffffffff",
            INIT_5B => X"ffffffdbfffffffffffffff5ffffffffffffffd0fffffffffffffffcffffffff",
            INIT_5C => X"0000000f000000000000000f00000000ffffffebffffffffffffffb2ffffffff",
            INIT_5D => X"000000120000000000000000000000000000000f000000000000000000000000",
            INIT_5E => X"0000003700000000fffffff2ffffffffffffffe3ffffffff0000001400000000",
            INIT_5F => X"0000001d00000000ffffffcafffffffffffffff1fffffffffffffff0ffffffff",
            INIT_60 => X"00000000000000000000000f00000000ffffffcdfffffffffffffffaffffffff",
            INIT_61 => X"fffffff2ffffffff00000007000000000000001800000000ffffffccffffffff",
            INIT_62 => X"00000001000000000000003b000000000000001500000000fffffffeffffffff",
            INIT_63 => X"ffffffe8ffffffffffffffd6ffffffff0000003c00000000fffffff2ffffffff",
            INIT_64 => X"000000220000000000000023000000000000001b00000000fffffffcffffffff",
            INIT_65 => X"00000010000000000000000b000000000000001e000000000000001b00000000",
            INIT_66 => X"0000000000000000ffffffe3ffffffff0000001c000000000000002900000000",
            INIT_67 => X"ffffffe8ffffffffffffffeeffffffffffffffccffffffff0000000b00000000",
            INIT_68 => X"0000000e000000000000001a0000000000000006000000000000000c00000000",
            INIT_69 => X"00000002000000000000001500000000fffffffcfffffffffffffff4ffffffff",
            INIT_6A => X"0000002a000000000000004b000000000000003300000000fffffff9ffffffff",
            INIT_6B => X"00000042000000000000003e0000000000000040000000000000004300000000",
            INIT_6C => X"ffffffbafffffffffffffff0ffffffff0000003a000000000000003800000000",
            INIT_6D => X"ffffffbcffffffffffffff8affffffffffffffbcfffffffffffffff5ffffffff",
            INIT_6E => X"ffffffdeffffffffffffffdaffffffffffffff94ffffffffffffffbeffffffff",
            INIT_6F => X"ffffffc0ffffffffffffffdeffffffffffffffe3ffffffffffffffdfffffffff",
            INIT_70 => X"ffffffe5ffffffffffffffe4ffffffffffffffa2ffffffffffffffefffffffff",
            INIT_71 => X"ffffffc4ffffffffffffffe6ffffffffffffffe2fffffffffffffff7ffffffff",
            INIT_72 => X"ffffffbeffffffffffffff86ffffffff0000000c00000000ffffffbbffffffff",
            INIT_73 => X"ffffffd9ffffffffffffffe9fffffffffffffffaffffffffffffffe1ffffffff",
            INIT_74 => X"0000003700000000ffffffffffffffff00000000000000000000000c00000000",
            INIT_75 => X"0000004200000000fffffffeffffffff00000042000000000000002f00000000",
            INIT_76 => X"0000000d00000000ffffffebfffffffffffffff7ffffffff0000002700000000",
            INIT_77 => X"0000000e00000000ffffffefffffffffffffffe0ffffffffffffffdcffffffff",
            INIT_78 => X"00000021000000000000001000000000fffffffbffffffff0000000100000000",
            INIT_79 => X"0000000800000000000000150000000000000027000000000000000500000000",
            INIT_7A => X"0000001e00000000000000220000000000000015000000000000000a00000000",
            INIT_7B => X"00000010000000000000000c000000000000000a00000000fffffff1ffffffff",
            INIT_7C => X"0000001b000000000000000b0000000000000014000000000000003800000000",
            INIT_7D => X"ffffffcbffffffff00000002000000000000000500000000ffffffdbffffffff",
            INIT_7E => X"000000100000000000000021000000000000000300000000ffffffdbffffffff",
            INIT_7F => X"0000002900000000fffffff5ffffffff00000022000000000000000d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE10;


    MEM_IWGHT_LAYER2_INSTANCE11 : if BRAM_NAME = "iwght_layer2_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff8ffffffff0000001700000000fffffffdffffffffffffffeeffffffff",
            INIT_01 => X"fffffff7fffffffffffffff0ffffffffffffffd8fffffffffffffff0ffffffff",
            INIT_02 => X"0000000a000000000000001e00000000ffffffe4ffffffffffffffe7ffffffff",
            INIT_03 => X"ffffffefffffffffffffffebffffffffffffffe9ffffffff0000000b00000000",
            INIT_04 => X"0000000c00000000fffffffffffffffffffffff1fffffffffffffff3ffffffff",
            INIT_05 => X"000000160000000000000021000000000000001300000000fffffff2ffffffff",
            INIT_06 => X"ffffffedffffffff000000320000000000000031000000000000001400000000",
            INIT_07 => X"ffffffe9ffffffff0000000c0000000000000009000000000000000700000000",
            INIT_08 => X"fffffffbffffffff0000000000000000ffffffedfffffffffffffffeffffffff",
            INIT_09 => X"ffffffe4ffffffff000000060000000000000010000000000000001e00000000",
            INIT_0A => X"0000000000000000ffffffdaffffffffffffffe9fffffffffffffffcffffffff",
            INIT_0B => X"00000009000000000000001000000000fffffffaffffffff0000000300000000",
            INIT_0C => X"fffffff9ffffffff0000005e000000000000005d000000000000003300000000",
            INIT_0D => X"000000130000000000000020000000000000003a000000000000004800000000",
            INIT_0E => X"fffffffdffffffff0000001e000000000000000e000000000000002500000000",
            INIT_0F => X"fffffff7ffffffff000000000000000000000005000000000000000a00000000",
            INIT_10 => X"0000000000000000ffffffeaffffffff0000000d000000000000000e00000000",
            INIT_11 => X"ffffffe6ffffffff0000000d00000000ffffffe3ffffffffffffffe8ffffffff",
            INIT_12 => X"0000001d00000000ffffffe4fffffffffffffff8ffffffffffffffe8ffffffff",
            INIT_13 => X"fffffff6ffffffff00000001000000000000001f000000000000000f00000000",
            INIT_14 => X"0000001900000000000000140000000000000014000000000000000800000000",
            INIT_15 => X"0000000f00000000ffffffeafffffffffffffff5ffffffffffffffd2ffffffff",
            INIT_16 => X"00000002000000000000001a00000000ffffffe7ffffffff0000001800000000",
            INIT_17 => X"0000000300000000000000190000000000000011000000000000000700000000",
            INIT_18 => X"0000000b00000000ffffffe6ffffffff0000000f00000000fffffffcffffffff",
            INIT_19 => X"00000012000000000000001c0000000000000011000000000000000700000000",
            INIT_1A => X"0000001c00000000000000110000000000000003000000000000002900000000",
            INIT_1B => X"00000003000000000000000300000000fffffff6fffffffffffffff4ffffffff",
            INIT_1C => X"0000000d00000000fffffff9ffffffff0000000400000000fffffff1ffffffff",
            INIT_1D => X"fffffff3ffffffff0000000400000000ffffffd3ffffffff0000000600000000",
            INIT_1E => X"ffffffb7fffffffffffffff7ffffffffffffffdeffffffffffffffbbffffffff",
            INIT_1F => X"ffffff70ffffffffffffff97ffffffffffffffc3ffffffffffffff94ffffffff",
            INIT_20 => X"000000240000000000000021000000000000000a00000000ffffffc0ffffffff",
            INIT_21 => X"000000040000000000000023000000000000000f000000000000001000000000",
            INIT_22 => X"0000001300000000000000030000000000000019000000000000001100000000",
            INIT_23 => X"00000009000000000000002d00000000ffffffd8ffffffff0000002100000000",
            INIT_24 => X"000000320000000000000006000000000000000a00000000ffffffe6ffffffff",
            INIT_25 => X"fffffffbffffffff0000000a0000000000000009000000000000001800000000",
            INIT_26 => X"ffffffecffffffff00000010000000000000002500000000ffffffedffffffff",
            INIT_27 => X"ffffffd2fffffffffffffff4ffffffffffffffd4fffffffffffffff6ffffffff",
            INIT_28 => X"ffffffe7ffffffffffffffc8ffffffff0000000900000000ffffffd5ffffffff",
            INIT_29 => X"0000000100000000ffffffe9ffffffffffffffefffffffff0000000800000000",
            INIT_2A => X"0000000400000000ffffffeaffffffff00000008000000000000000900000000",
            INIT_2B => X"ffffffe8fffffffffffffff1ffffffffffffffdfffffffffffffffeaffffffff",
            INIT_2C => X"000000030000000000000012000000000000001800000000ffffffe6ffffffff",
            INIT_2D => X"fffffff0ffffffff000000000000000000000015000000000000000d00000000",
            INIT_2E => X"0000000e000000000000000300000000fffffffcffffffff0000000f00000000",
            INIT_2F => X"00000009000000000000000000000000fffffffbffffffff0000000300000000",
            INIT_30 => X"ffffffeaffffffff0000000000000000ffffffeaffffffffffffffebffffffff",
            INIT_31 => X"0000000a00000000000000030000000000000003000000000000000b00000000",
            INIT_32 => X"fffffffcffffffff000000040000000000000011000000000000000a00000000",
            INIT_33 => X"ffffffd4ffffffffffffffe2ffffffffffffffc7ffffffffffffffefffffffff",
            INIT_34 => X"ffffffc1ffffffffffffffc2ffffffffffffffdeffffffffffffffd8ffffffff",
            INIT_35 => X"ffffffedffffffffffffff9affffffffffffffabffffffffffffffccffffffff",
            INIT_36 => X"00000009000000000000001500000000fffffffbffffffff0000000b00000000",
            INIT_37 => X"00000003000000000000002900000000ffffffd6fffffffffffffff7ffffffff",
            INIT_38 => X"fffffffeffffffff00000035000000000000003600000000ffffffe5ffffffff",
            INIT_39 => X"ffffffb2ffffffffffffffb3ffffffffffffffc1ffffffffffffff96ffffffff",
            INIT_3A => X"00000024000000000000000500000000ffffffe9ffffffffffffffd6ffffffff",
            INIT_3B => X"000000330000000000000042000000000000001a000000000000000500000000",
            INIT_3C => X"ffffffcfffffffff000000270000000000000016000000000000000000000000",
            INIT_3D => X"ffffffe9ffffffffffffffd8ffffffffffffffd6fffffffffffffff1ffffffff",
            INIT_3E => X"ffffffe5ffffffffffffffdeffffffffffffffa3ffffffffffffffbfffffffff",
            INIT_3F => X"0000001b000000000000002c00000000ffffffebffffffff0000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000fffffff7ffffffff0000000f000000000000000e00000000",
            INIT_41 => X"00000034000000000000000a000000000000001c000000000000001e00000000",
            INIT_42 => X"ffffffdafffffffffffffff9fffffffffffffffdfffffffffffffffaffffffff",
            INIT_43 => X"ffffffe7ffffffffffffffcbfffffffffffffff6ffffffffffffffcaffffffff",
            INIT_44 => X"fffffffcffffffff00000014000000000000001000000000ffffffeeffffffff",
            INIT_45 => X"fffffff8ffffffff0000000700000000ffffffedffffffff0000000100000000",
            INIT_46 => X"0000000700000000fffffff2ffffffffffffffeeffffffff0000000a00000000",
            INIT_47 => X"ffffffedfffffffffffffff3ffffffffffffffd8fffffffffffffff5ffffffff",
            INIT_48 => X"000000140000000000000024000000000000002900000000fffffff3ffffffff",
            INIT_49 => X"0000000c00000000000000080000000000000007000000000000001d00000000",
            INIT_4A => X"ffffffc6ffffffff0000001e00000000fffffffafffffffffffffff2ffffffff",
            INIT_4B => X"000000020000000000000018000000000000000300000000fffffffcffffffff",
            INIT_4C => X"000000010000000000000000000000000000000500000000fffffff9ffffffff",
            INIT_4D => X"ffffffd3ffffffffffffffd6ffffffffffffffdbffffffffffffffdaffffffff",
            INIT_4E => X"0000004d00000000fffffff2fffffffffffffff9ffffffff0000000300000000",
            INIT_4F => X"00000036000000000000000e000000000000003b000000000000003000000000",
            INIT_50 => X"ffffffecffffffff0000000e00000000ffffffe7ffffffff0000001800000000",
            INIT_51 => X"ffffffe9ffffffffffffffe3ffffffffffffffedffffffffffffffc4ffffffff",
            INIT_52 => X"fffffffdfffffffffffffffdfffffffffffffff1ffffffff0000000100000000",
            INIT_53 => X"0000000000000000ffffffedffffffffffffffd8ffffffffffffffebffffffff",
            INIT_54 => X"0000000b00000000ffffffd5ffffffff00000007000000000000000400000000",
            INIT_55 => X"0000003600000000000000170000000000000034000000000000001000000000",
            INIT_56 => X"0000000600000000fffffff5fffffffffffffff4ffffffff0000001600000000",
            INIT_57 => X"0000000800000000fffffffffffffffffffffff1ffffffff0000001b00000000",
            INIT_58 => X"fffffff9ffffffffffffffd6ffffffff0000000b000000000000001400000000",
            INIT_59 => X"ffffffffffffffff0000000500000000fffffff0ffffffffffffffd2ffffffff",
            INIT_5A => X"fffffffbffffffffffffffe4ffffffff0000000a000000000000002a00000000",
            INIT_5B => X"0000001500000000ffffffedffffffff0000001b000000000000000c00000000",
            INIT_5C => X"00000013000000000000000500000000ffffffeffffffffffffffff6ffffffff",
            INIT_5D => X"0000001f00000000fffffff4ffffffff0000000d000000000000000c00000000",
            INIT_5E => X"0000000400000000fffffff7fffffffffffffff6ffffffff0000001c00000000",
            INIT_5F => X"ffffffffffffffff00000010000000000000003100000000ffffffebffffffff",
            INIT_60 => X"ffffffd2ffffffffffffffe7ffffffff0000000e00000000fffffffaffffffff",
            INIT_61 => X"0000001a00000000fffffffdffffffff0000001400000000ffffffeeffffffff",
            INIT_62 => X"0000002800000000000000150000000000000002000000000000000c00000000",
            INIT_63 => X"0000000300000000fffffff7ffffffff0000000600000000ffffffebffffffff",
            INIT_64 => X"fffffff6ffffffff000000060000000000000012000000000000000f00000000",
            INIT_65 => X"00000011000000000000001a000000000000000d00000000ffffffecffffffff",
            INIT_66 => X"ffffffcfffffffff0000002d000000000000001d00000000ffffffc4ffffffff",
            INIT_67 => X"0000000e00000000ffffffc6ffffffff00000050000000000000003400000000",
            INIT_68 => X"ffffffcbffffffffffffffcdffffffffffffffc9ffffffff0000008d00000000",
            INIT_69 => X"0000002a00000000ffffffe6ffffffff0000000000000000ffffffe2ffffffff",
            INIT_6A => X"fffffff3ffffffff00000001000000000000002e000000000000003a00000000",
            INIT_6B => X"fffffff3ffffffffffffffeffffffffffffffff4ffffffff0000000400000000",
            INIT_6C => X"ffffffe4ffffffff000000010000000000000020000000000000003100000000",
            INIT_6D => X"fffffff1ffffffffffffffe5ffffffff0000000a000000000000000800000000",
            INIT_6E => X"00000016000000000000001500000000ffffffbffffffffffffffff9ffffffff",
            INIT_6F => X"0000002a00000000ffffffd9fffffffffffffff4fffffffffffffff0ffffffff",
            INIT_70 => X"00000036000000000000003700000000ffffffe7ffffffff0000000900000000",
            INIT_71 => X"00000016000000000000002e000000000000001100000000ffffffebffffffff",
            INIT_72 => X"ffffffd8ffffffff0000000d000000000000000600000000ffffffeaffffffff",
            INIT_73 => X"0000000e0000000000000022000000000000001d00000000ffffffe9ffffffff",
            INIT_74 => X"fffffffdffffffff0000001e000000000000002500000000fffffff3ffffffff",
            INIT_75 => X"0000002500000000fffffff8ffffffff00000010000000000000001b00000000",
            INIT_76 => X"0000001600000000000000360000000000000028000000000000001700000000",
            INIT_77 => X"fffffffaffffffff00000022000000000000001c00000000ffffffd9ffffffff",
            INIT_78 => X"00000006000000000000000c000000000000000800000000fffffffeffffffff",
            INIT_79 => X"000000170000000000000004000000000000001a000000000000000a00000000",
            INIT_7A => X"fffffff3ffffffff0000000400000000fffffff7fffffffffffffff5ffffffff",
            INIT_7B => X"0000000500000000000000180000000000000006000000000000000300000000",
            INIT_7C => X"fffffffaffffffff0000000f00000000ffffffedffffffff0000003000000000",
            INIT_7D => X"ffffffe9ffffffffffffffeafffffffffffffff0fffffffffffffff3ffffffff",
            INIT_7E => X"fffffff7fffffffffffffffbffffffffffffffd9ffffffff0000001500000000",
            INIT_7F => X"ffffffeaffffffff0000000600000000ffffffd1ffffffffffffffe2ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE11;


    MEM_IWGHT_LAYER2_INSTANCE12 : if BRAM_NAME = "iwght_layer2_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004d000000000000001a0000000000000002000000000000002c00000000",
            INIT_01 => X"ffffffdefffffffffffffffaffffffffffffffbfffffffffffffffe2ffffffff",
            INIT_02 => X"ffffffa3fffffffffffffffeffffffffffffffffffffffffffffffd2ffffffff",
            INIT_03 => X"0000000f00000000ffffffecfffffffffffffff4ffffffffffffffaaffffffff",
            INIT_04 => X"ffffffecfffffffffffffffbfffffffffffffff3ffffffff0000000000000000",
            INIT_05 => X"00000025000000000000002100000000fffffff1ffffffffffffffe2ffffffff",
            INIT_06 => X"ffffffd6ffffffffffffffa8ffffffffffffffa2fffffffffffffff1ffffffff",
            INIT_07 => X"ffffffecffffffff0000000000000000ffffffc5ffffffffffffffc5ffffffff",
            INIT_08 => X"fffffff0ffffffffffffffcaffffffff00000007000000000000001b00000000",
            INIT_09 => X"0000002e000000000000000e00000000ffffffe0ffffffff0000000a00000000",
            INIT_0A => X"0000000400000000000000110000000000000015000000000000002200000000",
            INIT_0B => X"fffffff3fffffffffffffffbffffffffffffffeaffffffff0000000600000000",
            INIT_0C => X"ffffffc9ffffffffffffffe5ffffffff0000000a00000000ffffffe9ffffffff",
            INIT_0D => X"0000001100000000ffffffd5ffffffff00000006000000000000001600000000",
            INIT_0E => X"00000016000000000000000a00000000ffffffacfffffffffffffff2ffffffff",
            INIT_0F => X"ffffffe4ffffffff00000022000000000000001d000000000000001f00000000",
            INIT_10 => X"0000000000000000ffffffd5ffffffffffffffecffffffffffffffeaffffffff",
            INIT_11 => X"00000008000000000000000700000000fffffff9fffffffffffffff6ffffffff",
            INIT_12 => X"00000009000000000000000a000000000000002200000000ffffffefffffffff",
            INIT_13 => X"ffffffd8ffffffffffffffe4ffffffffffffffe9ffffffffffffffe1ffffffff",
            INIT_14 => X"0000000200000000ffffffe1ffffffff0000000100000000fffffff9ffffffff",
            INIT_15 => X"fffffff5ffffffff000000230000000000000018000000000000000600000000",
            INIT_16 => X"00000016000000000000000b000000000000001d00000000fffffffdffffffff",
            INIT_17 => X"00000005000000000000000b000000000000000e000000000000000600000000",
            INIT_18 => X"ffffffeeffffffff000000150000000000000006000000000000000100000000",
            INIT_19 => X"fffffff8ffffffffffffffd1ffffffffffffffabffffffffffffffc6ffffffff",
            INIT_1A => X"fffffffcffffffff0000002800000000ffffffedfffffffffffffffdffffffff",
            INIT_1B => X"fffffff4ffffffff0000000300000000fffffff5fffffffffffffff2ffffffff",
            INIT_1C => X"0000004700000000000000210000000000000026000000000000003600000000",
            INIT_1D => X"0000000d000000000000000c0000000000000002000000000000003b00000000",
            INIT_1E => X"00000000000000000000000f00000000fffffff7ffffffff0000000200000000",
            INIT_1F => X"fffffff9fffffffffffffff8ffffffff00000021000000000000000500000000",
            INIT_20 => X"000000270000000000000023000000000000000600000000ffffffe2ffffffff",
            INIT_21 => X"fffffff5ffffffff0000002600000000ffffffdffffffffffffffffbffffffff",
            INIT_22 => X"0000000e00000000ffffffc7fffffffffffffff3ffffffffffffffb5ffffffff",
            INIT_23 => X"ffffffedfffffffffffffff1ffffffff00000014000000000000000d00000000",
            INIT_24 => X"ffffffffffffffffffffffd1ffffffffffffffbbffffffff0000000700000000",
            INIT_25 => X"ffffffe1ffffffff0000001c000000000000002f000000000000003300000000",
            INIT_26 => X"ffffffdeffffffffffffffc2ffffffff0000001500000000ffffffcfffffffff",
            INIT_27 => X"00000021000000000000001d0000000000000033000000000000000200000000",
            INIT_28 => X"ffffffe0ffffffff0000000d00000000fffffff8ffffffff0000000e00000000",
            INIT_29 => X"ffffffd9ffffffffffffffecffffffff0000002300000000ffffffcbffffffff",
            INIT_2A => X"ffffffd9ffffffff00000007000000000000000600000000ffffffffffffffff",
            INIT_2B => X"fffffffdffffffffffffffffffffffff00000009000000000000001000000000",
            INIT_2C => X"00000010000000000000000c0000000000000020000000000000002400000000",
            INIT_2D => X"ffffffdaffffffffffffffc3ffffffffffffff9dffffffff0000000f00000000",
            INIT_2E => X"0000002800000000fffffff7ffffffffffffffe8ffffffff0000003600000000",
            INIT_2F => X"ffffffc2ffffffff00000024000000000000000600000000ffffffb1ffffffff",
            INIT_30 => X"000000050000000000000003000000000000000400000000ffffffd8ffffffff",
            INIT_31 => X"ffffffeeffffffff0000000f00000000fffffff4ffffffff0000000900000000",
            INIT_32 => X"0000002600000000000000220000000000000019000000000000000100000000",
            INIT_33 => X"fffffff2ffffffff0000002a000000000000000f00000000fffffff1ffffffff",
            INIT_34 => X"ffffffe7ffffffffffffffccffffffff00000024000000000000000b00000000",
            INIT_35 => X"fffffff6fffffffffffffffbffffffffffffffd0ffffffffffffffe4ffffffff",
            INIT_36 => X"fffffff9ffffffffffffffd4ffffffffffffffeaffffffffffffffedffffffff",
            INIT_37 => X"ffffffe1ffffffffffffffe9ffffffffffffffd8ffffffff0000000600000000",
            INIT_38 => X"000000030000000000000007000000000000001200000000ffffffefffffffff",
            INIT_39 => X"fffffff2fffffffffffffffbffffffffffffffeeffffffff0000003400000000",
            INIT_3A => X"0000000c00000000fffffff8ffffffffffffffecffffffffffffffe9ffffffff",
            INIT_3B => X"0000000b000000000000001d00000000ffffffe8ffffffffffffffdeffffffff",
            INIT_3C => X"fffffffcffffffffffffffffffffffffffffffd9ffffffff0000000200000000",
            INIT_3D => X"0000000a000000000000002700000000ffffffd4ffffffffffffffadffffffff",
            INIT_3E => X"0000002c000000000000002200000000ffffffe0ffffffff0000001300000000",
            INIT_3F => X"fffffffbffffffff0000001d000000000000002900000000fffffff3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001300000000000000040000000000000018000000000000000100000000",
            INIT_41 => X"0000000a0000000000000016000000000000000d00000000fffffff6ffffffff",
            INIT_42 => X"0000001b00000000fffffffaffffffff00000000000000000000000100000000",
            INIT_43 => X"0000001000000000000000350000000000000028000000000000001300000000",
            INIT_44 => X"00000021000000000000003b00000000ffffffefffffffff0000003100000000",
            INIT_45 => X"00000012000000000000002d000000000000001f00000000fffffff4ffffffff",
            INIT_46 => X"0000001300000000fffffff9ffffffff0000000100000000ffffffd9ffffffff",
            INIT_47 => X"ffffffe3ffffffffffffffc9ffffffffffffffeffffffffffffffff8ffffffff",
            INIT_48 => X"fffffff1ffffffffffffffd6ffffffff0000000400000000ffffffedffffffff",
            INIT_49 => X"0000000000000000000000130000000000000006000000000000002800000000",
            INIT_4A => X"0000000d00000000000000070000000000000004000000000000002300000000",
            INIT_4B => X"fffffff8ffffffffffffffd4ffffffffffffffe6ffffffffffffffffffffffff",
            INIT_4C => X"fffffff3ffffffffffffffd9ffffffffffffffbeffffffffffffffe2ffffffff",
            INIT_4D => X"fffffff6ffffffffffffffe4ffffffffffffffd5ffffffffffffffb9ffffffff",
            INIT_4E => X"0000000c000000000000001f00000000fffffff8ffffffff0000000900000000",
            INIT_4F => X"fffffffdffffffff00000009000000000000001100000000ffffffe2ffffffff",
            INIT_50 => X"000000200000000000000004000000000000000000000000fffffff6ffffffff",
            INIT_51 => X"00000029000000000000001f00000000ffffffe4ffffffff0000000e00000000",
            INIT_52 => X"fffffff9fffffffffffffff6fffffffffffffff6ffffffff0000001100000000",
            INIT_53 => X"fffffff3ffffffffffffffe0ffffffff0000000a00000000ffffffedffffffff",
            INIT_54 => X"fffffffffffffffffffffffcfffffffffffffffeffffffff0000000e00000000",
            INIT_55 => X"fffffffeffffffffffffffebffffffff00000006000000000000002d00000000",
            INIT_56 => X"00000020000000000000002700000000ffffffd7fffffffffffffff6ffffffff",
            INIT_57 => X"0000001000000000000000200000000000000019000000000000001a00000000",
            INIT_58 => X"00000005000000000000001e00000000fffffff7fffffffffffffffaffffffff",
            INIT_59 => X"fffffffeffffffffffffffc4ffffffff00000018000000000000000300000000",
            INIT_5A => X"ffffffe0ffffffffffffffd4fffffffffffffff7ffffffff0000000000000000",
            INIT_5B => X"ffffffe4ffffffff0000000e000000000000001c000000000000000600000000",
            INIT_5C => X"fffffff6ffffffff0000000600000000fffffff6fffffffffffffff8ffffffff",
            INIT_5D => X"ffffffe7ffffffffffffffd9ffffffffffffffedffffffffffffffd8ffffffff",
            INIT_5E => X"fffffffdffffffff0000000c000000000000001d00000000ffffffe8ffffffff",
            INIT_5F => X"ffffffd2fffffffffffffff0ffffffffffffffe7ffffffff0000000400000000",
            INIT_60 => X"ffffffe9ffffffffffffffbdffffffffffffffe8fffffffffffffff0ffffffff",
            INIT_61 => X"0000001100000000fffffff4ffffffffffffffcefffffffffffffff2ffffffff",
            INIT_62 => X"ffffffddffffffff00000025000000000000000a000000000000000800000000",
            INIT_63 => X"ffffffd8fffffffffffffffdffffffff0000003200000000fffffff0ffffffff",
            INIT_64 => X"ffffffcbffffffff00000010000000000000003000000000fffffff3ffffffff",
            INIT_65 => X"0000001800000000ffffffdaffffffffffffffceffffffff0000001700000000",
            INIT_66 => X"fffffff8ffffffff0000002c000000000000001d000000000000000100000000",
            INIT_67 => X"ffffffd8ffffffff0000002f000000000000001200000000fffffffeffffffff",
            INIT_68 => X"ffffffe6ffffffff0000001200000000ffffffe9ffffffff0000001700000000",
            INIT_69 => X"fffffff9ffffffff0000002b0000000000000036000000000000001e00000000",
            INIT_6A => X"0000001200000000ffffffe1ffffffffffffffd9ffffffff0000003900000000",
            INIT_6B => X"ffffffd1fffffffffffffffdffffffff0000000b000000000000001000000000",
            INIT_6C => X"fffffffaffffffffffffffe2fffffffffffffffcffffffff0000000000000000",
            INIT_6D => X"00000012000000000000000e0000000000000010000000000000000800000000",
            INIT_6E => X"ffffffdeffffffffffffffebfffffffffffffff6ffffffffffffffe7ffffffff",
            INIT_6F => X"0000000a0000000000000011000000000000000b00000000ffffffe6ffffffff",
            INIT_70 => X"00000005000000000000000d00000000ffffffd4fffffffffffffff4ffffffff",
            INIT_71 => X"fffffff1ffffffffffffffdefffffffffffffff4ffffffffffffffe9ffffffff",
            INIT_72 => X"0000000d00000000fffffff8fffffffffffffffaffffffff0000001500000000",
            INIT_73 => X"0000002000000000fffffff4fffffffffffffff3ffffffff0000000800000000",
            INIT_74 => X"fffffff0fffffffffffffffeffffffff0000000c000000000000000000000000",
            INIT_75 => X"0000003300000000fffffffbfffffffffffffff1ffffffff0000000d00000000",
            INIT_76 => X"0000000900000000fffffff7ffffffffffffffd6ffffffff0000001100000000",
            INIT_77 => X"00000001000000000000001a00000000fffffff8ffffffff0000000400000000",
            INIT_78 => X"0000000c00000000000000220000000000000010000000000000000300000000",
            INIT_79 => X"ffffffd7ffffffff00000029000000000000003c000000000000001100000000",
            INIT_7A => X"0000000200000000fffffffaffffffff0000001d000000000000002900000000",
            INIT_7B => X"000000000000000000000008000000000000000f000000000000000000000000",
            INIT_7C => X"0000000300000000ffffffd6ffffffff00000005000000000000004500000000",
            INIT_7D => X"0000000600000000ffffffc8ffffffff0000001d00000000fffffff6ffffffff",
            INIT_7E => X"ffffffd1fffffffffffffffcfffffffffffffff1ffffffffffffffe7ffffffff",
            INIT_7F => X"ffffffd1ffffffff0000000100000000ffffffecfffffffffffffff2ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE12;


    MEM_IWGHT_LAYER2_INSTANCE13 : if BRAM_NAME = "iwght_layer2_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffa9ffffffffffffffe7ffffffffffffffdcffffffffffffffbeffffffff",
            INIT_01 => X"0000000000000000ffffffe5fffffffffffffff8ffffffffffffffd5ffffffff",
            INIT_02 => X"0000000300000000ffffffc1ffffffffffffffcdffffffffffffffe1ffffffff",
            INIT_03 => X"00000000000000000000000400000000ffffffd8ffffffff0000002b00000000",
            INIT_04 => X"0000000100000000fffffffdfffffffffffffff7fffffffffffffffaffffffff",
            INIT_05 => X"000000050000000000000009000000000000000200000000ffffffeeffffffff",
            INIT_06 => X"fffffffbffffffff000000200000000000000005000000000000000e00000000",
            INIT_07 => X"ffffffe0fffffffffffffff1ffffffff0000001c000000000000001900000000",
            INIT_08 => X"0000000a000000000000001000000000fffffff6fffffffffffffff6ffffffff",
            INIT_09 => X"fffffff0ffffffff0000000a00000000fffffff2fffffffffffffffeffffffff",
            INIT_0A => X"ffffffdbffffffffffffffc9ffffffffffffffdefffffffffffffff5ffffffff",
            INIT_0B => X"0000002800000000ffffffc4ffffffffffffffebffffffff0000002500000000",
            INIT_0C => X"ffffffc7ffffffffffffffe3ffffffffffffffecffffffff0000000400000000",
            INIT_0D => X"0000000d00000000fffffff0ffffffffffffffe6ffffffffffffffd6ffffffff",
            INIT_0E => X"fffffff4ffffffff00000029000000000000000a00000000ffffffdbffffffff",
            INIT_0F => X"fffffffbffffffffffffffe6ffffffffffffffd8ffffffffffffffb8ffffffff",
            INIT_10 => X"0000003300000000fffffff0ffffffffffffffe8ffffffff0000002800000000",
            INIT_11 => X"ffffffeeffffffffffffffc8ffffffffffffffb7ffffffffffffffeaffffffff",
            INIT_12 => X"0000005400000000fffffff2ffffffff0000001000000000ffffffeaffffffff",
            INIT_13 => X"ffffffeefffffffffffffffbffffffffffffffdaffffffff0000004d00000000",
            INIT_14 => X"0000002900000000ffffffe6ffffffff0000000e00000000ffffffe2ffffffff",
            INIT_15 => X"00000017000000000000001b000000000000002f000000000000002900000000",
            INIT_16 => X"0000001a0000000000000031000000000000001e00000000ffffffffffffffff",
            INIT_17 => X"0000002800000000ffffffc2ffffffffffffffc7ffffffffffffffd9ffffffff",
            INIT_18 => X"0000003a000000000000003f0000000000000013000000000000001800000000",
            INIT_19 => X"0000001100000000ffffffedfffffffffffffff0ffffffff0000001800000000",
            INIT_1A => X"fffffff1ffffffffffffffecfffffffffffffff5ffffffffffffffcfffffffff",
            INIT_1B => X"00000049000000000000002e00000000ffffffeefffffffffffffffaffffffff",
            INIT_1C => X"00000024000000000000001a0000000000000018000000000000001000000000",
            INIT_1D => X"ffffffc8ffffffff0000003a0000000000000020000000000000002800000000",
            INIT_1E => X"ffffffddffffffffffffffcffffffffffffffff5ffffffffffffffd7ffffffff",
            INIT_1F => X"00000003000000000000000700000000fffffff9ffffffffffffffd9ffffffff",
            INIT_20 => X"ffffffdcffffffff000000000000000000000021000000000000000c00000000",
            INIT_21 => X"00000028000000000000000000000000fffffff4ffffffffffffffdcffffffff",
            INIT_22 => X"00000035000000000000000c00000000ffffffe4ffffffff0000000a00000000",
            INIT_23 => X"0000000600000000ffffffedfffffffffffffffbffffffff0000000900000000",
            INIT_24 => X"fffffff7fffffffffffffff9fffffffffffffff8ffffffff0000001500000000",
            INIT_25 => X"00000025000000000000000e0000000000000042000000000000001200000000",
            INIT_26 => X"ffffffeeffffffff000000190000000000000028000000000000006e00000000",
            INIT_27 => X"ffffffe5ffffffffffffffa2fffffffffffffff0ffffffffffffffc3ffffffff",
            INIT_28 => X"00000009000000000000003c000000000000000000000000ffffffbcffffffff",
            INIT_29 => X"00000005000000000000000d000000000000003f000000000000002300000000",
            INIT_2A => X"ffffffe5ffffffffffffffedfffffffffffffffaffffffff0000001400000000",
            INIT_2B => X"ffffffedffffffffffffffdbffffffff0000000d00000000fffffff5ffffffff",
            INIT_2C => X"0000005100000000000000310000000000000030000000000000002c00000000",
            INIT_2D => X"0000003500000000000000150000000000000046000000000000003000000000",
            INIT_2E => X"fffffff2fffffffffffffffdffffffff00000005000000000000000e00000000",
            INIT_2F => X"ffffffdcfffffffffffffffcffffffff0000000000000000ffffffffffffffff",
            INIT_30 => X"0000000400000000fffffff1ffffffffffffffeeffffffffffffffcdffffffff",
            INIT_31 => X"0000000100000000ffffffeeffffffffffffffe1ffffffff0000000d00000000",
            INIT_32 => X"ffffffd2ffffffffffffffd5ffffffff0000000600000000ffffffd7ffffffff",
            INIT_33 => X"ffffffffffffffff0000000000000000ffffffc0ffffffffffffffecffffffff",
            INIT_34 => X"000000020000000000000035000000000000001900000000ffffffdfffffffff",
            INIT_35 => X"0000001700000000ffffffccffffffffffffffe0ffffffffffffffdcffffffff",
            INIT_36 => X"0000003b000000000000003b00000000fffffff7ffffffff0000001a00000000",
            INIT_37 => X"ffffffbefffffffffffffff9ffffffffffffffebfffffffffffffff9ffffffff",
            INIT_38 => X"0000004200000000ffffffdefffffffffffffffaffffffff0000000f00000000",
            INIT_39 => X"0000000700000000000000240000000000000003000000000000003500000000",
            INIT_3A => X"0000000100000000fffffffbffffffff00000013000000000000001200000000",
            INIT_3B => X"ffffffcbffffffffffffffeeffffffffffffffcbffffffffffffffdcffffffff",
            INIT_3C => X"0000002d000000000000000100000000ffffffecffffffffffffffd5ffffffff",
            INIT_3D => X"ffffffcfffffffff0000000c000000000000000a00000000ffffffedffffffff",
            INIT_3E => X"ffffffd8ffffffff00000000000000000000003400000000ffffffb9ffffffff",
            INIT_3F => X"0000001800000000ffffffccffffffff00000018000000000000004000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe2ffffffffffffffc9ffffffff00000023000000000000004b00000000",
            INIT_41 => X"fffffffcffffffff000000040000000000000005000000000000004500000000",
            INIT_42 => X"0000002d00000000fffffff8ffffffffffffffe1ffffffffffffffe5ffffffff",
            INIT_43 => X"0000003c00000000fffffffafffffffffffffff3ffffffff0000001a00000000",
            INIT_44 => X"0000001e00000000fffffffaffffffffffffffbeffffffffffffffe1ffffffff",
            INIT_45 => X"000000230000000000000014000000000000002d000000000000004400000000",
            INIT_46 => X"fffffff1ffffffff0000000800000000ffffffefffffffff0000001c00000000",
            INIT_47 => X"0000000d000000000000000a00000000ffffffd5ffffffffffffffefffffffff",
            INIT_48 => X"fffffffdfffffffffffffff1ffffffff0000001300000000ffffffdaffffffff",
            INIT_49 => X"000000480000000000000043000000000000000c000000000000003a00000000",
            INIT_4A => X"ffffffbdffffffff0000002f000000000000001d000000000000000d00000000",
            INIT_4B => X"ffffffe8ffffffff0000000200000000ffffffd5ffffffffffffffd7ffffffff",
            INIT_4C => X"00000010000000000000002a000000000000002200000000ffffffecffffffff",
            INIT_4D => X"0000000300000000fffffff7ffffffff0000000d000000000000002a00000000",
            INIT_4E => X"ffffffe7fffffffffffffffdffffffff0000002c000000000000001800000000",
            INIT_4F => X"0000000100000000ffffffefffffffffffffffeaffffffff0000001300000000",
            INIT_50 => X"00000008000000000000000000000000fffffffaffffffff0000000000000000",
            INIT_51 => X"0000000700000000fffffff7fffffffffffffff2ffffffff0000000a00000000",
            INIT_52 => X"fffffff4ffffffff0000001300000000ffffffedffffffff0000001200000000",
            INIT_53 => X"fffffff5fffffffffffffff5fffffffffffffff6ffffffff0000000200000000",
            INIT_54 => X"0000000700000000fffffffcfffffffffffffffafffffffffffffff3ffffffff",
            INIT_55 => X"fffffff0fffffffffffffff3fffffffffffffff9ffffffff0000000a00000000",
            INIT_56 => X"0000000000000000fffffffbfffffffffffffff9ffffffff0000001000000000",
            INIT_57 => X"ffffffffffffffff0000000000000000fffffff5ffffffff0000000e00000000",
            INIT_58 => X"0000000b00000000fffffff4ffffffff00000007000000000000000200000000",
            INIT_59 => X"0000000000000000ffffffe6ffffffffffffffedfffffffffffffffdffffffff",
            INIT_5A => X"ffffffffffffffffffffffeeffffffff0000000000000000fffffffcffffffff",
            INIT_5B => X"000000030000000000000000000000000000000500000000fffffff9ffffffff",
            INIT_5C => X"ffffffebfffffffffffffff4fffffffffffffff4fffffffffffffff7ffffffff",
            INIT_5D => X"fffffff6fffffffffffffffefffffffffffffff1fffffffffffffffcffffffff",
            INIT_5E => X"0000000000000000ffffffecfffffffffffffffdffffffff0000001000000000",
            INIT_5F => X"fffffff3fffffffffffffff6ffffffff00000004000000000000000000000000",
            INIT_60 => X"ffffffe9ffffffff00000001000000000000000d00000000fffffff4ffffffff",
            INIT_61 => X"fffffffaffffffff000000030000000000000010000000000000000400000000",
            INIT_62 => X"fffffffdffffffffffffffefffffffff0000000900000000fffffff1ffffffff",
            INIT_63 => X"0000000000000000fffffffcfffffffffffffffbfffffffffffffff0ffffffff",
            INIT_64 => X"0000000a0000000000000000000000000000000a00000000fffffffbffffffff",
            INIT_65 => X"0000000300000000000000110000000000000003000000000000000a00000000",
            INIT_66 => X"0000001300000000fffffffdfffffffffffffff5fffffffffffffff6ffffffff",
            INIT_67 => X"0000000400000000fffffffeffffffff0000000200000000fffffffbffffffff",
            INIT_68 => X"fffffff9fffffffffffffffdfffffffffffffff1ffffffff0000001700000000",
            INIT_69 => X"fffffff5ffffffff0000000c0000000000000007000000000000000600000000",
            INIT_6A => X"000000070000000000000000000000000000000000000000fffffff3ffffffff",
            INIT_6B => X"fffffff7ffffffff0000000200000000ffffffecffffffff0000000f00000000",
            INIT_6C => X"0000000d00000000000000000000000000000001000000000000000300000000",
            INIT_6D => X"0000000b00000000ffffffebffffffff0000000600000000fffffffdffffffff",
            INIT_6E => X"fffffff5fffffffffffffff0ffffffff0000000200000000ffffffefffffffff",
            INIT_6F => X"0000000e00000000fffffffdfffffffffffffffbfffffffffffffff7ffffffff",
            INIT_70 => X"0000000b00000000fffffff9ffffffff00000000000000000000000000000000",
            INIT_71 => X"0000000300000000fffffff4ffffffffffffffecfffffffffffffff1ffffffff",
            INIT_72 => X"0000000600000000ffffffeaffffffffffffffeaffffffff0000000000000000",
            INIT_73 => X"ffffffeaffffffff0000001100000000ffffffecffffffffffffffffffffffff",
            INIT_74 => X"fffffff0ffffffffffffffeeffffffff00000011000000000000001000000000",
            INIT_75 => X"0000000500000000fffffff5ffffffff0000000f000000000000000c00000000",
            INIT_76 => X"fffffff6fffffffffffffff8ffffffffffffffebffffffff0000000e00000000",
            INIT_77 => X"00000004000000000000000700000000fffffff5ffffffff0000000000000000",
            INIT_78 => X"000000110000000000000015000000000000000a00000000fffffff1ffffffff",
            INIT_79 => X"fffffffbffffffff0000000700000000fffffff3ffffffff0000000200000000",
            INIT_7A => X"0000000300000000fffffff0fffffffffffffff9fffffffffffffffaffffffff",
            INIT_7B => X"0000000c00000000fffffff3ffffffffffffffedffffffff0000000e00000000",
            INIT_7C => X"0000000200000000ffffffffffffffff0000000e00000000fffffff3ffffffff",
            INIT_7D => X"0000000400000000ffffffe8fffffffffffffffffffffffffffffff9ffffffff",
            INIT_7E => X"0000000300000000fffffff5ffffffff00000002000000000000000d00000000",
            INIT_7F => X"fffffff4ffffffff0000000b000000000000000600000000fffffffdffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE13;


    MEM_IWGHT_LAYER2_INSTANCE14 : if BRAM_NAME = "iwght_layer2_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000009000000000000000a00000000fffffff4ffffffffffffffe9ffffffff",
            INIT_01 => X"0000000d00000000fffffff0ffffffff0000000a00000000ffffffebffffffff",
            INIT_02 => X"ffffffe9ffffffff0000000500000000fffffffafffffffffffffffcffffffff",
            INIT_03 => X"fffffffdfffffffffffffff9ffffffff0000001200000000ffffffeeffffffff",
            INIT_04 => X"fffffff0fffffffffffffff2fffffffffffffff4fffffffffffffff1ffffffff",
            INIT_05 => X"ffffffeaffffffffffffffedfffffffffffffff3ffffffff0000000400000000",
            INIT_06 => X"0000000300000000fffffff6fffffffffffffff8fffffffffffffff0ffffffff",
            INIT_07 => X"fffffffeffffffff00000005000000000000000a00000000fffffffeffffffff",
            INIT_08 => X"ffffffe8fffffffffffffffefffffffffffffff4ffffffffffffffe8ffffffff",
            INIT_09 => X"0000000300000000fffffff9fffffffffffffff3ffffffff0000000400000000",
            INIT_0A => X"fffffff6fffffffffffffffeffffffff0000000000000000fffffffeffffffff",
            INIT_0B => X"fffffff6ffffffff0000000f0000000000000005000000000000000b00000000",
            INIT_0C => X"fffffff6ffffffff0000000d0000000000000007000000000000001100000000",
            INIT_0D => X"fffffffbffffffffffffffeffffffffffffffff5ffffffff0000000900000000",
            INIT_0E => X"ffffffeeffffffff0000000400000000ffffffebfffffffffffffffaffffffff",
            INIT_0F => X"fffffff8ffffffff00000004000000000000000000000000fffffff6ffffffff",
            INIT_10 => X"0000000300000000fffffff6fffffffffffffff5ffffffff0000000100000000",
            INIT_11 => X"fffffff2fffffffffffffff8ffffffff0000000000000000fffffff5ffffffff",
            INIT_12 => X"0000000000000000fffffffcfffffffffffffff9ffffffffffffffebffffffff",
            INIT_13 => X"0000000900000000ffffffeaffffffffffffffecffffffff0000000700000000",
            INIT_14 => X"fffffff9ffffffff0000000000000000ffffffeefffffffffffffff3ffffffff",
            INIT_15 => X"00000006000000000000000300000000fffffffbfffffffffffffff7ffffffff",
            INIT_16 => X"fffffffbfffffffffffffff9ffffffffffffffffffffffff0000000800000000",
            INIT_17 => X"ffffffe9fffffffffffffff4fffffffffffffff3ffffffffffffffeeffffffff",
            INIT_18 => X"fffffff8fffffffffffffffefffffffffffffffafffffffffffffff8ffffffff",
            INIT_19 => X"ffffffe9ffffffff0000000600000000ffffffe7ffffffff0000000800000000",
            INIT_1A => X"00000002000000000000001500000000fffffffdffffffffffffffeeffffffff",
            INIT_1B => X"fffffffaffffffffffffffd5ffffffffffffffe9fffffffffffffffdffffffff",
            INIT_1C => X"fffffffcffffffffffffffddfffffffffffffff3ffffffffffffffe4ffffffff",
            INIT_1D => X"0000001f000000000000001400000000fffffffcffffffffffffffdfffffffff",
            INIT_1E => X"0000001d00000000000000280000000000000043000000000000002e00000000",
            INIT_1F => X"00000018000000000000003a0000000000000040000000000000004800000000",
            INIT_20 => X"ffffffe6ffffffff00000002000000000000000b000000000000001e00000000",
            INIT_21 => X"0000003000000000ffffffdafffffffffffffff2fffffffffffffff9ffffffff",
            INIT_22 => X"00000031000000000000002c00000000fffffff0ffffffff0000000b00000000",
            INIT_23 => X"fffffff7ffffffffffffffe0fffffffffffffffbffffffff0000003300000000",
            INIT_24 => X"ffffffe9ffffffffffffffeefffffffffffffffdffffffffffffffe0ffffffff",
            INIT_25 => X"0000000a00000000ffffffeaffffffffffffffe1ffffffff0000001700000000",
            INIT_26 => X"fffffff7ffffffffffffffd7fffffffffffffffefffffffffffffffeffffffff",
            INIT_27 => X"0000000500000000ffffffe9fffffffffffffff6fffffffffffffff4ffffffff",
            INIT_28 => X"0000002200000000000000130000000000000004000000000000001800000000",
            INIT_29 => X"0000000000000000000000270000000000000020000000000000002600000000",
            INIT_2A => X"0000001b0000000000000019000000000000001c000000000000001600000000",
            INIT_2B => X"ffffffe9ffffffff0000000d000000000000000100000000fffffff4ffffffff",
            INIT_2C => X"ffffffe8ffffffffffffff9affffffffffffffb2ffffffff0000000600000000",
            INIT_2D => X"0000002200000000ffffffe5ffffffffffffffc3ffffffffffffffdbffffffff",
            INIT_2E => X"0000002f00000000000000080000000000000024000000000000000000000000",
            INIT_2F => X"ffffffefffffffffffffffdbfffffffffffffff2ffffffff0000000200000000",
            INIT_30 => X"ffffffc9ffffffffffffffe0ffffffffffffffe8ffffffff0000000c00000000",
            INIT_31 => X"ffffffc4ffffffffffffffd2ffffffffffffffe6ffffffffffffffc1ffffffff",
            INIT_32 => X"ffffffcfffffffffffffffbfffffffffffffffeeffffffffffffffd5ffffffff",
            INIT_33 => X"fffffffcffffffffffffffe5ffffffffffffffceffffffff0000000100000000",
            INIT_34 => X"00000021000000000000001300000000fffffff5ffffffff0000000300000000",
            INIT_35 => X"00000002000000000000000c00000000ffffffedffffffff0000001000000000",
            INIT_36 => X"0000001700000000fffffffeffffffff00000005000000000000000200000000",
            INIT_37 => X"ffffffeeffffffff00000016000000000000002e000000000000000d00000000",
            INIT_38 => X"0000001500000000fffffff2ffffffff0000001000000000fffffff6ffffffff",
            INIT_39 => X"ffffffeaffffffffffffffeffffffffffffffff9ffffffff0000000100000000",
            INIT_3A => X"fffffff2ffffffffffffffddfffffffffffffff2ffffffffffffffd1ffffffff",
            INIT_3B => X"0000001e0000000000000009000000000000000700000000fffffff9ffffffff",
            INIT_3C => X"ffffffafffffffffffffffefffffffffffffffc6ffffffffffffffcfffffffff",
            INIT_3D => X"ffffffe0ffffffffffffffe5ffffffffffffffddffffffffffffffaeffffffff",
            INIT_3E => X"fffffffffffffffffffffff7ffffffffffffffc7ffffffffffffffcdffffffff",
            INIT_3F => X"fffffffdffffffff0000000900000000ffffffc3ffffffff0000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001b0000000000000001000000000000000700000000fffffff8ffffffff",
            INIT_41 => X"ffffffb1ffffffffffffffb1ffffffffffffffb8fffffffffffffff4ffffffff",
            INIT_42 => X"0000002800000000ffffffc7ffffffffffffffa3ffffffffffffffbaffffffff",
            INIT_43 => X"0000002c000000000000002600000000ffffffecffffffff0000000900000000",
            INIT_44 => X"0000001f00000000000000130000000000000025000000000000000600000000",
            INIT_45 => X"0000001300000000fffffff4ffffffff00000001000000000000001500000000",
            INIT_46 => X"ffffffecffffffffffffffdefffffffffffffff1ffffffffffffffebffffffff",
            INIT_47 => X"ffffffecffffffff0000000b000000000000002700000000fffffff5ffffffff",
            INIT_48 => X"0000000900000000000000040000000000000013000000000000002b00000000",
            INIT_49 => X"ffffffebffffffffffffffd5ffffffff0000000900000000fffffffaffffffff",
            INIT_4A => X"0000000600000000ffffffd1fffffffffffffff2fffffffffffffff6ffffffff",
            INIT_4B => X"fffffffeffffffff0000001c000000000000000a000000000000001600000000",
            INIT_4C => X"fffffffffffffffffffffff3ffffffff00000014000000000000000700000000",
            INIT_4D => X"ffffffffffffffff0000000700000000fffffff9ffffffff0000000400000000",
            INIT_4E => X"0000002c00000000000000190000000000000030000000000000002000000000",
            INIT_4F => X"fffffffbffffffff0000000000000000fffffffdffffffff0000002900000000",
            INIT_50 => X"0000002000000000000000420000000000000024000000000000000b00000000",
            INIT_51 => X"0000002300000000000000240000000000000007000000000000002300000000",
            INIT_52 => X"ffffffbdffffffffffffffb7ffffffff00000017000000000000000100000000",
            INIT_53 => X"0000000700000000fffffffcffffffffffffffc7fffffffffffffff7ffffffff",
            INIT_54 => X"000000170000000000000020000000000000000b00000000fffffffdffffffff",
            INIT_55 => X"0000002800000000fffffffcfffffffffffffffbffffffffffffffe2ffffffff",
            INIT_56 => X"000000130000000000000006000000000000000a000000000000001f00000000",
            INIT_57 => X"000000240000000000000024000000000000002e000000000000004100000000",
            INIT_58 => X"ffffffeeffffffff0000000b0000000000000014000000000000001400000000",
            INIT_59 => X"0000000c00000000ffffffcaffffffffffffffdcfffffffffffffff0ffffffff",
            INIT_5A => X"0000000d000000000000000300000000ffffffdaffffffff0000000400000000",
            INIT_5B => X"00000010000000000000000f0000000000000001000000000000000800000000",
            INIT_5C => X"0000001d000000000000000b0000000000000028000000000000001300000000",
            INIT_5D => X"ffffffedfffffffffffffff2ffffffffffffffeffffffffffffffff5ffffffff",
            INIT_5E => X"ffffffdcffffffffffffffbeffffffff0000000200000000ffffffb8ffffffff",
            INIT_5F => X"000000220000000000000014000000000000000b000000000000001000000000",
            INIT_60 => X"00000007000000000000001500000000fffffff9ffffffff0000000000000000",
            INIT_61 => X"0000000600000000fffffffdfffffffffffffff7fffffffffffffff6ffffffff",
            INIT_62 => X"000000280000000000000013000000000000003500000000ffffffe9ffffffff",
            INIT_63 => X"00000003000000000000002300000000fffffff9ffffffff0000000300000000",
            INIT_64 => X"fffffffcffffffff0000002a0000000000000002000000000000000000000000",
            INIT_65 => X"00000015000000000000002e000000000000002d000000000000003c00000000",
            INIT_66 => X"ffffffc8ffffffff000000160000000000000030000000000000002c00000000",
            INIT_67 => X"ffffffdffffffffffffffff7ffffffffffffffe9fffffffffffffff1ffffffff",
            INIT_68 => X"ffffffcfffffffff0000000c000000000000001200000000ffffffeeffffffff",
            INIT_69 => X"0000003700000000ffffffccffffffff0000001900000000ffffffefffffffff",
            INIT_6A => X"0000001d00000000000000140000000000000014000000000000003500000000",
            INIT_6B => X"ffffffd8ffffffffffffffddffffffffffffffdbffffffff0000000200000000",
            INIT_6C => X"0000000e00000000000000230000000000000027000000000000000e00000000",
            INIT_6D => X"00000038000000000000004d0000000000000007000000000000001e00000000",
            INIT_6E => X"00000020000000000000001c000000000000000e000000000000003300000000",
            INIT_6F => X"0000001c00000000ffffffc3ffffffffffffffc7fffffffffffffff5ffffffff",
            INIT_70 => X"fffffff7ffffffffffffffe9ffffffff00000016000000000000003300000000",
            INIT_71 => X"fffffffbffffffffffffffc9ffffffffffffffe8ffffffffffffffd3ffffffff",
            INIT_72 => X"00000001000000000000000700000000fffffff8ffffffff0000002e00000000",
            INIT_73 => X"0000001b0000000000000012000000000000002a000000000000002c00000000",
            INIT_74 => X"fffffffeffffffff00000011000000000000002c000000000000001700000000",
            INIT_75 => X"0000002600000000ffffffe7ffffffffffffffdfffffffff0000002b00000000",
            INIT_76 => X"ffffffebffffffff0000000100000000ffffffefffffffff0000000000000000",
            INIT_77 => X"00000033000000000000000000000000ffffffddffffffff0000000600000000",
            INIT_78 => X"fffffff6fffffffffffffff3fffffffffffffff2ffffffffffffffe9ffffffff",
            INIT_79 => X"0000001f00000000ffffffe2ffffffff0000000e000000000000002d00000000",
            INIT_7A => X"ffffffe0ffffffffffffffdcffffffff00000007000000000000001e00000000",
            INIT_7B => X"0000000a00000000000000040000000000000004000000000000001b00000000",
            INIT_7C => X"fffffff8ffffffff0000000600000000ffffffdfffffffff0000001100000000",
            INIT_7D => X"000000350000000000000012000000000000003000000000ffffffe3ffffffff",
            INIT_7E => X"fffffff2ffffffffffffffddffffffffffffffe2ffffffff0000000200000000",
            INIT_7F => X"0000000d000000000000000c00000000ffffffe9ffffffffffffffe5ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE14;


    MEM_IWGHT_LAYER2_INSTANCE15 : if BRAM_NAME = "iwght_layer2_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000021000000000000003f000000000000001000000000ffffffedffffffff",
            INIT_01 => X"000000060000000000000018000000000000003e000000000000001000000000",
            INIT_02 => X"fffffffaffffffff0000001d0000000000000003000000000000000800000000",
            INIT_03 => X"0000000100000000ffffffe7fffffffffffffff6ffffffffffffffe5ffffffff",
            INIT_04 => X"0000000b000000000000001300000000fffffffbffffffffffffffe4ffffffff",
            INIT_05 => X"ffffffd6ffffffffffffffd1ffffffff0000002900000000ffffffefffffffff",
            INIT_06 => X"000000280000000000000010000000000000001a00000000fffffff9ffffffff",
            INIT_07 => X"fffffff6ffffffff0000002700000000fffffff4ffffffff0000000500000000",
            INIT_08 => X"0000000600000000fffffff6ffffffffffffffe9ffffffffffffffdeffffffff",
            INIT_09 => X"000000090000000000000004000000000000001800000000fffffff5ffffffff",
            INIT_0A => X"0000000e00000000fffffff1ffffffff00000007000000000000002400000000",
            INIT_0B => X"00000035000000000000000800000000fffffff4fffffffffffffffdffffffff",
            INIT_0C => X"fffffff6ffffffff0000000800000000fffffff2ffffffff0000000000000000",
            INIT_0D => X"0000000a00000000fffffff4fffffffffffffff2fffffffffffffffdffffffff",
            INIT_0E => X"0000000e00000000fffffff6ffffffffffffffdeffffffff0000000300000000",
            INIT_0F => X"ffffffe9ffffffff000000010000000000000000000000000000000600000000",
            INIT_10 => X"0000001c00000000000000100000000000000013000000000000000f00000000",
            INIT_11 => X"0000002a000000000000004a000000000000000f000000000000000b00000000",
            INIT_12 => X"00000017000000000000000b0000000000000015000000000000002800000000",
            INIT_13 => X"ffffffe3fffffffffffffff7ffffffffffffffefffffffff0000002800000000",
            INIT_14 => X"0000000a000000000000000500000000ffffffd7fffffffffffffff2ffffffff",
            INIT_15 => X"ffffffe0fffffffffffffffbffffffff0000000d00000000fffffff5ffffffff",
            INIT_16 => X"00000012000000000000000000000000ffffffcfffffffff0000000100000000",
            INIT_17 => X"0000000100000000ffffffdcffffffff0000003f00000000fffffff8ffffffff",
            INIT_18 => X"fffffffaffffffff0000000b00000000fffffffeffffffff0000002200000000",
            INIT_19 => X"ffffffbcffffffffffffffdcffffffffffffffe7ffffffffffffffefffffffff",
            INIT_1A => X"fffffffdffffffff0000001300000000ffffffb5ffffffffffffffc7ffffffff",
            INIT_1B => X"0000000100000000ffffffe1ffffffff0000001100000000ffffffffffffffff",
            INIT_1C => X"0000004800000000fffffffeffffffffffffffd8ffffffff0000001900000000",
            INIT_1D => X"000000030000000000000019000000000000001e000000000000001300000000",
            INIT_1E => X"fffffff3fffffffffffffff4fffffffffffffffeffffffff0000001100000000",
            INIT_1F => X"0000000100000000fffffff4fffffffffffffff6fffffffffffffff1ffffffff",
            INIT_20 => X"0000003a000000000000001a000000000000001f000000000000000400000000",
            INIT_21 => X"000000190000000000000025000000000000002000000000fffffff1ffffffff",
            INIT_22 => X"fffffffbfffffffffffffff8ffffffff00000002000000000000001b00000000",
            INIT_23 => X"fffffffaffffffffffffffe1ffffffff0000001300000000ffffffdbffffffff",
            INIT_24 => X"fffffff1fffffffffffffff5fffffffffffffff7ffffffffffffffddffffffff",
            INIT_25 => X"0000001e00000000ffffffebffffffff0000000100000000ffffffe9ffffffff",
            INIT_26 => X"ffffffd7fffffffffffffff5fffffffffffffffbffffffff0000001000000000",
            INIT_27 => X"ffffffedffffffff00000001000000000000001900000000fffffff6ffffffff",
            INIT_28 => X"0000001400000000ffffffebffffffffffffffeeffffffff0000000a00000000",
            INIT_29 => X"0000000a00000000000000150000000000000008000000000000000300000000",
            INIT_2A => X"ffffffeffffffffffffffff0ffffffffffffffe7ffffffff0000000000000000",
            INIT_2B => X"0000000800000000fffffffeffffffffffffffeaffffffff0000000100000000",
            INIT_2C => X"0000000a00000000000000020000000000000000000000000000000200000000",
            INIT_2D => X"0000000800000000fffffff5ffffffffffffffedffffffff0000000500000000",
            INIT_2E => X"ffffffe8ffffffffffffffedffffffffffffffebfffffffffffffffdffffffff",
            INIT_2F => X"00000004000000000000000d00000000fffffff4ffffffff0000000b00000000",
            INIT_30 => X"fffffffdffffffff00000002000000000000001100000000fffffff3ffffffff",
            INIT_31 => X"0000000700000000fffffff6fffffffffffffffdffffffff0000000200000000",
            INIT_32 => X"0000000a000000000000000c00000000fffffff6ffffffff0000001500000000",
            INIT_33 => X"fffffffcfffffffffffffff8fffffffffffffffeffffffff0000000200000000",
            INIT_34 => X"0000000500000000ffffffe6ffffffff0000000b00000000fffffffeffffffff",
            INIT_35 => X"00000007000000000000000b000000000000000300000000ffffffffffffffff",
            INIT_36 => X"fffffff4fffffffffffffff4ffffffff0000000000000000ffffffffffffffff",
            INIT_37 => X"00000007000000000000000600000000ffffffe5fffffffffffffff1ffffffff",
            INIT_38 => X"ffffffeafffffffffffffffcffffffff0000000100000000ffffffebffffffff",
            INIT_39 => X"0000000100000000fffffff6fffffffffffffffbfffffffffffffff8ffffffff",
            INIT_3A => X"ffffffefffffffff00000005000000000000000900000000fffffff1ffffffff",
            INIT_3B => X"fffffff2fffffffffffffff5ffffffffffffffe7fffffffffffffff0ffffffff",
            INIT_3C => X"ffffffebfffffffffffffff1ffffffff0000000c00000000ffffffedffffffff",
            INIT_3D => X"ffffffe8ffffffffffffffe7ffffffff00000000000000000000000900000000",
            INIT_3E => X"0000000500000000ffffffe7fffffffffffffff9ffffffffffffffe5ffffffff",
            INIT_3F => X"ffffffeeffffffff0000000a0000000000000001000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000a00000000ffffffeefffffffffffffff9fffffffffffffffdffffffff",
            INIT_41 => X"fffffff5ffffffff0000000f00000000fffffffdfffffffffffffff9ffffffff",
            INIT_42 => X"fffffffdffffffff00000000000000000000000000000000fffffff9ffffffff",
            INIT_43 => X"fffffff1fffffffffffffffcffffffffffffffebffffffffffffffecffffffff",
            INIT_44 => X"fffffffaffffffff00000009000000000000000b00000000ffffffe5ffffffff",
            INIT_45 => X"fffffff4ffffffff0000000900000000ffffffefffffffffffffffffffffffff",
            INIT_46 => X"fffffffcfffffffffffffffeffffffff0000000200000000fffffff5ffffffff",
            INIT_47 => X"fffffff5ffffffffffffffe6ffffffffffffffe6ffffffff0000000000000000",
            INIT_48 => X"fffffff1ffffffff00000000000000000000000100000000ffffffe9ffffffff",
            INIT_49 => X"fffffff0ffffffff000000020000000000000004000000000000000400000000",
            INIT_4A => X"0000000f000000000000000f0000000000000007000000000000000400000000",
            INIT_4B => X"0000000100000000fffffff9fffffffffffffff1fffffffffffffff1ffffffff",
            INIT_4C => X"0000000000000000fffffff5fffffffffffffff3fffffffffffffffcffffffff",
            INIT_4D => X"0000000700000000fffffff1ffffffff00000000000000000000000b00000000",
            INIT_4E => X"00000001000000000000000b000000000000000300000000fffffffcffffffff",
            INIT_4F => X"ffffffeafffffffffffffff9ffffffff0000000200000000ffffffebffffffff",
            INIT_50 => X"0000000d00000000fffffff5ffffffffffffffeeffffffff0000000900000000",
            INIT_51 => X"00000000000000000000000200000000ffffffecffffffff0000000800000000",
            INIT_52 => X"00000007000000000000000f000000000000000f00000000ffffffecffffffff",
            INIT_53 => X"fffffff3fffffffffffffffffffffffffffffff2fffffffffffffffcffffffff",
            INIT_54 => X"fffffff6ffffffffffffffe3fffffffffffffffefffffffffffffff6ffffffff",
            INIT_55 => X"ffffffecffffffff0000000b00000000fffffff9fffffffffffffff2ffffffff",
            INIT_56 => X"fffffff0ffffffffffffffe3ffffffffffffffedfffffffffffffff8ffffffff",
            INIT_57 => X"00000005000000000000000e00000000ffffffebffffffff0000000000000000",
            INIT_58 => X"ffffffeefffffffffffffff6ffffffff0000000d000000000000000700000000",
            INIT_59 => X"0000000d000000000000000000000000ffffffecffffffff0000000e00000000",
            INIT_5A => X"fffffff8ffffffffffffffefffffffff0000000400000000ffffffffffffffff",
            INIT_5B => X"fffffff0ffffffff0000000700000000ffffffedfffffffffffffff4ffffffff",
            INIT_5C => X"ffffffeafffffffffffffff0ffffffff00000000000000000000000400000000",
            INIT_5D => X"0000000500000000ffffffeeffffffff0000000700000000fffffff9ffffffff",
            INIT_5E => X"fffffff2ffffffffffffffe7ffffffff00000002000000000000000000000000",
            INIT_5F => X"0000000b000000000000000700000000ffffffe4ffffffff0000000400000000",
            INIT_60 => X"00000003000000000000000000000000ffffffe1ffffffffffffffedffffffff",
            INIT_61 => X"fffffff4ffffffffffffffdeffffffffffffffdfffffffffffffffe6ffffffff",
            INIT_62 => X"0000000600000000fffffff8ffffffffffffffefffffffffffffffe0ffffffff",
            INIT_63 => X"fffffffdfffffffffffffff3fffffffffffffff6ffffffff0000001300000000",
            INIT_64 => X"ffffffe9fffffffffffffff0ffffffff0000000000000000fffffff6ffffffff",
            INIT_65 => X"fffffff8fffffffffffffffaffffffff0000000100000000fffffff3ffffffff",
            INIT_66 => X"ffffffe7ffffffff0000000500000000ffffffecffffffffffffffebffffffff",
            INIT_67 => X"fffffffdffffffffffffffe6ffffffff0000000700000000fffffff4ffffffff",
            INIT_68 => X"00000005000000000000001300000000fffffff2ffffffff0000000700000000",
            INIT_69 => X"0000000b00000000ffffffecffffffffffffffffffffffffffffffe3ffffffff",
            INIT_6A => X"fffffff3ffffffff0000000500000000fffffff4ffffffff0000001000000000",
            INIT_6B => X"ffffffe7fffffffffffffffbfffffffffffffffcffffffffffffffe5ffffffff",
            INIT_6C => X"fffffffefffffffffffffff2fffffffffffffff5ffffffff0000000000000000",
            INIT_6D => X"fffffff4fffffffffffffffdffffffff0000000600000000ffffffebffffffff",
            INIT_6E => X"ffffffecfffffffffffffff9fffffffffffffffdfffffffffffffff4ffffffff",
            INIT_6F => X"0000000500000000ffffffe8ffffffff0000000f000000000000000600000000",
            INIT_70 => X"ffffffedffffffff0000001200000000fffffffdfffffffffffffff6ffffffff",
            INIT_71 => X"0000000600000000fffffffdfffffffffffffffeffffffff0000001400000000",
            INIT_72 => X"ffffffebfffffffffffffffdffffffff0000000400000000ffffffefffffffff",
            INIT_73 => X"00000003000000000000000a0000000000000003000000000000000900000000",
            INIT_74 => X"fffffff7ffffffffffffffedffffffff0000000000000000ffffffffffffffff",
            INIT_75 => X"000000110000000000000004000000000000000500000000fffffffdffffffff",
            INIT_76 => X"0000000000000000ffffffe9ffffffff00000005000000000000000100000000",
            INIT_77 => X"fffffff7ffffffffffffffefffffffffffffffecffffffffffffffebffffffff",
            INIT_78 => X"fffffff2fffffffffffffff7ffffffff0000000900000000ffffffecffffffff",
            INIT_79 => X"fffffffcffffffff0000000300000000fffffff3ffffffffffffffeeffffffff",
            INIT_7A => X"fffffff4fffffffffffffff0ffffffff00000006000000000000000900000000",
            INIT_7B => X"0000000200000000ffffffe4ffffffffffffffe9ffffffffffffffeeffffffff",
            INIT_7C => X"0000000900000000ffffffe2ffffffffffffffefffffffffffffffe4ffffffff",
            INIT_7D => X"ffffffe8fffffffffffffff4fffffffffffffff4ffffffff0000000b00000000",
            INIT_7E => X"00000002000000000000000200000000fffffff5fffffffffffffffeffffffff",
            INIT_7F => X"ffffffeafffffffffffffffeffffffffffffffecfffffffffffffffaffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE15;


    MEM_IWGHT_LAYER2_INSTANCE16 : if BRAM_NAME = "iwght_layer2_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff6ffffffff0000000500000000fffffff9fffffffffffffff3ffffffff",
            INIT_01 => X"ffffffecffffffffffffffe7fffffffffffffff5fffffffffffffff1ffffffff",
            INIT_02 => X"0000000000000000ffffffe7ffffffffffffffefffffffff0000000700000000",
            INIT_03 => X"0000000b000000000000000000000000fffffffeffffffff0000000000000000",
            INIT_04 => X"fffffff6fffffffffffffff0ffffffff00000006000000000000000300000000",
            INIT_05 => X"00000008000000000000000800000000fffffffeffffffffffffffedffffffff",
            INIT_06 => X"0000000500000000000000000000000000000005000000000000000800000000",
            INIT_07 => X"0000000500000000ffffffe3fffffffffffffffcfffffffffffffffcffffffff",
            INIT_08 => X"ffffffebffffffff0000000000000000fffffff7fffffffffffffff5ffffffff",
            INIT_09 => X"ffffffe9ffffffffffffffeaffffffff0000000b00000000fffffff9ffffffff",
            INIT_0A => X"0000000300000000ffffffe9fffffffffffffffcffffffff0000000e00000000",
            INIT_0B => X"0000000500000000fffffffaffffffff0000000f000000000000000800000000",
            INIT_0C => X"0000000b000000000000000f0000000000000008000000000000000900000000",
            INIT_0D => X"0000000c00000000000000040000000000000002000000000000000400000000",
            INIT_0E => X"0000000a00000000ffffffecfffffffffffffffdffffffffffffffe9ffffffff",
            INIT_0F => X"0000000a00000000ffffffe9fffffffffffffffffffffffffffffff6ffffffff",
            INIT_10 => X"00000000000000000000000600000000fffffff2fffffffffffffffeffffffff",
            INIT_11 => X"fffffffaffffffffffffffebffffffff00000006000000000000000800000000",
            INIT_12 => X"fffffff8ffffffff0000000000000000fffffff6ffffffff0000000e00000000",
            INIT_13 => X"fffffffcfffffffffffffff7fffffffffffffff3ffffffff0000000100000000",
            INIT_14 => X"fffffff6ffffffff0000000c0000000000000012000000000000000e00000000",
            INIT_15 => X"ffffffedffffffff0000000000000000fffffff1fffffffffffffffeffffffff",
            INIT_16 => X"fffffff4ffffffff0000000600000000fffffff8ffffffff0000000400000000",
            INIT_17 => X"0000000800000000ffffffedffffffffffffffeafffffffffffffffdffffffff",
            INIT_18 => X"0000000500000000fffffffcfffffffffffffff7fffffffffffffffcffffffff",
            INIT_19 => X"fffffffbffffffff0000000500000000fffffff6ffffffff0000000a00000000",
            INIT_1A => X"0000000d00000000fffffffaffffffffffffffefffffffff0000001300000000",
            INIT_1B => X"fffffff9fffffffffffffffcfffffffffffffff9ffffffffffffffeaffffffff",
            INIT_1C => X"ffffffe5ffffffff0000000a00000000ffffffe9fffffffffffffff1ffffffff",
            INIT_1D => X"ffffffffffffffff0000000a00000000ffffffecffffffff0000000200000000",
            INIT_1E => X"fffffff2ffffffff0000000300000000fffffff5fffffffffffffff0ffffffff",
            INIT_1F => X"0000000700000000fffffff4ffffffff0000000200000000ffffffefffffffff",
            INIT_20 => X"ffffffecfffffffffffffff2ffffffff0000000500000000fffffff9ffffffff",
            INIT_21 => X"fffffffbffffffffffffffeffffffffffffffff2ffffffffffffffebffffffff",
            INIT_22 => X"fffffff6fffffffffffffffeffffffff0000000000000000ffffffecffffffff",
            INIT_23 => X"0000000600000000ffffffedffffffff0000000000000000fffffff1ffffffff",
            INIT_24 => X"ffffffffffffffff00000004000000000000000b000000000000000500000000",
            INIT_25 => X"fffffffafffffffffffffff9ffffffffffffffe7fffffffffffffffaffffffff",
            INIT_26 => X"fffffff6ffffffff0000000a000000000000000900000000fffffff4ffffffff",
            INIT_27 => X"ffffffebfffffffffffffffaffffffffffffffe6ffffffff0000000f00000000",
            INIT_28 => X"0000000300000000fffffff2ffffffffffffffebffffffff0000000c00000000",
            INIT_29 => X"ffffffeefffffffffffffff8ffffffffffffffe9ffffffffffffffebffffffff",
            INIT_2A => X"0000000f00000000fffffff9fffffffffffffff3ffffffff0000000400000000",
            INIT_2B => X"fffffff5ffffffffffffffeafffffffffffffff0ffffffff0000000000000000",
            INIT_2C => X"ffffffe9fffffffffffffffcffffffffffffffe4fffffffffffffff8ffffffff",
            INIT_2D => X"ffffffeaffffffffffffffecffffffff00000010000000000000000500000000",
            INIT_2E => X"ffffffeefffffffffffffff5fffffffffffffffafffffffffffffff1ffffffff",
            INIT_2F => X"fffffff5ffffffff0000000700000000fffffffbffffffffffffffeaffffffff",
            INIT_30 => X"fffffff9fffffffffffffff5ffffffff0000000900000000ffffffefffffffff",
            INIT_31 => X"fffffff5ffffffffffffffe5ffffffffffffffeefffffffffffffffaffffffff",
            INIT_32 => X"0000000e0000000000000002000000000000000300000000ffffffebffffffff",
            INIT_33 => X"fffffffaffffffffffffffecffffffff0000000300000000fffffff1ffffffff",
            INIT_34 => X"0000000000000000fffffff5ffffffff0000000500000000fffffffaffffffff",
            INIT_35 => X"ffffffeeffffffffffffffeefffffffffffffff3fffffffffffffffaffffffff",
            INIT_36 => X"fffffffffffffffffffffffeffffffffffffffffffffffff0000000600000000",
            INIT_37 => X"fffffff7ffffffffffffffeeffffffff0000000d00000000fffffff9ffffffff",
            INIT_38 => X"ffffffe9ffffffff000000110000000000000008000000000000000000000000",
            INIT_39 => X"ffffffedfffffffffffffffafffffffffffffff7ffffffff0000000800000000",
            INIT_3A => X"0000001e000000000000002d0000000000000002000000000000000000000000",
            INIT_3B => X"0000001600000000fffffff6ffffffffffffffeeffffffffffffffdcffffffff",
            INIT_3C => X"0000002e00000000000000220000000000000000000000000000000c00000000",
            INIT_3D => X"fffffff4ffffffff000000260000000000000032000000000000000500000000",
            INIT_3E => X"fffffffdfffffffffffffff9ffffffff00000031000000000000003500000000",
            INIT_3F => X"ffffffc9fffffffffffffff2ffffffffffffffd4ffffffffffffffe9ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffb3ffffffffffffffa7ffffffff0000001200000000ffffffa9ffffffff",
            INIT_41 => X"0000003e00000000ffffffd9fffffffffffffffbffffffff0000001e00000000",
            INIT_42 => X"0000000a000000000000003800000000fffffffcffffffff0000000b00000000",
            INIT_43 => X"fffffff2ffffffff0000000b000000000000000b000000000000000a00000000",
            INIT_44 => X"ffffffe9ffffffff000000170000000000000029000000000000001600000000",
            INIT_45 => X"00000022000000000000002a00000000ffffffe2ffffffffffffffe8ffffffff",
            INIT_46 => X"ffffffeaffffffff0000000300000000fffffffaffffffff0000000f00000000",
            INIT_47 => X"ffffffe1ffffffffffffffb7ffffffffffffffecffffffffffffffe4ffffffff",
            INIT_48 => X"0000001000000000ffffffdfffffffff0000001800000000ffffffffffffffff",
            INIT_49 => X"0000002d0000000000000015000000000000003a00000000fffffff3ffffffff",
            INIT_4A => X"0000000700000000fffffff2ffffffff0000001a000000000000003500000000",
            INIT_4B => X"0000000f000000000000000300000000fffffff0ffffffffffffffe1ffffffff",
            INIT_4C => X"0000002200000000ffffffd5ffffffff0000000d000000000000000e00000000",
            INIT_4D => X"00000016000000000000002600000000fffffffcffffffffffffffe9ffffffff",
            INIT_4E => X"0000002e0000000000000004000000000000002a00000000fffffff8ffffffff",
            INIT_4F => X"ffffffe4ffffffffffffffbeffffffffffffffd3ffffffff0000000100000000",
            INIT_50 => X"fffffffbffffffff0000000c00000000fffffff7ffffffff0000001300000000",
            INIT_51 => X"ffffffe0ffffffff00000018000000000000000e000000000000002600000000",
            INIT_52 => X"0000000600000000ffffffc9ffffffff0000001200000000fffffff5ffffffff",
            INIT_53 => X"fffffffdffffffffffffffddffffffffffffffeaffffffff0000000100000000",
            INIT_54 => X"0000000800000000000000150000000000000018000000000000000700000000",
            INIT_55 => X"00000013000000000000000000000000ffffffdcffffffff0000001300000000",
            INIT_56 => X"fffffffaffffffff0000000600000000ffffffffffffffffffffffd6ffffffff",
            INIT_57 => X"0000000c000000000000003800000000fffffff5ffffffff0000001500000000",
            INIT_58 => X"fffffffeffffffff0000001800000000ffffffffffffffff0000000400000000",
            INIT_59 => X"ffffffecffffffffffffffe7fffffffffffffff3fffffffffffffffcffffffff",
            INIT_5A => X"fffffff1ffffffffffffffe4ffffffff00000015000000000000000300000000",
            INIT_5B => X"00000020000000000000000500000000ffffffd1ffffffff0000002a00000000",
            INIT_5C => X"ffffffbdffffffff0000001400000000fffffff2ffffffffffffffc6ffffffff",
            INIT_5D => X"0000000e00000000fffffff4ffffffffffffffd9ffffffffffffffd2ffffffff",
            INIT_5E => X"00000023000000000000000100000000fffffffeffffffffffffffcbffffffff",
            INIT_5F => X"00000000000000000000001a00000000ffffffe9ffffffff0000000200000000",
            INIT_60 => X"fffffff7ffffffffffffffc6ffffffff00000005000000000000000c00000000",
            INIT_61 => X"0000003f00000000fffffffcffffffff0000000a000000000000001200000000",
            INIT_62 => X"0000001600000000ffffffe5ffffffffffffffdcffffffffffffffceffffffff",
            INIT_63 => X"00000009000000000000001d000000000000001a000000000000002e00000000",
            INIT_64 => X"fffffff1ffffffff0000000d00000000fffffff9ffffffff0000000b00000000",
            INIT_65 => X"fffffff0ffffffff0000002a000000000000001b00000000ffffffe3ffffffff",
            INIT_66 => X"0000001c00000000ffffffedffffffff00000013000000000000000000000000",
            INIT_67 => X"0000000a000000000000002d0000000000000031000000000000001900000000",
            INIT_68 => X"ffffffecffffffff00000003000000000000000d000000000000000500000000",
            INIT_69 => X"00000026000000000000001800000000fffffff7ffffffff0000000e00000000",
            INIT_6A => X"fffffffdffffffffffffffffffffffff00000017000000000000000a00000000",
            INIT_6B => X"0000003400000000fffffffcffffffff0000001c000000000000000c00000000",
            INIT_6C => X"00000008000000000000000600000000ffffffe6ffffffff0000001400000000",
            INIT_6D => X"ffffffeefffffffffffffff4ffffffffffffffeffffffffffffffffcffffffff",
            INIT_6E => X"ffffffe9ffffffff0000001e000000000000002d000000000000001600000000",
            INIT_6F => X"ffffffe4ffffffffffffffaafffffffffffffff4ffffffffffffffdbffffffff",
            INIT_70 => X"00000013000000000000000300000000fffffff2ffffffffffffffd3ffffffff",
            INIT_71 => X"0000000500000000ffffffebffffffff0000000d00000000fffffffeffffffff",
            INIT_72 => X"ffffffe6fffffffffffffff6ffffffffffffffe3fffffffffffffff8ffffffff",
            INIT_73 => X"00000035000000000000000800000000fffffff9ffffffff0000001800000000",
            INIT_74 => X"0000001f000000000000001900000000fffffffffffffffffffffff9ffffffff",
            INIT_75 => X"00000010000000000000001700000000fffffff1ffffffff0000001d00000000",
            INIT_76 => X"ffffffedffffffff0000001d00000000ffffffe9ffffffff0000000d00000000",
            INIT_77 => X"fffffff8ffffffffffffffaffffffffffffffff8fffffffffffffff8ffffffff",
            INIT_78 => X"ffffffcfffffffffffffffdaffffffffffffffcdfffffffffffffff0ffffffff",
            INIT_79 => X"00000000000000000000000600000000fffffff8ffffffffffffffbfffffffff",
            INIT_7A => X"00000009000000000000002b000000000000000d00000000ffffffebffffffff",
            INIT_7B => X"0000000300000000ffffffcfffffffffffffffefffffffffffffffffffffffff",
            INIT_7C => X"ffffffdaffffffff0000000000000000ffffffe8fffffffffffffff9ffffffff",
            INIT_7D => X"00000001000000000000000c0000000000000008000000000000001500000000",
            INIT_7E => X"fffffff3ffffffff0000000e000000000000001c00000000ffffffd7ffffffff",
            INIT_7F => X"00000007000000000000000100000000ffffffe1ffffffff0000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE16;


    MEM_IWGHT_LAYER2_INSTANCE17 : if BRAM_NAME = "iwght_layer2_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000fffffff9fffffffffffffffeffffffff0000000c00000000",
            INIT_01 => X"fffffff4ffffffff0000000c00000000ffffffefffffffff0000000d00000000",
            INIT_02 => X"ffffffe4ffffffffffffffe3ffffffff00000002000000000000000e00000000",
            INIT_03 => X"ffffffe1ffffffffffffffedfffffffffffffffeffffffffffffffdcffffffff",
            INIT_04 => X"0000000200000000ffffffeffffffffffffffff0ffffffff0000000a00000000",
            INIT_05 => X"ffffffedfffffffffffffff7ffffffffffffffe8ffffffffffffffdfffffffff",
            INIT_06 => X"0000000400000000fffffff9ffffffffffffffeeffffffff0000000d00000000",
            INIT_07 => X"0000000900000000fffffff9fffffffffffffffdffffffffffffffe9ffffffff",
            INIT_08 => X"ffffffebffffffffffffffd4ffffffffffffffedfffffffffffffff7ffffffff",
            INIT_09 => X"fffffff5fffffffffffffff0fffffffffffffff4ffffffffffffffe4ffffffff",
            INIT_0A => X"0000000300000000fffffffefffffffffffffffaffffffff0000000c00000000",
            INIT_0B => X"fffffff9ffffffff0000000f00000000ffffffedffffffff0000000000000000",
            INIT_0C => X"0000000000000000fffffff4ffffffff00000004000000000000000100000000",
            INIT_0D => X"0000000200000000ffffffedffffffffffffffe9ffffffff0000000100000000",
            INIT_0E => X"ffffffeefffffffffffffffbffffffffffffffe5ffffffff0000000300000000",
            INIT_0F => X"fffffff7fffffffffffffff2ffffffff0000000000000000ffffffebffffffff",
            INIT_10 => X"0000000600000000ffffffebfffffffffffffff0ffffffff0000000200000000",
            INIT_11 => X"fffffffdffffffff0000000700000000ffffffe9fffffffffffffff4ffffffff",
            INIT_12 => X"ffffffebffffffff0000000a000000000000000000000000fffffff6ffffffff",
            INIT_13 => X"0000000800000000ffffffe9ffffffffffffffecfffffffffffffffdffffffff",
            INIT_14 => X"fffffff2ffffffff00000003000000000000000900000000fffffff1ffffffff",
            INIT_15 => X"0000000d00000000ffffffe8fffffffffffffff8ffffffff0000000700000000",
            INIT_16 => X"fffffff5fffffffffffffff5ffffffff0000001600000000ffffffffffffffff",
            INIT_17 => X"fffffff3fffffffffffffff1fffffffffffffffeffffffff0000000d00000000",
            INIT_18 => X"00000000000000000000000400000000ffffffe8ffffffffffffffeaffffffff",
            INIT_19 => X"fffffff8ffffffffffffffe9ffffffff00000013000000000000001200000000",
            INIT_1A => X"0000000500000000ffffffe9fffffffffffffffdffffffffffffffe6ffffffff",
            INIT_1B => X"fffffff6ffffffffffffffeaffffffff0000000f000000000000000600000000",
            INIT_1C => X"fffffffefffffffffffffffeffffffffffffffedffffffffffffffe4ffffffff",
            INIT_1D => X"fffffff1ffffffffffffffe4ffffffff0000000500000000fffffff1ffffffff",
            INIT_1E => X"00000001000000000000000000000000ffffffe8ffffffff0000000200000000",
            INIT_1F => X"00000011000000000000000b000000000000000a00000000fffffff7ffffffff",
            INIT_20 => X"ffffffebfffffffffffffff3ffffffffffffffe9ffffffffffffffeeffffffff",
            INIT_21 => X"ffffffeefffffffffffffffdffffffffffffffe5fffffffffffffff4ffffffff",
            INIT_22 => X"fffffff7ffffffffffffffedffffffff0000000300000000fffffff9ffffffff",
            INIT_23 => X"fffffff8ffffffff00000000000000000000000c00000000fffffff9ffffffff",
            INIT_24 => X"fffffff7fffffffffffffffbffffffff00000010000000000000001600000000",
            INIT_25 => X"000000200000000000000008000000000000000c00000000fffffffeffffffff",
            INIT_26 => X"00000014000000000000001900000000fffffffdffffffff0000000000000000",
            INIT_27 => X"0000000100000000fffffffdffffffff00000000000000000000001100000000",
            INIT_28 => X"fffffff5ffffffff00000005000000000000000400000000fffffff6ffffffff",
            INIT_29 => X"fffffffafffffffffffffff9fffffffffffffffdffffffff0000001100000000",
            INIT_2A => X"ffffffe8ffffffff00000000000000000000000200000000fffffff6ffffffff",
            INIT_2B => X"ffffffe6fffffffffffffff1ffffffffffffffebffffffff0000000000000000",
            INIT_2C => X"0000000200000000fffffff7ffffffffffffffe8ffffffffffffffffffffffff",
            INIT_2D => X"ffffffefffffffffffffffefffffffffffffffecffffffffffffffe0ffffffff",
            INIT_2E => X"ffffffecffffffff0000000000000000fffffff4ffffffffffffffe0ffffffff",
            INIT_2F => X"0000000000000000ffffffe0fffffffffffffff5ffffffffffffffe3ffffffff",
            INIT_30 => X"fffffffdfffffffffffffff2ffffffffffffffebfffffffffffffff7ffffffff",
            INIT_31 => X"ffffffe6ffffffffffffffe0ffffffff00000008000000000000000200000000",
            INIT_32 => X"0000000c00000000fffffff9ffffffff0000000f00000000fffffff7ffffffff",
            INIT_33 => X"0000000b00000000fffffff3ffffffff0000002000000000fffffffdffffffff",
            INIT_34 => X"000000000000000000000009000000000000001200000000fffffffaffffffff",
            INIT_35 => X"0000000800000000ffffffedffffffff00000006000000000000000000000000",
            INIT_36 => X"ffffffe9ffffffffffffffdcfffffffffffffff4fffffffffffffff1ffffffff",
            INIT_37 => X"0000000c000000000000000000000000ffffffe6ffffffffffffffe8ffffffff",
            INIT_38 => X"ffffffd9fffffffffffffffcffffffff0000000b00000000ffffffdbffffffff",
            INIT_39 => X"ffffffebffffffffffffffeafffffffffffffff0ffffffffffffffe6ffffffff",
            INIT_3A => X"fffffffafffffffffffffff3ffffffffffffffedffffffffffffffedffffffff",
            INIT_3B => X"fffffffcffffffff0000000f0000000000000012000000000000001100000000",
            INIT_3C => X"0000000400000000ffffffe6ffffffff0000000e00000000ffffffe5ffffffff",
            INIT_3D => X"ffffffe3fffffffffffffff8fffffffffffffff0ffffffff0000000800000000",
            INIT_3E => X"fffffff0fffffffffffffffefffffffffffffff8fffffffffffffffaffffffff",
            INIT_3F => X"fffffff7fffffffffffffff4ffffffff0000000200000000ffffffe8ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffecffffffff00000003000000000000000100000000fffffffaffffffff",
            INIT_41 => X"fffffff1ffffffff0000000000000000fffffff6fffffffffffffff5ffffffff",
            INIT_42 => X"ffffffeaffffffff0000000900000000ffffffffffffffffffffffeaffffffff",
            INIT_43 => X"00000007000000000000000a00000000fffffff0fffffffffffffff1ffffffff",
            INIT_44 => X"fffffffaffffffff0000000800000000ffffffebfffffffffffffff0ffffffff",
            INIT_45 => X"ffffffe3fffffffffffffffefffffffffffffff9fffffffffffffff2ffffffff",
            INIT_46 => X"fffffffcffffffff0000000e00000000fffffff9fffffffffffffffaffffffff",
            INIT_47 => X"ffffffffffffffffffffffe9ffffffffffffffebfffffffffffffff9ffffffff",
            INIT_48 => X"0000000400000000ffffffeeffffffff0000001a000000000000001900000000",
            INIT_49 => X"0000001a0000000000000018000000000000000e000000000000000700000000",
            INIT_4A => X"00000042000000000000003c000000000000001c000000000000000500000000",
            INIT_4B => X"00000057000000000000003a0000000000000062000000000000004a00000000",
            INIT_4C => X"ffffffefffffffff0000000000000000ffffffc6ffffffff0000000600000000",
            INIT_4D => X"ffffffaeffffffffffffffb6ffffffffffffffc0fffffffffffffff7ffffffff",
            INIT_4E => X"ffffffe5ffffffffffffff74ffffffffffffffb8ffffffffffffff83ffffffff",
            INIT_4F => X"fffffff4ffffffffffffffe5ffffffff0000001200000000fffffff5ffffffff",
            INIT_50 => X"00000063000000000000000f000000000000001b000000000000001c00000000",
            INIT_51 => X"ffffffdcfffffffffffffffdffffffff0000000600000000fffffffdffffffff",
            INIT_52 => X"ffffff63ffffffffffffffebffffffffffffffc4ffffffffffffffbcffffffff",
            INIT_53 => X"fffffffaffffffff00000018000000000000001a00000000ffffffbeffffffff",
            INIT_54 => X"0000002a00000000ffffffedffffffffffffffe0ffffffff0000000400000000",
            INIT_55 => X"0000000a00000000fffffff6ffffffff00000054000000000000003400000000",
            INIT_56 => X"000000000000000000000008000000000000001200000000fffffff4ffffffff",
            INIT_57 => X"00000009000000000000000000000000ffffffe5ffffffff0000000000000000",
            INIT_58 => X"fffffff4fffffffffffffffcfffffffffffffffaffffffff0000001100000000",
            INIT_59 => X"00000007000000000000002d0000000000000016000000000000000600000000",
            INIT_5A => X"0000001900000000000000300000000000000014000000000000001600000000",
            INIT_5B => X"00000009000000000000002c0000000000000014000000000000003a00000000",
            INIT_5C => X"ffffffc3fffffffffffffff1ffffffffffffffe5ffffffffffffffbbffffffff",
            INIT_5D => X"0000000700000000ffffffb0ffffffffffffffe0fffffffffffffff5ffffffff",
            INIT_5E => X"00000024000000000000002500000000fffffff1fffffffffffffff5ffffffff",
            INIT_5F => X"ffffffffffffffff0000002a0000000000000047000000000000000200000000",
            INIT_60 => X"fffffffdffffffffffffff6effffffffffffff9effffffff0000002300000000",
            INIT_61 => X"ffffff84ffffffffffffffc9ffffffffffffffb5fffffffffffffff5ffffffff",
            INIT_62 => X"ffffffdfffffffffffffffc1fffffffffffffffeffffffffffffffcbffffffff",
            INIT_63 => X"00000004000000000000000e00000000ffffffeeffffffffffffffddffffffff",
            INIT_64 => X"00000031000000000000001d00000000fffffff9ffffffffffffffedffffffff",
            INIT_65 => X"ffffffdcffffffff00000023000000000000000f000000000000006500000000",
            INIT_66 => X"fffffffdfffffffffffffff9ffffffff0000001f000000000000003100000000",
            INIT_67 => X"ffffffd6ffffffff0000001200000000fffffff9fffffffffffffffbffffffff",
            INIT_68 => X"ffffffa8ffffffffffffffe4fffffffffffffff0ffffffffffffffd7ffffffff",
            INIT_69 => X"fffffffcffffffff00000031000000000000001f000000000000000a00000000",
            INIT_6A => X"ffffffdeffffffff0000001400000000ffffffd6ffffffffffffffe1ffffffff",
            INIT_6B => X"000000220000000000000016000000000000000300000000ffffffe7ffffffff",
            INIT_6C => X"0000002c00000000000000140000000000000049000000000000000a00000000",
            INIT_6D => X"0000000200000000fffffff6ffffffffffffffedffffffff0000000700000000",
            INIT_6E => X"0000000b000000000000000f000000000000002800000000ffffffeaffffffff",
            INIT_6F => X"0000000100000000000000170000000000000021000000000000002200000000",
            INIT_70 => X"ffffffdaffffffff00000002000000000000001500000000fffffffcffffffff",
            INIT_71 => X"ffffffe8ffffffff0000001600000000ffffffe1ffffffff0000000e00000000",
            INIT_72 => X"0000001b00000000fffffffbffffffff0000001800000000fffffff6ffffffff",
            INIT_73 => X"0000000200000000fffffff9ffffffff00000015000000000000000e00000000",
            INIT_74 => X"0000001300000000000000130000000000000009000000000000000200000000",
            INIT_75 => X"ffffffdcfffffffffffffffdfffffffffffffff9ffffffff0000000e00000000",
            INIT_76 => X"fffffff6fffffffffffffff8fffffffffffffff6ffffffffffffffeaffffffff",
            INIT_77 => X"fffffffdffffffff00000000000000000000001d000000000000000100000000",
            INIT_78 => X"fffffff8ffffffff0000000a000000000000000000000000fffffff1ffffffff",
            INIT_79 => X"0000000c00000000ffffffe8ffffffff0000000900000000fffffffbffffffff",
            INIT_7A => X"ffffffeeffffffff0000000f00000000fffffffdffffffff0000000f00000000",
            INIT_7B => X"000000210000000000000000000000000000000900000000fffffff3ffffffff",
            INIT_7C => X"ffffffe6ffffffff0000001e00000000fffffff3ffffffff0000000100000000",
            INIT_7D => X"ffffffc7ffffffffffffffcdffffffffffffffebffffffffffffffe4ffffffff",
            INIT_7E => X"ffffffb8ffffffffffffffffffffffffffffffb8ffffffffffffffe6ffffffff",
            INIT_7F => X"ffffffb5fffffffffffffff5ffffffffffffff9bffffffffffffffd6ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE17;


    MEM_IWGHT_LAYER2_INSTANCE18 : if BRAM_NAME = "iwght_layer2_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000320000000000000024000000000000002f00000000ffffffa2ffffffff",
            INIT_01 => X"0000000c0000000000000007000000000000002a000000000000002000000000",
            INIT_02 => X"fffffff9ffffffff0000002e00000000ffffffe9fffffffffffffff4ffffffff",
            INIT_03 => X"ffffffdefffffffffffffffbfffffffffffffffaffffffffffffffecffffffff",
            INIT_04 => X"fffffff3ffffffff0000000f00000000fffffffffffffffffffffff7ffffffff",
            INIT_05 => X"fffffff8ffffffff0000000e00000000ffffffeafffffffffffffffeffffffff",
            INIT_06 => X"0000000e000000000000000f000000000000000c00000000fffffff0ffffffff",
            INIT_07 => X"ffffffe4ffffffff0000001d00000000ffffffd0fffffffffffffff0ffffffff",
            INIT_08 => X"00000019000000000000003b00000000fffffffafffffffffffffff3ffffffff",
            INIT_09 => X"ffffffd3ffffffffffffffd2ffffffffffffffe0ffffffff0000000e00000000",
            INIT_0A => X"0000001300000000ffffffcfffffffffffffffc0ffffffffffffffbbffffffff",
            INIT_0B => X"0000000f00000000fffffff1ffffffff00000014000000000000000b00000000",
            INIT_0C => X"0000001700000000ffffffe6fffffffffffffff9ffffffff0000000100000000",
            INIT_0D => X"0000000e000000000000001a000000000000000b000000000000000900000000",
            INIT_0E => X"ffffffffffffffff0000000500000000fffffff6ffffffffffffffe5ffffffff",
            INIT_0F => X"0000001b000000000000001a00000000fffffffdfffffffffffffffeffffffff",
            INIT_10 => X"000000040000000000000014000000000000001800000000fffffffcffffffff",
            INIT_11 => X"00000010000000000000000e000000000000000800000000fffffffcffffffff",
            INIT_12 => X"fffffffdffffffff000000210000000000000012000000000000000200000000",
            INIT_13 => X"ffffffefffffffffffffffeffffffffffffffff7ffffffff0000001700000000",
            INIT_14 => X"ffffffedfffffffffffffff9ffffffff0000000c00000000ffffffd0ffffffff",
            INIT_15 => X"ffffffc4ffffffffffffffd2ffffffffffffffeeffffffffffffffccffffffff",
            INIT_16 => X"0000001a00000000ffffffcbffffffffffffffd5ffffffff0000000300000000",
            INIT_17 => X"00000019000000000000002f0000000000000007000000000000000000000000",
            INIT_18 => X"fffffff0ffffffff00000021000000000000003b000000000000002c00000000",
            INIT_19 => X"ffffffe5ffffffffffffffe0ffffffffffffff96fffffffffffffff3ffffffff",
            INIT_1A => X"ffffffeaffffffffffffffd9ffffffffffffffcfffffffffffffff94ffffffff",
            INIT_1B => X"ffffffc4fffffffffffffff2ffffffffffffffcaffffffffffffffe6ffffffff",
            INIT_1C => X"ffffffdffffffffffffffff5ffffffff0000000900000000ffffffe9ffffffff",
            INIT_1D => X"0000000000000000000000160000000000000031000000000000004000000000",
            INIT_1E => X"0000001d00000000ffffffeeffffffff00000009000000000000001300000000",
            INIT_1F => X"ffffffdbffffffffffffffeeffffffffffffffedffffffffffffffe2ffffffff",
            INIT_20 => X"0000001300000000fffffff6ffffffff0000000500000000ffffffd3ffffffff",
            INIT_21 => X"0000001f00000000fffffffcffffffff0000000f000000000000002900000000",
            INIT_22 => X"0000004d000000000000000f0000000000000032000000000000004d00000000",
            INIT_23 => X"fffffffffffffffffffffff9ffffffffffffffeaffffffff0000000500000000",
            INIT_24 => X"fffffff5ffffffffffffffeaffffffff0000000200000000fffffff6ffffffff",
            INIT_25 => X"ffffffe9ffffffffffffffdafffffffffffffff4ffffffff0000000a00000000",
            INIT_26 => X"00000021000000000000002500000000ffffffe3fffffffffffffff6ffffffff",
            INIT_27 => X"ffffffe0ffffffffffffffd7ffffffff0000002400000000ffffffffffffffff",
            INIT_28 => X"0000000000000000ffffffe1ffffffff0000000000000000fffffff5ffffffff",
            INIT_29 => X"0000001d00000000fffffffeffffffffffffffecffffffffffffffebffffffff",
            INIT_2A => X"fffffffefffffffffffffffbfffffffffffffff2ffffffff0000000200000000",
            INIT_2B => X"fffffff3fffffffffffffffbffffffffffffffdffffffffffffffff3ffffffff",
            INIT_2C => X"0000001800000000000000150000000000000029000000000000001600000000",
            INIT_2D => X"ffffffdeffffffffffffffe7ffffffffffffffdeffffffff0000001700000000",
            INIT_2E => X"0000002200000000000000370000000000000005000000000000001500000000",
            INIT_2F => X"ffffffefffffffff00000011000000000000000100000000fffffff9ffffffff",
            INIT_30 => X"0000000b00000000fffffff6ffffffffffffffe4ffffffffffffffd8ffffffff",
            INIT_31 => X"000000010000000000000008000000000000001200000000fffffff4ffffffff",
            INIT_32 => X"0000001900000000ffffffe9ffffffffffffffe0ffffffffffffffdaffffffff",
            INIT_33 => X"00000012000000000000000d0000000000000001000000000000001900000000",
            INIT_34 => X"0000002e00000000000000260000000000000039000000000000005f00000000",
            INIT_35 => X"0000000600000000fffffff4ffffffff00000026000000000000002800000000",
            INIT_36 => X"00000011000000000000000b0000000000000009000000000000002400000000",
            INIT_37 => X"00000008000000000000002600000000fffffffcffffffff0000001200000000",
            INIT_38 => X"ffffffd0fffffffffffffff6ffffffffffffffe8ffffffffffffffebffffffff",
            INIT_39 => X"fffffff0fffffffffffffff8ffffffffffffffecffffffffffffffb4ffffffff",
            INIT_3A => X"00000000000000000000001900000000ffffffeeffffffffffffffeaffffffff",
            INIT_3B => X"ffffffe1ffffffff0000000e00000000ffffffe5ffffffffffffffeeffffffff",
            INIT_3C => X"0000002e000000000000002200000000ffffffe5fffffffffffffffdffffffff",
            INIT_3D => X"ffffffbfffffffffffffffd8ffffffffffffffe7ffffffffffffffe7ffffffff",
            INIT_3E => X"0000001c00000000ffffffd8ffffffffffffffe8ffffffffffffffe6ffffffff",
            INIT_3F => X"ffffffdeffffffffffffffeffffffffffffffff6ffffffff0000002a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff8ffffffffffffffd8ffffffffffffffdcffffffffffffffc1ffffffff",
            INIT_41 => X"ffffffeafffffffffffffffeffffffff00000042000000000000004000000000",
            INIT_42 => X"0000000400000000ffffffeefffffffffffffff2ffffffffffffffd1ffffffff",
            INIT_43 => X"0000004000000000fffffff7ffffffffffffffeaffffffffffffffd3ffffffff",
            INIT_44 => X"ffffffe5ffffffff00000017000000000000000a000000000000001900000000",
            INIT_45 => X"fffffff6fffffffffffffff6fffffffffffffffefffffffffffffffdffffffff",
            INIT_46 => X"0000004c00000000ffffffbfffffffffffffffdbfffffffffffffffaffffffff",
            INIT_47 => X"0000001e000000000000000000000000ffffffd2fffffffffffffffeffffffff",
            INIT_48 => X"fffffff1ffffffffffffffe5ffffffff00000005000000000000001700000000",
            INIT_49 => X"000000010000000000000008000000000000000d00000000fffffff0ffffffff",
            INIT_4A => X"0000000e00000000ffffffffffffffff0000000a000000000000000500000000",
            INIT_4B => X"0000000500000000000000050000000000000022000000000000001300000000",
            INIT_4C => X"ffffffddfffffffffffffff3fffffffffffffff8ffffffff0000000700000000",
            INIT_4D => X"ffffffeefffffffffffffffaffffffffffffffcdffffffffffffffd8ffffffff",
            INIT_4E => X"0000000400000000fffffff4ffffffffffffffebffffffff0000000900000000",
            INIT_4F => X"0000003000000000000000210000000000000019000000000000000600000000",
            INIT_50 => X"00000001000000000000001f000000000000000f000000000000000800000000",
            INIT_51 => X"fffffff6fffffffffffffffcfffffffffffffff3ffffffffffffffdeffffffff",
            INIT_52 => X"fffffff6ffffffffffffffe6ffffffff0000000d00000000fffffff4ffffffff",
            INIT_53 => X"ffffffeeffffffffffffffdbffffffff0000001200000000ffffffe7ffffffff",
            INIT_54 => X"fffffff4ffffffffffffffe5ffffffffffffffb0ffffffffffffffd4ffffffff",
            INIT_55 => X"ffffffe3ffffffff00000018000000000000000c00000000fffffff4ffffffff",
            INIT_56 => X"0000001100000000fffffffbffffffff00000017000000000000000200000000",
            INIT_57 => X"0000001200000000fffffff9ffffffff00000018000000000000002f00000000",
            INIT_58 => X"ffffffdfffffffffffffffedffffffff0000000100000000fffffff7ffffffff",
            INIT_59 => X"ffffffe8ffffffffffffffe3ffffffff0000000a00000000fffffff6ffffffff",
            INIT_5A => X"ffffffebfffffffffffffff6ffffffff0000001a00000000ffffffe8ffffffff",
            INIT_5B => X"ffffff78ffffffffffffffb9ffffffffffffff9affffffffffffff9bffffffff",
            INIT_5C => X"00000019000000000000001800000000ffffffc6ffffffffffffff87ffffffff",
            INIT_5D => X"fffffffcffffffff0000000600000000ffffffe0ffffffffffffffeaffffffff",
            INIT_5E => X"00000002000000000000000e000000000000001b000000000000002600000000",
            INIT_5F => X"ffffffc1ffffffff0000000a00000000ffffffdcffffffffffffffb3ffffffff",
            INIT_60 => X"ffffffd6ffffffffffffffe9ffffffff0000001100000000ffffffccffffffff",
            INIT_61 => X"00000027000000000000000000000000ffffffeeffffffff0000000a00000000",
            INIT_62 => X"0000002c000000000000002b00000000ffffffefffffffff0000001400000000",
            INIT_63 => X"ffffffffffffffff000000220000000000000029000000000000000a00000000",
            INIT_64 => X"0000000c00000000fffffff6ffffffff00000027000000000000003900000000",
            INIT_65 => X"0000000800000000ffffffeffffffffffffffff6ffffffff0000001700000000",
            INIT_66 => X"ffffffe0fffffffffffffff5fffffffffffffff9ffffffffffffffebffffffff",
            INIT_67 => X"0000000c00000000fffffff3fffffffffffffff2fffffffffffffffdffffffff",
            INIT_68 => X"0000001b00000000fffffff4ffffffff00000001000000000000002000000000",
            INIT_69 => X"00000019000000000000001a0000000000000026000000000000003800000000",
            INIT_6A => X"ffffffb8fffffffffffffff6ffffffffffffffe4fffffffffffffff4ffffffff",
            INIT_6B => X"fffffff0ffffffffffffffcaffffffffffffffeeffffffffffffffc9ffffffff",
            INIT_6C => X"0000000500000000000000110000000000000001000000000000000300000000",
            INIT_6D => X"0000000c00000000ffffffe9fffffffffffffff7ffffffffffffffffffffffff",
            INIT_6E => X"00000009000000000000000100000000fffffffefffffffffffffff9ffffffff",
            INIT_6F => X"ffffffc7ffffffffffffffc3ffffffffffffffdcfffffffffffffffdffffffff",
            INIT_70 => X"0000000a000000000000000e00000000fffffff1ffffffffffffffdaffffffff",
            INIT_71 => X"ffffffd0ffffffff0000001e00000000ffffffedffffffff0000000b00000000",
            INIT_72 => X"ffffffe3ffffffffffffffd8ffffffff0000002f00000000ffffffddffffffff",
            INIT_73 => X"0000000500000000ffffffe1fffffffffffffff4fffffffffffffffaffffffff",
            INIT_74 => X"00000010000000000000002000000000fffffff1fffffffffffffffdffffffff",
            INIT_75 => X"000000280000000000000022000000000000000d00000000ffffffc8ffffffff",
            INIT_76 => X"0000000600000000fffffffffffffffffffffffaffffffffffffffe3ffffffff",
            INIT_77 => X"fffffff2ffffffff000000030000000000000002000000000000000300000000",
            INIT_78 => X"fffffff2ffffffff0000000e000000000000003f00000000ffffffe9ffffffff",
            INIT_79 => X"fffffff0fffffffffffffff0ffffffff00000012000000000000001300000000",
            INIT_7A => X"0000001b000000000000000f000000000000000d00000000fffffff5ffffffff",
            INIT_7B => X"fffffffaffffffff0000000e000000000000001900000000fffffff1ffffffff",
            INIT_7C => X"ffffffb4ffffffffffffffc4ffffffffffffffe2ffffffffffffffccffffffff",
            INIT_7D => X"ffffffb0ffffffff0000000400000000ffffffbbffffffffffffffe0ffffffff",
            INIT_7E => X"000000110000000000000014000000000000001e00000000ffffffc2ffffffff",
            INIT_7F => X"0000000200000000ffffffe4ffffffff00000011000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE18;


    MEM_IWGHT_LAYER2_INSTANCE19 : if BRAM_NAME = "iwght_layer2_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004a000000000000002c00000000ffffffcefffffffffffffffaffffffff",
            INIT_01 => X"ffffffedffffffffffffffdaffffffff00000007000000000000004c00000000",
            INIT_02 => X"fffffffbffffffffffffffdaffffffffffffffbbfffffffffffffffcffffffff",
            INIT_03 => X"0000000d0000000000000017000000000000000000000000ffffffe7ffffffff",
            INIT_04 => X"000000190000000000000023000000000000000f000000000000000b00000000",
            INIT_05 => X"00000022000000000000001c00000000fffffff8ffffffff0000000400000000",
            INIT_06 => X"fffffff2fffffffffffffff9fffffffffffffff8ffffffff0000000400000000",
            INIT_07 => X"fffffff9fffffffffffffff7ffffffff00000007000000000000000000000000",
            INIT_08 => X"000000070000000000000000000000000000000b000000000000001900000000",
            INIT_09 => X"fffffff7ffffffff00000000000000000000001a000000000000000800000000",
            INIT_0A => X"fffffff5ffffffff00000007000000000000000500000000fffffffcffffffff",
            INIT_0B => X"0000002000000000ffffffefffffffff00000022000000000000000000000000",
            INIT_0C => X"0000000d000000000000001300000000fffffffdfffffffffffffff7ffffffff",
            INIT_0D => X"0000000b00000000000000190000000000000020000000000000000800000000",
            INIT_0E => X"ffffffebffffffffffffffd9ffffffff0000001000000000fffffff3ffffffff",
            INIT_0F => X"0000002100000000fffffff1ffffffff00000030000000000000000300000000",
            INIT_10 => X"0000000d00000000000000110000000000000000000000000000004200000000",
            INIT_11 => X"0000001700000000ffffffe1fffffffffffffff5ffffffffffffffdbffffffff",
            INIT_12 => X"0000002600000000fffffffaffffffff0000000e00000000ffffffedffffffff",
            INIT_13 => X"ffffffefffffffff0000000e0000000000000000000000000000002900000000",
            INIT_14 => X"fffffffcffffffffffffffe3fffffffffffffff6ffffffff0000002600000000",
            INIT_15 => X"0000000000000000ffffffe8ffffffffffffffccffffffffffffffebffffffff",
            INIT_16 => X"0000000500000000000000210000000000000006000000000000000900000000",
            INIT_17 => X"0000001900000000ffffffe6ffffffff00000000000000000000001d00000000",
            INIT_18 => X"0000003a00000000fffffffbffffffffffffffd9ffffffff0000000800000000",
            INIT_19 => X"ffffffccffffffff0000002100000000fffffff4ffffffffffffffe8ffffffff",
            INIT_1A => X"0000002900000000ffffffffffffffff0000002c000000000000000700000000",
            INIT_1B => X"ffffffe6ffffffffffffffffffffffffffffffecfffffffffffffffbffffffff",
            INIT_1C => X"0000000e00000000ffffffecffffffff0000000e000000000000000100000000",
            INIT_1D => X"00000021000000000000000c0000000000000006000000000000001400000000",
            INIT_1E => X"0000001b000000000000000e0000000000000032000000000000001b00000000",
            INIT_1F => X"ffffffceffffffff000000230000000000000010000000000000000200000000",
            INIT_20 => X"fffffffcffffffffffffffe3fffffffffffffff5ffffffffffffffedffffffff",
            INIT_21 => X"fffffffaffffffff00000001000000000000000e000000000000001000000000",
            INIT_22 => X"0000000e000000000000001500000000fffffffdfffffffffffffff0ffffffff",
            INIT_23 => X"0000000e00000000000000320000000000000016000000000000003600000000",
            INIT_24 => X"00000011000000000000002f0000000000000020000000000000002000000000",
            INIT_25 => X"0000000c000000000000001100000000ffffffddffffffff0000001a00000000",
            INIT_26 => X"ffffffe8ffffffff00000042000000000000001c000000000000001500000000",
            INIT_27 => X"0000003b00000000000000180000000000000007000000000000001500000000",
            INIT_28 => X"0000000b00000000ffffffeaffffffffffffffd6ffffffff0000000700000000",
            INIT_29 => X"00000010000000000000001500000000ffffffdaffffffff0000001c00000000",
            INIT_2A => X"0000000800000000ffffffe8ffffffff00000029000000000000000f00000000",
            INIT_2B => X"ffffffebffffffffffffffd8ffffffffffffffcdffffffff0000002700000000",
            INIT_2C => X"ffffffb8ffffffffffffffeeffffffffffffffe4ffffffffffffffe7ffffffff",
            INIT_2D => X"fffffff9ffffffffffffffeaffffffffffffffe7ffffffffffffffc7ffffffff",
            INIT_2E => X"ffffffb5ffffffffffffffb9ffffffffffffffafffffffffffffffd5ffffffff",
            INIT_2F => X"0000002200000000fffffffcfffffffffffffff2fffffffffffffffeffffffff",
            INIT_30 => X"fffffff1ffffffff0000001200000000fffffff5ffffffff0000003a00000000",
            INIT_31 => X"0000001500000000fffffff9ffffffff0000001100000000ffffffe5ffffffff",
            INIT_32 => X"ffffffe8ffffffff0000000200000000fffffffbffffffffffffffecffffffff",
            INIT_33 => X"0000000100000000ffffffc8ffffffff00000011000000000000000900000000",
            INIT_34 => X"00000018000000000000000b00000000ffffffeeffffffff0000003e00000000",
            INIT_35 => X"00000006000000000000000200000000fffffff7ffffffff0000000900000000",
            INIT_36 => X"0000000d00000000ffffffe9ffffffff0000000d000000000000000b00000000",
            INIT_37 => X"0000001a00000000fffffffeffffffff00000009000000000000001a00000000",
            INIT_38 => X"ffffffe5ffffffff000000130000000000000029000000000000000300000000",
            INIT_39 => X"fffffff1ffffffffffffffb7ffffffff0000000e00000000ffffffa8ffffffff",
            INIT_3A => X"ffffffcfffffffffffffffe2ffffffffffffffc0ffffffffffffffe7ffffffff",
            INIT_3B => X"ffffffc9fffffffffffffffbfffffffffffffff4ffffffffffffffeaffffffff",
            INIT_3C => X"ffffffc2fffffffffffffffaffffffff0000000f00000000fffffff2ffffffff",
            INIT_3D => X"ffffffd5fffffffffffffffaffffffffffffffdeffffffffffffffbbffffffff",
            INIT_3E => X"fffffffdffffffffffffffe3ffffffffffffffccffffffffffffffd8ffffffff",
            INIT_3F => X"ffffffbfffffffffffffffdfffffffffffffffecffffffff0000001200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffbffffffffffffff9affffffffffffffc0fffffffffffffff0ffffffff",
            INIT_41 => X"fffffff0ffffffffffffffc9ffffffffffffffa5ffffffffffffff97ffffffff",
            INIT_42 => X"ffffffeaffffffffffffffeaffffffff0000001e000000000000000000000000",
            INIT_43 => X"ffffffbfffffffffffffffd7fffffffffffffff2ffffffff0000000100000000",
            INIT_44 => X"ffffffbbffffffffffffffe7ffffffffffffffeaffffffffffffffccffffffff",
            INIT_45 => X"ffffff82ffffffffffffffcaffffffffffffffa9ffffffffffffffabffffffff",
            INIT_46 => X"0000001a000000000000000000000000ffffffd1ffffffffffffffd7ffffffff",
            INIT_47 => X"ffffffd9ffffffffffffffe1ffffffffffffffabfffffffffffffff0ffffffff",
            INIT_48 => X"fffffffcffffffffffffffffffffffffffffffe6fffffffffffffffdffffffff",
            INIT_49 => X"00000000000000000000000000000000ffffffe1ffffffff0000002400000000",
            INIT_4A => X"0000000e000000000000001c00000000ffffffcfffffffffffffffddffffffff",
            INIT_4B => X"000000140000000000000002000000000000001b000000000000001800000000",
            INIT_4C => X"ffffffd7ffffffffffffffdfffffffff00000013000000000000000300000000",
            INIT_4D => X"0000001700000000000000300000000000000045000000000000000f00000000",
            INIT_4E => X"ffffffe3fffffffffffffffaffffffff0000003e000000000000003600000000",
            INIT_4F => X"000000330000000000000033000000000000000e00000000ffffffedffffffff",
            INIT_50 => X"ffffffe0ffffffff000000140000000000000035000000000000001100000000",
            INIT_51 => X"ffffffefffffffffffffffe2ffffffffffffffedffffffffffffffedffffffff",
            INIT_52 => X"00000007000000000000000b00000000ffffffe9ffffffff0000000200000000",
            INIT_53 => X"ffffffefffffffff0000000e000000000000000100000000ffffffebffffffff",
            INIT_54 => X"ffffffe3ffffffffffffffe2ffffffff0000001b00000000fffffff7ffffffff",
            INIT_55 => X"ffffffe5ffffffffffffffcaffffffffffffffddffffffff0000001500000000",
            INIT_56 => X"0000002400000000ffffffecffffffff0000001d000000000000000800000000",
            INIT_57 => X"0000001a00000000000000310000000000000016000000000000003200000000",
            INIT_58 => X"ffffffe7ffffffff00000013000000000000002b00000000fffffff3ffffffff",
            INIT_59 => X"0000000500000000000000060000000000000016000000000000000000000000",
            INIT_5A => X"00000015000000000000000000000000fffffff0fffffffffffffff3ffffffff",
            INIT_5B => X"0000004300000000000000210000000000000000000000000000003900000000",
            INIT_5C => X"ffffffdbffffffff00000038000000000000001a00000000fffffff8ffffffff",
            INIT_5D => X"ffffffb0ffffffffffffffeeffffffffffffffdeffffffffffffffd2ffffffff",
            INIT_5E => X"ffffff9effffffffffffffb6ffffffff0000002f00000000ffffffd1ffffffff",
            INIT_5F => X"00000030000000000000002c0000000000000000000000000000000800000000",
            INIT_60 => X"0000000d000000000000000c0000000000000031000000000000000400000000",
            INIT_61 => X"ffffffc3ffffffffffffff95ffffffffffffff97ffffffff0000001100000000",
            INIT_62 => X"0000002200000000ffffff76ffffffffffffff90ffffffffffffffc5ffffffff",
            INIT_63 => X"00000015000000000000000800000000ffffffcdffffffff0000000400000000",
            INIT_64 => X"0000000d00000000000000310000000000000015000000000000003200000000",
            INIT_65 => X"fffffff4ffffffffffffffcfffffffffffffffe3ffffffff0000000400000000",
            INIT_66 => X"0000002b00000000000000110000000000000044000000000000000c00000000",
            INIT_67 => X"0000001f00000000fffffff4fffffffffffffffbffffffff0000001a00000000",
            INIT_68 => X"ffffffe1ffffffffffffffefffffffff00000013000000000000001300000000",
            INIT_69 => X"00000000000000000000000100000000fffffff3ffffffff0000000200000000",
            INIT_6A => X"ffffff9affffffffffffffceffffffffffffffe6ffffffff0000000000000000",
            INIT_6B => X"ffffffeaffffffffffffffa7ffffffffffffffbcffffffffffffffd0ffffffff",
            INIT_6C => X"ffffffeaffffffff0000000400000000fffffff6ffffffffffffffe0ffffffff",
            INIT_6D => X"0000000300000000ffffffdeffffffff0000000b00000000ffffffcaffffffff",
            INIT_6E => X"ffffffeeffffffffffffffe1fffffffffffffffeffffffff0000000200000000",
            INIT_6F => X"0000001100000000ffffffe4fffffffffffffff1fffffffffffffffbffffffff",
            INIT_70 => X"fffffffaffffffff0000000500000000ffffffe2ffffffff0000001600000000",
            INIT_71 => X"0000000400000000ffffffc9ffffffffffffffd8fffffffffffffff1ffffffff",
            INIT_72 => X"ffffffdaffffffffffffffd6ffffffffffffffe5fffffffffffffff0ffffffff",
            INIT_73 => X"0000002e000000000000002d000000000000000f00000000ffffffe5ffffffff",
            INIT_74 => X"000000250000000000000020000000000000001c000000000000001f00000000",
            INIT_75 => X"ffffffddffffffff0000001400000000fffffffdfffffffffffffffcffffffff",
            INIT_76 => X"0000000500000000ffffffecffffffff0000000e00000000ffffffcaffffffff",
            INIT_77 => X"fffffffbffffffff0000001400000000fffffffbffffffff0000002200000000",
            INIT_78 => X"0000000f000000000000002900000000ffffffdfffffffff0000001700000000",
            INIT_79 => X"ffffffe3ffffffff0000000e0000000000000012000000000000001800000000",
            INIT_7A => X"0000000000000000fffffffaffffffffffffffe4ffffffff0000001900000000",
            INIT_7B => X"ffffffeeffffffffffffffe9fffffffffffffff7ffffffffffffffdfffffffff",
            INIT_7C => X"fffffff3ffffffffffffffe0ffffffffffffffedffffffff0000000c00000000",
            INIT_7D => X"00000011000000000000000200000000ffffffffffffffffffffffedffffffff",
            INIT_7E => X"ffffffe9ffffffff000000130000000000000015000000000000002400000000",
            INIT_7F => X"fffffff9fffffffffffffff1ffffffff0000001c00000000ffffffcbffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE19;


    MEM_IWGHT_LAYER2_INSTANCE20 : if BRAM_NAME = "iwght_layer2_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000005000000000000001a000000000000000c000000000000000400000000",
            INIT_01 => X"0000001c0000000000000017000000000000003700000000fffffff9ffffffff",
            INIT_02 => X"00000004000000000000000a000000000000001f000000000000002600000000",
            INIT_03 => X"fffffff8ffffffff0000002e000000000000000900000000ffffffe3ffffffff",
            INIT_04 => X"0000000400000000fffffff9ffffffff0000001e000000000000000100000000",
            INIT_05 => X"ffffffccfffffffffffffff1fffffffffffffffeffffffff0000000900000000",
            INIT_06 => X"ffffffd6ffffffffffffffdfffffffffffffffc7ffffffffffffffecffffffff",
            INIT_07 => X"0000002a000000000000001900000000fffffff2ffffffff0000000a00000000",
            INIT_08 => X"00000008000000000000001c0000000000000021000000000000002100000000",
            INIT_09 => X"ffffffeaffffffffffffffdaffffffff00000007000000000000002400000000",
            INIT_0A => X"ffffffe6ffffffffffffffdaffffffff0000001000000000ffffffd6ffffffff",
            INIT_0B => X"0000000a00000000fffffffdffffffffffffffe1ffffffff0000000000000000",
            INIT_0C => X"fffffffbffffffffffffffd7ffffffffffffffcaffffffffffffffe6ffffffff",
            INIT_0D => X"fffffff3ffffffffffffffe1ffffffffffffffc4ffffffffffffffd6ffffffff",
            INIT_0E => X"0000000d00000000ffffffeafffffffffffffffeffffffffffffffdaffffffff",
            INIT_0F => X"0000000d00000000000000130000000000000000000000000000001900000000",
            INIT_10 => X"0000000400000000000000330000000000000017000000000000003800000000",
            INIT_11 => X"00000004000000000000000400000000ffffffd1ffffffff0000002c00000000",
            INIT_12 => X"fffffffbffffffff00000047000000000000000000000000fffffff4ffffffff",
            INIT_13 => X"0000001c00000000000000110000000000000012000000000000001d00000000",
            INIT_14 => X"ffffffecfffffffffffffffcffffffff00000029000000000000000600000000",
            INIT_15 => X"0000001100000000000000040000000000000011000000000000001e00000000",
            INIT_16 => X"00000019000000000000001100000000fffffff7ffffffff0000001200000000",
            INIT_17 => X"000000150000000000000016000000000000000e000000000000000d00000000",
            INIT_18 => X"fffffffdffffffff0000000b000000000000000400000000fffffff5ffffffff",
            INIT_19 => X"fffffff1fffffffffffffff7ffffffff0000000900000000fffffff2ffffffff",
            INIT_1A => X"0000001a0000000000000008000000000000000c00000000fffffff0ffffffff",
            INIT_1B => X"000000090000000000000015000000000000001b000000000000001100000000",
            INIT_1C => X"fffffff5ffffffff0000001800000000fffffff1ffffffff0000001e00000000",
            INIT_1D => X"ffffffdbffffffffffffffe5ffffffff0000002100000000fffffffdffffffff",
            INIT_1E => X"0000002d0000000000000047000000000000003d000000000000006300000000",
            INIT_1F => X"00000022000000000000005b0000000000000069000000000000004c00000000",
            INIT_20 => X"ffffffbdffffffffffffffd9fffffffffffffffaffffffff0000001100000000",
            INIT_21 => X"0000000400000000ffffffdcffffffffffffffbfffffffffffffffeeffffffff",
            INIT_22 => X"0000000500000000fffffff6fffffffffffffff9ffffffffffffffdeffffffff",
            INIT_23 => X"0000001c0000000000000016000000000000000500000000fffffff3ffffffff",
            INIT_24 => X"000000010000000000000024000000000000003c000000000000001400000000",
            INIT_25 => X"fffffff9ffffffff0000002200000000fffffffefffffffffffffffbffffffff",
            INIT_26 => X"0000000c0000000000000028000000000000002f00000000fffffffaffffffff",
            INIT_27 => X"000000020000000000000014000000000000000b000000000000001100000000",
            INIT_28 => X"fffffff2ffffffffffffffdeffffffff0000001a000000000000000100000000",
            INIT_29 => X"fffffff9ffffffff000000000000000000000007000000000000002300000000",
            INIT_2A => X"0000004100000000000000150000000000000026000000000000001100000000",
            INIT_2B => X"0000001400000000000000140000000000000003000000000000002100000000",
            INIT_2C => X"ffffffeaffffffff0000000e0000000000000012000000000000001100000000",
            INIT_2D => X"ffffffeffffffffffffffffafffffffffffffff0ffffffff0000000d00000000",
            INIT_2E => X"ffffffedffffffff00000000000000000000000600000000fffffff5ffffffff",
            INIT_2F => X"0000001a00000000000000270000000000000006000000000000000f00000000",
            INIT_30 => X"fffffff3fffffffffffffff0ffffffff0000000800000000ffffffffffffffff",
            INIT_31 => X"00000016000000000000001400000000fffffff3ffffffff0000000e00000000",
            INIT_32 => X"ffffffd7fffffffffffffffeffffffff0000000800000000fffffffeffffffff",
            INIT_33 => X"ffffffddffffffffffffffebfffffffffffffff6ffffffffffffffceffffffff",
            INIT_34 => X"0000004b00000000ffffffffffffffffffffffc0ffffffffffffffc0ffffffff",
            INIT_35 => X"0000000c00000000000000470000000000000034000000000000001900000000",
            INIT_36 => X"fffffffcffffffff000000000000000000000007000000000000002000000000",
            INIT_37 => X"ffffffdaffffffff00000009000000000000001f00000000fffffff1ffffffff",
            INIT_38 => X"000000260000000000000005000000000000002d00000000ffffffeaffffffff",
            INIT_39 => X"fffffffeffffffff0000003d0000000000000024000000000000002c00000000",
            INIT_3A => X"00000005000000000000004a00000000ffffffe6fffffffffffffff5ffffffff",
            INIT_3B => X"000000060000000000000000000000000000000c000000000000003c00000000",
            INIT_3C => X"0000000000000000ffffffeaffffffff0000001d000000000000003200000000",
            INIT_3D => X"ffffffe7ffffffffffffffd4ffffffffffffffd1fffffffffffffffbffffffff",
            INIT_3E => X"00000016000000000000000200000000ffffffd8fffffffffffffff3ffffffff",
            INIT_3F => X"ffffffe8fffffffffffffffdfffffffffffffff6ffffffffffffffc3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffd1fffffffffffffffaffffffff0000000b000000000000001100000000",
            INIT_41 => X"0000001f000000000000000d000000000000000200000000ffffffecffffffff",
            INIT_42 => X"00000001000000000000000a0000000000000014000000000000001b00000000",
            INIT_43 => X"fffffffaffffffff000000020000000000000024000000000000000000000000",
            INIT_44 => X"ffffffe4fffffffffffffff5ffffffffffffffdfffffffff0000001a00000000",
            INIT_45 => X"ffffffd9fffffffffffffffeffffffff00000037000000000000001f00000000",
            INIT_46 => X"ffffffecffffffff00000011000000000000000a00000000fffffffaffffffff",
            INIT_47 => X"0000001e000000000000000600000000fffffffbfffffffffffffff7ffffffff",
            INIT_48 => X"ffffffdfffffffff0000001f000000000000001c00000000fffffff4ffffffff",
            INIT_49 => X"ffffffcfffffffff00000017000000000000000700000000fffffff2ffffffff",
            INIT_4A => X"ffffffe1ffffffffffffffc9ffffffffffffffe2ffffffff0000000f00000000",
            INIT_4B => X"ffffffceffffffffffffffddffffffffffffffc4ffffffffffffffa2ffffffff",
            INIT_4C => X"ffffffdffffffffffffffffaffffffffffffffc7ffffffffffffffcaffffffff",
            INIT_4D => X"fffffff0ffffffff00000004000000000000000200000000ffffffd5ffffffff",
            INIT_4E => X"ffffffd8fffffffffffffff2ffffffffffffffe6ffffffff0000001200000000",
            INIT_4F => X"ffffffd7ffffffff0000000000000000ffffffd6fffffffffffffff0ffffffff",
            INIT_50 => X"ffffffecfffffffffffffffbffffffffffffffe9ffffffffffffffffffffffff",
            INIT_51 => X"ffffff91ffffffffffffffeaffffffffffffffe8fffffffffffffff9ffffffff",
            INIT_52 => X"ffffffc6ffffffffffffffbfffffffffffffffd7ffffffffffffff95ffffffff",
            INIT_53 => X"ffffffffffffffff00000003000000000000001200000000ffffffdaffffffff",
            INIT_54 => X"ffffffe2ffffffffffffff9dffffffffffffffb9ffffffffffffffddffffffff",
            INIT_55 => X"0000000300000000000000160000000000000016000000000000000e00000000",
            INIT_56 => X"ffffffcdffffffffffffffedffffffffffffffbcffffffffffffffdfffffffff",
            INIT_57 => X"ffffffe5ffffffff0000001300000000ffffffdffffffffffffffff2ffffffff",
            INIT_58 => X"0000001b0000000000000026000000000000000c000000000000001500000000",
            INIT_59 => X"0000000c00000000ffffffffffffffff00000037000000000000002a00000000",
            INIT_5A => X"ffffffecffffffff0000002900000000fffffff8ffffffff0000002400000000",
            INIT_5B => X"fffffffaffffffffffffffffffffffffffffffffffffffffffffffe5ffffffff",
            INIT_5C => X"0000001700000000fffffff2fffffffffffffff3fffffffffffffffcffffffff",
            INIT_5D => X"0000000d00000000fffffff2ffffffff00000005000000000000000900000000",
            INIT_5E => X"00000001000000000000000f000000000000000900000000fffffffaffffffff",
            INIT_5F => X"fffffffeffffffffffffffe8ffffffffffffffe9ffffffff0000001d00000000",
            INIT_60 => X"ffffffefffffffff0000000c000000000000000a000000000000000700000000",
            INIT_61 => X"ffffffc4ffffffffffffffa5fffffffffffffffeffffffffffffffebffffffff",
            INIT_62 => X"ffffffd9ffffffffffffffdffffffffffffffff3ffffffffffffffdcffffffff",
            INIT_63 => X"fffffff2fffffffffffffffcffffffffffffffe8fffffffffffffffbffffffff",
            INIT_64 => X"00000011000000000000001600000000ffffffffffffffffffffffe9ffffffff",
            INIT_65 => X"000000290000000000000007000000000000000c000000000000001900000000",
            INIT_66 => X"ffffffc6ffffffffffffffffffffffff0000001c00000000ffffffe2ffffffff",
            INIT_67 => X"0000002400000000ffffffdbffffffffffffffd2ffffffffffffffeaffffffff",
            INIT_68 => X"0000000000000000000000030000000000000029000000000000001000000000",
            INIT_69 => X"0000002000000000000000330000000000000025000000000000001400000000",
            INIT_6A => X"fffffff7ffffffffffffffffffffffff0000001e000000000000003100000000",
            INIT_6B => X"ffffffddfffffffffffffffdffffffff0000001800000000ffffffecffffffff",
            INIT_6C => X"ffffffb9ffffffff0000000100000000ffffffe9fffffffffffffffdffffffff",
            INIT_6D => X"ffffffe7ffffffffffffffc6ffffffffffffffd1fffffffffffffff4ffffffff",
            INIT_6E => X"ffffffdcffffffff0000001700000000ffffffb2fffffffffffffff1ffffffff",
            INIT_6F => X"000000110000000000000025000000000000002e000000000000002700000000",
            INIT_70 => X"0000001c000000000000002f00000000fffffff9fffffffffffffff2ffffffff",
            INIT_71 => X"ffffffb1ffffffffffffffd2ffffffffffffffe9ffffffff0000000400000000",
            INIT_72 => X"ffffffe4ffffffff0000001300000000ffffffefffffffffffffffe8ffffffff",
            INIT_73 => X"0000000300000000000000110000000000000017000000000000000b00000000",
            INIT_74 => X"0000001b00000000000000020000000000000019000000000000000500000000",
            INIT_75 => X"0000000c00000000000000150000000000000019000000000000000d00000000",
            INIT_76 => X"ffffffaafffffffffffffff3ffffffffffffffe2ffffffffffffffeeffffffff",
            INIT_77 => X"ffffffeefffffffffffffff1ffffffffffffffdcffffffffffffffcdffffffff",
            INIT_78 => X"0000000200000000fffffff4fffffffffffffff1fffffffffffffff5ffffffff",
            INIT_79 => X"0000001000000000fffffffcfffffffffffffff7ffffffff0000000500000000",
            INIT_7A => X"ffffffe7ffffffff00000001000000000000000f000000000000000d00000000",
            INIT_7B => X"ffffffe1ffffffffffffffe6ffffffff0000000900000000ffffffe9ffffffff",
            INIT_7C => X"0000001a000000000000000f00000000ffffffe5fffffffffffffff2ffffffff",
            INIT_7D => X"0000002a000000000000002d0000000000000005000000000000003600000000",
            INIT_7E => X"0000005f00000000000000160000000000000036000000000000001100000000",
            INIT_7F => X"00000015000000000000001700000000ffffffe5ffffffff0000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE20;


    MEM_IWGHT_LAYER2_INSTANCE21 : if BRAM_NAME = "iwght_layer2_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000014000000000000000d00000000ffffffe6ffffffffffffffe8ffffffff",
            INIT_01 => X"0000001e00000000000000050000000000000025000000000000002b00000000",
            INIT_02 => X"fffffff9ffffffff0000000100000000fffffff4ffffffff0000003100000000",
            INIT_03 => X"0000000200000000ffffffacffffffffffffffb1ffffffff0000001000000000",
            INIT_04 => X"ffffffc9ffffffff0000001a00000000ffffffe8ffffffffffffffd0ffffffff",
            INIT_05 => X"ffffffcbffffffffffffffeafffffffffffffff6ffffffffffffffe7ffffffff",
            INIT_06 => X"0000000b00000000ffffffeaffffffffffffffe4ffffffffffffffd1ffffffff",
            INIT_07 => X"fffffff5ffffffff00000027000000000000000c000000000000002500000000",
            INIT_08 => X"0000000900000000000000360000000000000000000000000000001900000000",
            INIT_09 => X"0000000d000000000000000a000000000000002c000000000000003a00000000",
            INIT_0A => X"ffffffa9ffffffffffffffd6ffffffff0000000800000000ffffffdeffffffff",
            INIT_0B => X"fffffff6ffffffffffffffcdffffffffffffffeffffffffffffffff9ffffffff",
            INIT_0C => X"ffffffdeffffffffffffffccffffffffffffffbefffffffffffffff4ffffffff",
            INIT_0D => X"0000000800000000ffffffdbffffffffffffffeaffffffffffffffeeffffffff",
            INIT_0E => X"ffffffe3ffffffffffffffeeffffffffffffffe6fffffffffffffff1ffffffff",
            INIT_0F => X"0000001300000000fffffffaffffffffffffffd6ffffffff0000001100000000",
            INIT_10 => X"fffffff4fffffffffffffff7ffffffffffffffdffffffffffffffff6ffffffff",
            INIT_11 => X"ffffffbbfffffffffffffff2ffffffff0000001d00000000fffffff5ffffffff",
            INIT_12 => X"ffffffd0ffffffffffffffd3ffffffffffffffcafffffffffffffffbffffffff",
            INIT_13 => X"fffffff7fffffffffffffff3ffffffffffffffeaffffffffffffffd1ffffffff",
            INIT_14 => X"0000001100000000fffffffaffffffff00000003000000000000001600000000",
            INIT_15 => X"ffffffebffffffff00000011000000000000001c000000000000002000000000",
            INIT_16 => X"0000002f000000000000000d000000000000001f000000000000005900000000",
            INIT_17 => X"ffffffdbffffffffffffffaafffffffffffffff2fffffffffffffffbffffffff",
            INIT_18 => X"0000000200000000fffffffdffffffffffffffc7ffffffffffffffe6ffffffff",
            INIT_19 => X"fffffff7ffffffffffffffdfffffffffffffffdcffffffff0000000200000000",
            INIT_1A => X"0000000700000000fffffff1ffffffff00000000000000000000000a00000000",
            INIT_1B => X"0000000200000000000000230000000000000001000000000000001100000000",
            INIT_1C => X"00000048000000000000000300000000fffffff5ffffffff0000004200000000",
            INIT_1D => X"ffffffbfffffffff0000001600000000ffffffc5fffffffffffffff9ffffffff",
            INIT_1E => X"fffffff2ffffffffffffffe4ffffffffffffffd6fffffffffffffffaffffffff",
            INIT_1F => X"00000007000000000000001000000000ffffffecffffffffffffffefffffffff",
            INIT_20 => X"ffffffc0ffffffffffffffdfffffffff00000024000000000000001100000000",
            INIT_21 => X"ffffffc7ffffffffffffffebfffffffffffffff5ffffffffffffffd1ffffffff",
            INIT_22 => X"ffffffedffffffff0000000b00000000ffffffe3ffffffff0000001100000000",
            INIT_23 => X"0000000200000000fffffff0ffffffff00000015000000000000000c00000000",
            INIT_24 => X"0000002100000000000000020000000000000001000000000000001000000000",
            INIT_25 => X"fffffffeffffffff0000000300000000fffffffefffffffffffffff1ffffffff",
            INIT_26 => X"0000000700000000fffffffdfffffffffffffff9fffffffffffffff9ffffffff",
            INIT_27 => X"00000004000000000000002300000000fffffffbffffffffffffffe6ffffffff",
            INIT_28 => X"fffffffcffffffff0000001b000000000000002000000000fffffffeffffffff",
            INIT_29 => X"fffffffbffffffffffffffecffffffffffffffe8ffffffffffffffeeffffffff",
            INIT_2A => X"0000001300000000ffffffe6ffffffffffffffffffffffff0000001300000000",
            INIT_2B => X"ffffffeeffffffff000000360000000000000013000000000000000700000000",
            INIT_2C => X"0000000000000000fffffff2ffffffff0000001800000000ffffffd7ffffffff",
            INIT_2D => X"0000002d000000000000000e000000000000000e00000000fffffff5ffffffff",
            INIT_2E => X"ffffffd4ffffffff0000002c000000000000003400000000fffffff9ffffffff",
            INIT_2F => X"ffffffccffffffffffffffd9ffffffff0000002f000000000000001400000000",
            INIT_30 => X"000000120000000000000020000000000000003700000000ffffffe9ffffffff",
            INIT_31 => X"0000002e00000000000000060000000000000013000000000000002f00000000",
            INIT_32 => X"fffffffbffffffffffffffedffffffff00000004000000000000000600000000",
            INIT_33 => X"fffffffcffffffff00000025000000000000002e00000000fffffff3ffffffff",
            INIT_34 => X"ffffffc4ffffffff00000007000000000000000c00000000fffffff9ffffffff",
            INIT_35 => X"ffffffe7ffffffff0000000400000000ffffffd1ffffffffffffffdcffffffff",
            INIT_36 => X"00000020000000000000001e0000000000000000000000000000001600000000",
            INIT_37 => X"0000000d00000000ffffffd3ffffffffffffffe0ffffffff0000001200000000",
            INIT_38 => X"0000002000000000ffffffe0ffffffffffffffcefffffffffffffffdffffffff",
            INIT_39 => X"0000001a00000000ffffffd3ffffffffffffffbaffffffffffffffe9ffffffff",
            INIT_3A => X"0000000400000000fffffffaffffffffffffffe7ffffffffffffffe7ffffffff",
            INIT_3B => X"0000001400000000ffffffebffffffff0000003300000000fffffff5ffffffff",
            INIT_3C => X"0000001200000000000000070000000000000011000000000000001900000000",
            INIT_3D => X"fffffff0ffffffff000000040000000000000001000000000000000a00000000",
            INIT_3E => X"00000016000000000000000c00000000fffffffcffffffff0000000c00000000",
            INIT_3F => X"fffffffcffffffff000000230000000000000019000000000000001300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffebffffffffffffffe9fffffffffffffff6ffffffffffffffecffffffff",
            INIT_41 => X"0000001000000000fffffff9ffffffffffffffdffffffffffffffff6ffffffff",
            INIT_42 => X"0000001500000000fffffff6fffffffffffffff4ffffffff0000000300000000",
            INIT_43 => X"ffffffb2ffffffff0000001d000000000000000300000000fffffff6ffffffff",
            INIT_44 => X"ffffffedffffffffffffffdfffffffff00000010000000000000000200000000",
            INIT_45 => X"0000000900000000fffffffaffffffff0000001700000000ffffffebffffffff",
            INIT_46 => X"fffffffeffffffff00000018000000000000003700000000ffffffffffffffff",
            INIT_47 => X"0000000900000000000000010000000000000028000000000000001f00000000",
            INIT_48 => X"ffffffd2fffffffffffffff8ffffffff0000000d00000000ffffffe9ffffffff",
            INIT_49 => X"0000000900000000ffffffd4ffffffffffffffcfffffffffffffffd4ffffffff",
            INIT_4A => X"0000004d00000000000000240000000000000006000000000000002c00000000",
            INIT_4B => X"fffffffdfffffffffffffffeffffffff00000000000000000000000000000000",
            INIT_4C => X"0000003400000000ffffffddffffffff00000010000000000000002300000000",
            INIT_4D => X"0000000f000000000000000300000000fffffff4ffffffff0000001e00000000",
            INIT_4E => X"00000009000000000000001200000000fffffff0ffffffff0000002300000000",
            INIT_4F => X"ffffffe1ffffffff0000000e0000000000000000000000000000000900000000",
            INIT_50 => X"fffffff0fffffffffffffff2ffffffff00000020000000000000000200000000",
            INIT_51 => X"000000030000000000000007000000000000001a000000000000000c00000000",
            INIT_52 => X"0000003500000000fffffff3ffffffff00000024000000000000001300000000",
            INIT_53 => X"0000000000000000000000120000000000000002000000000000002500000000",
            INIT_54 => X"00000016000000000000001400000000ffffffaeffffffffffffffd9ffffffff",
            INIT_55 => X"ffffffaeffffffff00000031000000000000003600000000ffffffb3ffffffff",
            INIT_56 => X"0000001300000000000000030000000000000046000000000000000a00000000",
            INIT_57 => X"ffffffedffffffff00000006000000000000002100000000fffffff4ffffffff",
            INIT_58 => X"ffffffe3ffffffffffffffdafffffffffffffff1fffffffffffffffaffffffff",
            INIT_59 => X"fffffffbffffffffffffffc9ffffffff0000000000000000fffffffcffffffff",
            INIT_5A => X"00000000000000000000001d00000000fffffff6ffffffff0000000b00000000",
            INIT_5B => X"ffffffe8fffffffffffffff8ffffffff00000009000000000000000000000000",
            INIT_5C => X"ffffffd1ffffffff0000001500000000fffffff6fffffffffffffff7ffffffff",
            INIT_5D => X"00000015000000000000001900000000ffffffbbffffffffffffffdeffffffff",
            INIT_5E => X"ffffff9bffffffff00000006000000000000002000000000ffffffc1ffffffff",
            INIT_5F => X"0000000700000000000000040000000000000039000000000000000500000000",
            INIT_60 => X"fffffffaffffffff0000000b000000000000003600000000ffffffdbffffffff",
            INIT_61 => X"0000000000000000ffffffefffffffff00000039000000000000002b00000000",
            INIT_62 => X"0000000900000000fffffff2ffffffff0000001c00000000fffffff5ffffffff",
            INIT_63 => X"0000001200000000fffffffcffffffff0000000d000000000000002000000000",
            INIT_64 => X"00000019000000000000004a000000000000004a00000000fffffffaffffffff",
            INIT_65 => X"fffffffbffffffffffffffc2ffffffff00000052000000000000004500000000",
            INIT_66 => X"0000002d00000000fffffff4ffffffffffffffc6ffffffff0000001600000000",
            INIT_67 => X"ffffffdaffffffff0000001d000000000000002600000000ffffffdfffffffff",
            INIT_68 => X"0000000500000000000000390000000000000017000000000000001700000000",
            INIT_69 => X"0000001400000000ffffffceffffffffffffffffffffffffffffffe9ffffffff",
            INIT_6A => X"000000270000000000000017000000000000000a000000000000000500000000",
            INIT_6B => X"fffffff2ffffffff0000002c00000000ffffffdaffffffffffffffe2ffffffff",
            INIT_6C => X"ffffffd4ffffffff00000000000000000000002a00000000ffffffd2ffffffff",
            INIT_6D => X"0000002c00000000ffffffdbffffffffffffffefffffffff0000003700000000",
            INIT_6E => X"00000000000000000000003f00000000ffffffd1fffffffffffffff1ffffffff",
            INIT_6F => X"ffffffd0ffffffffffffffcfffffffff0000002f00000000ffffffd9ffffffff",
            INIT_70 => X"0000002c00000000ffffffc9fffffffffffffff6ffffffff0000001000000000",
            INIT_71 => X"0000001800000000ffffffeeffffffffffffffe5fffffffffffffff5ffffffff",
            INIT_72 => X"0000002d000000000000000e00000000ffffffccffffffff0000000600000000",
            INIT_73 => X"00000002000000000000002b00000000ffffffe8ffffffffffffffe1ffffffff",
            INIT_74 => X"00000002000000000000003000000000ffffffccffffffffffffffe2ffffffff",
            INIT_75 => X"ffffffacffffffff00000003000000000000001c00000000ffffffdcffffffff",
            INIT_76 => X"0000001500000000000000010000000000000031000000000000003f00000000",
            INIT_77 => X"fffffff1ffffffff000000190000000000000007000000000000001a00000000",
            INIT_78 => X"fffffffdffffffff0000000d00000000ffffffd4ffffffff0000000d00000000",
            INIT_79 => X"ffffffdefffffffffffffff4ffffffff00000015000000000000000a00000000",
            INIT_7A => X"fffffff2ffffffffffffff9fffffffff0000000100000000fffffffbffffffff",
            INIT_7B => X"0000004b000000000000002300000000ffffffd0ffffffff0000003300000000",
            INIT_7C => X"fffffffaffffffff0000003f000000000000000c00000000ffffffb6ffffffff",
            INIT_7D => X"fffffff8ffffffffffffffe9fffffffffffffff7fffffffffffffff3ffffffff",
            INIT_7E => X"0000001200000000fffffff5ffffffff00000014000000000000000500000000",
            INIT_7F => X"0000000f00000000fffffffeffffffff0000001c00000000ffffffe9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE21;


    MEM_IWGHT_LAYER2_INSTANCE22 : if BRAM_NAME = "iwght_layer2_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff8fffffffffffffff3ffffffff00000015000000000000001600000000",
            INIT_01 => X"0000000b00000000fffffff6ffffffffffffffcdffffffffffffffe3ffffffff",
            INIT_02 => X"ffffffe8ffffffff0000001c00000000fffffffcffffffffffffffcbffffffff",
            INIT_03 => X"fffffff5ffffffff0000002b000000000000001a00000000ffffffefffffffff",
            INIT_04 => X"ffffffddffffffffffffffe9ffffffff0000002300000000ffffffebffffffff",
            INIT_05 => X"ffffffdcffffffffffffffccffffffff0000000a000000000000005000000000",
            INIT_06 => X"0000000000000000ffffffc8ffffffff0000003b00000000ffffffffffffffff",
            INIT_07 => X"0000001500000000fffffff6ffffffffffffffc1ffffffff0000002e00000000",
            INIT_08 => X"ffffffe4fffffffffffffff6ffffffff00000002000000000000001400000000",
            INIT_09 => X"fffffff1ffffffff0000000500000000ffffffe8ffffffff0000000100000000",
            INIT_0A => X"00000027000000000000000a000000000000002300000000ffffffeaffffffff",
            INIT_0B => X"0000000300000000ffffffedfffffffffffffffcffffffff0000002f00000000",
            INIT_0C => X"fffffff0ffffffffffffffe9ffffffffffffffcaffffffffffffffe4ffffffff",
            INIT_0D => X"ffffffd2ffffffffffffffc6ffffffff0000000d00000000fffffff7ffffffff",
            INIT_0E => X"ffffffcffffffffffffffff9ffffffff00000016000000000000003300000000",
            INIT_0F => X"ffffffc9ffffffff00000020000000000000001600000000ffffffcdffffffff",
            INIT_10 => X"ffffffeeffffffffffffffcbffffffff0000002d00000000ffffffbbffffffff",
            INIT_11 => X"0000001500000000ffffffaeffffffffffffffc7fffffffffffffff3ffffffff",
            INIT_12 => X"00000025000000000000005f00000000ffffffc0ffffffffffffffc7ffffffff",
            INIT_13 => X"ffffffe8fffffffffffffffbffffffff0000003300000000fffffff3ffffffff",
            INIT_14 => X"ffffffe7ffffffffffffffeffffffffffffffff6ffffffff0000001000000000",
            INIT_15 => X"00000008000000000000003700000000ffffffd6fffffffffffffff3ffffffff",
            INIT_16 => X"ffffffeaffffffff00000000000000000000000d00000000fffffff2ffffffff",
            INIT_17 => X"ffffffe8ffffffffffffffecffffffff00000007000000000000000500000000",
            INIT_18 => X"fffffff0ffffffffffffffc9ffffffff00000052000000000000001100000000",
            INIT_19 => X"0000001b00000000ffffffedffffffffffffffceffffffff0000001100000000",
            INIT_1A => X"0000001f00000000ffffffedffffffff0000001c000000000000000e00000000",
            INIT_1B => X"ffffffffffffffff0000000400000000ffffffd3fffffffffffffffbffffffff",
            INIT_1C => X"ffffffd6ffffffffffffffc0ffffffff0000000e00000000ffffffd4ffffffff",
            INIT_1D => X"0000001500000000fffffff5fffffffffffffffcffffffff0000002800000000",
            INIT_1E => X"00000001000000000000000f00000000ffffffc1fffffffffffffffdffffffff",
            INIT_1F => X"0000000000000000ffffffeffffffffffffffffcffffffff0000000a00000000",
            INIT_20 => X"ffffffedfffffffffffffffeffffffff0000000b00000000ffffffebffffffff",
            INIT_21 => X"ffffffdbffffffffffffffe1ffffffff0000002a00000000ffffffebffffffff",
            INIT_22 => X"ffffffd9ffffffffffffffbeffffffffffffffe9fffffffffffffff3ffffffff",
            INIT_23 => X"0000000b000000000000000900000000ffffffe3ffffffff0000003100000000",
            INIT_24 => X"ffffffe1ffffffffffffffe4ffffffffffffffceffffffffffffffe8ffffffff",
            INIT_25 => X"0000002600000000ffffffe9ffffffff0000000200000000ffffffcdffffffff",
            INIT_26 => X"0000001f00000000000000080000000000000013000000000000004c00000000",
            INIT_27 => X"00000005000000000000000300000000ffffffedffffffff0000000a00000000",
            INIT_28 => X"ffffffe0ffffffffffffffe0ffffffff00000004000000000000000700000000",
            INIT_29 => X"0000003100000000ffffffc6ffffffffffffffddffffffffffffffd2ffffffff",
            INIT_2A => X"00000003000000000000002b00000000fffffffbfffffffffffffff3ffffffff",
            INIT_2B => X"0000000d0000000000000027000000000000002100000000fffffff7ffffffff",
            INIT_2C => X"00000043000000000000000f0000000000000029000000000000000800000000",
            INIT_2D => X"00000014000000000000003d000000000000004b000000000000005100000000",
            INIT_2E => X"0000000900000000fffffff0ffffffff0000001000000000fffffff9ffffffff",
            INIT_2F => X"0000000800000000ffffffddffffffff0000000b000000000000001200000000",
            INIT_30 => X"ffffffe1ffffffffffffffccffffffffffffffc7fffffffffffffffbffffffff",
            INIT_31 => X"000000060000000000000005000000000000000800000000ffffffe5ffffffff",
            INIT_32 => X"0000000100000000fffffff1ffffffff00000021000000000000000c00000000",
            INIT_33 => X"fffffffcfffffffffffffff6ffffffff0000000a000000000000000300000000",
            INIT_34 => X"00000008000000000000000b00000000fffffff4ffffffff0000000200000000",
            INIT_35 => X"ffffffedffffffff0000001800000000fffffffefffffffffffffff6ffffffff",
            INIT_36 => X"0000000600000000fffffff5ffffffff0000000f000000000000001700000000",
            INIT_37 => X"00000003000000000000001100000000fffffff9ffffffff0000001500000000",
            INIT_38 => X"0000000c000000000000001300000000ffffffe8fffffffffffffffeffffffff",
            INIT_39 => X"0000000200000000000000220000000000000011000000000000003e00000000",
            INIT_3A => X"ffffffdcfffffffffffffffbffffffff0000003600000000ffffffd2ffffffff",
            INIT_3B => X"0000001400000000ffffffc4fffffffffffffffbfffffffffffffff4ffffffff",
            INIT_3C => X"00000001000000000000000000000000ffffffc7ffffffffffffffd9ffffffff",
            INIT_3D => X"000000160000000000000004000000000000000800000000ffffffffffffffff",
            INIT_3E => X"0000000f000000000000004d0000000000000070000000000000004b00000000",
            INIT_3F => X"0000001500000000ffffffeeffffffff0000003e000000000000004a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000002000000000000000b00000000ffffffecffffffff0000003300000000",
            INIT_41 => X"00000027000000000000001900000000fffffffcffffffff0000002600000000",
            INIT_42 => X"ffffffd3ffffffff0000001b000000000000001e000000000000000700000000",
            INIT_43 => X"fffffffaffffffff00000007000000000000002e00000000ffffffdbffffffff",
            INIT_44 => X"0000000c00000000ffffffd8fffffffffffffff8ffffffff0000002e00000000",
            INIT_45 => X"00000000000000000000000600000000fffffffbffffffff0000002d00000000",
            INIT_46 => X"ffffffd6ffffffff0000000000000000ffffffe6ffffffff0000000400000000",
            INIT_47 => X"fffffff2fffffffffffffff6ffffffffffffffb1ffffffffffffffe0ffffffff",
            INIT_48 => X"fffffff8ffffffff0000003900000000ffffffb3ffffffffffffffd8ffffffff",
            INIT_49 => X"0000000e000000000000000e000000000000001700000000ffffffe2ffffffff",
            INIT_4A => X"ffffffd1ffffffff0000001d00000000fffffff8ffffffffffffffdfffffffff",
            INIT_4B => X"ffffffe0fffffffffffffff1ffffffffffffffc4ffffffffffffffe8ffffffff",
            INIT_4C => X"0000001600000000fffffff7ffffffffffffffe6ffffffff0000000f00000000",
            INIT_4D => X"0000001e000000000000000100000000ffffffdfffffffffffffffbfffffffff",
            INIT_4E => X"fffffffeffffffff0000003300000000ffffffe7ffffffffffffffe1ffffffff",
            INIT_4F => X"ffffffecffffffff00000031000000000000001100000000ffffffe7ffffffff",
            INIT_50 => X"fffffffbfffffffffffffffbffffffff0000001900000000ffffffffffffffff",
            INIT_51 => X"0000001c000000000000001c000000000000001f000000000000001400000000",
            INIT_52 => X"0000003900000000ffffffc0ffffffffffffffbdffffffff0000000f00000000",
            INIT_53 => X"00000008000000000000002900000000ffffffeeffffffffffffffc9ffffffff",
            INIT_54 => X"ffffffa3ffffffffffffffa8fffffffffffffff6ffffffff0000000800000000",
            INIT_55 => X"ffffff9fffffffffffffffaaffffffffffffffbdffffffffffffffcbffffffff",
            INIT_56 => X"00000011000000000000000800000000ffffffe2ffffffff0000000300000000",
            INIT_57 => X"00000020000000000000000f0000000000000041000000000000003100000000",
            INIT_58 => X"0000000e000000000000001f0000000000000015000000000000000c00000000",
            INIT_59 => X"ffffff9cffffffffffffffb0ffffffffffffff7dffffffffffffffdaffffffff",
            INIT_5A => X"fffffffefffffffffffffff4ffffffffffffffeeffffffffffffffbeffffffff",
            INIT_5B => X"0000001b0000000000000033000000000000004100000000ffffffffffffffff",
            INIT_5C => X"000000070000000000000010000000000000001f000000000000001800000000",
            INIT_5D => X"ffffffe9fffffffffffffff4ffffffff0000000500000000ffffffe8ffffffff",
            INIT_5E => X"0000000000000000fffffff9fffffffffffffff4fffffffffffffff9ffffffff",
            INIT_5F => X"fffffff6ffffffff0000001e000000000000001800000000fffffffdffffffff",
            INIT_60 => X"ffffffd9ffffffff000000090000000000000001000000000000000300000000",
            INIT_61 => X"ffffffebffffffff0000000900000000ffffffe3ffffffffffffffe3ffffffff",
            INIT_62 => X"ffffffe1ffffffff0000003d00000000ffffffdeffffffffffffffddffffffff",
            INIT_63 => X"fffffff9ffffffffffffffdfffffffff00000020000000000000000000000000",
            INIT_64 => X"0000001500000000fffffffafffffffffffffff1ffffffff0000000d00000000",
            INIT_65 => X"ffffffebffffffff0000000c00000000fffffffeffffffffffffffe9ffffffff",
            INIT_66 => X"ffffffd7ffffffffffffffcfffffffff00000022000000000000001500000000",
            INIT_67 => X"0000001200000000fffffff0fffffffffffffff9fffffffffffffff8ffffffff",
            INIT_68 => X"00000010000000000000000800000000fffffffbffffffff0000001100000000",
            INIT_69 => X"0000000b000000000000000400000000ffffffffffffffff0000000900000000",
            INIT_6A => X"fffffff0fffffffffffffff8ffffffff0000000800000000ffffffc5ffffffff",
            INIT_6B => X"000000170000000000000008000000000000000c000000000000002d00000000",
            INIT_6C => X"0000000d000000000000000b0000000000000021000000000000001f00000000",
            INIT_6D => X"0000001e00000000ffffffe6ffffffffffffffbfffffffff0000001d00000000",
            INIT_6E => X"ffffffe3ffffffff00000017000000000000000300000000ffffffd1ffffffff",
            INIT_6F => X"0000002c0000000000000033000000000000000b000000000000001300000000",
            INIT_70 => X"fffffff4ffffffff000000280000000000000011000000000000001500000000",
            INIT_71 => X"00000016000000000000000f00000000fffffff9ffffffff0000001800000000",
            INIT_72 => X"0000002400000000ffffffe5ffffffff0000000b000000000000000c00000000",
            INIT_73 => X"0000000c0000000000000028000000000000000300000000fffffff9ffffffff",
            INIT_74 => X"000000020000000000000044000000000000002b00000000ffffffc7ffffffff",
            INIT_75 => X"0000005500000000000000170000000000000048000000000000003400000000",
            INIT_76 => X"fffffffcffffffffffffffdaffffffffffffffdeffffffff0000003900000000",
            INIT_77 => X"0000001e000000000000000300000000ffffffefffffffff0000000000000000",
            INIT_78 => X"0000002d00000000fffffffcffffffff00000024000000000000000300000000",
            INIT_79 => X"fffffffaffffffff0000002200000000fffffffafffffffffffffff3ffffffff",
            INIT_7A => X"0000001e00000000fffffff1ffffffff0000001b00000000fffffff2ffffffff",
            INIT_7B => X"0000000e000000000000001400000000fffffff6ffffffff0000002400000000",
            INIT_7C => X"0000001c000000000000000b0000000000000019000000000000000c00000000",
            INIT_7D => X"0000001c00000000ffffffdfffffffff0000001a000000000000000300000000",
            INIT_7E => X"0000000f00000000fffffff1ffffffffffffffe3fffffffffffffffbffffffff",
            INIT_7F => X"ffffffeeffffffff00000000000000000000000400000000ffffffd9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE22;


    MEM_IWGHT_LAYER2_INSTANCE23 : if BRAM_NAME = "iwght_layer2_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000fffffff5ffffffff00000018000000000000002a00000000",
            INIT_01 => X"fffffff4ffffffff0000000b00000000fffffff8ffffffff0000000300000000",
            INIT_02 => X"00000003000000000000002600000000ffffffe4ffffffff0000002d00000000",
            INIT_03 => X"0000000b0000000000000007000000000000001e00000000fffffff0ffffffff",
            INIT_04 => X"00000011000000000000000c00000000ffffffdbffffffff0000000400000000",
            INIT_05 => X"0000001500000000fffffff4ffffffff0000001a000000000000000300000000",
            INIT_06 => X"ffffffefffffffff0000000b00000000ffffffb2ffffffff0000000a00000000",
            INIT_07 => X"0000002900000000ffffffecffffffffffffffd9fffffffffffffff8ffffffff",
            INIT_08 => X"0000001600000000ffffffd6ffffffffffffffc6ffffffff0000000100000000",
            INIT_09 => X"0000003a000000000000003400000000ffffffeffffffffffffffff9ffffffff",
            INIT_0A => X"0000001200000000ffffffe0ffffffff00000009000000000000002900000000",
            INIT_0B => X"00000015000000000000000600000000ffffffd5ffffffff0000001700000000",
            INIT_0C => X"ffffffffffffffff00000025000000000000000700000000ffffffe7ffffffff",
            INIT_0D => X"0000001c000000000000000d0000000000000014000000000000001100000000",
            INIT_0E => X"0000000100000000fffffff8fffffffffffffff9ffffffff0000001500000000",
            INIT_0F => X"00000006000000000000001a00000000ffffffe8fffffffffffffff1ffffffff",
            INIT_10 => X"0000000b000000000000000f000000000000000c000000000000000c00000000",
            INIT_11 => X"00000006000000000000000900000000ffffffefffffffff0000002b00000000",
            INIT_12 => X"ffffffeeffffffff0000000b00000000fffffff7fffffffffffffffaffffffff",
            INIT_13 => X"00000016000000000000000000000000fffffffdffffffff0000000200000000",
            INIT_14 => X"fffffff4ffffffff00000004000000000000001700000000ffffffe0ffffffff",
            INIT_15 => X"fffffff2ffffffffffffffecfffffffffffffff8ffffffff0000001400000000",
            INIT_16 => X"0000001000000000ffffffe5ffffffff0000000200000000fffffff0ffffffff",
            INIT_17 => X"00000004000000000000000000000000ffffffe6ffffffff0000001100000000",
            INIT_18 => X"0000000600000000fffffff9fffffffffffffff6ffffffff0000000f00000000",
            INIT_19 => X"ffffffefffffffffffffffe9ffffffffffffffe9ffffffffffffffe7ffffffff",
            INIT_1A => X"0000003200000000fffffffcffffffffffffffdffffffffffffffff9ffffffff",
            INIT_1B => X"0000001f0000000000000016000000000000001200000000fffffffbffffffff",
            INIT_1C => X"ffffffe8ffffffffffffffccfffffffffffffff0ffffffff0000003c00000000",
            INIT_1D => X"0000000900000000ffffffd1ffffffffffffffe6ffffffffffffffe1ffffffff",
            INIT_1E => X"ffffffeefffffffffffffffaffffffffffffffbdffffffffffffffe0ffffffff",
            INIT_1F => X"0000005200000000000000130000000000000012000000000000003500000000",
            INIT_20 => X"00000038000000000000001e0000000000000032000000000000005300000000",
            INIT_21 => X"fffffff5ffffffffffffffffffffffff0000002200000000ffffffd9ffffffff",
            INIT_22 => X"fffffff7ffffffffffffffddffffffff00000039000000000000000200000000",
            INIT_23 => X"fffffff5ffffffff0000001e000000000000001000000000ffffffe8ffffffff",
            INIT_24 => X"ffffffdafffffffffffffff5ffffffff00000000000000000000001500000000",
            INIT_25 => X"ffffffefffffffffffffffe9fffffffffffffff4fffffffffffffff5ffffffff",
            INIT_26 => X"0000002c00000000000000210000000000000016000000000000002000000000",
            INIT_27 => X"fffffff9ffffffff0000004500000000ffffffffffffffff0000000500000000",
            INIT_28 => X"ffffffefffffffffffffffe7ffffffff0000002a000000000000001500000000",
            INIT_29 => X"0000000700000000ffffffdeffffffff0000000f00000000ffffffeeffffffff",
            INIT_2A => X"ffffffa4ffffffff0000001500000000ffffffe8ffffffffffffffc0ffffffff",
            INIT_2B => X"0000003600000000ffffffc5ffffffff00000028000000000000001900000000",
            INIT_2C => X"ffffffebffffffffffffffeeffffffff0000002200000000ffffffe1ffffffff",
            INIT_2D => X"ffffffffffffffffffffffbdffffffffffffffe2ffffffff0000001300000000",
            INIT_2E => X"ffffffdeffffffffffffffc5ffffffffffffffeeffffffff0000000300000000",
            INIT_2F => X"00000025000000000000000900000000ffffffabffffffff0000003300000000",
            INIT_30 => X"fffffff3ffffffffffffffd1ffffffffffffffe1ffffffffffffffeeffffffff",
            INIT_31 => X"ffffffb1ffffffffffffffbcffffffffffffffd7ffffffffffffffddffffffff",
            INIT_32 => X"ffffff97ffffffffffffffaefffffffffffffff0ffffffffffffffb2ffffffff",
            INIT_33 => X"00000000000000000000000b0000000000000001000000000000001c00000000",
            INIT_34 => X"00000018000000000000001e00000000ffffffe2fffffffffffffff4ffffffff",
            INIT_35 => X"fffffff2fffffffffffffff7ffffffff00000001000000000000000c00000000",
            INIT_36 => X"0000002700000000ffffffdfffffffff00000011000000000000001d00000000",
            INIT_37 => X"0000000500000000ffffffedfffffffffffffffefffffffffffffff8ffffffff",
            INIT_38 => X"0000000200000000ffffffddffffffffffffffe7fffffffffffffffeffffffff",
            INIT_39 => X"0000002300000000fffffff9ffffffffffffffcdffffffffffffffecffffffff",
            INIT_3A => X"ffffffe7ffffffff0000002000000000ffffffe3fffffffffffffff7ffffffff",
            INIT_3B => X"ffffffeeffffffff00000009000000000000000d00000000ffffffefffffffff",
            INIT_3C => X"fffffff2ffffffffffffffd4ffffffffffffffe9ffffffffffffffe4ffffffff",
            INIT_3D => X"0000000b00000000000000100000000000000034000000000000000200000000",
            INIT_3E => X"fffffffcffffffffffffffedfffffffffffffff7ffffffff0000001300000000",
            INIT_3F => X"0000002800000000000000170000000000000008000000000000001400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003400000000000000250000000000000008000000000000000400000000",
            INIT_41 => X"00000017000000000000003c000000000000002b000000000000000b00000000",
            INIT_42 => X"0000002500000000ffffffd3ffffffff00000003000000000000002f00000000",
            INIT_43 => X"fffffffcffffffff000000120000000000000025000000000000002000000000",
            INIT_44 => X"00000027000000000000001200000000ffffffeaffffffff0000000e00000000",
            INIT_45 => X"fffffff9ffffffffffffffdfffffffff00000013000000000000001600000000",
            INIT_46 => X"ffffffe3ffffffffffffffd1fffffffffffffffcffffffffffffffedffffffff",
            INIT_47 => X"0000001b0000000000000016000000000000000200000000ffffffe7ffffffff",
            INIT_48 => X"00000013000000000000000f000000000000000b000000000000001200000000",
            INIT_49 => X"000000070000000000000001000000000000000b000000000000000a00000000",
            INIT_4A => X"00000006000000000000001b0000000000000026000000000000002100000000",
            INIT_4B => X"ffffffb9ffffffff0000000e000000000000002e000000000000001a00000000",
            INIT_4C => X"0000001500000000ffffffd7ffffffff0000001800000000fffffff7ffffffff",
            INIT_4D => X"0000002e000000000000000300000000fffffff3ffffffff0000000b00000000",
            INIT_4E => X"ffffffc3fffffffffffffff2ffffffffffffffc4ffffffffffffffd3ffffffff",
            INIT_4F => X"ffffffabffffffffffffffaeffffffffffffffeffffffffffffffff0ffffffff",
            INIT_50 => X"00000028000000000000000900000000ffffffc7ffffffffffffffc7ffffffff",
            INIT_51 => X"0000001000000000000000270000000000000030000000000000000300000000",
            INIT_52 => X"ffffffeaffffffff0000002500000000fffffffdffffffff0000001d00000000",
            INIT_53 => X"ffffffcaffffffff00000007000000000000002d00000000ffffffd8ffffffff",
            INIT_54 => X"0000001000000000ffffffedffffffff00000000000000000000000f00000000",
            INIT_55 => X"fffffffeffffffff0000000900000000fffffffdfffffffffffffff6ffffffff",
            INIT_56 => X"ffffffecffffffff0000000800000000fffffffbffffffffffffffe1ffffffff",
            INIT_57 => X"0000001600000000fffffffafffffffffffffffdffffffff0000000300000000",
            INIT_58 => X"0000001500000000000000000000000000000048000000000000006000000000",
            INIT_59 => X"ffffffe0ffffffffffffffd7ffffffff0000000b000000000000002b00000000",
            INIT_5A => X"ffffffe5ffffffffffffffbcffffffffffffffb8ffffffff0000000400000000",
            INIT_5B => X"00000015000000000000000800000000ffffffeeffffffffffffffd6ffffffff",
            INIT_5C => X"00000009000000000000000600000000ffffffd4fffffffffffffff8ffffffff",
            INIT_5D => X"0000000900000000fffffff0ffffffff0000000600000000ffffffeaffffffff",
            INIT_5E => X"00000002000000000000001a0000000000000003000000000000001200000000",
            INIT_5F => X"fffffff1ffffffff00000007000000000000002200000000fffffffbffffffff",
            INIT_60 => X"0000000800000000ffffffe8ffffffff0000000900000000ffffffffffffffff",
            INIT_61 => X"00000013000000000000000000000000fffffff8ffffffffffffffecffffffff",
            INIT_62 => X"00000001000000000000002a00000000ffffffebffffffff0000001900000000",
            INIT_63 => X"0000003600000000ffffffe4ffffffffffffffbeffffffffffffffe9ffffffff",
            INIT_64 => X"00000037000000000000001700000000ffffffebffffffff0000001e00000000",
            INIT_65 => X"0000004d00000000000000470000000000000013000000000000004200000000",
            INIT_66 => X"0000002800000000000000280000000000000041000000000000001100000000",
            INIT_67 => X"00000018000000000000004500000000ffffffe8ffffffff0000000e00000000",
            INIT_68 => X"00000022000000000000001700000000fffffff9ffffffff0000000800000000",
            INIT_69 => X"0000004a000000000000001a000000000000004b000000000000003800000000",
            INIT_6A => X"0000002e0000000000000017000000000000003e000000000000003700000000",
            INIT_6B => X"0000002c0000000000000026000000000000001f000000000000002e00000000",
            INIT_6C => X"ffffffe7ffffffff00000035000000000000003e000000000000002100000000",
            INIT_6D => X"00000016000000000000002f00000000fffffffffffffffffffffffcffffffff",
            INIT_6E => X"ffffffe6fffffffffffffffcffffffffffffffc9ffffffff0000001000000000",
            INIT_6F => X"fffffff0ffffffff0000000b000000000000000400000000fffffff5ffffffff",
            INIT_70 => X"ffffffdaffffffffffffffc8ffffffff0000000b000000000000000b00000000",
            INIT_71 => X"fffffff0fffffffffffffff3fffffffffffffff0ffffffffffffffc7ffffffff",
            INIT_72 => X"ffffffd9ffffffff000000000000000000000009000000000000000a00000000",
            INIT_73 => X"000000030000000000000012000000000000000000000000ffffffdfffffffff",
            INIT_74 => X"00000018000000000000002e0000000000000023000000000000001900000000",
            INIT_75 => X"ffffffeafffffffffffffff7ffffffff0000001300000000fffffff2ffffffff",
            INIT_76 => X"000000260000000000000000000000000000000a00000000fffffff9ffffffff",
            INIT_77 => X"ffffffeafffffffffffffff0fffffffffffffff1ffffffffffffffd1ffffffff",
            INIT_78 => X"0000001d000000000000000e000000000000001b000000000000000800000000",
            INIT_79 => X"00000006000000000000002100000000ffffffd5ffffffffffffffe4ffffffff",
            INIT_7A => X"fffffffbfffffffffffffff9ffffffff0000002700000000ffffffe9ffffffff",
            INIT_7B => X"fffffff0fffffffffffffffbfffffffffffffff6ffffffff0000002200000000",
            INIT_7C => X"ffffffe1ffffffffffffffdfffffffffffffffecffffffff0000000000000000",
            INIT_7D => X"fffffff4fffffffffffffff8ffffffffffffffd8fffffffffffffff1ffffffff",
            INIT_7E => X"fffffffcffffffffffffffc9ffffffffffffffbbffffffffffffffbaffffffff",
            INIT_7F => X"0000002400000000fffffffcffffffff00000029000000000000002a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE23;


    MEM_IWGHT_LAYER2_INSTANCE24 : if BRAM_NAME = "iwght_layer2_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000b0000000000000023000000000000000700000000fffffff1ffffffff",
            INIT_01 => X"0000003400000000ffffffe2ffffffffffffffc7ffffffffffffffdbffffffff",
            INIT_02 => X"0000000d000000000000002200000000fffffff5ffffffff0000001100000000",
            INIT_03 => X"ffffffc3ffffffff0000000000000000ffffffefffffffff0000000600000000",
            INIT_04 => X"fffffff1ffffffff000000290000000000000008000000000000000000000000",
            INIT_05 => X"0000002b000000000000001700000000fffffff4ffffffff0000000a00000000",
            INIT_06 => X"ffffffebfffffffffffffff6ffffffff0000001900000000fffffffeffffffff",
            INIT_07 => X"0000000a000000000000000000000000fffffffefffffffffffffff5ffffffff",
            INIT_08 => X"ffffffdcfffffffffffffff5ffffffffffffffdaffffffff0000000700000000",
            INIT_09 => X"0000000e00000000ffffffc4ffffffff0000001200000000fffffff7ffffffff",
            INIT_0A => X"fffffffdffffffff0000000400000000fffffffbfffffffffffffffdffffffff",
            INIT_0B => X"ffffffedffffffff0000001100000000ffffffe0ffffffff0000000700000000",
            INIT_0C => X"ffffffefffffffffffffffe0ffffffffffffffd2ffffffff0000000000000000",
            INIT_0D => X"0000000600000000fffffff0ffffffffffffffdbffffffffffffffebffffffff",
            INIT_0E => X"ffffffefffffffffffffffe7ffffffff0000001800000000ffffffeeffffffff",
            INIT_0F => X"fffffffbfffffffffffffff8ffffffff0000002400000000ffffffdcffffffff",
            INIT_10 => X"ffffffe4ffffffff0000000d0000000000000017000000000000000e00000000",
            INIT_11 => X"00000023000000000000003300000000ffffffccffffffffffffffddffffffff",
            INIT_12 => X"fffffff1fffffffffffffffcfffffffffffffffdffffffff0000000c00000000",
            INIT_13 => X"fffffff9ffffffffffffffe1fffffffffffffff3ffffffffffffffcbffffffff",
            INIT_14 => X"fffffff9ffffffff0000000e00000000ffffffccffffffffffffffd4ffffffff",
            INIT_15 => X"0000002c000000000000000b00000000fffffff9ffffffffffffffe9ffffffff",
            INIT_16 => X"0000001200000000000000120000000000000040000000000000003d00000000",
            INIT_17 => X"ffffffecffffffffffffffe5ffffffff00000049000000000000005300000000",
            INIT_18 => X"ffffffebffffffff0000001800000000ffffffdcffffffff0000002f00000000",
            INIT_19 => X"ffffffe3ffffffffffffffd7ffffffffffffffd8ffffffffffffffd8ffffffff",
            INIT_1A => X"0000000c000000000000000300000000fffffffdffffffff0000000c00000000",
            INIT_1B => X"ffffffe2fffffffffffffffdfffffffffffffffffffffffffffffff6ffffffff",
            INIT_1C => X"0000002400000000fffffff1ffffffffffffffebffffffffffffffdfffffffff",
            INIT_1D => X"0000001a00000000ffffffdaffffffffffffffddffffffff0000003100000000",
            INIT_1E => X"fffffff8fffffffffffffff1fffffffffffffff3ffffffffffffffeaffffffff",
            INIT_1F => X"0000003900000000fffffff8ffffffff0000001a000000000000003900000000",
            INIT_20 => X"0000002900000000ffffffe4ffffffff00000015000000000000005700000000",
            INIT_21 => X"ffffffc6ffffffffffffffcaffffffffffffffe0ffffffffffffffe7ffffffff",
            INIT_22 => X"ffffffe6ffffffffffffffd5fffffffffffffffeffffffffffffffdcffffffff",
            INIT_23 => X"ffffffd5fffffffffffffff6ffffffffffffffdbffffffffffffffdaffffffff",
            INIT_24 => X"ffffffeeffffffff00000000000000000000000500000000fffffff1ffffffff",
            INIT_25 => X"0000001b000000000000000400000000ffffffffffffffff0000000600000000",
            INIT_26 => X"0000000a00000000ffffffffffffffff0000001200000000fffffffaffffffff",
            INIT_27 => X"ffffffeeffffffff00000000000000000000000900000000ffffffeeffffffff",
            INIT_28 => X"0000002200000000000000240000000000000013000000000000000400000000",
            INIT_29 => X"00000013000000000000000d0000000000000009000000000000001000000000",
            INIT_2A => X"fffffffeffffffffffffffd4fffffffffffffff8fffffffffffffff9ffffffff",
            INIT_2B => X"0000003600000000000000220000000000000013000000000000001400000000",
            INIT_2C => X"000000210000000000000000000000000000003d000000000000003600000000",
            INIT_2D => X"00000027000000000000004c000000000000002900000000fffffff4ffffffff",
            INIT_2E => X"ffffffffffffffff000000510000000000000065000000000000005600000000",
            INIT_2F => X"fffffff9ffffffff0000001200000000fffffff7ffffffffffffffddffffffff",
            INIT_30 => X"0000001800000000fffffffdffffffffffffffc3ffffffffffffffd6ffffffff",
            INIT_31 => X"0000005200000000fffffff9ffffffff0000001400000000fffffffcffffffff",
            INIT_32 => X"0000004000000000000000440000000000000033000000000000006c00000000",
            INIT_33 => X"000000420000000000000048000000000000002f000000000000005700000000",
            INIT_34 => X"ffffff83ffffffff00000000000000000000001100000000ffffffddffffffff",
            INIT_35 => X"00000016000000000000000800000000ffffffb9ffffffffffffff98ffffffff",
            INIT_36 => X"ffffffafffffffffffffffcaffffffff00000000000000000000001400000000",
            INIT_37 => X"fffffffbffffffffffffffe0ffffffffffffffc5ffffffffffffffc2ffffffff",
            INIT_38 => X"ffffffd6ffffffff0000002c00000000ffffffe5ffffffffffffffe1ffffffff",
            INIT_39 => X"000000100000000000000010000000000000000c00000000fffffff3ffffffff",
            INIT_3A => X"ffffffebffffffff0000000e0000000000000017000000000000000a00000000",
            INIT_3B => X"000000190000000000000003000000000000001300000000fffffff9ffffffff",
            INIT_3C => X"fffffff8ffffffff0000000500000000fffffff6ffffffff0000002000000000",
            INIT_3D => X"fffffffbffffffff0000000c00000000fffffff8ffffffff0000000100000000",
            INIT_3E => X"00000009000000000000001b00000000ffffffdafffffffffffffff8ffffffff",
            INIT_3F => X"0000001e000000000000000d000000000000000d000000000000002300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000000000010000000000000004000000000000001400000000",
            INIT_41 => X"fffffff4fffffffffffffffdffffffff00000027000000000000002000000000",
            INIT_42 => X"ffffffe3ffffffff0000000000000000ffffffc3ffffffffffffffdfffffffff",
            INIT_43 => X"ffffffeeffffffff000000170000000000000029000000000000000e00000000",
            INIT_44 => X"0000000400000000ffffffcbffffffffffffffdbffffffff0000001e00000000",
            INIT_45 => X"ffffffe3ffffffff0000000300000000ffffffffffffffffffffffe7ffffffff",
            INIT_46 => X"fffffff1fffffffffffffff0ffffffffffffffc6fffffffffffffff0ffffffff",
            INIT_47 => X"00000027000000000000001f0000000000000013000000000000001600000000",
            INIT_48 => X"fffffffbffffffffffffffceffffffffffffffcaffffffff0000002300000000",
            INIT_49 => X"fffffff7ffffffffffffffd4ffffffffffffffbaffffffffffffff8cffffffff",
            INIT_4A => X"0000001300000000ffffffe0ffffffff0000001a000000000000000d00000000",
            INIT_4B => X"fffffff2ffffffffffffffeaffffffffffffffefffffffff0000000b00000000",
            INIT_4C => X"0000000b00000000000000400000000000000047000000000000003600000000",
            INIT_4D => X"0000000000000000fffffffdffffffff00000009000000000000002800000000",
            INIT_4E => X"00000006000000000000001c000000000000003200000000ffffffdeffffffff",
            INIT_4F => X"ffffffe6ffffffffffffffe7fffffffffffffffefffffffffffffffaffffffff",
            INIT_50 => X"000000420000000000000038000000000000000d000000000000000600000000",
            INIT_51 => X"fffffff5ffffffff0000000600000000fffffffbffffffff0000004b00000000",
            INIT_52 => X"0000001100000000ffffffe5ffffffffffffffa1ffffffffffffffb8ffffffff",
            INIT_53 => X"0000001800000000fffffff6ffffffff00000023000000000000003000000000",
            INIT_54 => X"ffffffc8ffffffffffffffbfffffffffffffffe9ffffffff0000001300000000",
            INIT_55 => X"fffffff2ffffffff0000001c0000000000000014000000000000001000000000",
            INIT_56 => X"ffffffa1ffffffffffffffd5fffffffffffffffcfffffffffffffffbffffffff",
            INIT_57 => X"000000180000000000000039000000000000002a00000000ffffffdeffffffff",
            INIT_58 => X"ffffffbdffffffff00000018000000000000001200000000fffffff5ffffffff",
            INIT_59 => X"0000000400000000ffffffffffffffffffffffe7ffffffffffffffd7ffffffff",
            INIT_5A => X"fffffffafffffffffffffff6fffffffffffffffcffffffff0000001400000000",
            INIT_5B => X"0000002700000000ffffffe8fffffffffffffffefffffffffffffff6ffffffff",
            INIT_5C => X"0000000f00000000fffffff0ffffffff00000044000000000000003300000000",
            INIT_5D => X"ffffffc1ffffffffffffff96ffffffffffffff9dffffffff0000000000000000",
            INIT_5E => X"ffffffdcffffffffffffffccffffffffffffffebffffffffffffffeeffffffff",
            INIT_5F => X"000000060000000000000012000000000000000000000000ffffffd6ffffffff",
            INIT_60 => X"fffffffdfffffffffffffff0ffffffff00000000000000000000000f00000000",
            INIT_61 => X"00000003000000000000001b00000000ffffffebffffffff0000001a00000000",
            INIT_62 => X"0000000a000000000000000e00000000fffffff2ffffffffffffffeeffffffff",
            INIT_63 => X"fffffff2ffffffff0000000100000000ffffffe7fffffffffffffff6ffffffff",
            INIT_64 => X"0000000100000000ffffffe1fffffffffffffff4ffffffff0000000400000000",
            INIT_65 => X"fffffff4ffffffffffffffddffffffff0000000c00000000fffffff7ffffffff",
            INIT_66 => X"ffffffeeffffffffffffffe7fffffffffffffff9ffffffff0000001200000000",
            INIT_67 => X"fffffff6ffffffffffffffc7ffffffffffffffdcffffffffffffffeaffffffff",
            INIT_68 => X"ffffffe6ffffffffffffffc6ffffffffffffffe0ffffffff0000000100000000",
            INIT_69 => X"fffffffaffffffff000000050000000000000001000000000000002100000000",
            INIT_6A => X"0000000b00000000ffffffd3fffffffffffffffcffffffffffffffccffffffff",
            INIT_6B => X"00000016000000000000000f00000000fffffff2ffffffff0000001b00000000",
            INIT_6C => X"ffffffe3ffffffffffffffeeffffffffffffffeaffffffff0000002000000000",
            INIT_6D => X"0000001c00000000ffffffcdffffffffffffffcaffffffffffffffc7ffffffff",
            INIT_6E => X"0000001100000000fffffff2ffffffff00000021000000000000002500000000",
            INIT_6F => X"ffffffecffffffff0000001400000000fffffff1ffffffff0000000500000000",
            INIT_70 => X"fffffffeffffffff00000005000000000000000300000000ffffffefffffffff",
            INIT_71 => X"0000000e00000000000000120000000000000001000000000000000e00000000",
            INIT_72 => X"ffffffeeffffffffffffffecffffffffffffffe5ffffffff0000001a00000000",
            INIT_73 => X"fffffff7ffffffffffffffeaffffffffffffffdbffffffffffffffe5ffffffff",
            INIT_74 => X"00000045000000000000000000000000ffffffd3ffffffffffffffe3ffffffff",
            INIT_75 => X"0000007000000000000000510000000000000014000000000000003d00000000",
            INIT_76 => X"fffffffeffffffff0000001500000000fffffff3fffffffffffffff7ffffffff",
            INIT_77 => X"0000004700000000ffffffe6fffffffffffffffeffffffff0000001100000000",
            INIT_78 => X"00000013000000000000002900000000ffffffd9ffffffff0000002900000000",
            INIT_79 => X"0000002000000000fffffffcffffffff0000003b000000000000003e00000000",
            INIT_7A => X"0000002100000000ffffffdbffffffff00000045000000000000004400000000",
            INIT_7B => X"000000020000000000000001000000000000000700000000ffffffffffffffff",
            INIT_7C => X"0000002900000000000000130000000000000003000000000000000c00000000",
            INIT_7D => X"0000000e00000000ffffffe6ffffffff00000012000000000000001e00000000",
            INIT_7E => X"ffffffddffffffff0000000800000000fffffff7ffffffffffffffe7ffffffff",
            INIT_7F => X"00000001000000000000000c000000000000000500000000fffffff1ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE24;


    MEM_IWGHT_LAYER2_INSTANCE25 : if BRAM_NAME = "iwght_layer2_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff9ffffffffffffffebfffffffffffffff8ffffffff0000000000000000",
            INIT_01 => X"00000019000000000000000c000000000000000b00000000fffffff6ffffffff",
            INIT_02 => X"0000000a00000000000000210000000000000031000000000000001000000000",
            INIT_03 => X"ffffffdbfffffffffffffffaffffffff0000000100000000fffffff6ffffffff",
            INIT_04 => X"fffffff5ffffffffffffffe2fffffffffffffff0ffffffff0000000800000000",
            INIT_05 => X"00000025000000000000000100000000fffffff6ffffffff0000001000000000",
            INIT_06 => X"0000000a00000000ffffffebfffffffffffffffaffffffffffffffeeffffffff",
            INIT_07 => X"0000000a00000000000000000000000000000007000000000000001a00000000",
            INIT_08 => X"0000000500000000ffffffccffffffffffffffb8ffffffffffffffc9ffffffff",
            INIT_09 => X"0000002500000000000000140000000000000019000000000000000200000000",
            INIT_0A => X"ffffffceffffffff0000001d00000000fffffff7ffffffff0000000700000000",
            INIT_0B => X"0000001700000000fffffff4fffffffffffffff2fffffffffffffff4ffffffff",
            INIT_0C => X"0000002a000000000000002000000000ffffffdffffffffffffffffaffffffff",
            INIT_0D => X"ffffffebffffffffffffffe2ffffffff0000000b000000000000000700000000",
            INIT_0E => X"0000002800000000000000110000000000000005000000000000000600000000",
            INIT_0F => X"0000000f000000000000000000000000fffffffbfffffffffffffffeffffffff",
            INIT_10 => X"00000026000000000000001a000000000000002e000000000000002000000000",
            INIT_11 => X"0000001800000000fffffffdffffffff00000031000000000000000e00000000",
            INIT_12 => X"ffffffd7ffffffff0000001900000000ffffffd5ffffffffffffffceffffffff",
            INIT_13 => X"000000340000000000000036000000000000004f00000000ffffffd7ffffffff",
            INIT_14 => X"ffffffe3ffffffffffffffd7fffffffffffffffafffffffffffffff2ffffffff",
            INIT_15 => X"00000024000000000000004c00000000ffffffd9ffffffffffffffe6ffffffff",
            INIT_16 => X"ffffffd2ffffffffffffffdcffffffffffffffdcffffffff0000002b00000000",
            INIT_17 => X"0000000500000000fffffff7ffffffffffffffe5ffffffffffffffe6ffffffff",
            INIT_18 => X"00000016000000000000000c0000000000000003000000000000002400000000",
            INIT_19 => X"00000016000000000000001a0000000000000028000000000000000b00000000",
            INIT_1A => X"ffffffe8ffffffff000000160000000000000033000000000000000900000000",
            INIT_1B => X"fffffffeffffffff0000001000000000ffffffebfffffffffffffff1ffffffff",
            INIT_1C => X"0000001a0000000000000000000000000000000300000000ffffffdeffffffff",
            INIT_1D => X"ffffffe4ffffffff0000000400000000ffffffdfffffffff0000000900000000",
            INIT_1E => X"0000001f000000000000001e00000000ffffffd1ffffffffffffffebffffffff",
            INIT_1F => X"fffffff7ffffffffffffffe4fffffffffffffff8fffffffffffffff1ffffffff",
            INIT_20 => X"0000000000000000ffffffe9fffffffffffffffdffffffff0000000800000000",
            INIT_21 => X"ffffffccffffffffffffffd9fffffffffffffffdffffffff0000001700000000",
            INIT_22 => X"000000190000000000000000000000000000000800000000ffffffe6ffffffff",
            INIT_23 => X"0000000c000000000000002b0000000000000031000000000000002800000000",
            INIT_24 => X"00000005000000000000000500000000ffffffecffffffff0000002300000000",
            INIT_25 => X"0000000300000000ffffffecffffffff0000000100000000ffffffebffffffff",
            INIT_26 => X"0000001200000000000000580000000000000043000000000000000b00000000",
            INIT_27 => X"ffffffd8ffffffffffffffe2ffffffff00000047000000000000002f00000000",
            INIT_28 => X"fffffff7ffffffffffffffe4ffffffff0000000a000000000000001100000000",
            INIT_29 => X"00000015000000000000000d000000000000000400000000ffffffffffffffff",
            INIT_2A => X"ffffffe6fffffffffffffffcffffffff00000010000000000000000900000000",
            INIT_2B => X"ffffffffffffffffffffffe5fffffffffffffffffffffffffffffffeffffffff",
            INIT_2C => X"ffffffe4ffffffff0000001d000000000000000d000000000000002a00000000",
            INIT_2D => X"0000000400000000fffffff5ffffffffffffffcfffffffffffffffd9ffffffff",
            INIT_2E => X"00000022000000000000001b0000000000000029000000000000000700000000",
            INIT_2F => X"fffffff5fffffffffffffffbffffffff0000002e000000000000002900000000",
            INIT_30 => X"0000001e00000000ffffffdaffffffff0000003e000000000000005100000000",
            INIT_31 => X"0000001200000000fffffffbfffffffffffffff1ffffffff0000001700000000",
            INIT_32 => X"0000001a000000000000000a000000000000000400000000fffffff1ffffffff",
            INIT_33 => X"00000000000000000000000d000000000000002a000000000000000900000000",
            INIT_34 => X"ffffffe4ffffffffffffffeeffffffffffffffe6ffffffffffffffecffffffff",
            INIT_35 => X"ffffffe7ffffffff000000160000000000000026000000000000002300000000",
            INIT_36 => X"ffffffe5ffffffff0000000300000000ffffffebffffffffffffffddffffffff",
            INIT_37 => X"000000050000000000000024000000000000001e000000000000000000000000",
            INIT_38 => X"ffffffecffffffff0000000800000000fffffffffffffffffffffffbffffffff",
            INIT_39 => X"fffffff0ffffffff0000000800000000fffffffbfffffffffffffff6ffffffff",
            INIT_3A => X"0000000600000000fffffffbfffffffffffffffaffffffff0000000f00000000",
            INIT_3B => X"0000000000000000ffffffe0fffffffffffffff0ffffffff0000000000000000",
            INIT_3C => X"0000000600000000ffffffe8ffffffff00000004000000000000000400000000",
            INIT_3D => X"ffffffecffffffff0000000000000000ffffffeffffffffffffffff7ffffffff",
            INIT_3E => X"ffffffebffffffff0000001000000000fffffffffffffffffffffff7ffffffff",
            INIT_3F => X"0000000d000000000000001200000000fffffffcfffffffffffffff2ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe8ffffffffffffffe8fffffffffffffff6ffffffff0000001a00000000",
            INIT_41 => X"0000001e00000000000000060000000000000002000000000000000c00000000",
            INIT_42 => X"ffffffefffffffff0000000c00000000fffffffbfffffffffffffffdffffffff",
            INIT_43 => X"0000000b0000000000000000000000000000001a00000000fffffff9ffffffff",
            INIT_44 => X"fffffffefffffffffffffff8ffffffff0000000700000000fffffff5ffffffff",
            INIT_45 => X"ffffffe9fffffffffffffff5ffffffffffffffedfffffffffffffff1ffffffff",
            INIT_46 => X"ffffffecffffffffffffffe5ffffffffffffffdaffffffff0000000700000000",
            INIT_47 => X"ffffffe4ffffffffffffffe9ffffffffffffffebffffffffffffffe4ffffffff",
            INIT_48 => X"000000000000000000000007000000000000000d00000000ffffffe5ffffffff",
            INIT_49 => X"00000000000000000000000b0000000000000008000000000000000c00000000",
            INIT_4A => X"fffffff6ffffffffffffffeafffffffffffffff2ffffffffffffffedffffffff",
            INIT_4B => X"ffffffdffffffffffffffffbffffffffffffffffffffffffffffffe8ffffffff",
            INIT_4C => X"ffffffe5ffffffffffffffe3ffffffff00000006000000000000001400000000",
            INIT_4D => X"ffffffedffffffff0000000b00000000ffffffebffffffffffffffebffffffff",
            INIT_4E => X"0000000800000000ffffffeefffffffffffffff0ffffffffffffffedffffffff",
            INIT_4F => X"0000000400000000fffffffbffffffffffffffeaffffffffffffffe7ffffffff",
            INIT_50 => X"ffffffe8ffffffff0000000000000000ffffffecfffffffffffffff8ffffffff",
            INIT_51 => X"ffffffe8fffffffffffffffaffffffffffffffedfffffffffffffff3ffffffff",
            INIT_52 => X"ffffffebfffffffffffffff3fffffffffffffff2fffffffffffffff3ffffffff",
            INIT_53 => X"ffffffe6ffffffff0000000400000000fffffff5ffffffffffffffedffffffff",
            INIT_54 => X"ffffffe2ffffffffffffffedffffffffffffffeeffffffff0000000a00000000",
            INIT_55 => X"ffffffdfffffffffffffffe1ffffffffffffffefffffffffffffffeeffffffff",
            INIT_56 => X"fffffff0ffffffff000000090000000000000006000000000000000000000000",
            INIT_57 => X"ffffffe5ffffffff00000001000000000000000500000000ffffffecffffffff",
            INIT_58 => X"0000000a00000000ffffffdcffffffffffffffebffffffff0000000800000000",
            INIT_59 => X"ffffffebfffffffffffffffbfffffffffffffff8fffffffffffffff0ffffffff",
            INIT_5A => X"0000000400000000ffffffe3ffffffff0000000a000000000000000100000000",
            INIT_5B => X"fffffff0ffffffff00000001000000000000000000000000ffffffe8ffffffff",
            INIT_5C => X"fffffffaffffffffffffffeefffffffffffffffbffffffffffffffe6ffffffff",
            INIT_5D => X"0000000d000000000000000500000000fffffff6fffffffffffffff4ffffffff",
            INIT_5E => X"fffffff4ffffffffffffffd9ffffffffffffffddfffffffffffffffdffffffff",
            INIT_5F => X"0000000c0000000000000000000000000000000100000000fffffffeffffffff",
            INIT_60 => X"fffffffcfffffffffffffff5fffffffffffffff8ffffffffffffffe5ffffffff",
            INIT_61 => X"fffffff1fffffffffffffff0fffffffffffffff1ffffffff0000000300000000",
            INIT_62 => X"ffffffe5ffffffff00000000000000000000000c000000000000000b00000000",
            INIT_63 => X"0000000000000000fffffffeffffffffffffffffffffffffffffffe1ffffffff",
            INIT_64 => X"fffffff0ffffffff0000000300000000ffffffeeffffffffffffffecffffffff",
            INIT_65 => X"fffffff5ffffffff0000000800000000ffffffe7ffffffff0000000f00000000",
            INIT_66 => X"ffffffe4ffffffff0000000000000000ffffffecffffffff0000000600000000",
            INIT_67 => X"0000000700000000fffffffaffffffff0000000a000000000000000d00000000",
            INIT_68 => X"ffffffeaffffffffffffffe9ffffffffffffffe1ffffffffffffffe3ffffffff",
            INIT_69 => X"ffffffe2fffffffffffffffaffffffffffffffeeffffffffffffffe8ffffffff",
            INIT_6A => X"00000005000000000000000500000000ffffffdfffffffff0000000100000000",
            INIT_6B => X"ffffffe4fffffffffffffff5fffffffffffffffcfffffffffffffff0ffffffff",
            INIT_6C => X"ffffffe5ffffffffffffffecffffffff00000003000000000000000300000000",
            INIT_6D => X"ffffffeaffffffffffffffe7ffffffffffffffffffffffff0000000a00000000",
            INIT_6E => X"ffffffe9ffffffffffffffffffffffffffffffe6fffffffffffffff6ffffffff",
            INIT_6F => X"0000000d00000000ffffffe6fffffffffffffff4ffffffffffffffe9ffffffff",
            INIT_70 => X"fffffff5ffffffffffffffedffffffffffffffe7fffffffffffffff8ffffffff",
            INIT_71 => X"ffffffefffffffffffffffe9ffffffff00000000000000000000000800000000",
            INIT_72 => X"ffffffe9ffffffffffffffecffffffff0000000700000000fffffffbffffffff",
            INIT_73 => X"fffffffcffffffffffffffeeffffffff0000000400000000ffffffe7ffffffff",
            INIT_74 => X"fffffffffffffffffffffffcffffffffffffffedffffffff0000000100000000",
            INIT_75 => X"fffffffcffffffff00000007000000000000000a00000000ffffffe9ffffffff",
            INIT_76 => X"fffffff7ffffffff00000002000000000000000200000000ffffffe2ffffffff",
            INIT_77 => X"00000002000000000000000e00000000fffffff5fffffffffffffff3ffffffff",
            INIT_78 => X"000000080000000000000001000000000000000200000000ffffffe7ffffffff",
            INIT_79 => X"fffffff8ffffffff0000000000000000fffffffbffffffffffffffe2ffffffff",
            INIT_7A => X"0000000000000000fffffff7ffffffffffffffefffffffff0000000500000000",
            INIT_7B => X"0000000a00000000ffffffeafffffffffffffff2fffffffffffffffaffffffff",
            INIT_7C => X"ffffffecffffffffffffffedffffffff00000000000000000000000200000000",
            INIT_7D => X"0000000a00000000fffffffbffffffff00000009000000000000000900000000",
            INIT_7E => X"fffffff9ffffffff0000000800000000fffffffcfffffffffffffff2ffffffff",
            INIT_7F => X"00000008000000000000001600000000fffffffffffffffffffffff1ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE25;


    MEM_IWGHT_LAYER2_INSTANCE26 : if BRAM_NAME = "iwght_layer2_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000008000000000000000000000000ffffffecfffffffffffffff6ffffffff",
            INIT_01 => X"0000000b000000000000000a000000000000000700000000ffffffe8ffffffff",
            INIT_02 => X"ffffffd3fffffffffffffff2ffffffffffffffefffffffffffffffebffffffff",
            INIT_03 => X"0000001500000000ffffffedfffffffffffffff8ffffffff0000001400000000",
            INIT_04 => X"0000000a000000000000001800000000ffffffdbffffffff0000000100000000",
            INIT_05 => X"000000100000000000000031000000000000003c000000000000000a00000000",
            INIT_06 => X"ffffffdbffffffff0000002b0000000000000037000000000000002f00000000",
            INIT_07 => X"ffffffe5ffffffffffffffc1ffffffffffffffd8ffffffff0000000b00000000",
            INIT_08 => X"ffffffc7ffffffffffffffb6ffffffffffffffd8ffffffffffffffb8ffffffff",
            INIT_09 => X"0000001a000000000000001c00000000fffffff9fffffffffffffffcffffffff",
            INIT_0A => X"000000550000000000000023000000000000004d000000000000003b00000000",
            INIT_0B => X"00000017000000000000002200000000fffffffaffffffff0000003000000000",
            INIT_0C => X"fffffff0fffffffffffffffbffffffff0000000a00000000ffffffeaffffffff",
            INIT_0D => X"0000001b000000000000002100000000fffffffdffffffffffffffdeffffffff",
            INIT_0E => X"fffffff1ffffffffffffffd2ffffffffffffffd8ffffffff0000001700000000",
            INIT_0F => X"fffffffcffffffffffffffe6ffffffffffffffcbffffffffffffffe2ffffffff",
            INIT_10 => X"ffffffffffffffff0000001600000000ffffffedffffffffffffffe7ffffffff",
            INIT_11 => X"00000005000000000000000b000000000000000b00000000fffffff8ffffffff",
            INIT_12 => X"fffffff3ffffffff00000023000000000000000d000000000000002a00000000",
            INIT_13 => X"ffffff95ffffffffffffffb9fffffffffffffff2ffffffff0000001a00000000",
            INIT_14 => X"000000140000000000000000000000000000000200000000ffffffb0ffffffff",
            INIT_15 => X"fffffff4ffffffff00000000000000000000001700000000ffffffc9ffffffff",
            INIT_16 => X"ffffffe2fffffffffffffff4ffffffff0000000300000000fffffffeffffffff",
            INIT_17 => X"ffffffdfffffffffffffffdafffffffffffffff6ffffffff0000000800000000",
            INIT_18 => X"fffffff7ffffffffffffffceffffffffffffffcbffffffffffffffd1ffffffff",
            INIT_19 => X"0000000c00000000fffffffbffffffff00000000000000000000001000000000",
            INIT_1A => X"0000001d00000000ffffffeaffffffffffffffc4fffffffffffffff9ffffffff",
            INIT_1B => X"ffffffe9fffffffffffffff1ffffffff0000000f000000000000001300000000",
            INIT_1C => X"0000000200000000ffffffe3ffffffff0000000e000000000000001000000000",
            INIT_1D => X"fffffffcffffffff0000000600000000ffffffccffffffff0000001400000000",
            INIT_1E => X"00000015000000000000000f000000000000000f00000000fffffffbffffffff",
            INIT_1F => X"00000011000000000000001b0000000000000022000000000000001600000000",
            INIT_20 => X"00000000000000000000000100000000ffffffd9ffffffff0000001900000000",
            INIT_21 => X"fffffff2ffffffffffffffd0ffffffffffffffabffffffffffffffa8ffffffff",
            INIT_22 => X"00000030000000000000001000000000ffffffd0ffffffff0000000b00000000",
            INIT_23 => X"0000003500000000000000440000000000000021000000000000000c00000000",
            INIT_24 => X"fffffff9ffffffff0000000d000000000000000100000000ffffffe9ffffffff",
            INIT_25 => X"000000210000000000000002000000000000001a000000000000000700000000",
            INIT_26 => X"0000001f00000000000000190000000000000006000000000000001400000000",
            INIT_27 => X"ffffffb7fffffffffffffff4ffffffffffffffefffffffffffffffefffffffff",
            INIT_28 => X"ffffffedffffffffffffffd6ffffffffffffffe9ffffffffffffffdfffffffff",
            INIT_29 => X"ffffffc1ffffffffffffffb6ffffffffffffffc1ffffffffffffffbdffffffff",
            INIT_2A => X"0000000e00000000ffffffe2ffffffff0000000200000000ffffffd5ffffffff",
            INIT_2B => X"fffffff0ffffffff000000040000000000000005000000000000000e00000000",
            INIT_2C => X"0000000e00000000000000190000000000000005000000000000000800000000",
            INIT_2D => X"0000002700000000ffffffd6ffffffffffffffeeffffffffffffffe3ffffffff",
            INIT_2E => X"00000019000000000000003b00000000ffffffdcfffffffffffffff5ffffffff",
            INIT_2F => X"ffffffe6fffffffffffffff0fffffffffffffffcfffffffffffffff8ffffffff",
            INIT_30 => X"0000002300000000ffffffebffffffff00000015000000000000001500000000",
            INIT_31 => X"0000002200000000000000100000000000000006000000000000001900000000",
            INIT_32 => X"0000000a000000000000000500000000ffffffeeffffffff0000001500000000",
            INIT_33 => X"0000001d00000000ffffffddffffffffffffffccffffffffffffffd4ffffffff",
            INIT_34 => X"fffffffcffffffffffffffdaffffffff00000027000000000000001600000000",
            INIT_35 => X"ffffffe5ffffffffffffffbdffffffffffffff9dffffffff0000000700000000",
            INIT_36 => X"ffffffd0ffffffffffffffeeffffffff0000003200000000ffffffecffffffff",
            INIT_37 => X"ffffff9afffffffffffffffbffffffffffffffd9ffffffffffffffccffffffff",
            INIT_38 => X"000000180000000000000005000000000000001500000000ffffffceffffffff",
            INIT_39 => X"0000002700000000fffffffdffffffff0000001e000000000000002000000000",
            INIT_3A => X"0000000100000000ffffffe7ffffffff00000007000000000000001f00000000",
            INIT_3B => X"0000001500000000fffffffdfffffffffffffff2ffffffff0000002300000000",
            INIT_3C => X"0000000a0000000000000017000000000000001500000000fffffff8ffffffff",
            INIT_3D => X"ffffffeeffffffffffffffe3ffffffff00000003000000000000000900000000",
            INIT_3E => X"fffffffbffffffffffffffe0ffffffff0000000e000000000000000c00000000",
            INIT_3F => X"ffffffc1ffffffff0000000900000000ffffffffffffffffffffffe6ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffc9ffffffffffffffc5ffffffffffffffccffffffffffffffb8ffffffff",
            INIT_41 => X"0000001700000000fffffff2ffffffffffffffdeffffffffffffffecffffffff",
            INIT_42 => X"ffffffbeffffffff0000000100000000fffffff7ffffffffffffffebffffffff",
            INIT_43 => X"0000000b000000000000000700000000fffffffbffffffffffffffd5ffffffff",
            INIT_44 => X"ffffffedffffffff000000210000000000000019000000000000000500000000",
            INIT_45 => X"fffffff3ffffffff000000120000000000000035000000000000003900000000",
            INIT_46 => X"000000170000000000000004000000000000001a000000000000000b00000000",
            INIT_47 => X"fffffff7fffffffffffffffcffffffffffffffd8ffffffff0000002f00000000",
            INIT_48 => X"0000000d000000000000000f000000000000000c00000000fffffffeffffffff",
            INIT_49 => X"ffffffffffffffff000000240000000000000012000000000000000100000000",
            INIT_4A => X"fffffff5ffffffffffffffe9fffffffffffffff7fffffffffffffffbffffffff",
            INIT_4B => X"ffffffb9ffffffffffffffd0ffffffffffffff98ffffffffffffffc9ffffffff",
            INIT_4C => X"0000000900000000fffffff0ffffffffffffffdeffffffffffffff8affffffff",
            INIT_4D => X"0000004e00000000000000350000000000000033000000000000000c00000000",
            INIT_4E => X"0000002600000000000000260000000000000055000000000000004300000000",
            INIT_4F => X"0000004300000000000000340000000000000026000000000000005900000000",
            INIT_50 => X"000000080000000000000018000000000000002c000000000000003100000000",
            INIT_51 => X"0000002a00000000ffffffe2ffffffffffffffecfffffffffffffffdffffffff",
            INIT_52 => X"00000018000000000000003100000000ffffffe6ffffffff0000002600000000",
            INIT_53 => X"ffffffe6ffffffff00000008000000000000000a00000000fffffffaffffffff",
            INIT_54 => X"0000002c000000000000000f000000000000001b000000000000001b00000000",
            INIT_55 => X"ffffffe4ffffffffffffffefffffffff00000022000000000000002800000000",
            INIT_56 => X"ffffffedfffffffffffffff7fffffffffffffffeffffffffffffffcdffffffff",
            INIT_57 => X"ffffffdfffffffffffffffffffffffff00000000000000000000002500000000",
            INIT_58 => X"fffffffdffffffffffffffeeffffffffffffffe0ffffffff0000000000000000",
            INIT_59 => X"fffffff0ffffffffffffffd9ffffffffffffffc7ffffffffffffffedffffffff",
            INIT_5A => X"0000001a00000000ffffffffffffffff0000000a000000000000003900000000",
            INIT_5B => X"fffffff6fffffffffffffffbfffffffffffffffcfffffffffffffff4ffffffff",
            INIT_5C => X"ffffffeeffffffffffffffdeffffffffffffffe8ffffffff0000000000000000",
            INIT_5D => X"0000001e00000000ffffffebfffffffffffffff6ffffffff0000002300000000",
            INIT_5E => X"00000006000000000000001600000000fffffffdfffffffffffffffcffffffff",
            INIT_5F => X"ffffffe1ffffffffffffffedffffffff0000001b000000000000001000000000",
            INIT_60 => X"fffffff0fffffffffffffff1fffffffffffffff1ffffffffffffffecffffffff",
            INIT_61 => X"0000002300000000fffffff9ffffffff0000002000000000fffffffcffffffff",
            INIT_62 => X"000000220000000000000006000000000000002c000000000000001b00000000",
            INIT_63 => X"00000018000000000000000000000000fffffff7ffffffffffffffedffffffff",
            INIT_64 => X"0000002800000000000000150000000000000013000000000000000b00000000",
            INIT_65 => X"ffffffe7ffffffffffffffccfffffffffffffffcffffffff0000000300000000",
            INIT_66 => X"ffffffebffffffffffffffe1ffffffffffffffcfffffffff0000001a00000000",
            INIT_67 => X"fffffffdffffffff0000000e00000000ffffffe1ffffffffffffffcfffffffff",
            INIT_68 => X"0000000000000000000000220000000000000004000000000000000a00000000",
            INIT_69 => X"fffffffffffffffffffffff9ffffffff00000034000000000000001700000000",
            INIT_6A => X"00000018000000000000001200000000ffffffe5fffffffffffffffeffffffff",
            INIT_6B => X"0000000a0000000000000006000000000000000b000000000000001200000000",
            INIT_6C => X"0000002a00000000ffffffedffffffffffffffe3ffffffff0000000600000000",
            INIT_6D => X"ffffffd3ffffffffffffffe2ffffffffffffffdbffffffffffffffabffffffff",
            INIT_6E => X"ffffffe3fffffffffffffff5ffffffff0000001800000000ffffffd2ffffffff",
            INIT_6F => X"0000001a00000000ffffffd7ffffffff00000009000000000000005100000000",
            INIT_70 => X"ffffffccffffffffffffffd1ffffffffffffffd2fffffffffffffff3ffffffff",
            INIT_71 => X"fffffffaffffffffffffffdcffffffffffffffe5ffffffffffffffbbffffffff",
            INIT_72 => X"ffffffdcfffffffffffffff5fffffffffffffff0ffffffffffffffeaffffffff",
            INIT_73 => X"ffffffeaffffffffffffffddffffffff0000001400000000fffffff1ffffffff",
            INIT_74 => X"0000001600000000fffffff5fffffffffffffff0ffffffff0000001700000000",
            INIT_75 => X"ffffffe7ffffffff0000000c000000000000000d00000000ffffffe0ffffffff",
            INIT_76 => X"ffffffe8ffffffffffffffdbffffffff00000022000000000000000900000000",
            INIT_77 => X"0000000600000000ffffffe1ffffffffffffffc9ffffffff0000000700000000",
            INIT_78 => X"ffffffe9ffffffff0000001d000000000000000a00000000ffffffe9ffffffff",
            INIT_79 => X"0000000000000000ffffffeeffffffff00000022000000000000000000000000",
            INIT_7A => X"ffffffe0ffffffff000000020000000000000034000000000000000500000000",
            INIT_7B => X"0000001100000000fffffff1ffffffff00000005000000000000003500000000",
            INIT_7C => X"0000001600000000fffffff8fffffffffffffff9fffffffffffffff1ffffffff",
            INIT_7D => X"000000040000000000000003000000000000001600000000fffffff5ffffffff",
            INIT_7E => X"0000003f00000000000000200000000000000045000000000000003600000000",
            INIT_7F => X"00000045000000000000005a000000000000001d000000000000006f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE26;


    MEM_IWGHT_LAYER2_INSTANCE27 : if BRAM_NAME = "iwght_layer2_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffff2ffffffffffffffe2ffffffff00000001000000000000003500000000",
            INIT_01 => X"ffffffd2fffffffffffffffbffffffffffffffe5ffffffffffffffe1ffffffff",
            INIT_02 => X"fffffffcffffffff0000000800000000ffffffd3ffffffffffffffaeffffffff",
            INIT_03 => X"ffffffd5fffffffffffffffaffffffff0000003100000000fffffff4ffffffff",
            INIT_04 => X"ffffffdaffffffffffffffe0fffffffffffffff9ffffffff0000003400000000",
            INIT_05 => X"ffffffe0ffffffffffffffdbffffffff0000001400000000ffffffe7ffffffff",
            INIT_06 => X"0000001b00000000fffffff2ffffffffffffffe1fffffffffffffffeffffffff",
            INIT_07 => X"0000007b00000000000000170000000000000049000000000000003500000000",
            INIT_08 => X"0000002700000000000000690000000000000038000000000000005b00000000",
            INIT_09 => X"0000001100000000ffffffdcffffffffffffffd6ffffffff0000003600000000",
            INIT_0A => X"ffffffe5ffffffffffffffe8ffffffff0000000500000000fffffffeffffffff",
            INIT_0B => X"ffffffefffffffffffffffe6ffffffff0000000f00000000ffffffe6ffffffff",
            INIT_0C => X"00000022000000000000001c00000000ffffffe7ffffffff0000001200000000",
            INIT_0D => X"fffffff7ffffffff0000001600000000fffffff1ffffffffffffffecffffffff",
            INIT_0E => X"ffffffe5ffffffff0000001e00000000fffffff1ffffffff0000000000000000",
            INIT_0F => X"ffffffc8fffffffffffffffbffffffff0000003500000000fffffff1ffffffff",
            INIT_10 => X"00000016000000000000000400000000fffffff7ffffffff0000001400000000",
            INIT_11 => X"0000000000000000ffffffe1ffffffff0000000000000000fffffff9ffffffff",
            INIT_12 => X"ffffffbdffffffff0000001e000000000000003f000000000000000800000000",
            INIT_13 => X"fffffff0ffffffff0000002600000000fffffff9ffffffffffffffd7ffffffff",
            INIT_14 => X"00000001000000000000001a00000000fffffff9ffffffffffffffd8ffffffff",
            INIT_15 => X"00000021000000000000000a000000000000000a00000000ffffffd8ffffffff",
            INIT_16 => X"ffffffd4ffffffff0000000900000000ffffffecffffffffffffffefffffffff",
            INIT_17 => X"fffffff0ffffffffffffffd1ffffffff0000000100000000ffffffdfffffffff",
            INIT_18 => X"fffffff0fffffffffffffff6ffffffffffffffcaffffffff0000001000000000",
            INIT_19 => X"0000000f0000000000000028000000000000000c000000000000001a00000000",
            INIT_1A => X"0000000600000000fffffffeffffffff0000002800000000fffffffcffffffff",
            INIT_1B => X"0000000b000000000000001900000000ffffffe9ffffffffffffffd8ffffffff",
            INIT_1C => X"000000180000000000000014000000000000000e00000000fffffff7ffffffff",
            INIT_1D => X"ffffffd6ffffffffffffffb0ffffffff00000015000000000000002300000000",
            INIT_1E => X"ffffffd4ffffffffffffffe6ffffffffffffffd7ffffffff0000000300000000",
            INIT_1F => X"ffffffccffffffffffffffd5fffffffffffffff8fffffffffffffff0ffffffff",
            INIT_20 => X"0000000200000000ffffffd8ffffffffffffffc2ffffffffffffffcbffffffff",
            INIT_21 => X"0000000600000000ffffffd1ffffffffffffffeaffffffffffffffe2ffffffff",
            INIT_22 => X"ffffffdfffffffff000000350000000000000033000000000000003100000000",
            INIT_23 => X"fffffff8ffffffffffffffd9ffffffff0000003300000000fffffff7ffffffff",
            INIT_24 => X"ffffffd3fffffffffffffff9ffffffffffffffe5ffffffff0000002300000000",
            INIT_25 => X"fffffffcffffffffffffffc1fffffffffffffff2ffffffffffffffd0ffffffff",
            INIT_26 => X"00000016000000000000000f00000000fffffff9fffffffffffffff4ffffffff",
            INIT_27 => X"0000004400000000ffffffddffffffffffffffc5ffffffff0000000d00000000",
            INIT_28 => X"ffffffdbffffffff0000002000000000ffffffe3ffffffffffffffd9ffffffff",
            INIT_29 => X"ffffffc2fffffffffffffff0fffffffffffffff1ffffffffffffffebffffffff",
            INIT_2A => X"fffffff0ffffffffffffffddffffffff00000010000000000000000100000000",
            INIT_2B => X"ffffffddffffffffffffffeaffffffffffffffceffffffffffffffd7ffffffff",
            INIT_2C => X"ffffffcbffffffff0000000300000000fffffffeffffffffffffff9fffffffff",
            INIT_2D => X"fffffff9ffffffffffffffccffffffffffffffe2ffffffffffffffc5ffffffff",
            INIT_2E => X"ffffffe8fffffffffffffffaffffffffffffffdfffffffff0000000100000000",
            INIT_2F => X"0000002200000000ffffffbeffffffff0000000200000000fffffffaffffffff",
            INIT_30 => X"0000000300000000ffffffdfffffffffffffffd9ffffffff0000004800000000",
            INIT_31 => X"ffffffd2ffffffffffffffe4ffffffffffffffddfffffffffffffff8ffffffff",
            INIT_32 => X"ffffffdafffffffffffffffaffffffffffffffd7fffffffffffffff4ffffffff",
            INIT_33 => X"ffffffcdffffffff00000016000000000000001700000000ffffff9cffffffff",
            INIT_34 => X"ffffffc4fffffffffffffff8ffffffff00000036000000000000000700000000",
            INIT_35 => X"0000000b00000000ffffffd0ffffffff00000030000000000000000500000000",
            INIT_36 => X"0000000b000000000000000e00000000fffffff3ffffffff0000002b00000000",
            INIT_37 => X"fffffffcffffffff0000002800000000fffffff2ffffffffffffffb4ffffffff",
            INIT_38 => X"00000038000000000000000600000000fffffff7fffffffffffffff1ffffffff",
            INIT_39 => X"0000003c000000000000004e0000000000000069000000000000003900000000",
            INIT_3A => X"ffffffe0ffffffff000000230000000000000066000000000000005500000000",
            INIT_3B => X"ffffffc4ffffffffffffffdaffffffff0000000000000000fffffffaffffffff",
            INIT_3C => X"ffffffaaffffffffffffffcaffffffffffffffdbffffffffffffffb1ffffffff",
            INIT_3D => X"fffffffcfffffffffffffff9ffffffffffffffd6ffffffffffffffdfffffffff",
            INIT_3E => X"fffffffdfffffffffffffffaffffffffffffffb4fffffffffffffff2ffffffff",
            INIT_3F => X"fffffffcffffffff0000000d000000000000000400000000ffffffd0ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffffbffffffffffffffe4ffffffffffffffeafffffffffffffff7ffffffff",
            INIT_41 => X"ffffffeffffffffffffffff1ffffffffffffffdbffffffff0000001800000000",
            INIT_42 => X"ffffffebffffffffffffffdcffffffffffffffe5fffffffffffffff2ffffffff",
            INIT_43 => X"0000000100000000ffffffe4ffffffff00000047000000000000001300000000",
            INIT_44 => X"ffffffeeffffffffffffffd0ffffffff0000003d000000000000002e00000000",
            INIT_45 => X"0000001c00000000ffffffdbffffffffffffffd5ffffffff0000002300000000",
            INIT_46 => X"ffffffdefffffffffffffff2ffffffff0000000b00000000fffffff0ffffffff",
            INIT_47 => X"ffffffd6ffffffff000000070000000000000027000000000000000b00000000",
            INIT_48 => X"0000000c00000000ffffffe9ffffffff00000021000000000000000300000000",
            INIT_49 => X"ffffffdfffffffff0000000a00000000fffffff9ffffffffffffffe9ffffffff",
            INIT_4A => X"fffffff2ffffffffffffffe9ffffffff0000001500000000ffffffe1ffffffff",
            INIT_4B => X"ffffffe6fffffffffffffff5fffffffffffffff7fffffffffffffffbffffffff",
            INIT_4C => X"ffffffd1ffffffff00000032000000000000000700000000ffffffedffffffff",
            INIT_4D => X"ffffffe3ffffffffffffffd6fffffffffffffffcffffffffffffffe7ffffffff",
            INIT_4E => X"ffffffd7ffffffff0000000e00000000ffffffdcfffffffffffffffbffffffff",
            INIT_4F => X"fffffff8ffffffff00000028000000000000001400000000ffffffd6ffffffff",
            INIT_50 => X"000000110000000000000003000000000000003a000000000000000e00000000",
            INIT_51 => X"ffffffecffffffffffffffcbffffffffffffffd8ffffffff0000002900000000",
            INIT_52 => X"ffffffefffffffff0000000700000000fffffff4ffffffffffffffeaffffffff",
            INIT_53 => X"ffffffccffffffffffffffdcffffffff00000043000000000000001700000000",
            INIT_54 => X"ffffffe2ffffffffffffffe1ffffffff00000004000000000000000500000000",
            INIT_55 => X"0000001400000000ffffffd2ffffffffffffffefffffffff0000000c00000000",
            INIT_56 => X"fffffff9ffffffff0000000a0000000000000012000000000000002400000000",
            INIT_57 => X"00000023000000000000001a0000000000000021000000000000001100000000",
            INIT_58 => X"0000000c00000000fffffffcfffffffffffffffcffffffff0000001200000000",
            INIT_59 => X"fffffff2fffffffffffffff0fffffffffffffff0ffffffff0000001400000000",
            INIT_5A => X"fffffff1ffffffff000000370000000000000036000000000000001900000000",
            INIT_5B => X"fffffff2ffffffff000000090000000000000013000000000000000300000000",
            INIT_5C => X"0000001500000000ffffffceffffffff0000000f00000000fffffffcffffffff",
            INIT_5D => X"fffffffbffffffff0000004100000000fffffffcffffffff0000000a00000000",
            INIT_5E => X"ffffffd6ffffffff0000000900000000fffffffbffffffffffffffe6ffffffff",
            INIT_5F => X"0000002c000000000000001000000000ffffffd2fffffffffffffff8ffffffff",
            INIT_60 => X"0000003a0000000000000023000000000000000c000000000000001100000000",
            INIT_61 => X"0000001e000000000000003100000000fffffffeffffffffffffffd5ffffffff",
            INIT_62 => X"ffffffc9ffffffff0000003400000000fffffffcffffffffffffffdcffffffff",
            INIT_63 => X"0000000c0000000000000019000000000000000600000000fffffff6ffffffff",
            INIT_64 => X"fffffff3fffffffffffffff9ffffffff00000008000000000000000000000000",
            INIT_65 => X"0000001000000000fffffffaffffffffffffffdaffffffff0000000100000000",
            INIT_66 => X"00000006000000000000000e000000000000000000000000ffffffc4ffffffff",
            INIT_67 => X"ffffffebffffffffffffffe0fffffffffffffffffffffffffffffffaffffffff",
            INIT_68 => X"0000000700000000fffffff5ffffffff0000000000000000ffffffe0ffffffff",
            INIT_69 => X"00000013000000000000000d00000000fffffff4ffffffff0000001f00000000",
            INIT_6A => X"fffffff1ffffffff00000007000000000000002a000000000000000a00000000",
            INIT_6B => X"0000000600000000fffffff9fffffffffffffff7ffffffff0000001500000000",
            INIT_6C => X"ffffffecfffffffffffffff0ffffffff0000000a000000000000003600000000",
            INIT_6D => X"fffffff0ffffffffffffffb7ffffffffffffffc4ffffffffffffffffffffffff",
            INIT_6E => X"0000001c00000000fffffff1ffffffffffffffedffffffffffffffe5ffffffff",
            INIT_6F => X"000000170000000000000007000000000000001d00000000ffffffebffffffff",
            INIT_70 => X"fffffffcffffffff0000002400000000fffffff6ffffffff0000001c00000000",
            INIT_71 => X"ffffffddfffffffffffffffdfffffffffffffff1ffffffffffffffd2ffffffff",
            INIT_72 => X"ffffffa8ffffffffffffffdbffffffffffffffc4ffffffffffffffe7ffffffff",
            INIT_73 => X"fffffff8ffffffff0000001000000000ffffffeaffffffff0000000000000000",
            INIT_74 => X"ffffffd9ffffffffffffffd0ffffffffffffffebffffffffffffffe5ffffffff",
            INIT_75 => X"ffffffddffffffff0000000700000000fffffff3ffffffffffffffd3ffffffff",
            INIT_76 => X"00000001000000000000000000000000fffffff4ffffffff0000000b00000000",
            INIT_77 => X"ffffffd4fffffffffffffffbffffffff00000019000000000000000600000000",
            INIT_78 => X"ffffffddfffffffffffffff0ffffffff0000000700000000ffffffefffffffff",
            INIT_79 => X"0000000700000000ffffffb7ffffffffffffffcdffffffffffffffccffffffff",
            INIT_7A => X"ffffffe3ffffffffffffffe1ffffffffffffffd9ffffffffffffffdaffffffff",
            INIT_7B => X"fffffff1ffffffffffffffebffffffffffffffe4ffffffffffffffc4ffffffff",
            INIT_7C => X"ffffff93ffffffffffffffbdffffffffffffffa4ffffffffffffffcdffffffff",
            INIT_7D => X"0000000600000000ffffffdfffffffffffffffe0ffffffffffffffc8ffffffff",
            INIT_7E => X"ffffffe7ffffffff00000011000000000000001f00000000ffffffdbffffffff",
            INIT_7F => X"0000001000000000fffffffaffffffff00000004000000000000002d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE27;


    MEM_IWGHT_LAYER2_INSTANCE28 : if BRAM_NAME = "iwght_layer2_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004a0000000000000010000000000000000a000000000000000a00000000",
            INIT_01 => X"0000005b0000000000000066000000000000000d000000000000004800000000",
            INIT_02 => X"ffffffeeffffffff000000380000000000000090000000000000005300000000",
            INIT_03 => X"ffffffe0ffffffffffffffd9ffffffff0000000700000000fffffff3ffffffff",
            INIT_04 => X"fffffff3ffffffffffffffcaffffffffffffffdefffffffffffffffcffffffff",
            INIT_05 => X"ffffffe7fffffffffffffffdfffffffffffffff1ffffffffffffffdbffffffff",
            INIT_06 => X"fffffffbfffffffffffffff4ffffffff0000001000000000fffffff0ffffffff",
            INIT_07 => X"ffffffedfffffffffffffffbfffffffffffffff9ffffffffffffffefffffffff",
            INIT_08 => X"ffffffecfffffffffffffffeffffffff0000000900000000ffffffd0ffffffff",
            INIT_09 => X"00000000000000000000001d00000000ffffffddffffffffffffffedffffffff",
            INIT_0A => X"fffffffefffffffffffffff9ffffffff0000002300000000ffffffe2ffffffff",
            INIT_0B => X"0000000800000000ffffffedfffffffffffffffefffffffffffffff6ffffffff",
            INIT_0C => X"ffffffd2ffffffff0000000f00000000ffffffcdffffffffffffffcaffffffff",
            INIT_0D => X"ffffffffffffffffffffffc8ffffffffffffffdaffffffffffffffcfffffffff",
            INIT_0E => X"000000180000000000000012000000000000003e000000000000000900000000",
            INIT_0F => X"ffffffe9fffffffffffffffefffffffffffffffbffffffff0000003b00000000",
            INIT_10 => X"00000007000000000000000000000000fffffffcffffffff0000000d00000000",
            INIT_11 => X"ffffffedffffffff0000000b000000000000000600000000ffffffebffffffff",
            INIT_12 => X"00000000000000000000003b0000000000000045000000000000000f00000000",
            INIT_13 => X"ffffffc6ffffffff00000001000000000000000b00000000ffffffe2ffffffff",
            INIT_14 => X"fffffff7ffffffffffffffd9ffffffffffffffdaffffffffffffffe7ffffffff",
            INIT_15 => X"ffffffffffffffffffffffe6ffffffffffffffffffffffff0000003a00000000",
            INIT_16 => X"ffffffdfffffffffffffffceffffffffffffffddffffffffffffffcaffffffff",
            INIT_17 => X"0000002500000000fffffff1ffffffff0000001200000000fffffff4ffffffff",
            INIT_18 => X"00000034000000000000002a0000000000000018000000000000004e00000000",
            INIT_19 => X"0000001300000000fffffff5ffffffff00000002000000000000003e00000000",
            INIT_1A => X"ffffffe3ffffffffffffffbfffffffff0000000600000000fffffff7ffffffff",
            INIT_1B => X"fffffffaffffffffffffffc6ffffffffffffffe3fffffffffffffff3ffffffff",
            INIT_1C => X"0000001000000000fffffff6ffffffffffffffdaffffffff0000000800000000",
            INIT_1D => X"000000370000000000000007000000000000001200000000fffffff0ffffffff",
            INIT_1E => X"0000000d000000000000001e00000000ffffffecffffffff0000000e00000000",
            INIT_1F => X"fffffff2ffffffff0000000a00000000fffffffcffffffffffffffdaffffffff",
            INIT_20 => X"00000012000000000000002400000000fffffffdfffffffffffffff8ffffffff",
            INIT_21 => X"fffffffeffffffffffffffe0ffffffff0000001b000000000000000400000000",
            INIT_22 => X"00000000000000000000000a000000000000001100000000fffffff5ffffffff",
            INIT_23 => X"0000000c000000000000002200000000fffffff0fffffffffffffffdffffffff",
            INIT_24 => X"ffffffbcffffffffffffffc4ffffffff00000016000000000000001700000000",
            INIT_25 => X"ffffffccffffffffffffffcfffffffffffffffd6ffffffffffffffdaffffffff",
            INIT_26 => X"ffffffc5ffffffffffffffeeffffffffffffffddfffffffffffffff8ffffffff",
            INIT_27 => X"0000002500000000ffffffa1ffffffff0000001c000000000000001200000000",
            INIT_28 => X"00000010000000000000001600000000fffffff0ffffffff0000000000000000",
            INIT_29 => X"ffffffa5ffffffffffffffe1ffffffffffffffa0ffffffffffffff76ffffffff",
            INIT_2A => X"ffffffc1ffffffff00000003000000000000000b00000000ffffff7bffffffff",
            INIT_2B => X"0000001f000000000000000d000000000000000f000000000000000100000000",
            INIT_2C => X"0000000100000000000000160000000000000028000000000000000000000000",
            INIT_2D => X"000000210000000000000004000000000000002c000000000000002200000000",
            INIT_2E => X"0000002500000000ffffffe8ffffffffffffffe2ffffffff0000001100000000",
            INIT_2F => X"0000003900000000fffffff7ffffffffffffffbeffffffffffffffaaffffffff",
            INIT_30 => X"00000029000000000000002800000000fffffff2ffffffff0000000600000000",
            INIT_31 => X"0000001e000000000000001a000000000000002000000000fffffff2ffffffff",
            INIT_32 => X"ffffffe8fffffffffffffff9ffffffffffffffe5ffffffff0000003700000000",
            INIT_33 => X"ffffffcfffffffffffffffdbffffffffffffffeeffffffffffffffdeffffffff",
            INIT_34 => X"00000028000000000000001c000000000000002700000000ffffffd6ffffffff",
            INIT_35 => X"ffffffe8ffffffff00000010000000000000002100000000ffffffedffffffff",
            INIT_36 => X"0000001a000000000000001200000000fffffffbfffffffffffffff9ffffffff",
            INIT_37 => X"0000000f00000000fffffff8ffffffff0000000000000000fffffff9ffffffff",
            INIT_38 => X"0000000d00000000ffffffd8ffffffffffffffe5ffffffff0000001a00000000",
            INIT_39 => X"0000001700000000ffffffd6ffffffff0000002d000000000000002c00000000",
            INIT_3A => X"0000000d000000000000001300000000ffffffe7ffffffff0000001500000000",
            INIT_3B => X"ffffffeaffffffff00000019000000000000000f000000000000001000000000",
            INIT_3C => X"0000000b00000000000000000000000000000011000000000000002000000000",
            INIT_3D => X"000000020000000000000010000000000000001b000000000000002000000000",
            INIT_3E => X"ffffffdffffffffffffffffcffffffff0000002300000000ffffffffffffffff",
            INIT_3F => X"0000002a00000000fffffff8ffffffff00000025000000000000000600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002000000000fffffffeffffffffffffffe8ffffffff0000002e00000000",
            INIT_41 => X"ffffffe0ffffffff0000000b00000000ffffffecffffffffffffffe3ffffffff",
            INIT_42 => X"0000000600000000ffffffe0ffffffff0000000f00000000fffffff2ffffffff",
            INIT_43 => X"00000023000000000000000c0000000000000012000000000000000300000000",
            INIT_44 => X"ffffffc9fffffffffffffff6ffffffffffffffdeffffffffffffffb6ffffffff",
            INIT_45 => X"0000003900000000ffffffc4ffffffffffffffdaffffffffffffffc3ffffffff",
            INIT_46 => X"00000038000000000000002800000000fffffffcffffffff0000000300000000",
            INIT_47 => X"ffffffc1ffffffff0000002300000000fffffff3fffffffffffffffdffffffff",
            INIT_48 => X"fffffff0ffffffff0000001c000000000000000500000000ffffffffffffffff",
            INIT_49 => X"0000001900000000ffffffd6fffffffffffffff7ffffffffffffffe7ffffffff",
            INIT_4A => X"ffffffe0ffffffffffffffeeffffffff0000001100000000fffffff7ffffffff",
            INIT_4B => X"ffffffe1ffffffff0000001600000000ffffffecffffffffffffffc3ffffffff",
            INIT_4C => X"0000000500000000fffffffbffffffff0000003300000000ffffffe7ffffffff",
            INIT_4D => X"0000003500000000ffffffdaffffffffffffffc7fffffffffffffff9ffffffff",
            INIT_4E => X"0000001c000000000000005900000000ffffffb7fffffffffffffffaffffffff",
            INIT_4F => X"ffffffe1ffffffffffffffe3ffffffffffffffeeffffffffffffffecffffffff",
            INIT_50 => X"0000003b00000000ffffffe8ffffffffffffffdfffffffff0000002200000000",
            INIT_51 => X"0000000200000000fffffffbffffffffffffffe3ffffffff0000000100000000",
            INIT_52 => X"fffffffaffffffff0000000d00000000fffffffdffffffff0000002700000000",
            INIT_53 => X"ffffffdfffffffff0000001900000000fffffff4ffffffffffffffd3ffffffff",
            INIT_54 => X"ffffffebffffffffffffffe0ffffffff0000001b00000000fffffff3ffffffff",
            INIT_55 => X"fffffff2ffffffffffffffe9ffffffffffffffe8ffffffff0000001600000000",
            INIT_56 => X"0000001600000000ffffffd5ffffffffffffffdfffffffffffffffc0ffffffff",
            INIT_57 => X"0000002a000000000000002300000000ffffffcfffffffff0000002a00000000",
            INIT_58 => X"ffffffe3ffffffff0000000300000000ffffffe4ffffffff0000000000000000",
            INIT_59 => X"0000003a00000000000000040000000000000012000000000000000600000000",
            INIT_5A => X"0000000c00000000ffffffebffffffff00000016000000000000001700000000",
            INIT_5B => X"00000013000000000000000c00000000ffffffc5ffffffff0000001600000000",
            INIT_5C => X"fffffff4ffffffff0000000800000000fffffff4ffffffffffffffb8ffffffff",
            INIT_5D => X"fffffff1fffffffffffffff2ffffffff0000000a00000000fffffff4ffffffff",
            INIT_5E => X"0000002500000000ffffffc7fffffffffffffff8ffffffff0000000e00000000",
            INIT_5F => X"ffffffa8fffffffffffffffeffffffffffffffe2fffffffffffffffeffffffff",
            INIT_60 => X"fffffffeffffffffffffffc1ffffffffffffffecfffffffffffffff3ffffffff",
            INIT_61 => X"00000027000000000000002000000000ffffffe5ffffffff0000001b00000000",
            INIT_62 => X"fffffffaffffffff000000090000000000000025000000000000000c00000000",
            INIT_63 => X"fffffff7ffffffff000000020000000000000000000000000000000d00000000",
            INIT_64 => X"ffffffdcfffffffffffffff0ffffffff0000002d00000000ffffffedffffffff",
            INIT_65 => X"fffffff0ffffffffffffffefffffffff00000016000000000000004d00000000",
            INIT_66 => X"0000000e00000000ffffffadffffffff00000026000000000000001300000000",
            INIT_67 => X"0000001c00000000fffffffdffffffffffffffd4ffffffff0000000d00000000",
            INIT_68 => X"00000012000000000000000400000000fffffff8ffffffff0000000000000000",
            INIT_69 => X"0000001200000000fffffffefffffffffffffffbffffffff0000000600000000",
            INIT_6A => X"fffffff9ffffffff0000000700000000fffffff2fffffffffffffff7ffffffff",
            INIT_6B => X"0000000500000000ffffffeafffffffffffffff9fffffffffffffff9ffffffff",
            INIT_6C => X"fffffff8fffffffffffffff1ffffffff0000000300000000ffffffeeffffffff",
            INIT_6D => X"fffffff0ffffffff0000000100000000fffffffefffffffffffffff6ffffffff",
            INIT_6E => X"fffffff4fffffffffffffff6ffffffff0000000b000000000000000600000000",
            INIT_6F => X"00000000000000000000000600000000ffffffffffffffff0000000000000000",
            INIT_70 => X"fffffff3ffffffff0000000500000000ffffffe8ffffffff0000000000000000",
            INIT_71 => X"fffffffeffffffff0000000d00000000ffffffffffffffff0000000600000000",
            INIT_72 => X"ffffffe9fffffffffffffff6ffffffff0000000e00000000fffffff2ffffffff",
            INIT_73 => X"fffffff6fffffffffffffff2ffffffff0000000600000000fffffffdffffffff",
            INIT_74 => X"ffffffefffffffffffffffeaffffffffffffffeaffffffff0000000700000000",
            INIT_75 => X"0000000a00000000fffffffcffffffff0000000600000000ffffffffffffffff",
            INIT_76 => X"fffffffaffffffff0000000c000000000000000c00000000fffffff1ffffffff",
            INIT_77 => X"fffffffafffffffffffffffbffffffffffffffe9fffffffffffffff5ffffffff",
            INIT_78 => X"0000000600000000fffffff2ffffffffffffffe7ffffffff0000000400000000",
            INIT_79 => X"000000000000000000000000000000000000000600000000fffffff4ffffffff",
            INIT_7A => X"ffffffefffffffff0000000b00000000fffffff9fffffffffffffffeffffffff",
            INIT_7B => X"ffffffe7ffffffff0000000900000000fffffff7ffffffff0000000200000000",
            INIT_7C => X"00000012000000000000000200000000fffffffbfffffffffffffff2ffffffff",
            INIT_7D => X"00000008000000000000000a00000000fffffff4ffffffffffffffecffffffff",
            INIT_7E => X"fffffff2ffffffffffffffedffffffff0000000000000000fffffff9ffffffff",
            INIT_7F => X"00000000000000000000000000000000fffffff1ffffffff0000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE28;


    MEM_IWGHT_LAYER2_INSTANCE29 : if BRAM_NAME = "iwght_layer2_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffecffffffff0000000d00000000ffffffe7ffffffff0000000e00000000",
            INIT_01 => X"0000000a000000000000000a00000000ffffffecffffffff0000000000000000",
            INIT_02 => X"ffffffedffffffff0000001000000000fffffffbffffffffffffffecffffffff",
            INIT_03 => X"0000000f00000000fffffff3fffffffffffffff5ffffffff0000000f00000000",
            INIT_04 => X"fffffff0ffffffff0000000d00000000fffffff4ffffffff0000000a00000000",
            INIT_05 => X"fffffff2fffffffffffffffffffffffffffffffbffffffff0000001100000000",
            INIT_06 => X"00000001000000000000000000000000ffffffeefffffffffffffffcffffffff",
            INIT_07 => X"0000000100000000fffffff8ffffffff0000000000000000ffffffe6ffffffff",
            INIT_08 => X"fffffff7ffffffffffffffeafffffffffffffff1fffffffffffffff0ffffffff",
            INIT_09 => X"0000000600000000fffffff8ffffffff0000000700000000fffffffdffffffff",
            INIT_0A => X"ffffffebfffffffffffffffbfffffffffffffff9fffffffffffffffdffffffff",
            INIT_0B => X"ffffffeeffffffffffffffefffffffffffffffefffffffffffffffedffffffff",
            INIT_0C => X"fffffffcfffffffffffffff8ffffffff0000000200000000fffffffdffffffff",
            INIT_0D => X"ffffffeffffffffffffffff1ffffffffffffffeefffffffffffffff4ffffffff",
            INIT_0E => X"0000000f00000000ffffffeaffffffff0000000b000000000000000900000000",
            INIT_0F => X"ffffffecfffffffffffffffbffffffff0000000e00000000fffffff2ffffffff",
            INIT_10 => X"00000007000000000000001200000000fffffff3ffffffffffffffebffffffff",
            INIT_11 => X"0000000900000000fffffff4ffffffff0000000d000000000000000f00000000",
            INIT_12 => X"ffffffe8fffffffffffffff9ffffffff00000001000000000000000d00000000",
            INIT_13 => X"00000000000000000000000600000000ffffffe9ffffffffffffffebffffffff",
            INIT_14 => X"0000000c000000000000000800000000ffffffe5ffffffffffffffe7ffffffff",
            INIT_15 => X"fffffff0fffffffffffffff3ffffffff0000000e00000000ffffffedffffffff",
            INIT_16 => X"0000000a00000000ffffffe7ffffffffffffffecfffffffffffffff3ffffffff",
            INIT_17 => X"fffffff8ffffffff00000005000000000000000600000000ffffffe9ffffffff",
            INIT_18 => X"0000000400000000fffffff9ffffffff0000000b000000000000000300000000",
            INIT_19 => X"ffffffecfffffffffffffff9ffffffff00000006000000000000000100000000",
            INIT_1A => X"ffffffeefffffffffffffff7fffffffffffffff6ffffffffffffffedffffffff",
            INIT_1B => X"00000005000000000000000100000000fffffff0ffffffff0000000d00000000",
            INIT_1C => X"0000000000000000ffffffeffffffffffffffff4ffffffffffffffecffffffff",
            INIT_1D => X"0000000600000000fffffffcffffffffffffffe9fffffffffffffff3ffffffff",
            INIT_1E => X"0000000a00000000fffffffcffffffff0000000500000000ffffffecffffffff",
            INIT_1F => X"ffffffeafffffffffffffffdffffffffffffffecffffffffffffffefffffffff",
            INIT_20 => X"fffffffdffffffffffffffe9fffffffffffffffdfffffffffffffffeffffffff",
            INIT_21 => X"0000000900000000fffffff8ffffffff0000000a00000000fffffff3ffffffff",
            INIT_22 => X"ffffffe7ffffffff00000001000000000000000000000000ffffffe2ffffffff",
            INIT_23 => X"ffffffeaffffffff0000000100000000fffffffeffffffff0000000700000000",
            INIT_24 => X"ffffffeefffffffffffffffbfffffffffffffff5fffffffffffffff4ffffffff",
            INIT_25 => X"0000000d000000000000000300000000fffffff0ffffffff0000000800000000",
            INIT_26 => X"0000000700000000ffffffeffffffffffffffffeffffffff0000000f00000000",
            INIT_27 => X"0000000e000000000000000c00000000fffffff0ffffffff0000000500000000",
            INIT_28 => X"fffffffbfffffffffffffff3ffffffffffffffedffffffff0000001500000000",
            INIT_29 => X"0000000b000000000000000c00000000fffffff0ffffffffffffffe4ffffffff",
            INIT_2A => X"0000000d0000000000000012000000000000000500000000fffffff1ffffffff",
            INIT_2B => X"ffffffedfffffffffffffffbfffffffffffffff4ffffffffffffffe9ffffffff",
            INIT_2C => X"ffffffebffffffffffffffe8ffffffff0000000b00000000fffffff0ffffffff",
            INIT_2D => X"fffffff0ffffffff0000000a000000000000000d000000000000000f00000000",
            INIT_2E => X"00000007000000000000000c0000000000000002000000000000000700000000",
            INIT_2F => X"0000000d000000000000000400000000fffffff3fffffffffffffffcffffffff",
            INIT_30 => X"0000001000000000ffffffeaffffffff0000000000000000fffffff0ffffffff",
            INIT_31 => X"00000015000000000000000c0000000000000004000000000000001100000000",
            INIT_32 => X"fffffff5ffffffffffffffe4fffffffffffffffdfffffffffffffff7ffffffff",
            INIT_33 => X"ffffffffffffffff0000000a00000000ffffffe6fffffffffffffffcffffffff",
            INIT_34 => X"00000032000000000000001d000000000000001900000000fffffffeffffffff",
            INIT_35 => X"fffffffbffffffff000000260000000000000005000000000000000b00000000",
            INIT_36 => X"ffffffdfffffffff000000020000000000000024000000000000001a00000000",
            INIT_37 => X"fffffff9ffffffff0000000000000000fffffffaffffffffffffffd5ffffffff",
            INIT_38 => X"fffffffaffffffff000000080000000000000014000000000000001100000000",
            INIT_39 => X"fffffffcfffffffffffffff9ffffffff0000001500000000fffffff3ffffffff",
            INIT_3A => X"0000000f00000000000000030000000000000013000000000000002d00000000",
            INIT_3B => X"0000000f00000000fffffffeffffffffffffffe6ffffffff0000000a00000000",
            INIT_3C => X"fffffff1fffffffffffffffdffffffff0000000100000000ffffffceffffffff",
            INIT_3D => X"ffffffe1fffffffffffffff7fffffffffffffff4ffffffffffffffc7ffffffff",
            INIT_3E => X"fffffffcffffffff00000002000000000000000400000000ffffffedffffffff",
            INIT_3F => X"fffffffdffffffffffffffcdffffffffffffffd3ffffffff0000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000013000000000000002b00000000ffffffe6fffffffffffffff5ffffffff",
            INIT_41 => X"ffffffe7ffffffff000000180000000000000025000000000000000500000000",
            INIT_42 => X"ffffffecffffffff0000000b0000000000000006000000000000000000000000",
            INIT_43 => X"0000000700000000000000050000000000000025000000000000000f00000000",
            INIT_44 => X"fffffffdffffffffffffffbfffffffffffffffe6fffffffffffffffbffffffff",
            INIT_45 => X"fffffffaffffffffffffffa2ffffffffffffffc2ffffffff0000000900000000",
            INIT_46 => X"00000018000000000000000700000000fffffff7fffffffffffffff3ffffffff",
            INIT_47 => X"0000001400000000fffffff8ffffffff0000000d000000000000001c00000000",
            INIT_48 => X"0000001f000000000000002d000000000000001400000000fffffff6ffffffff",
            INIT_49 => X"fffffffffffffffffffffff2fffffffffffffff2ffffffff0000000a00000000",
            INIT_4A => X"0000000000000000fffffff4ffffffffffffffdeffffffff0000000300000000",
            INIT_4B => X"00000004000000000000001a0000000000000016000000000000000100000000",
            INIT_4C => X"0000000c000000000000000f000000000000000b000000000000000100000000",
            INIT_4D => X"ffffffc6ffffffffffffffc3ffffffff0000000d000000000000000f00000000",
            INIT_4E => X"fffffff4ffffffffffffffc2ffffffffffffffc0ffffffff0000000f00000000",
            INIT_4F => X"0000000800000000ffffffe9ffffffff0000000400000000fffffff3ffffffff",
            INIT_50 => X"0000000600000000fffffffbffffffffffffffd8ffffffff0000000500000000",
            INIT_51 => X"0000000f000000000000000e00000000ffffffe9ffffffffffffffc5ffffffff",
            INIT_52 => X"00000005000000000000000b0000000000000000000000000000000600000000",
            INIT_53 => X"ffffffcafffffffffffffff4ffffffff0000003300000000fffffffaffffffff",
            INIT_54 => X"0000000000000000fffffffcffffffffffffffe0ffffffff0000001300000000",
            INIT_55 => X"ffffffb4ffffffffffffffe7ffffffffffffffafffffffffffffffc5ffffffff",
            INIT_56 => X"fffffff0fffffffffffffffafffffffffffffff1fffffffffffffff0ffffffff",
            INIT_57 => X"fffffffeffffffffffffffc6ffffffffffffffe3ffffffff0000002000000000",
            INIT_58 => X"0000003b000000000000002500000000ffffffcfffffffffffffffcaffffffff",
            INIT_59 => X"ffffffd2ffffffffffffffe4fffffffffffffff3ffffffff0000000000000000",
            INIT_5A => X"fffffff0ffffffffffffffc8ffffffffffffffc8fffffffffffffff7ffffffff",
            INIT_5B => X"0000000900000000ffffffdcffffffff0000001d000000000000000b00000000",
            INIT_5C => X"00000008000000000000000000000000ffffffeffffffffffffffffeffffffff",
            INIT_5D => X"fffffffaffffffff00000011000000000000000000000000ffffffd6ffffffff",
            INIT_5E => X"ffffffe9ffffffffffffffd7ffffffffffffffe5fffffffffffffffaffffffff",
            INIT_5F => X"0000000c000000000000001000000000fffffff0fffffffffffffff4ffffffff",
            INIT_60 => X"fffffff3ffffffff0000000600000000fffffffcffffffffffffffe4ffffffff",
            INIT_61 => X"0000000400000000ffffffeffffffffffffffffffffffffffffffff4ffffffff",
            INIT_62 => X"ffffffeeffffffffffffffdcffffffff0000000b00000000ffffffe5ffffffff",
            INIT_63 => X"0000000a00000000ffffffe8ffffffffffffffbcffffffff0000002900000000",
            INIT_64 => X"0000000b0000000000000004000000000000002600000000fffffffaffffffff",
            INIT_65 => X"fffffff8ffffffff0000000d00000000ffffffffffffffff0000001700000000",
            INIT_66 => X"0000004d0000000000000019000000000000001700000000fffffff6ffffffff",
            INIT_67 => X"0000005300000000000000340000000000000001000000000000001200000000",
            INIT_68 => X"0000000000000000ffffffe7ffffffff0000001000000000ffffffffffffffff",
            INIT_69 => X"0000000b000000000000000000000000ffffffffffffffff0000000e00000000",
            INIT_6A => X"ffffffe7fffffffffffffff3ffffffff0000002b00000000fffffff5ffffffff",
            INIT_6B => X"ffffffe9ffffffffffffffddffffffff0000003b00000000fffffff7ffffffff",
            INIT_6C => X"fffffff6ffffffffffffffe4ffffffffffffffe7ffffffff0000000e00000000",
            INIT_6D => X"fffffffaffffffff0000000600000000ffffffe6ffffffffffffffebffffffff",
            INIT_6E => X"ffffffd4ffffffffffffffedffffffffffffffefffffffff0000000c00000000",
            INIT_6F => X"ffffffffffffffffffffffecffffffffffffffd0ffffffffffffffe4ffffffff",
            INIT_70 => X"fffffffdffffffff0000001200000000fffffff0ffffffffffffffdbffffffff",
            INIT_71 => X"000000310000000000000020000000000000000900000000fffffff6ffffffff",
            INIT_72 => X"ffffffe8ffffffffffffffe2ffffffffffffffe3ffffffff0000001800000000",
            INIT_73 => X"0000001200000000ffffffd2fffffffffffffff0ffffffff0000000c00000000",
            INIT_74 => X"00000018000000000000000300000000fffffff1ffffffff0000002300000000",
            INIT_75 => X"000000290000000000000024000000000000001e00000000fffffff0ffffffff",
            INIT_76 => X"fffffff5ffffffff0000002800000000ffffffe3ffffffff0000000000000000",
            INIT_77 => X"ffffffc6fffffffffffffff5ffffffff0000001c00000000ffffffb8ffffffff",
            INIT_78 => X"000000080000000000000006000000000000000000000000ffffffffffffffff",
            INIT_79 => X"fffffffeffffffff0000000000000000fffffff3ffffffff0000000100000000",
            INIT_7A => X"0000001300000000000000060000000000000023000000000000000700000000",
            INIT_7B => X"ffffffdcffffffff000000290000000000000038000000000000000e00000000",
            INIT_7C => X"fffffffdfffffffffffffff8ffffffff00000010000000000000000700000000",
            INIT_7D => X"ffffffd9ffffffffffffffd1fffffffffffffffdffffffff0000001900000000",
            INIT_7E => X"ffffffb9ffffffffffffffafffffffffffffffbefffffffffffffff2ffffffff",
            INIT_7F => X"ffffff99ffffffffffffffb7ffffffffffffffd8ffffffffffffffd0ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE29;


    MEM_IWGHT_LAYER2_INSTANCE30 : if BRAM_NAME = "iwght_layer2_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffff9dffffffffffffff86ffffffffffffffafffffffffffffffc5ffffffff",
            INIT_01 => X"ffffffb7ffffffff00000026000000000000004600000000ffffffe7ffffffff",
            INIT_02 => X"ffffffc0fffffffffffffff5fffffffffffffffbffffffffffffffefffffffff",
            INIT_03 => X"000000130000000000000028000000000000003d000000000000000100000000",
            INIT_04 => X"0000003400000000000000230000000000000000000000000000000000000000",
            INIT_05 => X"fffffff6fffffffffffffffcffffffff00000023000000000000001000000000",
            INIT_06 => X"000000000000000000000005000000000000000300000000fffffffeffffffff",
            INIT_07 => X"fffffff8fffffffffffffffdffffffff0000000000000000fffffff8ffffffff",
            INIT_08 => X"0000001f000000000000001e000000000000000f000000000000001400000000",
            INIT_09 => X"0000001c000000000000000f0000000000000022000000000000002200000000",
            INIT_0A => X"ffffffdffffffffffffffffcffffffffffffffebffffffffffffffdcffffffff",
            INIT_0B => X"0000000a00000000fffffff0ffffffffffffffd0ffffffff0000001200000000",
            INIT_0C => X"ffffffedffffffffffffffebffffffff0000000a00000000ffffffefffffffff",
            INIT_0D => X"ffffffedffffffff0000000a00000000fffffffcfffffffffffffff3ffffffff",
            INIT_0E => X"fffffff1ffffffffffffffeafffffffffffffff9fffffffffffffff5ffffffff",
            INIT_0F => X"fffffff2ffffffffffffffecffffffff0000000a00000000ffffffe2ffffffff",
            INIT_10 => X"fffffff8ffffffff000000010000000000000008000000000000000c00000000",
            INIT_11 => X"0000000100000000fffffffdffffffff0000000100000000fffffffcffffffff",
            INIT_12 => X"fffffff3ffffffff000000020000000000000014000000000000000400000000",
            INIT_13 => X"fffffffbffffffff000000120000000000000000000000000000000b00000000",
            INIT_14 => X"00000014000000000000001b000000000000001500000000ffffffefffffffff",
            INIT_15 => X"000000090000000000000002000000000000000a000000000000001200000000",
            INIT_16 => X"0000000000000000000000370000000000000047000000000000001200000000",
            INIT_17 => X"0000001400000000000000250000000000000018000000000000001200000000",
            INIT_18 => X"0000001600000000000000150000000000000007000000000000003300000000",
            INIT_19 => X"00000010000000000000002a0000000000000027000000000000002100000000",
            INIT_1A => X"0000000300000000ffffffe5fffffffffffffff9ffffffff0000000c00000000",
            INIT_1B => X"00000014000000000000000500000000ffffffedfffffffffffffffcffffffff",
            INIT_1C => X"ffffffecffffffff00000018000000000000000c00000000ffffffd3ffffffff",
            INIT_1D => X"0000002400000000ffffffe6ffffffff00000010000000000000002800000000",
            INIT_1E => X"0000000500000000fffffffefffffffffffffffefffffffffffffff5ffffffff",
            INIT_1F => X"fffffffcffffffff00000005000000000000000e000000000000000900000000",
            INIT_20 => X"ffffffeaffffffff0000001800000000fffffffaffffffff0000001600000000",
            INIT_21 => X"ffffffecffffffffffffffceffffffff0000001400000000ffffffe7ffffffff",
            INIT_22 => X"fffffff7fffffffffffffff9ffffffff0000001d00000000fffffff9ffffffff",
            INIT_23 => X"ffffffecfffffffffffffff3ffffffff00000001000000000000000d00000000",
            INIT_24 => X"000000080000000000000013000000000000002600000000fffffffbffffffff",
            INIT_25 => X"fffffff2fffffffffffffff8ffffffffffffffffffffffffffffffe4ffffffff",
            INIT_26 => X"fffffff8ffffffff0000000000000000fffffff6ffffffffffffffedffffffff",
            INIT_27 => X"00000008000000000000000900000000fffffff9ffffffff0000001400000000",
            INIT_28 => X"fffffffffffffffffffffffbfffffffffffffff2fffffffffffffff1ffffffff",
            INIT_29 => X"fffffffefffffffffffffff9ffffffff0000001f00000000ffffffffffffffff",
            INIT_2A => X"ffffffe6ffffffff0000001b000000000000000e00000000ffffffe8ffffffff",
            INIT_2B => X"fffffffcfffffffffffffffcffffffff00000005000000000000000f00000000",
            INIT_2C => X"ffffffdcfffffffffffffff1fffffffffffffffdffffffffffffffe1ffffffff",
            INIT_2D => X"fffffff1ffffffff000000080000000000000019000000000000000500000000",
            INIT_2E => X"ffffff6dffffffffffffff95ffffffffffffffe1ffffffffffffff84ffffffff",
            INIT_2F => X"ffffffa3ffffffffffffffdeffffffffffffff94ffffffffffffff6effffffff",
            INIT_30 => X"0000001d0000000000000031000000000000000f00000000ffffff84ffffffff",
            INIT_31 => X"0000000e00000000000000340000000000000032000000000000000800000000",
            INIT_32 => X"0000001d00000000fffffffafffffffffffffff2fffffffffffffff8ffffffff",
            INIT_33 => X"00000012000000000000001100000000fffffff8ffffffff0000000100000000",
            INIT_34 => X"fffffffafffffffffffffff1ffffffff00000002000000000000000c00000000",
            INIT_35 => X"00000008000000000000001a00000000fffffff0ffffffffffffffeeffffffff",
            INIT_36 => X"00000029000000000000002d000000000000002b000000000000002400000000",
            INIT_37 => X"ffffffb5ffffffffffffffdcffffffffffffffe4ffffffffffffffd3ffffffff",
            INIT_38 => X"ffffffa1ffffffffffffffaaffffffffffffffa7ffffffffffffffa5ffffffff",
            INIT_39 => X"0000000d00000000fffffffbffffffff0000000000000000ffffffa9ffffffff",
            INIT_3A => X"0000003000000000000000110000000000000017000000000000000600000000",
            INIT_3B => X"ffffffe7ffffffffffffffe9ffffffff0000002e000000000000002700000000",
            INIT_3C => X"fffffffdfffffffffffffff1fffffffffffffff3ffffffffffffffecffffffff",
            INIT_3D => X"0000001c000000000000001c00000000ffffffffffffffff0000002300000000",
            INIT_3E => X"0000000c00000000ffffffebffffffff00000014000000000000001b00000000",
            INIT_3F => X"fffffff3fffffffffffffffafffffffffffffff0fffffffffffffffeffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000ffffffffffffffff00000018000000000000000900000000",
            INIT_41 => X"0000001500000000000000030000000000000015000000000000001700000000",
            INIT_42 => X"0000000900000000000000220000000000000015000000000000000e00000000",
            INIT_43 => X"ffffffe9ffffffff0000001500000000ffffffedffffffff0000000a00000000",
            INIT_44 => X"000000180000000000000019000000000000000e000000000000000200000000",
            INIT_45 => X"0000004800000000000000570000000000000027000000000000000800000000",
            INIT_46 => X"000000220000000000000049000000000000000b000000000000003500000000",
            INIT_47 => X"ffffffe6ffffffff00000015000000000000000e000000000000000100000000",
            INIT_48 => X"ffffffc7ffffffffffffffe4ffffffffffffffebffffffff0000000800000000",
            INIT_49 => X"0000002300000000ffffffedfffffffffffffff1ffffffff0000001800000000",
            INIT_4A => X"0000000c000000000000001a0000000000000040000000000000002900000000",
            INIT_4B => X"fffffff2ffffffffffffffe4ffffffffffffffe2ffffffff0000002c00000000",
            INIT_4C => X"0000003c0000000000000004000000000000001300000000fffffff6ffffffff",
            INIT_4D => X"00000032000000000000000a00000000fffffff9ffffffff0000002600000000",
            INIT_4E => X"fffffff2ffffffff0000000800000000fffffff1ffffffff0000001f00000000",
            INIT_4F => X"fffffff9ffffffffffffffd1ffffffffffffffc9ffffffffffffffd3ffffffff",
            INIT_50 => X"0000000400000000ffffffe4ffffffff0000000f00000000ffffffffffffffff",
            INIT_51 => X"0000001b00000000fffffff3ffffffffffffffe8ffffffffffffffebffffffff",
            INIT_52 => X"00000037000000000000000a000000000000002b000000000000003300000000",
            INIT_53 => X"0000000200000000000000170000000000000006000000000000002100000000",
            INIT_54 => X"fffffffdffffffff000000270000000000000008000000000000000600000000",
            INIT_55 => X"0000000100000000ffffffdfffffffff0000001d00000000fffffffbffffffff",
            INIT_56 => X"00000036000000000000001400000000ffffffd5ffffffff0000000400000000",
            INIT_57 => X"0000000900000000000000150000000000000006000000000000000900000000",
            INIT_58 => X"ffffffe1ffffffff0000001800000000fffffff7ffffffff0000001700000000",
            INIT_59 => X"00000004000000000000000a000000000000002100000000fffffff1ffffffff",
            INIT_5A => X"ffffffe6ffffffff0000000b0000000000000007000000000000002400000000",
            INIT_5B => X"ffffffd7ffffffff0000001600000000fffffffeffffffffffffffdbffffffff",
            INIT_5C => X"fffffff1ffffffffffffffeaffffffffffffffdcffffffffffffffe2ffffffff",
            INIT_5D => X"0000002c000000000000003800000000fffffffcffffffffffffffc9ffffffff",
            INIT_5E => X"ffffffe3ffffffffffffffe3ffffffff0000000600000000ffffffd1ffffffff",
            INIT_5F => X"ffffffe0ffffffffffffffe6ffffffff00000012000000000000001200000000",
            INIT_60 => X"0000000700000000fffffff6ffffffff0000001e00000000fffffff9ffffffff",
            INIT_61 => X"ffffffdaffffffff000000160000000000000006000000000000004300000000",
            INIT_62 => X"ffffffe5ffffffffffffffbeffffffff00000032000000000000000d00000000",
            INIT_63 => X"00000007000000000000000400000000ffffffceffffffff0000001400000000",
            INIT_64 => X"fffffffdffffffffffffffd1ffffffff0000003a000000000000001300000000",
            INIT_65 => X"fffffff4ffffffffffffffc7ffffffffffffff81fffffffffffffff0ffffffff",
            INIT_66 => X"0000003c0000000000000037000000000000001800000000ffffffdaffffffff",
            INIT_67 => X"0000000800000000fffffff0fffffffffffffff1ffffffff0000000300000000",
            INIT_68 => X"fffffff7ffffffffffffffe4ffffffffffffffc0ffffffffffffffdfffffffff",
            INIT_69 => X"fffffff7ffffffffffffffedffffffffffffffbffffffffffffffff3ffffffff",
            INIT_6A => X"fffffff1ffffffffffffffc9ffffffff0000000300000000ffffffd4ffffffff",
            INIT_6B => X"ffffffebffffffffffffffe2ffffffff0000000800000000fffffff0ffffffff",
            INIT_6C => X"fffffffdffffffffffffffe7ffffffff0000000f00000000fffffff3ffffffff",
            INIT_6D => X"ffffffd9ffffffff00000011000000000000000000000000ffffffffffffffff",
            INIT_6E => X"0000000900000000ffffffe0ffffffff00000021000000000000000600000000",
            INIT_6F => X"0000002d00000000fffffff7fffffffffffffff8ffffffff0000002c00000000",
            INIT_70 => X"fffffff3ffffffff0000002f000000000000001800000000ffffffedffffffff",
            INIT_71 => X"0000001900000000fffffff6ffffffff00000024000000000000000200000000",
            INIT_72 => X"00000009000000000000000900000000ffffffe8ffffffff0000002300000000",
            INIT_73 => X"0000001700000000ffffffc5ffffffffffffffe8fffffffffffffff7ffffffff",
            INIT_74 => X"0000000f000000000000000800000000ffffffe5ffffffff0000000b00000000",
            INIT_75 => X"fffffff1ffffffff000000060000000000000018000000000000000800000000",
            INIT_76 => X"ffffffd0ffffffffffffffd0ffffffffffffffb5fffffffffffffff7ffffffff",
            INIT_77 => X"ffffffd0fffffffffffffff5ffffffff0000001400000000ffffffb3ffffffff",
            INIT_78 => X"ffffffe6ffffffff00000015000000000000001100000000ffffffe0ffffffff",
            INIT_79 => X"fffffff3ffffffffffffffe3ffffffffffffffe8ffffffffffffffeaffffffff",
            INIT_7A => X"0000002e0000000000000003000000000000000c000000000000001100000000",
            INIT_7B => X"fffffff1fffffffffffffffcffffffffffffffeaffffffff0000000b00000000",
            INIT_7C => X"fffffff7ffffffff000000070000000000000013000000000000000400000000",
            INIT_7D => X"fffffff8ffffffffffffffd0ffffffff0000001b00000000fffffff0ffffffff",
            INIT_7E => X"fffffff2ffffffffffffffd1ffffffff0000001300000000ffffffc1ffffffff",
            INIT_7F => X"fffffff7ffffffff0000002d000000000000001d00000000fffffffeffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE30;


    MEM_IWGHT_LAYER2_INSTANCE31 : if BRAM_NAME = "iwght_layer2_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe8fffffffffffffffbffffffff00000016000000000000001500000000",
            INIT_01 => X"fffffffcffffffffffffffe2ffffffffffffffdcffffffff0000001100000000",
            INIT_02 => X"ffffffe5ffffffffffffffbaffffffffffffffeaffffffffffffffa8ffffffff",
            INIT_03 => X"fffffffbffffffff0000000100000000fffffff3fffffffffffffff4ffffffff",
            INIT_04 => X"0000002100000000fffffff6ffffffffffffffebffffffffffffffeeffffffff",
            INIT_05 => X"000000080000000000000013000000000000000900000000fffffff8ffffffff",
            INIT_06 => X"0000000300000000ffffffd7ffffffff00000020000000000000000600000000",
            INIT_07 => X"fffffffafffffffffffffff2ffffffffffffffcfffffffff0000000200000000",
            INIT_08 => X"00000000000000000000000000000000fffffff2fffffffffffffff7ffffffff",
            INIT_09 => X"0000000200000000fffffff6fffffffffffffffdffffffff0000001000000000",
            INIT_0A => X"0000000f0000000000000014000000000000002600000000fffffff8ffffffff",
            INIT_0B => X"0000001800000000fffffff4ffffffff00000023000000000000004900000000",
            INIT_0C => X"00000004000000000000000e0000000000000059000000000000003300000000",
            INIT_0D => X"fffffffaffffffffffffffedffffffff00000000000000000000002000000000",
            INIT_0E => X"0000001300000000ffffffe9ffffffffffffffbfffffffff0000000600000000",
            INIT_0F => X"000000320000000000000028000000000000001700000000fffffffbffffffff",
            INIT_10 => X"0000003400000000000000360000000000000011000000000000003f00000000",
            INIT_11 => X"ffffffc9ffffffff0000002d000000000000002a00000000fffffff0ffffffff",
            INIT_12 => X"ffffffe6ffffffffffffffe2fffffffffffffffefffffffffffffff3ffffffff",
            INIT_13 => X"00000013000000000000002000000000fffffffcffffffffffffffe5ffffffff",
            INIT_14 => X"ffffffd1ffffffff0000001a00000000ffffffdbffffffffffffffd8ffffffff",
            INIT_15 => X"0000001e00000000fffffff9ffffffff0000000000000000ffffffeaffffffff",
            INIT_16 => X"0000003e000000000000000600000000ffffffd0ffffffff0000001800000000",
            INIT_17 => X"fffffff9ffffffff0000001300000000fffffff1fffffffffffffffaffffffff",
            INIT_18 => X"000000380000000000000003000000000000003b000000000000002e00000000",
            INIT_19 => X"ffffffe2ffffffffffffffeafffffffffffffff9ffffffff0000002400000000",
            INIT_1A => X"fffffff7fffffffffffffff8ffffffffffffffd4ffffffff0000000400000000",
            INIT_1B => X"0000001f000000000000000a00000000ffffffecffffffff0000001300000000",
            INIT_1C => X"ffffffffffffffffffffffe3ffffffff0000000a000000000000002a00000000",
            INIT_1D => X"0000000500000000ffffffe2ffffffffffffffc7ffffffffffffffd9ffffffff",
            INIT_1E => X"fffffffcffffffffffffffefffffffffffffffedffffffffffffffdbffffffff",
            INIT_1F => X"0000001000000000fffffffaffffffffffffffd8ffffffffffffffefffffffff",
            INIT_20 => X"00000018000000000000003b000000000000001200000000ffffffe0ffffffff",
            INIT_21 => X"0000000c00000000ffffffcaffffffff00000020000000000000002d00000000",
            INIT_22 => X"0000001900000000ffffffe5ffffffffffffffbeffffffff0000001b00000000",
            INIT_23 => X"ffffffefffffffff0000001a0000000000000028000000000000002600000000",
            INIT_24 => X"0000000c00000000ffffffffffffffff00000004000000000000000b00000000",
            INIT_25 => X"000000020000000000000001000000000000000d000000000000000200000000",
            INIT_26 => X"0000002600000000ffffffd2ffffffffffffffe8ffffffff0000000900000000",
            INIT_27 => X"0000002500000000fffffff0fffffffffffffff0fffffffffffffff2ffffffff",
            INIT_28 => X"0000000600000000ffffffedffffffffffffff84ffffffff0000002100000000",
            INIT_29 => X"00000031000000000000001900000000fffffff0ffffffffffffff88ffffffff",
            INIT_2A => X"ffffffe7ffffffff0000001600000000fffffffdffffffff0000001d00000000",
            INIT_2B => X"ffffffe3fffffffffffffff9ffffffff0000001a00000000ffffffdcffffffff",
            INIT_2C => X"0000000800000000ffffffdcffffffffffffffeeffffffff0000000300000000",
            INIT_2D => X"0000001b00000000000000220000000000000028000000000000005000000000",
            INIT_2E => X"0000000500000000000000170000000000000029000000000000003e00000000",
            INIT_2F => X"ffffffe6ffffffff00000030000000000000000f000000000000000400000000",
            INIT_30 => X"fffffffbffffffffffffffe1ffffffff0000001b000000000000001300000000",
            INIT_31 => X"00000017000000000000002e0000000000000013000000000000001a00000000",
            INIT_32 => X"fffffffcffffffff00000010000000000000001b000000000000001400000000",
            INIT_33 => X"ffffffffffffffffffffffdcffffffff0000000c000000000000002600000000",
            INIT_34 => X"fffffff5ffffffff0000000f00000000ffffffd7ffffffff0000003800000000",
            INIT_35 => X"fffffff2fffffffffffffff6ffffffffffffffffffffffffffffffd9ffffffff",
            INIT_36 => X"fffffffbffffffffffffffd6ffffffff00000016000000000000002e00000000",
            INIT_37 => X"0000000f000000000000001c000000000000002a00000000fffffff6ffffffff",
            INIT_38 => X"ffffffe0ffffffff000000180000000000000025000000000000001a00000000",
            INIT_39 => X"fffffff2ffffffff0000001700000000fffffffeffffffffffffffedffffffff",
            INIT_3A => X"0000001700000000ffffffd7ffffffffffffffdfffffffff0000000800000000",
            INIT_3B => X"ffffffddffffffffffffffeffffffffffffffff1ffffffffffffffe6ffffffff",
            INIT_3C => X"0000001a00000000ffffffc3ffffffff0000000400000000fffffff6ffffffff",
            INIT_3D => X"0000000e000000000000002400000000ffffffdeffffffff0000001f00000000",
            INIT_3E => X"ffffffe5ffffffff0000001200000000ffffffdeffffffffffffffe8ffffffff",
            INIT_3F => X"ffffffecffffffff00000029000000000000000200000000ffffffd5ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffffffffffffffffffeaffffffffffffffe9ffffffffffffffe2ffffffff",
            INIT_41 => X"ffffffe3fffffffffffffff6fffffffffffffffdffffffffffffffe3ffffffff",
            INIT_42 => X"ffffffd0fffffffffffffffefffffffffffffffeffffffffffffffecffffffff",
            INIT_43 => X"ffffffc9ffffffffffffffd8ffffffff0000000400000000ffffffefffffffff",
            INIT_44 => X"0000000700000000fffffffbffffffff00000000000000000000002f00000000",
            INIT_45 => X"ffffffccffffffffffffffb3ffffffff00000022000000000000001600000000",
            INIT_46 => X"fffffff7ffffffffffffffe5ffffffff00000006000000000000002000000000",
            INIT_47 => X"ffffffffffffffff0000000500000000fffffff1ffffffff0000000200000000",
            INIT_48 => X"0000001900000000000000090000000000000026000000000000000800000000",
            INIT_49 => X"0000001800000000fffffff9ffffffff00000009000000000000001900000000",
            INIT_4A => X"00000026000000000000001100000000ffffffe4ffffffffffffffcdffffffff",
            INIT_4B => X"0000000000000000ffffffd9ffffffffffffffd6ffffffffffffffdaffffffff",
            INIT_4C => X"00000006000000000000001c00000000ffffffdcffffffff0000001600000000",
            INIT_4D => X"00000012000000000000000b000000000000000a00000000ffffffc3ffffffff",
            INIT_4E => X"fffffff8ffffffff00000029000000000000001700000000fffffff7ffffffff",
            INIT_4F => X"000000130000000000000006000000000000003300000000ffffffd7ffffffff",
            INIT_50 => X"0000000c00000000000000100000000000000003000000000000001400000000",
            INIT_51 => X"0000000e00000000fffffff9ffffffff0000000e000000000000002200000000",
            INIT_52 => X"0000000200000000000000000000000000000017000000000000000200000000",
            INIT_53 => X"ffffffe4ffffffffffffffdcffffffff0000001f00000000fffffff4ffffffff",
            INIT_54 => X"0000002e000000000000003d000000000000002200000000ffffffe2ffffffff",
            INIT_55 => X"fffffffcffffffff00000038000000000000001700000000fffffffbffffffff",
            INIT_56 => X"00000037000000000000000a00000000fffffff0fffffffffffffffcffffffff",
            INIT_57 => X"00000006000000000000003d00000000fffffff4ffffffff0000001d00000000",
            INIT_58 => X"ffffffd6ffffffff00000007000000000000004000000000ffffffe0ffffffff",
            INIT_59 => X"0000003c00000000ffffffe4ffffffffffffffe4fffffffffffffff1ffffffff",
            INIT_5A => X"ffffffcfffffffff0000004300000000ffffffbbffffffffffffffe9ffffffff",
            INIT_5B => X"00000017000000000000000000000000ffffffd8fffffffffffffffdffffffff",
            INIT_5C => X"000000380000000000000013000000000000000b000000000000001000000000",
            INIT_5D => X"0000000400000000000000000000000000000029000000000000000400000000",
            INIT_5E => X"0000001f00000000fffffff6ffffffffffffffedffffffff0000002c00000000",
            INIT_5F => X"ffffffd1ffffffff0000000900000000ffffffddffffffff0000001a00000000",
            INIT_60 => X"fffffff3ffffffffffffffbbffffffffffffffcaffffffffffffffe6ffffffff",
            INIT_61 => X"fffffffbffffffffffffffceffffffffffffffefffffffffffffffcfffffffff",
            INIT_62 => X"ffffffecffffffffffffffe9fffffffffffffff8ffffffff0000000f00000000",
            INIT_63 => X"ffffffd9ffffffff0000000200000000fffffff6ffffffff0000000a00000000",
            INIT_64 => X"00000006000000000000000000000000fffffff1ffffffffffffffe9ffffffff",
            INIT_65 => X"000000010000000000000015000000000000001a000000000000000b00000000",
            INIT_66 => X"00000007000000000000000c0000000000000013000000000000001c00000000",
            INIT_67 => X"0000000d000000000000001600000000ffffffe9ffffffff0000000a00000000",
            INIT_68 => X"fffffff3ffffffff0000000900000000ffffffe0ffffffffffffffcdffffffff",
            INIT_69 => X"000000030000000000000000000000000000001a000000000000000900000000",
            INIT_6A => X"00000001000000000000000a0000000000000017000000000000003700000000",
            INIT_6B => X"ffffffdbffffffff0000001200000000fffffffbffffffffffffffebffffffff",
            INIT_6C => X"0000000a0000000000000015000000000000000600000000ffffffebffffffff",
            INIT_6D => X"fffffffaffffffff00000003000000000000001f000000000000002a00000000",
            INIT_6E => X"0000002200000000fffffff9ffffffff0000000f00000000ffffffe6ffffffff",
            INIT_6F => X"ffffffe4ffffffffffffffc6fffffffffffffff3ffffffff0000000800000000",
            INIT_70 => X"00000004000000000000000500000000fffffff7ffffffff0000001800000000",
            INIT_71 => X"ffffffd9fffffffffffffff6ffffffff0000001700000000ffffffe9ffffffff",
            INIT_72 => X"0000000600000000ffffffe3fffffffffffffffcffffffffffffffe6ffffffff",
            INIT_73 => X"000000090000000000000020000000000000001300000000fffffffaffffffff",
            INIT_74 => X"0000000b00000000fffffff4ffffffff00000006000000000000000000000000",
            INIT_75 => X"ffffffebfffffffffffffffcfffffffffffffff9ffffffff0000002000000000",
            INIT_76 => X"0000002e000000000000000e00000000ffffffe1ffffffffffffffefffffffff",
            INIT_77 => X"0000000c000000000000002b000000000000001b000000000000000100000000",
            INIT_78 => X"0000002a000000000000004700000000fffffffeffffffff0000000d00000000",
            INIT_79 => X"0000002800000000000000060000000000000050000000000000001000000000",
            INIT_7A => X"ffffffdeffffffff00000054000000000000006b000000000000004b00000000",
            INIT_7B => X"ffffffd8ffffffffffffffc8ffffffffffffffe9ffffffffffffffdbffffffff",
            INIT_7C => X"fffffff1fffffffffffffff2ffffffffffffffc7ffffffffffffffe6ffffffff",
            INIT_7D => X"ffffffedffffffffffffffccffffffff0000001200000000fffffff9ffffffff",
            INIT_7E => X"fffffff7ffffffffffffffc3ffffffffffffffd3ffffffff0000000900000000",
            INIT_7F => X"ffffffceffffffffffffffd7ffffffff00000008000000000000000900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE31;


    MEM_IWGHT_LAYER2_INSTANCE32 : if BRAM_NAME = "iwght_layer2_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffe0ffffffffffffffd0fffffffffffffff0ffffffffffffffefffffffff",
            INIT_01 => X"fffffffeffffffff0000000700000000fffffffaffffffffffffffe8ffffffff",
            INIT_02 => X"0000001700000000ffffffecfffffffffffffff8ffffffff0000001600000000",
            INIT_03 => X"ffffffe4fffffffffffffff3ffffffff00000006000000000000001f00000000",
            INIT_04 => X"fffffffbffffffff000000180000000000000009000000000000000c00000000",
            INIT_05 => X"ffffffe3ffffffffffffffe9ffffffff00000015000000000000001000000000",
            INIT_06 => X"0000001c00000000ffffffe1ffffffffffffffe3ffffffffffffffebffffffff",
            INIT_07 => X"0000000500000000ffffffd7ffffffffffffffe5ffffffff0000003000000000",
            INIT_08 => X"fffffff6ffffffff00000002000000000000000e000000000000000b00000000",
            INIT_09 => X"fffffff3ffffffffffffffddffffffff0000002400000000fffffffeffffffff",
            INIT_0A => X"ffffffeeffffffffffffffecfffffffffffffff9ffffffffffffffd1ffffffff",
            INIT_0B => X"fffffffeffffffff00000016000000000000000d000000000000000300000000",
            INIT_0C => X"ffffffe2ffffffff0000000b0000000000000027000000000000003100000000",
            INIT_0D => X"0000000500000000ffffffe8ffffffff0000001300000000ffffffecffffffff",
            INIT_0E => X"0000001d000000000000001b00000000fffffff7ffffffffffffffe9ffffffff",
            INIT_0F => X"0000003300000000fffffffdffffffff00000023000000000000000e00000000",
            INIT_10 => X"0000001c000000000000000a00000000ffffffdbfffffffffffffff0ffffffff",
            INIT_11 => X"ffffffe9ffffffff0000000000000000ffffffeaffffffff0000000300000000",
            INIT_12 => X"0000002300000000000000220000000000000022000000000000000100000000",
            INIT_13 => X"ffffffd2fffffffffffffffaffffffff0000003c000000000000003700000000",
            INIT_14 => X"ffffffe0ffffffff0000000200000000ffffffceffffffffffffffc2ffffffff",
            INIT_15 => X"0000001800000000fffffff7ffffffffffffffd6ffffffffffffffc1ffffffff",
            INIT_16 => X"0000000000000000fffffffeffffffff00000009000000000000000000000000",
            INIT_17 => X"0000002000000000000000160000000000000041000000000000000400000000",
            INIT_18 => X"fffffff7ffffffffffffffecffffffff0000000d00000000fffffff9ffffffff",
            INIT_19 => X"0000001d00000000fffffff7ffffffff0000000a000000000000001000000000",
            INIT_1A => X"00000026000000000000001b000000000000000d000000000000001800000000",
            INIT_1B => X"000000130000000000000017000000000000001a000000000000001900000000",
            INIT_1C => X"ffffffeeffffffff000000420000000000000021000000000000001100000000",
            INIT_1D => X"ffffffa4ffffffff00000028000000000000002d00000000ffffffc2ffffffff",
            INIT_1E => X"0000000400000000fffffffdffffffffffffffffffffffff0000002800000000",
            INIT_1F => X"ffffffc0ffffffffffffffefffffffffffffffd0ffffffffffffffe2ffffffff",
            INIT_20 => X"ffffffaeffffffffffffffe6fffffffffffffff5ffffffffffffff8fffffffff",
            INIT_21 => X"0000003600000000ffffffbfffffffffffffffb6ffffffff0000003f00000000",
            INIT_22 => X"00000009000000000000005500000000ffffffbeffffffffffffffb7ffffffff",
            INIT_23 => X"0000001d00000000ffffffecfffffffffffffff7ffffffffffffffacffffffff",
            INIT_24 => X"ffffffeaffffffff000000090000000000000022000000000000000600000000",
            INIT_25 => X"00000020000000000000000a000000000000000000000000fffffff2ffffffff",
            INIT_26 => X"0000000a00000000ffffffffffffffff0000000600000000fffffff2ffffffff",
            INIT_27 => X"000000240000000000000013000000000000000e000000000000000700000000",
            INIT_28 => X"0000000900000000000000230000000000000035000000000000004000000000",
            INIT_29 => X"00000005000000000000001e0000000000000019000000000000000d00000000",
            INIT_2A => X"ffffffedffffffffffffffbcffffffffffffffeefffffffffffffff2ffffffff",
            INIT_2B => X"ffffffe4ffffffff0000000200000000ffffffcdffffffff0000000000000000",
            INIT_2C => X"ffffffe8ffffffff0000000800000000ffffffe8ffffffffffffffdcffffffff",
            INIT_2D => X"fffffff8fffffffffffffffcffffffff0000002700000000ffffffd4ffffffff",
            INIT_2E => X"ffffffeeffffffff0000000200000000fffffffbffffffff0000000300000000",
            INIT_2F => X"fffffffbffffffff00000030000000000000001e00000000ffffffe7ffffffff",
            INIT_30 => X"ffffffe7ffffffff00000012000000000000000e000000000000000b00000000",
            INIT_31 => X"ffffffe1ffffffffffffffffffffffffffffffe3fffffffffffffff9ffffffff",
            INIT_32 => X"00000011000000000000000100000000ffffffceffffffff0000000000000000",
            INIT_33 => X"ffffffecffffffff0000000f00000000fffffffbffffffff0000000000000000",
            INIT_34 => X"ffffffeaffffffffffffffc1ffffffff0000002c00000000fffffff5ffffffff",
            INIT_35 => X"0000000e000000000000003600000000ffffffe0ffffffff0000001300000000",
            INIT_36 => X"fffffffeffffffff0000002c000000000000003b000000000000000100000000",
            INIT_37 => X"0000000c00000000fffffff5ffffffff0000000c000000000000001200000000",
            INIT_38 => X"0000002800000000fffffffcffffffffffffffe1fffffffffffffffbffffffff",
            INIT_39 => X"0000000d00000000fffffffcffffffff0000000300000000ffffffe1ffffffff",
            INIT_3A => X"0000001a00000000ffffffecffffffff0000000a000000000000000e00000000",
            INIT_3B => X"fffffff7ffffffffffffffeaffffffffffffffc2ffffffff0000000b00000000",
            INIT_3C => X"0000001e0000000000000032000000000000002800000000ffffffceffffffff",
            INIT_3D => X"000000040000000000000003000000000000001e000000000000004200000000",
            INIT_3E => X"0000000e000000000000001000000000ffffffcdffffffff0000001500000000",
            INIT_3F => X"fffffff7ffffffff00000014000000000000002900000000fffffff8ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffd0ffffffffffffffeefffffffffffffff1ffffffff0000001800000000",
            INIT_41 => X"0000000b000000000000000b00000000fffffff8ffffffffffffff97ffffffff",
            INIT_42 => X"0000001b000000000000000a000000000000000900000000ffffffe5ffffffff",
            INIT_43 => X"0000001b00000000ffffffe8ffffffff00000014000000000000000300000000",
            INIT_44 => X"00000015000000000000000000000000ffffffe4ffffffff0000001c00000000",
            INIT_45 => X"0000000000000000000000040000000000000013000000000000000f00000000",
            INIT_46 => X"0000000000000000fffffff7ffffffff0000003a000000000000002500000000",
            INIT_47 => X"0000001300000000000000210000000000000013000000000000001e00000000",
            INIT_48 => X"ffffffe5ffffffff000000140000000000000006000000000000000200000000",
            INIT_49 => X"000000090000000000000022000000000000000600000000ffffffe3ffffffff",
            INIT_4A => X"fffffff0ffffffffffffffdafffffffffffffffeffffffffffffffebffffffff",
            INIT_4B => X"ffffffedffffffff00000002000000000000000b00000000ffffffdcffffffff",
            INIT_4C => X"fffffffefffffffffffffff4ffffffffffffffdbffffffffffffffd2ffffffff",
            INIT_4D => X"00000016000000000000000100000000ffffffe1ffffffff0000000200000000",
            INIT_4E => X"0000000300000000ffffffaeffffffffffffff99ffffffff0000002800000000",
            INIT_4F => X"ffffffc4ffffffff0000003800000000ffffff8cffffffffffffff9dffffffff",
            INIT_50 => X"000000020000000000000026000000000000001200000000ffffff77ffffffff",
            INIT_51 => X"fffffffdffffffff0000000e0000000000000002000000000000001c00000000",
            INIT_52 => X"0000000000000000ffffffedffffffff0000001f000000000000001500000000",
            INIT_53 => X"0000000e000000000000001600000000ffffffffffffffff0000000a00000000",
            INIT_54 => X"fffffffcffffffff0000000e0000000000000019000000000000001a00000000",
            INIT_55 => X"ffffffeaffffffffffffffd3ffffffff0000002500000000fffffff9ffffffff",
            INIT_56 => X"0000000000000000fffffff2ffffffff0000001b000000000000000300000000",
            INIT_57 => X"ffffffc6ffffffffffffffbcffffffffffffff91ffffffffffffffdbffffffff",
            INIT_58 => X"ffffffcdffffffff0000000600000000ffffffb1ffffffffffffff9cffffffff",
            INIT_59 => X"ffffffedffffffffffffffe2ffffffffffffffcfffffffffffffffb7ffffffff",
            INIT_5A => X"ffffffecfffffffffffffffcffffffff0000000a00000000ffffffc8ffffffff",
            INIT_5B => X"000000000000000000000010000000000000000300000000fffffffeffffffff",
            INIT_5C => X"00000016000000000000002b0000000000000002000000000000001100000000",
            INIT_5D => X"00000004000000000000001800000000fffffffeffffffffffffffeeffffffff",
            INIT_5E => X"00000010000000000000000600000000ffffffe5ffffffffffffffeaffffffff",
            INIT_5F => X"000000010000000000000007000000000000000e000000000000001c00000000",
            INIT_60 => X"fffffff3ffffffff0000000e000000000000001f000000000000000c00000000",
            INIT_61 => X"ffffffeeffffffff0000000900000000ffffffffffffffff0000000500000000",
            INIT_62 => X"fffffff2ffffffff00000031000000000000001800000000fffffff9ffffffff",
            INIT_63 => X"fffffff1fffffffffffffff8ffffffff00000025000000000000004700000000",
            INIT_64 => X"ffffffc2fffffffffffffff1ffffffff00000012000000000000001f00000000",
            INIT_65 => X"ffffffefffffffffffffffa6fffffffffffffff3ffffffffffffffe2ffffffff",
            INIT_66 => X"0000001700000000ffffffd9ffffffffffffffd6ffffffff0000001700000000",
            INIT_67 => X"0000003100000000000000410000000000000028000000000000003b00000000",
            INIT_68 => X"ffffffffffffffff000000280000000000000038000000000000003d00000000",
            INIT_69 => X"ffffffd9ffffffffffffffdcffffffffffffffa7ffffffffffffffc9ffffffff",
            INIT_6A => X"fffffff2fffffffffffffff0ffffffffffffffd9ffffffffffffffb3ffffffff",
            INIT_6B => X"fffffff2ffffffffffffffcdffffffffffffffbdffffffffffffffe7ffffffff",
            INIT_6C => X"0000002c00000000ffffffdaffffffffffffffb1fffffffffffffff3ffffffff",
            INIT_6D => X"0000001a00000000fffffff4ffffffffffffffdafffffffffffffffeffffffff",
            INIT_6E => X"0000002f000000000000003e000000000000003a000000000000004500000000",
            INIT_6F => X"0000001200000000ffffffddffffffff00000004000000000000000000000000",
            INIT_70 => X"fffffffbffffffff000000110000000000000007000000000000000c00000000",
            INIT_71 => X"0000001500000000ffffffecffffffffffffffd8ffffffff0000001500000000",
            INIT_72 => X"0000005200000000fffffff7ffffffff0000004800000000fffffffdffffffff",
            INIT_73 => X"00000018000000000000002d0000000000000013000000000000002200000000",
            INIT_74 => X"fffffff6ffffffffffffffdcffffffff0000000100000000fffffff3ffffffff",
            INIT_75 => X"fffffffbfffffffffffffff8ffffffff0000000100000000fffffff5ffffffff",
            INIT_76 => X"00000016000000000000000f0000000000000003000000000000001500000000",
            INIT_77 => X"00000011000000000000000c0000000000000021000000000000001e00000000",
            INIT_78 => X"ffffffd6ffffffff000000180000000000000014000000000000000d00000000",
            INIT_79 => X"ffffffbbffffffffffffffbbffffffffffffffbfffffffffffffff96ffffffff",
            INIT_7A => X"0000000f00000000fffffff8fffffffffffffffaffffffff0000000000000000",
            INIT_7B => X"0000001400000000fffffffffffffffffffffff7ffffffff0000001400000000",
            INIT_7C => X"ffffffedffffffffffffffefffffffff00000010000000000000000400000000",
            INIT_7D => X"ffffffd2ffffffff00000012000000000000000600000000fffffff1ffffffff",
            INIT_7E => X"ffffffabffffffffffffffe5ffffffff00000015000000000000002300000000",
            INIT_7F => X"ffffffbbffffffffffffffe3ffffffffffffffd3ffffffffffffffdbffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE32;


    MEM_IWGHT_LAYER2_INSTANCE33 : if BRAM_NAME = "iwght_layer2_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002200000000ffffffe0ffffffffffffffd7ffffffffffffffdeffffffff",
            INIT_01 => X"0000004100000000ffffffffffffffff00000013000000000000001200000000",
            INIT_02 => X"fffffff0ffffffff0000001a000000000000000400000000fffffff2ffffffff",
            INIT_03 => X"ffffffe6ffffffffffffffe6ffffffff0000002400000000fffffff1ffffffff",
            INIT_04 => X"fffffffaffffffff0000002c0000000000000005000000000000000900000000",
            INIT_05 => X"0000001b00000000ffffffe6ffffffffffffffdbffffffff0000000400000000",
            INIT_06 => X"0000001000000000000000220000000000000017000000000000001000000000",
            INIT_07 => X"0000000c00000000000000020000000000000011000000000000000700000000",
            INIT_08 => X"000000170000000000000023000000000000000f000000000000000900000000",
            INIT_09 => X"fffffffdffffffff00000011000000000000004600000000ffffffd7ffffffff",
            INIT_0A => X"fffffff4fffffffffffffff1fffffffffffffff7ffffffff0000001e00000000",
            INIT_0B => X"0000001200000000000000090000000000000026000000000000000a00000000",
            INIT_0C => X"0000001000000000fffffffaffffffff00000007000000000000000b00000000",
            INIT_0D => X"ffffffe5fffffffffffffff7fffffffffffffff1ffffffff0000000a00000000",
            INIT_0E => X"0000002e000000000000000200000000ffffffe9ffffffffffffffe8ffffffff",
            INIT_0F => X"00000020000000000000000300000000fffffffcffffffff0000003000000000",
            INIT_10 => X"0000002500000000000000110000000000000010000000000000000400000000",
            INIT_11 => X"0000001100000000fffffffdffffffff0000001a000000000000000d00000000",
            INIT_12 => X"0000000a0000000000000001000000000000000c000000000000001500000000",
            INIT_13 => X"fffffffefffffffffffffff6ffffffff00000003000000000000000100000000",
            INIT_14 => X"0000001e000000000000001f0000000000000018000000000000000200000000",
            INIT_15 => X"ffffffe0ffffffff0000001b000000000000000b000000000000002900000000",
            INIT_16 => X"0000002900000000000000270000000000000016000000000000001d00000000",
            INIT_17 => X"00000045000000000000003500000000fffffff5ffffffff0000001f00000000",
            INIT_18 => X"ffffffe5ffffffff0000001700000000ffffffebffffffff0000001c00000000",
            INIT_19 => X"ffffffd8ffffffffffffffefffffffffffffffeffffffffffffffff9ffffffff",
            INIT_1A => X"00000006000000000000000f000000000000002300000000ffffffffffffffff",
            INIT_1B => X"ffffffe8ffffffff0000000a000000000000001000000000ffffffebffffffff",
            INIT_1C => X"00000000000000000000000400000000fffffff8ffffffff0000001a00000000",
            INIT_1D => X"0000000700000000ffffffe4ffffffff0000000900000000fffffff9ffffffff",
            INIT_1E => X"fffffffcffffffffffffffe9fffffffffffffff3ffffffff0000002400000000",
            INIT_1F => X"00000024000000000000003c000000000000000a000000000000001d00000000",
            INIT_20 => X"00000011000000000000001400000000fffffffcfffffffffffffff1ffffffff",
            INIT_21 => X"ffffffceffffffffffffffc2ffffffffffffffedffffffffffffffe1ffffffff",
            INIT_22 => X"ffffffd7fffffffffffffff8ffffffffffffffb7ffffffffffffffd7ffffffff",
            INIT_23 => X"0000000600000000fffffff0ffffffffffffffddffffffffffffffc9ffffffff",
            INIT_24 => X"00000025000000000000000300000000ffffffdbffffffffffffffeeffffffff",
            INIT_25 => X"0000001d00000000fffffff9ffffffff0000002a000000000000000500000000",
            INIT_26 => X"0000001a0000000000000026000000000000001500000000fffffff7ffffffff",
            INIT_27 => X"0000002d000000000000001d000000000000004900000000fffffff9ffffffff",
            INIT_28 => X"0000000300000000000000170000000000000008000000000000000b00000000",
            INIT_29 => X"000000100000000000000018000000000000000f00000000fffffff1ffffffff",
            INIT_2A => X"ffffffe2ffffffff00000006000000000000001400000000fffffff8ffffffff",
            INIT_2B => X"0000002d000000000000000e000000000000001c000000000000002500000000",
            INIT_2C => X"0000000c00000000000000030000000000000019000000000000002a00000000",
            INIT_2D => X"00000000000000000000000900000000ffffffeaffffffffffffffd9ffffffff",
            INIT_2E => X"ffffffe9ffffffffffffffe6ffffffff0000000c00000000ffffffe4ffffffff",
            INIT_2F => X"ffffffecffffffffffffffe4ffffffffffffffafffffffffffffffc3ffffffff",
            INIT_30 => X"ffffffbdffffffffffffffbbffffffffffffffc6ffffffffffffffbeffffffff",
            INIT_31 => X"00000002000000000000000a000000000000002a000000000000004f00000000",
            INIT_32 => X"0000001200000000ffffffe5ffffffff0000000a000000000000003e00000000",
            INIT_33 => X"fffffffffffffffffffffff3fffffffffffffff6ffffffff0000000600000000",
            INIT_34 => X"fffffff0ffffffff00000014000000000000002100000000fffffff9ffffffff",
            INIT_35 => X"00000014000000000000001800000000ffffffeeffffffff0000000800000000",
            INIT_36 => X"fffffff1fffffffffffffff2fffffffffffffffbffffffff0000000d00000000",
            INIT_37 => X"0000001700000000fffffff9ffffffffffffffceffffffffffffffc6ffffffff",
            INIT_38 => X"fffffff2ffffffff0000000c0000000000000011000000000000000100000000",
            INIT_39 => X"00000029000000000000000b0000000000000004000000000000000000000000",
            INIT_3A => X"0000000500000000000000050000000000000005000000000000000300000000",
            INIT_3B => X"000000000000000000000008000000000000001c00000000fffffffaffffffff",
            INIT_3C => X"0000001c000000000000002c0000000000000028000000000000001100000000",
            INIT_3D => X"ffffff92ffffffff00000002000000000000001c000000000000001600000000",
            INIT_3E => X"0000001b000000000000001500000000ffffffc6ffffffffffffffb7ffffffff",
            INIT_3F => X"0000002a00000000000000080000000000000020000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000100000000ffffffefffffffff00000006000000000000000400000000",
            INIT_41 => X"fffffff2ffffffff0000000900000000ffffffcaffffffffffffffd4ffffffff",
            INIT_42 => X"ffffffb9ffffffffffffffd8ffffffffffffffefffffffffffffffc9ffffffff",
            INIT_43 => X"0000001300000000fffffff5fffffffffffffff6fffffffffffffff4ffffffff",
            INIT_44 => X"ffffffe3ffffffffffffffedfffffffffffffffdfffffffffffffffeffffffff",
            INIT_45 => X"000000100000000000000016000000000000000f000000000000000300000000",
            INIT_46 => X"fffffffbffffffffffffffe5ffffffff00000000000000000000000500000000",
            INIT_47 => X"fffffffcffffffffffffffe7ffffffffffffffe4fffffffffffffffeffffffff",
            INIT_48 => X"fffffff7ffffffff0000000d0000000000000008000000000000000000000000",
            INIT_49 => X"0000000c00000000ffffffeaffffffffffffffe5fffffffffffffffbffffffff",
            INIT_4A => X"00000015000000000000001f00000000ffffffd5ffffffff0000001600000000",
            INIT_4B => X"ffffffd5fffffffffffffff5fffffffffffffffeffffffffffffffffffffffff",
            INIT_4C => X"ffffffbffffffffffffffffeffffffffffffffe0ffffffffffffffd4ffffffff",
            INIT_4D => X"ffffff8effffffffffffffc2ffffffffffffffabffffffffffffffbbffffffff",
            INIT_4E => X"0000001d0000000000000022000000000000001900000000ffffffabffffffff",
            INIT_4F => X"ffffffb6ffffffff0000000000000000fffffff0ffffffff0000000f00000000",
            INIT_50 => X"0000003f000000000000003100000000ffffffc3ffffffffffffffb8ffffffff",
            INIT_51 => X"ffffffeefffffffffffffffbffffffff0000004000000000ffffffefffffffff",
            INIT_52 => X"fffffff6ffffffff0000000a000000000000002e000000000000001c00000000",
            INIT_53 => X"000000160000000000000013000000000000000100000000fffffffeffffffff",
            INIT_54 => X"00000010000000000000002900000000fffffffcffffffff0000000100000000",
            INIT_55 => X"0000002e00000000fffffff4ffffffff00000002000000000000000100000000",
            INIT_56 => X"0000000d00000000000000380000000000000001000000000000002200000000",
            INIT_57 => X"00000005000000000000000a0000000000000007000000000000002400000000",
            INIT_58 => X"0000001e0000000000000018000000000000001f000000000000001200000000",
            INIT_59 => X"0000003d00000000ffffffe9ffffffff0000002a000000000000000500000000",
            INIT_5A => X"ffffffe0ffffffffffffffffffffffffffffffedffffffff0000001900000000",
            INIT_5B => X"fffffff5ffffffffffffff9cffffffffffffffcbffffffffffffff80ffffffff",
            INIT_5C => X"fffffffbffffffffffffffebffffffff0000001000000000ffffffffffffffff",
            INIT_5D => X"0000001a00000000ffffffd1ffffffffffffffd8ffffffff0000001200000000",
            INIT_5E => X"ffffffceffffffffffffffebffffffffffffffd1ffffffffffffffe1ffffffff",
            INIT_5F => X"ffffffd0ffffffffffffff9affffffffffffffb9ffffffffffffffbbffffffff",
            INIT_60 => X"000000230000000000000027000000000000001900000000ffffffc2ffffffff",
            INIT_61 => X"0000001800000000000000170000000000000012000000000000002300000000",
            INIT_62 => X"000000460000000000000044000000000000000e00000000fffffffdffffffff",
            INIT_63 => X"fffffffcfffffffffffffff3ffffffff0000001e000000000000001e00000000",
            INIT_64 => X"fffffffaffffffffffffffd7ffffffffffffffe9ffffffffffffffccffffffff",
            INIT_65 => X"ffffffd3ffffffffffffffd3fffffffffffffffeffffffffffffffe3ffffffff",
            INIT_66 => X"ffffffd1ffffffffffffffd7ffffffffffffffebfffffffffffffffaffffffff",
            INIT_67 => X"ffffffedffffffffffffffd6ffffffffffffffccffffffff0000001a00000000",
            INIT_68 => X"ffffffbbffffffffffffffedffffffffffffffefffffffffffffffedffffffff",
            INIT_69 => X"0000002100000000ffffffccffffffffffffffdaffffffffffffffebffffffff",
            INIT_6A => X"ffffffd3ffffffffffffffa6ffffffffffffff7bffffffffffffffa5ffffffff",
            INIT_6B => X"00000017000000000000000a00000000ffffffb1ffffffffffffff90ffffffff",
            INIT_6C => X"00000008000000000000000d0000000000000023000000000000000000000000",
            INIT_6D => X"0000001600000000000000090000000000000025000000000000001800000000",
            INIT_6E => X"0000000400000000fffffff5ffffffff00000004000000000000003d00000000",
            INIT_6F => X"ffffffb9ffffffffffffffe6ffffffffffffffbfffffffff0000002900000000",
            INIT_70 => X"0000001000000000fffffff4ffffffff00000004000000000000000d00000000",
            INIT_71 => X"0000000600000000fffffffdffffffffffffffefffffffff0000001400000000",
            INIT_72 => X"00000000000000000000000b0000000000000010000000000000000c00000000",
            INIT_73 => X"0000000600000000ffffffe4ffffffff00000003000000000000000900000000",
            INIT_74 => X"0000001100000000000000030000000000000024000000000000001800000000",
            INIT_75 => X"000000100000000000000010000000000000000f00000000fffffffeffffffff",
            INIT_76 => X"ffffffc5ffffffff00000020000000000000001d000000000000001100000000",
            INIT_77 => X"ffffffeaffffffffffffffb2ffffffffffffffefffffffffffffffe0ffffffff",
            INIT_78 => X"ffffffeaffffffffffffffe2ffffffffffffffcfffffffffffffffdeffffffff",
            INIT_79 => X"0000002200000000fffffff4fffffffffffffff6ffffffff0000000600000000",
            INIT_7A => X"0000004800000000000000010000000000000018000000000000002b00000000",
            INIT_7B => X"0000000f00000000ffffffdcffffffff00000004000000000000002d00000000",
            INIT_7C => X"0000000800000000fffffff8fffffffffffffffaffffffff0000001300000000",
            INIT_7D => X"fffffff4ffffffff0000001d00000000ffffffe5ffffffff0000001800000000",
            INIT_7E => X"ffffffe0fffffffffffffff4fffffffffffffffefffffffffffffffaffffffff",
            INIT_7F => X"ffffffecffffffffffffffeffffffffffffffff2fffffffffffffff6ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE33;


    MEM_IWGHT_LAYER2_INSTANCE34 : if BRAM_NAME = "iwght_layer2_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffffffffffff0000000400000000ffffffedfffffffffffffff3ffffffff",
            INIT_01 => X"0000002d000000000000002b0000000000000007000000000000000b00000000",
            INIT_02 => X"000000470000000000000008000000000000001a000000000000000c00000000",
            INIT_03 => X"fffffffcffffffff0000001500000000ffffffddffffffff0000001e00000000",
            INIT_04 => X"0000000800000000fffffffbffffffff00000016000000000000000c00000000",
            INIT_05 => X"ffffffdcffffffff0000002100000000ffffffefffffffffffffffdfffffffff",
            INIT_06 => X"0000001800000000fffffffeffffffff0000001c00000000ffffffd8ffffffff",
            INIT_07 => X"ffffffedffffffffffffffedffffffff0000000f00000000fffffff9ffffffff",
            INIT_08 => X"ffffffe7fffffffffffffffaffffffffffffffedffffffff0000002b00000000",
            INIT_09 => X"ffffffcfffffffffffffffd5ffffffffffffffe1ffffffffffffffe8ffffffff",
            INIT_0A => X"ffffffcdffffffffffffffe1ffffffffffffffd1fffffffffffffff0ffffffff",
            INIT_0B => X"fffffff9ffffffff0000000900000000fffffff4ffffffff0000000400000000",
            INIT_0C => X"fffffffaffffffff0000000d000000000000000900000000fffffffeffffffff",
            INIT_0D => X"000000000000000000000015000000000000000700000000ffffffeaffffffff",
            INIT_0E => X"ffffffebffffffff00000034000000000000001e000000000000000200000000",
            INIT_0F => X"ffffffeefffffffffffffff7ffffffff00000019000000000000002000000000",
            INIT_10 => X"ffffffeffffffffffffffffaffffffff0000000c00000000ffffffe6ffffffff",
            INIT_11 => X"0000000400000000ffffffccffffffff00000000000000000000001a00000000",
            INIT_12 => X"0000002b000000000000001b0000000000000000000000000000001e00000000",
            INIT_13 => X"0000001d000000000000000400000000ffffffedffffffff0000001300000000",
            INIT_14 => X"ffffffe0ffffffffffffffbeffffffffffffffd3ffffffffffffffafffffffff",
            INIT_15 => X"ffffff97ffffffffffffffb9fffffffffffffff3ffffffffffffffcaffffffff",
            INIT_16 => X"00000006000000000000000100000000fffffff4ffffffffffffffa8ffffffff",
            INIT_17 => X"fffffff0ffffffffffffffdaffffffffffffffdbffffffffffffffe5ffffffff",
            INIT_18 => X"0000000600000000fffffffcffffffffffffffdeffffffffffffffd8ffffffff",
            INIT_19 => X"ffffffdaffffffffffffffd0ffffffffffffffc6ffffffff0000002300000000",
            INIT_1A => X"0000001a00000000ffffffebffffffffffffffdfffffffffffffff8dffffffff",
            INIT_1B => X"0000001d000000000000001d0000000000000013000000000000001b00000000",
            INIT_1C => X"00000023000000000000002e000000000000001000000000fffffffcffffffff",
            INIT_1D => X"0000001a00000000fffffffaffffffff0000000a000000000000000b00000000",
            INIT_1E => X"ffffffeeffffffff000000040000000000000022000000000000001200000000",
            INIT_1F => X"fffffff8ffffffff00000000000000000000001d000000000000002100000000",
            INIT_20 => X"0000001900000000000000000000000000000010000000000000000800000000",
            INIT_21 => X"ffffffe5ffffffffffffffceffffffff0000000a000000000000000800000000",
            INIT_22 => X"ffffffb2ffffffffffffffe3ffffffffffffffcbffffffffffffffecffffffff",
            INIT_23 => X"0000000600000000ffffffd0ffffffffffffffc3ffffffffffffffc8ffffffff",
            INIT_24 => X"fffffff4ffffffff000000160000000000000022000000000000001300000000",
            INIT_25 => X"fffffff8fffffffffffffff3ffffffff0000000600000000ffffffeaffffffff",
            INIT_26 => X"ffffffceffffffffffffffdafffffffffffffff5ffffffffffffffcfffffffff",
            INIT_27 => X"ffffffddffffffff0000000600000000ffffffaeffffffffffffffd7ffffffff",
            INIT_28 => X"0000002c0000000000000010000000000000000d00000000ffffffd9ffffffff",
            INIT_29 => X"0000001d000000000000000f0000000000000016000000000000001b00000000",
            INIT_2A => X"fffffffcffffffff00000007000000000000001b000000000000001400000000",
            INIT_2B => X"00000009000000000000000f00000000fffffff7ffffffff0000001b00000000",
            INIT_2C => X"00000008000000000000001200000000ffffffe5ffffffffffffffd6ffffffff",
            INIT_2D => X"000000000000000000000015000000000000000900000000ffffffe8ffffffff",
            INIT_2E => X"0000000600000000000000000000000000000001000000000000000300000000",
            INIT_2F => X"ffffffe4ffffffff00000013000000000000000200000000fffffff9ffffffff",
            INIT_30 => X"0000000000000000fffffff8fffffffffffffffdfffffffffffffff1ffffffff",
            INIT_31 => X"0000002b000000000000001b000000000000000000000000ffffffd8ffffffff",
            INIT_32 => X"ffffffe2ffffffffffffffdaffffffffffffffc5ffffffffffffffdeffffffff",
            INIT_33 => X"fffffffeffffffff0000000200000000ffffffddffffffffffffffceffffffff",
            INIT_34 => X"0000000a00000000000000040000000000000003000000000000001600000000",
            INIT_35 => X"0000001200000000fffffffbffffffffffffffedffffffff0000000100000000",
            INIT_36 => X"0000000900000000ffffffe9ffffffff00000001000000000000000f00000000",
            INIT_37 => X"ffffffecffffffffffffffdeffffffffffffffcafffffffffffffffeffffffff",
            INIT_38 => X"fffffff7ffffffff00000005000000000000000e000000000000000800000000",
            INIT_39 => X"00000000000000000000000000000000fffffff9ffffffffffffffecffffffff",
            INIT_3A => X"ffffffdfffffffffffffffebffffffff0000001b00000000ffffffefffffffff",
            INIT_3B => X"ffffffbfffffffff0000001f000000000000002100000000ffffffdfffffffff",
            INIT_3C => X"fffffffbffffffff0000001900000000ffffffebffffffffffffffcfffffffff",
            INIT_3D => X"000000190000000000000010000000000000000c000000000000000000000000",
            INIT_3E => X"ffffffe6ffffffffffffffbbfffffffffffffff8ffffffffffffffd6ffffffff",
            INIT_3F => X"fffffffbffffffff0000000200000000ffffffffffffffffffffffe3ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000fffffffbffffffffffffffe5ffffffff0000002000000000",
            INIT_41 => X"fffffff8fffffffffffffff3fffffffffffffff0fffffffffffffff4ffffffff",
            INIT_42 => X"ffffffd6ffffffff0000000d00000000ffffffe1fffffffffffffffaffffffff",
            INIT_43 => X"fffffffaffffffffffffffcfffffffffffffffdafffffffffffffff4ffffffff",
            INIT_44 => X"0000002900000000fffffffdffffffffffffffcdffffffff0000000600000000",
            INIT_45 => X"0000000200000000ffffffeefffffffffffffff2ffffffff0000000b00000000",
            INIT_46 => X"ffffffc6ffffffff0000001f000000000000000d000000000000000b00000000",
            INIT_47 => X"0000000000000000fffffff1fffffffffffffffaffffffff0000000700000000",
            INIT_48 => X"0000001000000000ffffffe4ffffffff0000001f000000000000001f00000000",
            INIT_49 => X"0000003700000000fffffffbfffffffffffffff7ffffffff0000002a00000000",
            INIT_4A => X"fffffff3ffffffff00000008000000000000001100000000ffffffd9ffffffff",
            INIT_4B => X"ffffffe2ffffffffffffffd5ffffffff0000000000000000fffffffeffffffff",
            INIT_4C => X"ffffffc0fffffffffffffff1ffffffff0000001600000000ffffffedffffffff",
            INIT_4D => X"0000002a00000000ffffffc7ffffffffffffffe9ffffffff0000001500000000",
            INIT_4E => X"0000004400000000fffffff8fffffffffffffff7fffffffffffffff0ffffffff",
            INIT_4F => X"0000004e000000000000000300000000ffffffd9ffffffff0000002c00000000",
            INIT_50 => X"0000000e00000000ffffffdcfffffffffffffff8ffffffffffffffb6ffffffff",
            INIT_51 => X"000000070000000000000027000000000000000f000000000000000500000000",
            INIT_52 => X"ffffffebffffffff000000120000000000000029000000000000004700000000",
            INIT_53 => X"0000002300000000ffffffefffffffffffffffdbffffffff0000001c00000000",
            INIT_54 => X"00000025000000000000003600000000ffffffdbfffffffffffffff3ffffffff",
            INIT_55 => X"ffffffe6ffffffff00000019000000000000000f000000000000000c00000000",
            INIT_56 => X"fffffffbffffffff00000005000000000000000b00000000ffffffd4ffffffff",
            INIT_57 => X"fffffff7ffffffffffffffcfffffffff0000001300000000fffffff6ffffffff",
            INIT_58 => X"fffffff9ffffffffffffffdaffffffffffffffffffffffff0000001600000000",
            INIT_59 => X"0000003a00000000000000030000000000000027000000000000002f00000000",
            INIT_5A => X"ffffffe7ffffffff0000003c00000000ffffffdcffffffffffffffd0ffffffff",
            INIT_5B => X"0000000600000000fffffffcffffffff0000004000000000ffffffd8ffffffff",
            INIT_5C => X"ffffffd0ffffffffffffffe0ffffffff0000001c00000000fffffff4ffffffff",
            INIT_5D => X"ffffffecffffffffffffffbefffffffffffffff9ffffffff0000002a00000000",
            INIT_5E => X"ffffffeeffffffffffffffeffffffffffffffff5ffffffff0000002300000000",
            INIT_5F => X"0000001500000000ffffffd6ffffffff0000001a00000000ffffffe7ffffffff",
            INIT_60 => X"0000000600000000000000310000000000000008000000000000003200000000",
            INIT_61 => X"ffffffccffffffff0000000700000000fffffffdfffffffffffffffeffffffff",
            INIT_62 => X"fffffff4ffffffff0000000200000000fffffff8ffffffff0000002a00000000",
            INIT_63 => X"ffffffeefffffffffffffff0ffffffff0000000b00000000ffffffd7ffffffff",
            INIT_64 => X"ffffffedffffffff0000000100000000fffffff2fffffffffffffffeffffffff",
            INIT_65 => X"00000015000000000000001600000000fffffff8ffffffffffffffddffffffff",
            INIT_66 => X"0000000300000000ffffffebffffffff00000004000000000000000200000000",
            INIT_67 => X"0000002000000000ffffffefffffffffffffffe2ffffffff0000002700000000",
            INIT_68 => X"00000010000000000000001d00000000ffffffe0ffffffffffffffefffffffff",
            INIT_69 => X"ffffffe2fffffffffffffffafffffffffffffffdfffffffffffffff8ffffffff",
            INIT_6A => X"ffffffc0ffffffffffffffe8ffffffff0000000600000000ffffffbeffffffff",
            INIT_6B => X"ffffffe3fffffffffffffff7ffffffff00000019000000000000002200000000",
            INIT_6C => X"ffffffedffffffffffffffc1ffffffff00000040000000000000001900000000",
            INIT_6D => X"0000001100000000fffffff5ffffffffffffffeeffffffff0000005500000000",
            INIT_6E => X"00000050000000000000001b000000000000002e000000000000004200000000",
            INIT_6F => X"0000001e0000000000000006000000000000005e000000000000005200000000",
            INIT_70 => X"ffffffe1ffffffff0000001b00000000ffffffe2ffffffff0000002300000000",
            INIT_71 => X"ffffffc8ffffffff00000016000000000000001300000000ffffffdaffffffff",
            INIT_72 => X"00000001000000000000001a0000000000000028000000000000000300000000",
            INIT_73 => X"ffffffceffffffffffffffedffffffff0000000d00000000ffffffdeffffffff",
            INIT_74 => X"0000000000000000fffffff7ffffffff0000001c000000000000002d00000000",
            INIT_75 => X"ffffffeafffffffffffffff5fffffffffffffffdffffffffffffffe3ffffffff",
            INIT_76 => X"0000001d000000000000001c000000000000000a00000000ffffffe3ffffffff",
            INIT_77 => X"0000001e00000000000000050000000000000027000000000000001700000000",
            INIT_78 => X"0000001200000000000000180000000000000021000000000000001f00000000",
            INIT_79 => X"ffffffe6ffffffff000000080000000000000005000000000000001d00000000",
            INIT_7A => X"000000170000000000000032000000000000003e000000000000002900000000",
            INIT_7B => X"ffffffc3ffffffffffffffcaffffffff00000050000000000000003b00000000",
            INIT_7C => X"fffffffaffffffffffffffd3ffffffffffffffdcffffffff0000000800000000",
            INIT_7D => X"0000000800000000fffffffefffffffffffffff8ffffffffffffffefffffffff",
            INIT_7E => X"ffffffefffffffff0000003600000000ffffffcaffffffffffffffdaffffffff",
            INIT_7F => X"000000110000000000000022000000000000005400000000ffffffd6ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE34;


    MEM_IWGHT_LAYER2_INSTANCE35 : if BRAM_NAME = "iwght_layer2_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffffffffffffffffff2fffffffffffffffeffffffff0000000600000000",
            INIT_01 => X"fffffff0ffffffff0000000400000000ffffffe5fffffffffffffffeffffffff",
            INIT_02 => X"0000002e0000000000000029000000000000000400000000fffffff3ffffffff",
            INIT_03 => X"0000001d000000000000001d0000000000000005000000000000002500000000",
            INIT_04 => X"ffffffa7ffffffffffffffb4ffffffff00000007000000000000002900000000",
            INIT_05 => X"ffffff8fffffffffffffff89ffffffffffffffbbffffffffffffffb5ffffffff",
            INIT_06 => X"fffffff8ffffffffffffffa1ffffffffffffffbeffffffffffffff93ffffffff",
            INIT_07 => X"000000370000000000000028000000000000002f000000000000003700000000",
            INIT_08 => X"000000150000000000000029000000000000002700000000ffffffffffffffff",
            INIT_09 => X"ffffffb3ffffffffffffffaeffffffffffffffb7ffffffffffffffadffffffff",
            INIT_0A => X"ffffffafffffffffffffffa9ffffffffffffffcfffffffffffffff96ffffffff",
            INIT_0B => X"000000180000000000000027000000000000000000000000ffffffcaffffffff",
            INIT_0C => X"ffffffd7ffffffff00000034000000000000002b000000000000000200000000",
            INIT_0D => X"00000028000000000000000e0000000000000010000000000000001200000000",
            INIT_0E => X"fffffff3ffffffffffffffedffffffffffffffecffffffff0000003200000000",
            INIT_0F => X"0000002600000000fffffff6ffffffffffffffdcffffffffffffffc5ffffffff",
            INIT_10 => X"fffffff5ffffffff0000000d00000000ffffffefffffffff0000001c00000000",
            INIT_11 => X"fffffffcffffffff000000020000000000000002000000000000000700000000",
            INIT_12 => X"0000000400000000fffffff4ffffffffffffffdaffffffffffffffe7ffffffff",
            INIT_13 => X"fffffff5ffffffffffffffe4ffffffff0000001a00000000fffffff5ffffffff",
            INIT_14 => X"0000001700000000ffffffeffffffffffffffff0ffffffffffffffc7ffffffff",
            INIT_15 => X"0000000000000000fffffff7ffffffffffffffd2fffffffffffffff7ffffffff",
            INIT_16 => X"ffffffe9fffffffffffffff9ffffffff00000000000000000000000900000000",
            INIT_17 => X"0000001e000000000000000000000000fffffff9fffffffffffffffeffffffff",
            INIT_18 => X"ffffffecffffffffffffffcaffffffffffffffeeffffffffffffffddffffffff",
            INIT_19 => X"0000001c000000000000000400000000ffffffe5fffffffffffffff1ffffffff",
            INIT_1A => X"0000001400000000ffffffdafffffffffffffff7ffffffff0000000900000000",
            INIT_1B => X"00000002000000000000001e00000000fffffffeffffffff0000001d00000000",
            INIT_1C => X"0000000000000000ffffffecffffffff0000002a000000000000002800000000",
            INIT_1D => X"000000070000000000000006000000000000000f000000000000000a00000000",
            INIT_1E => X"0000000f00000000fffffff1ffffffffffffffebffffffff0000000e00000000",
            INIT_1F => X"000000190000000000000011000000000000001a000000000000000e00000000",
            INIT_20 => X"00000019000000000000001a0000000000000007000000000000000700000000",
            INIT_21 => X"ffffffffffffffffffffffeaffffffffffffffddffffffffffffffe2ffffffff",
            INIT_22 => X"0000001200000000fffffffeffffffff00000000000000000000000600000000",
            INIT_23 => X"00000011000000000000000f000000000000000e000000000000000a00000000",
            INIT_24 => X"00000016000000000000000700000000ffffffe4ffffffffffffffe4ffffffff",
            INIT_25 => X"0000000e000000000000002100000000fffffffaffffffff0000000000000000",
            INIT_26 => X"0000002700000000000000160000000000000026000000000000001900000000",
            INIT_27 => X"0000000b000000000000000f0000000000000005000000000000000c00000000",
            INIT_28 => X"ffffffeeffffffff0000001500000000fffffff3fffffffffffffff7ffffffff",
            INIT_29 => X"ffffffacffffffffffffffd8ffffffff0000001e00000000ffffffd2ffffffff",
            INIT_2A => X"fffffff6ffffffffffffffd6ffffffffffffffe3ffffffff0000000d00000000",
            INIT_2B => X"000000170000000000000002000000000000002b000000000000001e00000000",
            INIT_2C => X"0000000b00000000fffffff9fffffffffffffff7ffffffff0000002700000000",
            INIT_2D => X"fffffffdfffffffffffffff8ffffffff0000000b00000000fffffffeffffffff",
            INIT_2E => X"0000000500000000ffffffeeffffffffffffffebfffffffffffffffdffffffff",
            INIT_2F => X"0000000f0000000000000028000000000000001e000000000000000000000000",
            INIT_30 => X"00000013000000000000001700000000fffffffdffffffff0000000f00000000",
            INIT_31 => X"000000230000000000000010000000000000001f000000000000001a00000000",
            INIT_32 => X"0000000c00000000fffffffdffffffff00000007000000000000002900000000",
            INIT_33 => X"00000017000000000000000000000000fffffffbfffffffffffffff9ffffffff",
            INIT_34 => X"00000029000000000000000a000000000000001b000000000000000900000000",
            INIT_35 => X"fffffff2ffffffffffffffc7ffffffffffffffc4ffffffff0000001600000000",
            INIT_36 => X"ffffffa0ffffffffffffff99ffffffffffffffc5ffffffffffffff77ffffffff",
            INIT_37 => X"ffffffe3ffffffffffffffb2ffffffffffffffd5ffffffffffffffe3ffffffff",
            INIT_38 => X"00000009000000000000000700000000fffffff2ffffffff0000000b00000000",
            INIT_39 => X"0000001e00000000fffffffaffffffffffffffe5fffffffffffffff9ffffffff",
            INIT_3A => X"0000000a00000000fffffffeffffffff00000008000000000000000500000000",
            INIT_3B => X"fffffff3fffffffffffffff5fffffffffffffff1ffffffff0000000800000000",
            INIT_3C => X"00000013000000000000001300000000fffffff1fffffffffffffffbffffffff",
            INIT_3D => X"0000002300000000fffffff2ffffffff0000000a000000000000000300000000",
            INIT_3E => X"00000002000000000000000600000000ffffffdeffffffff0000002900000000",
            INIT_3F => X"0000001800000000fffffffcffffffff0000001700000000ffffffebffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000b00000000fffffff1ffffffffffffffc6fffffffffffffff4ffffffff",
            INIT_41 => X"fffffffaffffffff0000000700000000fffffff5ffffffffffffffcaffffffff",
            INIT_42 => X"ffffffedfffffffffffffff9ffffffffffffffe3fffffffffffffffeffffffff",
            INIT_43 => X"00000008000000000000000200000000ffffffecffffffffffffffdeffffffff",
            INIT_44 => X"000000000000000000000008000000000000000d000000000000000700000000",
            INIT_45 => X"0000001100000000fffffffdffffffffffffffe4ffffffffffffffe7ffffffff",
            INIT_46 => X"0000001b00000000000000190000000000000007000000000000001300000000",
            INIT_47 => X"0000000500000000000000240000000000000020000000000000001d00000000",
            INIT_48 => X"ffffffecffffffffffffffe5fffffffffffffff3fffffffffffffffdffffffff",
            INIT_49 => X"000000030000000000000009000000000000001200000000fffffffbffffffff",
            INIT_4A => X"000000000000000000000018000000000000000f000000000000000500000000",
            INIT_4B => X"0000004600000000000000180000000000000026000000000000001c00000000",
            INIT_4C => X"0000000700000000000000220000000000000023000000000000004700000000",
            INIT_4D => X"fffffffdffffffffffffffc7ffffffff0000000d00000000ffffffffffffffff",
            INIT_4E => X"fffffffeffffffff0000000200000000ffffffd7ffffffffffffffebffffffff",
            INIT_4F => X"ffffffe5ffffffffffffffe6ffffffff0000000f00000000fffffffcffffffff",
            INIT_50 => X"0000000b00000000ffffffc7ffffffffffffff97fffffffffffffffcffffffff",
            INIT_51 => X"ffffff96ffffffff0000000000000000ffffffe7ffffffffffffffffffffffff",
            INIT_52 => X"ffffffcfffffffffffffffa0ffffffffffffffd0ffffffffffffffbcffffffff",
            INIT_53 => X"000000130000000000000023000000000000000e00000000ffffffe7ffffffff",
            INIT_54 => X"0000004100000000fffffff1ffffffff0000000a000000000000000e00000000",
            INIT_55 => X"0000000800000000000000270000000000000023000000000000002500000000",
            INIT_56 => X"ffffffefffffffff0000001300000000ffffffe7ffffffff0000002700000000",
            INIT_57 => X"0000000600000000fffffff5ffffffffffffffeaffffffffffffffcaffffffff",
            INIT_58 => X"fffffff2fffffffffffffff8ffffffff00000005000000000000000400000000",
            INIT_59 => X"fffffff0ffffffff0000000a00000000ffffffecfffffffffffffffaffffffff",
            INIT_5A => X"ffffffffffffffffffffffedffffffff0000000400000000ffffffffffffffff",
            INIT_5B => X"ffffffeeffffffff000000090000000000000024000000000000001500000000",
            INIT_5C => X"00000004000000000000001b000000000000000a000000000000001d00000000",
            INIT_5D => X"fffffff9ffffffff000000170000000000000013000000000000000500000000",
            INIT_5E => X"00000006000000000000000000000000fffffff3ffffffff0000002000000000",
            INIT_5F => X"00000023000000000000000b000000000000000b00000000fffffffcffffffff",
            INIT_60 => X"ffffffd9ffffffff000000050000000000000016000000000000000b00000000",
            INIT_61 => X"ffffffd2fffffffffffffff7fffffffffffffffcffffffffffffffe2ffffffff",
            INIT_62 => X"fffffff4ffffffff00000004000000000000000600000000ffffffeeffffffff",
            INIT_63 => X"ffffffe3ffffffff0000000c00000000fffffff3ffffffffffffffefffffffff",
            INIT_64 => X"ffffffeeffffffff0000000c00000000ffffffe4ffffffffffffffe8ffffffff",
            INIT_65 => X"fffffffcffffffff0000002100000000ffffffdafffffffffffffff7ffffffff",
            INIT_66 => X"00000000000000000000000f000000000000002c00000000fffffff4ffffffff",
            INIT_67 => X"ffffffedffffffff00000003000000000000001b000000000000003a00000000",
            INIT_68 => X"fffffffdffffffffffffffdfffffffffffffffeafffffffffffffffdffffffff",
            INIT_69 => X"0000000900000000ffffffffffffffff0000000400000000fffffffeffffffff",
            INIT_6A => X"fffffff9ffffffffffffffecfffffffffffffff5fffffffffffffffcffffffff",
            INIT_6B => X"0000000c000000000000000a000000000000001500000000ffffffefffffffff",
            INIT_6C => X"0000001b0000000000000039000000000000001e000000000000000900000000",
            INIT_6D => X"0000000e00000000fffffff8ffffffff00000045000000000000004600000000",
            INIT_6E => X"000000170000000000000023000000000000000b000000000000003f00000000",
            INIT_6F => X"ffffffe4ffffffff00000001000000000000000b000000000000000600000000",
            INIT_70 => X"000000260000000000000046000000000000000f00000000fffffff9ffffffff",
            INIT_71 => X"ffffffb0ffffffffffffffd4fffffffffffffffcffffffffffffffe3ffffffff",
            INIT_72 => X"0000003900000000ffffffcaffffffffffffffd7ffffffffffffffd4ffffffff",
            INIT_73 => X"fffffff4ffffffff000000080000000000000012000000000000000800000000",
            INIT_74 => X"ffffffedffffffffffffffedffffffffffffffeeffffffff0000000300000000",
            INIT_75 => X"fffffffdffffffff0000000400000000fffffff6ffffffff0000000c00000000",
            INIT_76 => X"ffffffb8ffffffffffffffe8ffffffffffffffc1ffffffffffffffceffffffff",
            INIT_77 => X"0000000c0000000000000027000000000000001b00000000ffffffc7ffffffff",
            INIT_78 => X"ffffffe9ffffffffffffffe2ffffffffffffffe5fffffffffffffff4ffffffff",
            INIT_79 => X"0000001e000000000000000400000000ffffffdcfffffffffffffff9ffffffff",
            INIT_7A => X"ffffffffffffffff0000000e00000000ffffffe8ffffffff0000001400000000",
            INIT_7B => X"0000000b00000000ffffffd6ffffffff0000000d00000000ffffffe6ffffffff",
            INIT_7C => X"0000001800000000fffffff6ffffffff00000012000000000000001000000000",
            INIT_7D => X"ffffffeafffffffffffffffaffffffffffffffedffffffff0000001000000000",
            INIT_7E => X"ffffffcbffffffffffffffc6ffffffffffffffc4fffffffffffffff4ffffffff",
            INIT_7F => X"ffffffcaffffffff0000000b00000000ffffffdeffffffffffffffacffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE35;


    MEM_IWGHT_LAYER2_INSTANCE36 : if BRAM_NAME = "iwght_layer2_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000150000000000000006000000000000001f00000000ffffff9dffffffff",
            INIT_01 => X"ffffffedffffffff0000001b0000000000000022000000000000001200000000",
            INIT_02 => X"0000000800000000fffffff8ffffffff00000012000000000000001400000000",
            INIT_03 => X"00000016000000000000002800000000fffffff2ffffffff0000000c00000000",
            INIT_04 => X"00000006000000000000002d000000000000001600000000ffffffefffffffff",
            INIT_05 => X"fffffffdfffffffffffffff9ffffffff0000000500000000fffffffaffffffff",
            INIT_06 => X"ffffffe5ffffffffffffffebffffffff0000002500000000fffffff3ffffffff",
            INIT_07 => X"ffffffd7ffffffffffffffecffffffff0000000200000000fffffff1ffffffff",
            INIT_08 => X"ffffffc4ffffffffffffffadffffffffffffffe4ffffffffffffffd5ffffffff",
            INIT_09 => X"ffffffe3ffffffffffffffd5ffffffffffffffe0ffffffff0000001600000000",
            INIT_0A => X"0000001f00000000ffffffd3ffffffffffffffedffffffffffffffefffffffff",
            INIT_0B => X"00000004000000000000002d000000000000001300000000fffffffeffffffff",
            INIT_0C => X"ffffffd1ffffffffffffffe3ffffffff0000000000000000fffffff7ffffffff",
            INIT_0D => X"0000000200000000ffffffd5ffffffffffffffd4fffffffffffffff4ffffffff",
            INIT_0E => X"0000000c00000000ffffffd6ffffffff00000000000000000000000b00000000",
            INIT_0F => X"0000001f000000000000000f00000000fffffff0fffffffffffffff9ffffffff",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER2_INSTANCE36;


    MEM_IWGHT_LAYER3_INSTANCE0 : if BRAM_NAME = "iwght_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000158b00000000fffffc2bfffffffffffff30cffffffffffffd650ffffffff",
            INIT_01 => X"ffffda7effffffff0000391000000000ffffd632ffffffff00002ad400000000",
            INIT_02 => X"ffffffe5ffffffffffffffe4fffffffffffff0dfffffffff00001da200000000",
            INIT_03 => X"00000013000000000000000000000000fffffff3ffffffff0000002200000000",
            INIT_04 => X"0000000a00000000ffffffe8ffffffff0000000e000000000000000000000000",
            INIT_05 => X"0000002a00000000ffffffa7ffffffff0000001d000000000000001900000000",
            INIT_06 => X"ffffffefffffffffffffffebffffffff0000002c00000000ffffffd0ffffffff",
            INIT_07 => X"ffffffd4ffffffff0000002800000000ffffffeeffffffff0000000400000000",
            INIT_08 => X"ffffffc8fffffffffffffff1ffffffff0000001e00000000fffffff4ffffffff",
            INIT_09 => X"ffffffedffffffff0000001600000000ffffffeeffffffff0000000b00000000",
            INIT_0A => X"fffffff7ffffffffffffffe4ffffffff0000000500000000ffffffe3ffffffff",
            INIT_0B => X"ffffff8affffffffffffffe2ffffffff0000002400000000ffffffb2ffffffff",
            INIT_0C => X"ffffffdbfffffffffffffff5fffffffffffffff7fffffffffffffff7ffffffff",
            INIT_0D => X"ffffffebffffffffffffffdfffffffff0000001700000000fffffff3ffffffff",
            INIT_0E => X"fffffffdfffffffffffffffcffffffff0000002f00000000fffffffaffffffff",
            INIT_0F => X"0000000700000000000000140000000000000008000000000000001100000000",
            INIT_10 => X"00000025000000000000001700000000fffffff8fffffffffffffff1ffffffff",
            INIT_11 => X"0000002700000000fffffff0ffffffffffffffe1ffffffffffffffeaffffffff",
            INIT_12 => X"0000000f00000000ffffffe6ffffffff0000002100000000ffffffddffffffff",
            INIT_13 => X"00000016000000000000000000000000ffffffe7ffffffffffffffe6ffffffff",
            INIT_14 => X"0000001a000000000000000c000000000000000d000000000000000400000000",
            INIT_15 => X"fffffff0ffffffffffffffdeffffffff0000002400000000fffffff7ffffffff",
            INIT_16 => X"fffffffeffffffff0000000300000000fffffff8ffffffff0000000a00000000",
            INIT_17 => X"ffffffe1ffffffff00000017000000000000000d00000000ffffffbdffffffff",
            INIT_18 => X"fffffff0ffffffff0000000000000000fffffff2ffffffffffffffdbffffffff",
            INIT_19 => X"0000000000000000ffffffecffffffff00000010000000000000000200000000",
            INIT_1A => X"0000002000000000ffffffdbffffffff0000002e00000000ffffffe6ffffffff",
            INIT_1B => X"ffffffc7ffffffffffffffe0ffffffff0000002500000000ffffffbdffffffff",
            INIT_1C => X"00000017000000000000001800000000ffffffe9fffffffffffffffdffffffff",
            INIT_1D => X"fffffff1ffffffff000000040000000000000009000000000000000d00000000",
            INIT_1E => X"0000001500000000fffffff1ffffffff00000036000000000000001300000000",
            INIT_1F => X"0000003c000000000000002000000000fffffffeffffffff0000002b00000000",
            INIT_20 => X"ffffffe7ffffffff0000001700000000ffffffecffffffff0000000a00000000",
            INIT_21 => X"0000002000000000ffffffe9fffffffffffffff2ffffffffffffffccffffffff",
            INIT_22 => X"00000009000000000000000b00000000ffffffecffffffff0000001800000000",
            INIT_23 => X"00000023000000000000002100000000ffffffe5fffffffffffffffdffffffff",
            INIT_24 => X"000000060000000000000008000000000000000a00000000fffffff7ffffffff",
            INIT_25 => X"fffffffaffffffffffffffdeffffffff00000000000000000000000f00000000",
            INIT_26 => X"fffffff8ffffffff000000050000000000000005000000000000000500000000",
            INIT_27 => X"fffffff5ffffffff000000220000000000000035000000000000001c00000000",
            INIT_28 => X"ffffffecffffffffffffffe9ffffffff0000000900000000ffffffe0ffffffff",
            INIT_29 => X"ffffffd9fffffffffffffff5ffffffffffffffe4ffffffffffffffe9ffffffff",
            INIT_2A => X"000000280000000000000017000000000000003900000000fffffff9ffffffff",
            INIT_2B => X"ffffffc3ffffffffffffffdbffffffffffffffeffffffffffffffff9ffffffff",
            INIT_2C => X"00000049000000000000001600000000ffffffd0ffffffffffffffdaffffffff",
            INIT_2D => X"ffffffd2ffffffffffffffedfffffffffffffffeffffffff0000002800000000",
            INIT_2E => X"0000000000000000ffffffc0ffffffff00000007000000000000001200000000",
            INIT_2F => X"fffffffefffffffffffffffaffffffff0000000200000000fffffff8ffffffff",
            INIT_30 => X"fffffff9ffffffff0000000e000000000000001b00000000ffffffc1ffffffff",
            INIT_31 => X"ffffffa6ffffffffffffffcafffffffffffffff8ffffffff0000000500000000",
            INIT_32 => X"ffffffedfffffffffffffffeffffffff0000002b000000000000000300000000",
            INIT_33 => X"ffffffe4ffffffffffffffedffffffff0000000a00000000fffffff8ffffffff",
            INIT_34 => X"0000003f000000000000003c000000000000000800000000ffffffbcffffffff",
            INIT_35 => X"fffffffdffffffff0000001900000000ffffffc7ffffffffffffffe2ffffffff",
            INIT_36 => X"ffffffbdffffffff00000017000000000000000c00000000fffffff8ffffffff",
            INIT_37 => X"ffffffd2fffffffffffffffbffffffff0000001e00000000ffffffd7ffffffff",
            INIT_38 => X"ffffffadffffffffffffffe4ffffffff00000007000000000000003800000000",
            INIT_39 => X"00000006000000000000000a00000000fffffff6fffffffffffffff0ffffffff",
            INIT_3A => X"ffffffd8ffffffffffffffe4ffffffff0000000800000000fffffff0ffffffff",
            INIT_3B => X"ffffffc4ffffffff00000012000000000000001100000000ffffffe0ffffffff",
            INIT_3C => X"0000000400000000000000140000000000000018000000000000000500000000",
            INIT_3D => X"ffffffdfffffffff0000001400000000ffffffeeffffffffffffffdeffffffff",
            INIT_3E => X"00000003000000000000000300000000ffffffe7ffffffff0000000200000000",
            INIT_3F => X"0000003400000000ffffffe7ffffffff0000000b000000000000000200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002d000000000000001a000000000000000300000000fffffff8ffffffff",
            INIT_41 => X"0000000800000000ffffffecfffffffffffffff6ffffffffffffffe0ffffffff",
            INIT_42 => X"00000010000000000000001500000000fffffffafffffffffffffffaffffffff",
            INIT_43 => X"00000011000000000000001300000000fffffffbffffffffffffffe2ffffffff",
            INIT_44 => X"ffffffeeffffffff00000007000000000000000200000000ffffffe7ffffffff",
            INIT_45 => X"0000001e000000000000001900000000ffffffc4ffffffffffffffeeffffffff",
            INIT_46 => X"ffffffadffffffff000000050000000000000000000000000000001500000000",
            INIT_47 => X"ffffffebffffffffffffffe1ffffffff0000001000000000ffffffeaffffffff",
            INIT_48 => X"ffffffbafffffffffffffffcffffffff00000033000000000000001500000000",
            INIT_49 => X"ffffffb7fffffffffffffffbffffffffffffffe5fffffffffffffff0ffffffff",
            INIT_4A => X"ffffffe3ffffffff0000000500000000ffffffecffffffff0000000000000000",
            INIT_4B => X"fffffff4ffffffff0000000700000000ffffffe5ffffffff0000002a00000000",
            INIT_4C => X"000000020000000000000013000000000000000a00000000ffffffe8ffffffff",
            INIT_4D => X"ffffffe8ffffffff0000000e0000000000000031000000000000000700000000",
            INIT_4E => X"0000000200000000ffffffdafffffffffffffff5ffffffff0000002200000000",
            INIT_4F => X"fffffffeffffffffffffffe5ffffffffffffffe9ffffffff0000001b00000000",
            INIT_50 => X"00000022000000000000000300000000ffffffeffffffffffffffff5ffffffff",
            INIT_51 => X"0000000800000000ffffffdffffffffffffffffaffffffffffffffe6ffffffff",
            INIT_52 => X"fffffff6ffffffff0000002800000000fffffff6ffffffff0000001000000000",
            INIT_53 => X"00000008000000000000000c000000000000001500000000ffffffe2ffffffff",
            INIT_54 => X"ffffffdeffffffff0000002800000000fffffff6ffffffffffffffc2ffffffff",
            INIT_55 => X"ffffffe5ffffffff0000002800000000ffffffc6ffffffff0000000800000000",
            INIT_56 => X"ffffffa1ffffffff0000004c000000000000000d000000000000000500000000",
            INIT_57 => X"ffffffedffffffff0000000a0000000000000034000000000000000600000000",
            INIT_58 => X"ffffffb9ffffffff0000000300000000ffffffd4ffffffff0000001000000000",
            INIT_59 => X"ffffffdaffffffff00000003000000000000000a00000000ffffffcfffffffff",
            INIT_5A => X"ffffffb6fffffffffffffff6ffffffff00000020000000000000000e00000000",
            INIT_5B => X"0000000300000000ffffffd8ffffffff0000000900000000ffffffd9ffffffff",
            INIT_5C => X"0000002a00000000fffffff9ffffffff0000000f00000000fffffff9ffffffff",
            INIT_5D => X"fffffff2ffffffffffffffccfffffffffffffff5ffffffff0000004300000000",
            INIT_5E => X"0000000700000000ffffffc2ffffffffffffffe6ffffffff0000002700000000",
            INIT_5F => X"0000001a00000000ffffffe2ffffffffffffffeeffffffffffffffdaffffffff",
            INIT_60 => X"000000160000000000000015000000000000002e00000000ffffffc8ffffffff",
            INIT_61 => X"ffffffe7ffffffffffffffe9fffffffffffffff6ffffffff0000004800000000",
            INIT_62 => X"ffffffcbfffffffffffffff2ffffffff0000000d000000000000002200000000",
            INIT_63 => X"fffffff5ffffffff00000011000000000000001300000000fffffffeffffffff",
            INIT_64 => X"0000002200000000000000090000000000000017000000000000002000000000",
            INIT_65 => X"fffffff4fffffffffffffff6ffffffffffffffe4ffffffffffffffb1ffffffff",
            INIT_66 => X"0000000900000000ffffffefffffffffffffffd0ffffffffffffffb3ffffffff",
            INIT_67 => X"ffffffe8ffffffffffffffd8ffffffff00000035000000000000001d00000000",
            INIT_68 => X"fffffff7ffffffff00000016000000000000001800000000ffffffd8ffffffff",
            INIT_69 => X"0000001500000000ffffffefffffffff0000000800000000fffffffeffffffff",
            INIT_6A => X"0000000400000000ffffffd3ffffffff0000005c00000000fffffff9ffffffff",
            INIT_6B => X"0000000400000000ffffffdeffffffff00000003000000000000000600000000",
            INIT_6C => X"0000002f000000000000003d00000000fffffffbffffffffffffffd5ffffffff",
            INIT_6D => X"fffffff9ffffffff0000000000000000ffffffefffffffff0000000200000000",
            INIT_6E => X"00000026000000000000000f000000000000000300000000ffffffc4ffffffff",
            INIT_6F => X"0000001800000000ffffffb7ffffffff0000000e00000000fffffff5ffffffff",
            INIT_70 => X"ffffffe5ffffffffffffffedffffffffffffffd3ffffffff0000002c00000000",
            INIT_71 => X"fffffff3ffffffff0000000200000000fffffffbfffffffffffffff4ffffffff",
            INIT_72 => X"0000000300000000ffffffd8ffffffff00000025000000000000002400000000",
            INIT_73 => X"ffffffebfffffffffffffffbffffffff0000000800000000ffffffe1ffffffff",
            INIT_74 => X"0000000d000000000000000e00000000ffffffe7ffffffff0000002400000000",
            INIT_75 => X"000000120000000000000011000000000000002700000000ffffffddffffffff",
            INIT_76 => X"fffffff0ffffffffffffffdbffffffff00000018000000000000000300000000",
            INIT_77 => X"0000000000000000ffffffe7ffffffff00000009000000000000004300000000",
            INIT_78 => X"ffffffdafffffffffffffffcfffffffffffffff7fffffffffffffff6ffffffff",
            INIT_79 => X"000000110000000000000010000000000000000c000000000000000700000000",
            INIT_7A => X"0000002300000000ffffffeaffffffff00000008000000000000000900000000",
            INIT_7B => X"0000001800000000ffffffc0ffffffff00000023000000000000000000000000",
            INIT_7C => X"00000003000000000000004b0000000000000004000000000000000700000000",
            INIT_7D => X"ffffffd4ffffffff0000002d000000000000003500000000ffffffe3ffffffff",
            INIT_7E => X"ffffffeafffffffffffffff5ffffffff0000002600000000fffffffaffffffff",
            INIT_7F => X"0000000100000000ffffffeffffffffffffffff8ffffffffffffffebffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE0;


    MEM_IWGHT_LAYER3_INSTANCE1 : if BRAM_NAME = "iwght_layer3_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000017000000000000001b00000000fffffffaffffffff0000000300000000",
            INIT_01 => X"0000002700000000000000200000000000000050000000000000000000000000",
            INIT_02 => X"ffffffb9ffffffff0000002100000000fffffff3ffffffffffffffefffffffff",
            INIT_03 => X"00000016000000000000001d000000000000001400000000ffffffddffffffff",
            INIT_04 => X"ffffffffffffffffffffffc2ffffffff00000013000000000000000e00000000",
            INIT_05 => X"0000004e00000000ffffffd7fffffffffffffff5ffffffffffffffc9ffffffff",
            INIT_06 => X"ffffffbdffffffff00000013000000000000000000000000fffffffbffffffff",
            INIT_07 => X"ffffffd4fffffffffffffff5ffffffff0000000e000000000000001e00000000",
            INIT_08 => X"fffffff7ffffffffffffffe9ffffffffffffffd4ffffffff0000000600000000",
            INIT_09 => X"0000001d00000000fffffff3ffffffff00000011000000000000000c00000000",
            INIT_0A => X"0000000a000000000000000800000000fffffff4ffffffffffffffe8ffffffff",
            INIT_0B => X"fffffff9ffffffffffffffc9ffffffff0000003400000000ffffffeeffffffff",
            INIT_0C => X"fffffffaffffffffffffffe4fffffffffffffff0ffffffff0000000e00000000",
            INIT_0D => X"fffffff5ffffffffffffffd8ffffffffffffffe7ffffffff0000000a00000000",
            INIT_0E => X"ffffffc5ffffffffffffffffffffffffffffffebffffffffffffffe1ffffffff",
            INIT_0F => X"0000000a00000000fffffffaffffffff0000000e00000000fffffffdffffffff",
            INIT_10 => X"000000340000000000000044000000000000001500000000ffffffdaffffffff",
            INIT_11 => X"ffffffdefffffffffffffff4ffffffff0000002f000000000000000200000000",
            INIT_12 => X"ffffffeeffffffff0000001000000000ffffffecffffffff0000002100000000",
            INIT_13 => X"ffffffc5ffffffffffffffd8fffffffffffffff0ffffffff0000000700000000",
            INIT_14 => X"0000000d00000000ffffffeefffffffffffffffdffffffffffffffefffffffff",
            INIT_15 => X"ffffffddffffffff0000000300000000fffffff5fffffffffffffffaffffffff",
            INIT_16 => X"0000002c000000000000001200000000ffffffdbffffffff0000002000000000",
            INIT_17 => X"ffffffe9fffffffffffffffaffffffff0000000600000000fffffffbffffffff",
            INIT_18 => X"fffffff9ffffffff00000000000000000000000c00000000fffffff4ffffffff",
            INIT_19 => X"fffffff4fffffffffffffff2ffffffff0000000a00000000ffffffe4ffffffff",
            INIT_1A => X"ffffffe6ffffffffffffffe7ffffffff0000001700000000ffffffdfffffffff",
            INIT_1B => X"0000001000000000000000140000000000000003000000000000000b00000000",
            INIT_1C => X"0000000200000000000000040000000000000006000000000000000200000000",
            INIT_1D => X"ffffffe9ffffffffffffffedffffffff0000002500000000fffffff7ffffffff",
            INIT_1E => X"ffffffe4ffffffffffffffedfffffffffffffff7fffffffffffffff6ffffffff",
            INIT_1F => X"fffffff7ffffffff000000000000000000000001000000000000001200000000",
            INIT_20 => X"fffffff5ffffffffffffffb8fffffffffffffffaffffffff0000000300000000",
            INIT_21 => X"ffffffa7fffffffffffffffcffffffff0000001700000000ffffffe2ffffffff",
            INIT_22 => X"ffffffefffffffffffffffd3ffffffff00000002000000000000000200000000",
            INIT_23 => X"ffffffdeffffffffffffffcbfffffffffffffff4ffffffffffffffe2ffffffff",
            INIT_24 => X"fffffff0ffffffff00000008000000000000000e00000000ffffffd6ffffffff",
            INIT_25 => X"00000023000000000000001700000000ffffffefffffffffffffffcfffffffff",
            INIT_26 => X"fffffff9ffffffff0000000200000000fffffff7ffffffff0000003300000000",
            INIT_27 => X"0000002200000000ffffffeeffffffff0000001100000000ffffffefffffffff",
            INIT_28 => X"00000007000000000000000200000000ffffffd6ffffffff0000001800000000",
            INIT_29 => X"000000020000000000000006000000000000000f00000000ffffffe4ffffffff",
            INIT_2A => X"ffffffcdffffffff0000000200000000ffffffdefffffffffffffffcffffffff",
            INIT_2B => X"0000002100000000ffffffeeffffffffffffffebffffffff0000001700000000",
            INIT_2C => X"ffffffd7ffffffff00000014000000000000003100000000ffffffe6ffffffff",
            INIT_2D => X"fffffffaffffffff000000160000000000000008000000000000003b00000000",
            INIT_2E => X"fffffff3ffffffffffffffe8ffffffffffffffddffffffff0000000200000000",
            INIT_2F => X"0000000500000000ffffffc3ffffffff0000001000000000ffffffffffffffff",
            INIT_30 => X"0000000300000000fffffff9ffffffff0000000e000000000000001300000000",
            INIT_31 => X"ffffffd1ffffffffffffffdefffffffffffffff8ffffffff0000000400000000",
            INIT_32 => X"ffffffe7ffffffff000000130000000000000030000000000000001d00000000",
            INIT_33 => X"ffffffffffffffffffffffd3ffffffff0000000f000000000000000600000000",
            INIT_34 => X"ffffffe8fffffffffffffff1ffffffffffffffecffffffff0000000e00000000",
            INIT_35 => X"0000001500000000ffffffe9ffffffffffffffe4fffffffffffffff3ffffffff",
            INIT_36 => X"0000002000000000ffffffedffffffff0000000d00000000fffffff0ffffffff",
            INIT_37 => X"000000310000000000000025000000000000000800000000ffffffd7ffffffff",
            INIT_38 => X"fffffffcffffffff000000130000000000000005000000000000002200000000",
            INIT_39 => X"0000001100000000fffffff7ffffffffffffffefffffffffffffffffffffffff",
            INIT_3A => X"ffffffd5ffffffffffffffe5ffffffffffffffcefffffffffffffffcffffffff",
            INIT_3B => X"0000002e00000000fffffffeffffffffffffffe3ffffffffffffffe7ffffffff",
            INIT_3C => X"ffffffedffffffff00000008000000000000001900000000ffffffc5ffffffff",
            INIT_3D => X"0000000200000000000000250000000000000001000000000000001b00000000",
            INIT_3E => X"ffffffd5ffffffffffffff83ffffffffffffffdffffffffffffffffcffffffff",
            INIT_3F => X"fffffff9ffffffff0000001e000000000000000700000000ffffffe6ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000200000000ffffffd9ffffffff0000001e000000000000000d00000000",
            INIT_41 => X"0000002300000000fffffff0fffffffffffffffeffffffff0000000000000000",
            INIT_42 => X"0000000500000000fffffff6ffffffffffffffe8ffffffff0000003000000000",
            INIT_43 => X"ffffffdeffffffff000000420000000000000006000000000000000500000000",
            INIT_44 => X"fffffff6ffffffffffffffe3ffffffffffffffecfffffffffffffff3ffffffff",
            INIT_45 => X"0000000600000000ffffffdfffffffffffffffe2ffffffffffffff94ffffffff",
            INIT_46 => X"0000002100000000ffffffe7ffffffff0000001000000000ffffffdbffffffff",
            INIT_47 => X"0000000e0000000000000016000000000000002e000000000000001600000000",
            INIT_48 => X"00000007000000000000001800000000ffffffe7ffffffff0000000e00000000",
            INIT_49 => X"00000015000000000000000600000000fffffff1ffffffff0000000100000000",
            INIT_4A => X"ffffffc1ffffffff0000003200000000ffffffd1ffffffff0000001400000000",
            INIT_4B => X"ffffffe4ffffffff0000001100000000ffffffdcffffffff0000000b00000000",
            INIT_4C => X"ffffffd6ffffffff0000002400000000ffffffe8ffffffff0000002300000000",
            INIT_4D => X"0000000200000000ffffffc2ffffffff0000003400000000ffffffd2ffffffff",
            INIT_4E => X"ffffffd0ffffffff0000004b00000000ffffffceffffffff0000000f00000000",
            INIT_4F => X"fffffff7ffffffffffffffbfffffffff00000003000000000000001c00000000",
            INIT_50 => X"00000030000000000000000200000000ffffffebffffffff0000000900000000",
            INIT_51 => X"ffffffd9ffffffffffffffdffffffffffffffff8ffffffff0000000d00000000",
            INIT_52 => X"0000000100000000000000080000000000000018000000000000000e00000000",
            INIT_53 => X"00000030000000000000002f00000000fffffffbffffffff0000001c00000000",
            INIT_54 => X"ffffffe3ffffffff0000000e00000000ffffffffffffffffffffffe0ffffffff",
            INIT_55 => X"00000029000000000000000700000000ffffffc6ffffffffffffff95ffffffff",
            INIT_56 => X"fffffffeffffffff00000000000000000000000800000000ffffffe5ffffffff",
            INIT_57 => X"00000005000000000000002a000000000000000b000000000000000400000000",
            INIT_58 => X"ffffffb3ffffffff00000015000000000000003800000000fffffff6ffffffff",
            INIT_59 => X"ffffffaffffffffffffffffaffffffff00000014000000000000002200000000",
            INIT_5A => X"ffffffd0ffffffff0000002c00000000ffffffc5ffffffff0000001900000000",
            INIT_5B => X"fffffffbfffffffffffffff5ffffffffffffffd4ffffffff0000000a00000000",
            INIT_5C => X"000000090000000000000000000000000000002b00000000fffffffaffffffff",
            INIT_5D => X"ffffffe3fffffffffffffff3fffffffffffffff4ffffffffffffffc5ffffffff",
            INIT_5E => X"ffffffe7ffffffff0000000200000000ffffffc3ffffffff0000000000000000",
            INIT_5F => X"0000001800000000ffffffb4fffffffffffffffaffffffffffffffdcffffffff",
            INIT_60 => X"00000019000000000000002400000000ffffffddffffffffffffffe5ffffffff",
            INIT_61 => X"0000001300000000ffffffe9ffffffff0000000a000000000000001100000000",
            INIT_62 => X"0000002c00000000ffffffccffffffff00000029000000000000000000000000",
            INIT_63 => X"000000320000000000000025000000000000001700000000ffffffeaffffffff",
            INIT_64 => X"ffffffcaffffffffffffffd3ffffffffffffffecffffffffffffffe5ffffffff",
            INIT_65 => X"0000003b00000000ffffff96ffffffffffffffc3ffffffffffffffe4ffffffff",
            INIT_66 => X"ffffffe8fffffffffffffffeffffffff0000000b00000000fffffff6ffffffff",
            INIT_67 => X"000000460000000000000028000000000000001500000000ffffffd3ffffffff",
            INIT_68 => X"ffffffceffffffffffffffeeffffffff0000000b00000000fffffff2ffffffff",
            INIT_69 => X"ffffffcdffffffff000000000000000000000014000000000000001600000000",
            INIT_6A => X"ffffff98ffffffff00000019000000000000001200000000ffffffefffffffff",
            INIT_6B => X"0000000800000000ffffffe0ffffffff0000000e00000000ffffffe5ffffffff",
            INIT_6C => X"0000002300000000ffffffe3ffffffff0000002600000000fffffff3ffffffff",
            INIT_6D => X"fffffffbfffffffffffffff6ffffffff0000000000000000ffffffebffffffff",
            INIT_6E => X"0000000c00000000ffffffe7ffffffffffffffb4fffffffffffffff8ffffffff",
            INIT_6F => X"ffffffeeffffffffffffffd1ffffffff0000000c00000000fffffff1ffffffff",
            INIT_70 => X"ffffffecffffffff0000000c00000000ffffffeaffffffff0000002100000000",
            INIT_71 => X"ffffffbcffffffffffffffe4ffffffff0000004a000000000000002800000000",
            INIT_72 => X"00000045000000000000000600000000fffffff0fffffffffffffffdffffffff",
            INIT_73 => X"ffffffedffffffff0000001a00000000fffffff7ffffffffffffffd7ffffffff",
            INIT_74 => X"fffffff8ffffffffffffffc4ffffffff0000000000000000ffffffe4ffffffff",
            INIT_75 => X"000000170000000000000036000000000000000400000000ffffffc6ffffffff",
            INIT_76 => X"000000150000000000000016000000000000004000000000fffffffeffffffff",
            INIT_77 => X"fffffff2ffffffffffffffbefffffffffffffffcfffffffffffffffbffffffff",
            INIT_78 => X"ffffffbeffffffff0000000500000000fffffff8ffffffff0000001d00000000",
            INIT_79 => X"ffffffccffffffff0000001900000000fffffffaffffffffffffffe8ffffffff",
            INIT_7A => X"0000003300000000ffffffe6fffffffffffffff2fffffffffffffffaffffffff",
            INIT_7B => X"ffffffafffffffffffffffbfffffffff00000016000000000000000c00000000",
            INIT_7C => X"ffffffadffffffffffffffcfffffffffffffffa4ffffffff0000002b00000000",
            INIT_7D => X"fffffff3ffffffff00000013000000000000002a00000000ffffffe7ffffffff",
            INIT_7E => X"ffffffc1ffffffff0000003c00000000ffffffd1fffffffffffffff6ffffffff",
            INIT_7F => X"0000002800000000ffffffeeffffffffffffffe9ffffffff0000001700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE1;


    MEM_IWGHT_LAYER3_INSTANCE2 : if BRAM_NAME = "iwght_layer3_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004000000000ffffffd3ffffffff0000002a000000000000003500000000",
            INIT_01 => X"0000004b00000000ffffffffffffffffffffffe9fffffffffffffff1ffffffff",
            INIT_02 => X"0000004d000000000000001b000000000000002300000000ffffffa3ffffffff",
            INIT_03 => X"0000001f000000000000000d0000000000000002000000000000001200000000",
            INIT_04 => X"ffffffbbffffffffffffffdaffffffffffffffe3ffffffffffffffb2ffffffff",
            INIT_05 => X"fffffffdffffffff0000000e00000000ffffffccffffffff0000003900000000",
            INIT_06 => X"fffffff4ffffffffffffffeaffffffff00000007000000000000004a00000000",
            INIT_07 => X"0000002200000000ffffffdcffffffff0000002900000000ffffffe1ffffffff",
            INIT_08 => X"ffffffe2ffffffff00000019000000000000001d000000000000000000000000",
            INIT_09 => X"000000120000000000000003000000000000000b000000000000000200000000",
            INIT_0A => X"ffffff9dffffffffffffffeefffffffffffffffbffffffff0000001b00000000",
            INIT_0B => X"00000006000000000000000000000000fffffff7ffffffff0000006a00000000",
            INIT_0C => X"fffffff3ffffffffffffffd5ffffffffffffffd8ffffffffffffffe1ffffffff",
            INIT_0D => X"0000001000000000000000270000000000000036000000000000004a00000000",
            INIT_0E => X"00000015000000000000000b0000000000000000000000000000000e00000000",
            INIT_0F => X"0000002f000000000000000a00000000ffffffe7ffffffffffffffd7ffffffff",
            INIT_10 => X"00000032000000000000000b0000000000000009000000000000000d00000000",
            INIT_11 => X"0000000b00000000ffffffd3ffffffff0000001d00000000ffffffe7ffffffff",
            INIT_12 => X"0000006e00000000fffffff7ffffffff0000001e00000000ffffffecffffffff",
            INIT_13 => X"ffffffc9ffffffff0000000b000000000000000000000000fffffffeffffffff",
            INIT_14 => X"ffffffbfffffffffffffffc3ffffffffffffffecffffffffffffffe8ffffffff",
            INIT_15 => X"ffffffe5ffffffff0000002b000000000000002100000000ffffffe9ffffffff",
            INIT_16 => X"0000002f00000000ffffffc1ffffffff0000000f00000000fffffffaffffffff",
            INIT_17 => X"0000004700000000fffffffaffffffff00000008000000000000003800000000",
            INIT_18 => X"ffffffbdffffffff00000001000000000000001a000000000000000a00000000",
            INIT_19 => X"ffffffdfffffffff0000000400000000fffffff8fffffffffffffff8ffffffff",
            INIT_1A => X"fffffffaffffffff0000000a000000000000005600000000fffffff7ffffffff",
            INIT_1B => X"ffffffe7ffffffffffffffcdffffffffffffffc0ffffffffffffffe0ffffffff",
            INIT_1C => X"0000004800000000ffffffe6ffffffffffffffc5ffffffffffffffc3ffffffff",
            INIT_1D => X"00000006000000000000001c0000000000000043000000000000000900000000",
            INIT_1E => X"0000000000000000ffffffceffffffffffffffe9fffffffffffffff0ffffffff",
            INIT_1F => X"0000001400000000ffffffd1ffffffff0000000200000000fffffffcffffffff",
            INIT_20 => X"ffffffd8ffffffff0000000500000000ffffffe0ffffffff0000002400000000",
            INIT_21 => X"ffffffefffffffffffffffeaffffffff0000000b00000000ffffffe5ffffffff",
            INIT_22 => X"ffffffdfffffffffffffffeeffffffff0000001800000000ffffffcbffffffff",
            INIT_23 => X"000000130000000000000006000000000000000900000000ffffffc5ffffffff",
            INIT_24 => X"0000002a00000000000000110000000000000011000000000000001b00000000",
            INIT_25 => X"fffffff5fffffffffffffff3ffffffff0000000300000000fffffff1ffffffff",
            INIT_26 => X"0000002700000000fffffff4ffffffff0000000a00000000ffffffe7ffffffff",
            INIT_27 => X"ffffffebffffffff0000000b000000000000000900000000ffffffccffffffff",
            INIT_28 => X"0000000800000000ffffffeaffffffffffffffc8ffffffff0000000900000000",
            INIT_29 => X"000000000000000000000013000000000000000300000000ffffffdbffffffff",
            INIT_2A => X"0000001000000000ffffffc2fffffffffffffff2ffffffff0000000400000000",
            INIT_2B => X"ffffffe4fffffffffffffff4ffffffff00000028000000000000001e00000000",
            INIT_2C => X"00000006000000000000001f00000000fffffffcffffffff0000002900000000",
            INIT_2D => X"ffffffe9ffffffff0000000200000000ffffffe7fffffffffffffff9ffffffff",
            INIT_2E => X"0000000800000000000000090000000000000019000000000000001400000000",
            INIT_2F => X"ffffffeeffffffffffffffe4ffffffff0000000900000000fffffffeffffffff",
            INIT_30 => X"fffffff8ffffffff0000001100000000ffffffd0ffffffffffffffe1ffffffff",
            INIT_31 => X"0000000c000000000000001f00000000ffffffffffffffff0000001700000000",
            INIT_32 => X"fffffff6fffffffffffffff2fffffffffffffffcffffffff0000000a00000000",
            INIT_33 => X"fffffffdffffffffffffffd5ffffffff00000004000000000000001300000000",
            INIT_34 => X"0000002b00000000ffffffdbfffffffffffffff7ffffffffffffffddffffffff",
            INIT_35 => X"0000001400000000fffffff2fffffffffffffff0ffffffff0000000300000000",
            INIT_36 => X"0000000c0000000000000019000000000000000b000000000000000400000000",
            INIT_37 => X"00000015000000000000000300000000fffffff3ffffffffffffffefffffffff",
            INIT_38 => X"ffffffebffffffff0000000b000000000000003d000000000000000000000000",
            INIT_39 => X"ffffffedffffffff00000000000000000000000300000000fffffffaffffffff",
            INIT_3A => X"fffffff3fffffffffffffffdffffffff00000024000000000000000000000000",
            INIT_3B => X"fffffffbffffffffffffffd9ffffffff0000000700000000fffffff2ffffffff",
            INIT_3C => X"0000001200000000000000080000000000000014000000000000004e00000000",
            INIT_3D => X"ffffffdbfffffffffffffffbffffffffffffffc3ffffffffffffffe5ffffffff",
            INIT_3E => X"000000130000000000000009000000000000003000000000ffffffebffffffff",
            INIT_3F => X"ffffffbdffffffff0000000a00000000fffffffaffffffff0000000e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff1fffffffffffffffaffffffff0000001d00000000ffffffefffffffff",
            INIT_41 => X"fffffff9ffffffffffffffd9fffffffffffffff6ffffffff0000001600000000",
            INIT_42 => X"fffffff3ffffffffffffffe7fffffffffffffff5ffffffff0000000b00000000",
            INIT_43 => X"000000240000000000000021000000000000000700000000ffffffffffffffff",
            INIT_44 => X"0000001b00000000fffffff2ffffffffffffffeefffffffffffffffcffffffff",
            INIT_45 => X"fffffffdffffffff0000001900000000ffffffe8ffffffff0000001500000000",
            INIT_46 => X"00000034000000000000000f00000000ffffffdffffffffffffffffeffffffff",
            INIT_47 => X"0000001d000000000000001900000000ffffffd0ffffffff0000000c00000000",
            INIT_48 => X"00000011000000000000001600000000fffffffbfffffffffffffff3ffffffff",
            INIT_49 => X"fffffff4fffffffffffffffbffffffff0000000200000000fffffff3ffffffff",
            INIT_4A => X"fffffff1fffffffffffffff5fffffffffffffff8ffffffff0000000900000000",
            INIT_4B => X"fffffff6ffffffffffffffe3fffffffffffffffaffffffff0000002e00000000",
            INIT_4C => X"0000001e00000000fffffff5ffffffffffffffefffffffff0000000800000000",
            INIT_4D => X"fffffff6ffffffff0000000d00000000ffffffcaffffffffffffffedffffffff",
            INIT_4E => X"ffffffe5ffffffffffffffdfffffffff0000001e00000000fffffff4ffffffff",
            INIT_4F => X"0000000e000000000000001600000000ffffffe6ffffffff0000002a00000000",
            INIT_50 => X"ffffffeaffffffffffffffe7ffffffffffffffd8ffffffffffffffffffffffff",
            INIT_51 => X"ffffffe9ffffffff0000000e0000000000000019000000000000000b00000000",
            INIT_52 => X"fffffff4ffffffffffffffe7ffffffffffffffdbffffffffffffffffffffffff",
            INIT_53 => X"0000003200000000ffffffdeffffffff0000000e00000000ffffffedffffffff",
            INIT_54 => X"fffffff2ffffffff0000002f000000000000001500000000fffffff3ffffffff",
            INIT_55 => X"ffffffeeffffffff0000000f000000000000001c000000000000000200000000",
            INIT_56 => X"0000000700000000ffffffe4ffffffffffffffe8ffffffff0000000600000000",
            INIT_57 => X"ffffffc7fffffffffffffff4ffffffff0000001f00000000ffffffc4ffffffff",
            INIT_58 => X"0000001700000000ffffffe4fffffffffffffff4fffffffffffffff7ffffffff",
            INIT_59 => X"ffffffefffffffffffffffeeffffffff0000000700000000ffffffeeffffffff",
            INIT_5A => X"0000002b00000000ffffffcffffffffffffffff3ffffffff0000000700000000",
            INIT_5B => X"ffffffdbffffffffffffffc6ffffffff0000002c000000000000003600000000",
            INIT_5C => X"0000000f000000000000001e0000000000000000000000000000001a00000000",
            INIT_5D => X"00000009000000000000001100000000ffffffe2ffffffff0000000b00000000",
            INIT_5E => X"ffffffc7ffffffffffffffd1ffffffff0000000e000000000000000300000000",
            INIT_5F => X"0000001500000000fffffff0ffffffffffffffeeffffffff0000004800000000",
            INIT_60 => X"ffffffcafffffffffffffffafffffffffffffff0ffffffffffffffe0ffffffff",
            INIT_61 => X"000000230000000000000021000000000000000500000000ffffffdcffffffff",
            INIT_62 => X"0000000a00000000ffffffdbffffffff00000016000000000000002c00000000",
            INIT_63 => X"ffffffe3ffffffffffffffe5ffffffff00000003000000000000002600000000",
            INIT_64 => X"ffffffe5fffffffffffffff1fffffffffffffffdffffffffffffffc3ffffffff",
            INIT_65 => X"ffffffe4ffffffff0000001200000000fffffff6fffffffffffffff5ffffffff",
            INIT_66 => X"fffffffafffffffffffffffcffffffffffffffc8ffffffff0000002900000000",
            INIT_67 => X"0000001b00000000fffffffbffffffff00000013000000000000000a00000000",
            INIT_68 => X"0000000200000000fffffff6ffffffff0000001100000000ffffffeeffffffff",
            INIT_69 => X"fffffff9ffffffffffffffe8ffffffff0000000e00000000ffffffd9ffffffff",
            INIT_6A => X"ffffffe5ffffffff0000003d000000000000002900000000fffffff0ffffffff",
            INIT_6B => X"fffffff1ffffffffffffffafffffffff0000003000000000fffffff2ffffffff",
            INIT_6C => X"0000000700000000ffffffe7ffffffff00000020000000000000002d00000000",
            INIT_6D => X"ffffffe7ffffffff0000002900000000ffffffe7ffffffff0000000400000000",
            INIT_6E => X"ffffffe2ffffffffffffffeaffffffffffffffebffffffffffffffc8ffffffff",
            INIT_6F => X"ffffffb7fffffffffffffffdffffffff00000000000000000000003400000000",
            INIT_70 => X"fffffff2ffffffff0000000b000000000000005900000000ffffffd9ffffffff",
            INIT_71 => X"0000003500000000ffffffebffffffffffffffd3ffffffff0000000c00000000",
            INIT_72 => X"0000000000000000ffffffdcffffffff0000001300000000ffffffe0ffffffff",
            INIT_73 => X"0000002900000000ffffffceffffffff0000000b000000000000001400000000",
            INIT_74 => X"0000000200000000fffffffbfffffffffffffff3fffffffffffffffcffffffff",
            INIT_75 => X"fffffffdffffffff000000250000000000000008000000000000000d00000000",
            INIT_76 => X"0000002800000000ffffffdeffffffffffffffd0ffffffff0000000c00000000",
            INIT_77 => X"00000002000000000000000300000000ffffffe0ffffffff0000001b00000000",
            INIT_78 => X"ffffffe0fffffffffffffff3ffffffffffffffd3ffffffffffffffd8ffffffff",
            INIT_79 => X"fffffffbfffffffffffffffeffffffff0000001200000000fffffff9ffffffff",
            INIT_7A => X"0000000500000000000000250000000000000011000000000000000800000000",
            INIT_7B => X"0000000c00000000ffffffcdffffffff0000001b00000000fffffff7ffffffff",
            INIT_7C => X"00000008000000000000001b00000000ffffffdfffffffff0000002b00000000",
            INIT_7D => X"0000000000000000ffffffddffffffffffffffe7ffffffff0000004100000000",
            INIT_7E => X"0000002c00000000ffffffedffffffff00000027000000000000001300000000",
            INIT_7F => X"00000009000000000000001a0000000000000010000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE2;


    MEM_IWGHT_LAYER3_INSTANCE3 : if BRAM_NAME = "iwght_layer3_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000fffffff0fffffffffffffff4ffffffffffffffe9ffffffff",
            INIT_01 => X"ffffffeffffffffffffffffcffffffff0000001500000000ffffffebffffffff",
            INIT_02 => X"ffffffdeffffffffffffffe3ffffffffffffffe5ffffffff0000003a00000000",
            INIT_03 => X"0000003200000000ffffffd9ffffffff0000000f000000000000002400000000",
            INIT_04 => X"ffffffe9ffffffff0000006900000000ffffffeefffffffffffffff9ffffffff",
            INIT_05 => X"fffffff1ffffffffffffffcdffffffff0000000400000000fffffffeffffffff",
            INIT_06 => X"ffffffd8fffffffffffffff2ffffffffffffffd8ffffffffffffffedffffffff",
            INIT_07 => X"ffffffe4ffffffff000000350000000000000019000000000000001c00000000",
            INIT_08 => X"0000001300000000ffffffebffffffff0000001f00000000ffffffe2ffffffff",
            INIT_09 => X"0000001e00000000fffffffdffffffff00000009000000000000001b00000000",
            INIT_0A => X"0000000c0000000000000001000000000000000600000000ffffffe9ffffffff",
            INIT_0B => X"fffffff3ffffffff0000003500000000ffffffe8ffffffff0000000600000000",
            INIT_0C => X"0000000e0000000000000009000000000000003700000000fffffff4ffffffff",
            INIT_0D => X"0000000e00000000ffffffc4ffffffffffffffbfffffffff0000001500000000",
            INIT_0E => X"0000000000000000ffffffd4ffffffffffffffffffffffff0000000900000000",
            INIT_0F => X"0000001700000000fffffff5fffffffffffffff8ffffffffffffffffffffffff",
            INIT_10 => X"0000000f000000000000002600000000ffffffc2ffffffffffffffe7ffffffff",
            INIT_11 => X"ffffffd8ffffffff00000032000000000000000400000000ffffffb6ffffffff",
            INIT_12 => X"ffffffdbffffffff0000001500000000ffffffeefffffffffffffffbffffffff",
            INIT_13 => X"ffffffeeffffffff0000000d00000000fffffff9ffffffff0000001a00000000",
            INIT_14 => X"000000240000000000000034000000000000000400000000fffffff4ffffffff",
            INIT_15 => X"00000006000000000000000200000000fffffffdffffffffffffffe4ffffffff",
            INIT_16 => X"ffffffe2fffffffffffffff7ffffffffffffffe8fffffffffffffff6ffffffff",
            INIT_17 => X"00000020000000000000004800000000ffffffeaffffffffffffffe6ffffffff",
            INIT_18 => X"0000000f0000000000000004000000000000000f00000000ffffffffffffffff",
            INIT_19 => X"ffffffdffffffffffffffff7ffffffff0000001300000000fffffffdffffffff",
            INIT_1A => X"0000003700000000fffffffafffffffffffffff2fffffffffffffffeffffffff",
            INIT_1B => X"fffffff0ffffffffffffffe6fffffffffffffff7ffffffffffffffd0ffffffff",
            INIT_1C => X"0000000200000000ffffffd4ffffffff00000026000000000000002800000000",
            INIT_1D => X"fffffffcffffffffffffffe0ffffffffffffffe5ffffffffffffffe6ffffffff",
            INIT_1E => X"0000000b00000000fffffff8ffffffff0000002500000000ffffffefffffffff",
            INIT_1F => X"ffffffbaffffffff0000000b00000000fffffff7fffffffffffffffbffffffff",
            INIT_20 => X"0000001300000000fffffff1ffffffffffffffebfffffffffffffffaffffffff",
            INIT_21 => X"00000003000000000000001000000000fffffff6ffffffff0000000a00000000",
            INIT_22 => X"ffffffbfffffffffffffffd2ffffffffffffffecffffffffffffffc1ffffffff",
            INIT_23 => X"0000002800000000ffffffe2ffffffff00000009000000000000000000000000",
            INIT_24 => X"0000001100000000000000110000000000000013000000000000000f00000000",
            INIT_25 => X"0000002d00000000ffffffd4ffffffff0000000100000000fffffffbffffffff",
            INIT_26 => X"0000001b000000000000000f00000000ffffffe7fffffffffffffffbffffffff",
            INIT_27 => X"ffffffddffffffff0000000b00000000ffffffeafffffffffffffff9ffffffff",
            INIT_28 => X"0000001700000000fffffff1ffffffffffffffc3fffffffffffffff3ffffffff",
            INIT_29 => X"ffffffeeffffffff0000000e00000000fffffff0ffffffffffffffebffffffff",
            INIT_2A => X"0000001700000000ffffffcfffffffffffffffc7fffffffffffffffdffffffff",
            INIT_2B => X"0000000600000000fffffffcffffffff0000000c000000000000001600000000",
            INIT_2C => X"ffffffefffffffff000000000000000000000010000000000000004a00000000",
            INIT_2D => X"0000000600000000ffffffb1ffffffffffffffaffffffffffffffffbffffffff",
            INIT_2E => X"00000035000000000000002a0000000000000037000000000000000d00000000",
            INIT_2F => X"00000028000000000000000c00000000ffffffe9ffffffff0000001f00000000",
            INIT_30 => X"0000003d000000000000000000000000ffffffcfffffffff0000000000000000",
            INIT_31 => X"ffffffd2ffffffff0000001c0000000000000008000000000000001b00000000",
            INIT_32 => X"0000001000000000000000020000000000000010000000000000000000000000",
            INIT_33 => X"fffffff6ffffffff0000000400000000fffffffcffffffff0000001b00000000",
            INIT_34 => X"fffffffbffffffffffffffe4ffffffffffffffe8fffffffffffffff5ffffffff",
            INIT_35 => X"0000001000000000000000300000000000000000000000000000001e00000000",
            INIT_36 => X"fffffff1ffffffffffffffedffffffffffffffeeffffffff0000000d00000000",
            INIT_37 => X"0000000700000000fffffff0ffffffffffffffefffffffffffffffccffffffff",
            INIT_38 => X"fffffff0ffffffff0000000e000000000000000c00000000fffffffcffffffff",
            INIT_39 => X"ffffffffffffffffffffffe6ffffffffffffffe9fffffffffffffffeffffffff",
            INIT_3A => X"0000000d00000000000000010000000000000018000000000000000a00000000",
            INIT_3B => X"00000018000000000000000700000000fffffffdffffffffffffffd9ffffffff",
            INIT_3C => X"fffffffdffffffff00000009000000000000000a000000000000001100000000",
            INIT_3D => X"fffffff8ffffffff0000000b000000000000000000000000ffffffedffffffff",
            INIT_3E => X"ffffffccffffffffffffffd2ffffffff0000003700000000ffffffebffffffff",
            INIT_3F => X"0000000a0000000000000007000000000000000200000000fffffff6ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffdbfffffffffffffff8ffffffff00000015000000000000001100000000",
            INIT_41 => X"0000002300000000fffffffbffffffffffffffd6ffffffffffffffeaffffffff",
            INIT_42 => X"00000026000000000000001a00000000ffffffd5ffffffffffffffe5ffffffff",
            INIT_43 => X"fffffff6ffffffff0000000e0000000000000014000000000000001200000000",
            INIT_44 => X"fffffff7ffffffff0000000600000000fffffff5ffffffffffffffefffffffff",
            INIT_45 => X"ffffffe4ffffffff00000007000000000000000e00000000fffffff5ffffffff",
            INIT_46 => X"0000000c00000000fffffff6ffffffffffffffefffffffff0000001000000000",
            INIT_47 => X"0000000500000000ffffffebfffffffffffffffbffffffff0000001300000000",
            INIT_48 => X"00000019000000000000001400000000fffffff4ffffffffffffffeeffffffff",
            INIT_49 => X"00000000000000000000000900000000fffffff7ffffffffffffffd4ffffffff",
            INIT_4A => X"0000001b00000000000000010000000000000018000000000000001300000000",
            INIT_4B => X"fffffff1ffffffff000000010000000000000015000000000000000100000000",
            INIT_4C => X"ffffffccfffffffffffffff7ffffffffffffffe3ffffffff0000000d00000000",
            INIT_4D => X"fffffff6ffffffff00000010000000000000001200000000ffffffc7ffffffff",
            INIT_4E => X"fffffff0fffffffffffffffefffffffffffffff8ffffffffffffffedffffffff",
            INIT_4F => X"00000000000000000000002800000000ffffffecffffffff0000001000000000",
            INIT_50 => X"fffffff8ffffffff0000000300000000fffffff1ffffffff0000000400000000",
            INIT_51 => X"00000028000000000000001c000000000000000c000000000000000a00000000",
            INIT_52 => X"00000005000000000000000e00000000ffffffd4ffffffff0000000900000000",
            INIT_53 => X"ffffffdaffffffff0000000f000000000000000600000000fffffff7ffffffff",
            INIT_54 => X"0000000000000000ffffffe7ffffffff0000000c000000000000001400000000",
            INIT_55 => X"fffffff3ffffffff0000000900000000fffffffeffffffff0000001200000000",
            INIT_56 => X"0000000a000000000000000200000000fffffffbffffffff0000001200000000",
            INIT_57 => X"0000001400000000fffffff0ffffffff0000001500000000ffffffeaffffffff",
            INIT_58 => X"0000001c000000000000001600000000ffffffeefffffffffffffff7ffffffff",
            INIT_59 => X"00000005000000000000000700000000fffffffcfffffffffffffffcffffffff",
            INIT_5A => X"ffffffddfffffffffffffff7fffffffffffffff5ffffffffffffffd7ffffffff",
            INIT_5B => X"fffffff5ffffffff0000000d000000000000000e00000000fffffffaffffffff",
            INIT_5C => X"ffffffefffffffff0000000000000000ffffffdeffffffff0000000e00000000",
            INIT_5D => X"fffffff2ffffffff0000000e000000000000001300000000fffffff4ffffffff",
            INIT_5E => X"0000000000000000fffffff2ffffffff0000000400000000fffffff4ffffffff",
            INIT_5F => X"fffffff7fffffffffffffffbffffffff0000000600000000ffffffd2ffffffff",
            INIT_60 => X"fffffff3ffffffffffffffdcfffffffffffffffffffffffffffffff4ffffffff",
            INIT_61 => X"0000001c00000000ffffffe2ffffffff0000000c000000000000001500000000",
            INIT_62 => X"ffffffe5ffffffffffffffe2ffffffffffffffddffffffffffffffffffffffff",
            INIT_63 => X"0000000a000000000000001400000000fffffffaffffffff0000000100000000",
            INIT_64 => X"0000001300000000fffffff2ffffffff0000000600000000fffffffeffffffff",
            INIT_65 => X"ffffffe9fffffffffffffff7ffffffff0000002700000000ffffffeeffffffff",
            INIT_66 => X"ffffffebfffffffffffffffefffffffffffffff6ffffffff0000001c00000000",
            INIT_67 => X"00000022000000000000001b00000000ffffffcefffffffffffffff1ffffffff",
            INIT_68 => X"00000023000000000000000300000000ffffffcdfffffffffffffff5ffffffff",
            INIT_69 => X"fffffff4ffffffff0000001700000000fffffff7fffffffffffffff6ffffffff",
            INIT_6A => X"0000000600000000ffffffefffffffff0000003a000000000000001d00000000",
            INIT_6B => X"0000000000000000ffffffe6fffffffffffffffdfffffffffffffffcffffffff",
            INIT_6C => X"ffffffeefffffffffffffff2fffffffffffffff1ffffffff0000000b00000000",
            INIT_6D => X"ffffffe8fffffffffffffff0ffffffffffffffe9ffffffff0000000900000000",
            INIT_6E => X"0000001c00000000ffffffbaffffffff0000003100000000ffffffc6ffffffff",
            INIT_6F => X"ffffffc1ffffffff00000010000000000000000700000000fffffffbffffffff",
            INIT_70 => X"ffffffeaffffffffffffffc5fffffffffffffff5ffffffff0000001800000000",
            INIT_71 => X"fffffffbfffffffffffffff7ffffffff00000005000000000000001a00000000",
            INIT_72 => X"ffffffc4ffffffffffffffebffffffffffffffe5ffffffff0000001100000000",
            INIT_73 => X"ffffffb0ffffffff0000000100000000fffffff4ffffffff0000000a00000000",
            INIT_74 => X"00000020000000000000000e00000000fffffff9ffffffff0000001500000000",
            INIT_75 => X"ffffffecffffffffffffffddffffffff00000032000000000000001e00000000",
            INIT_76 => X"00000030000000000000001a00000000ffffffbdffffffff0000001100000000",
            INIT_77 => X"ffffffb7ffffffff0000000500000000fffffff5fffffffffffffffdffffffff",
            INIT_78 => X"0000002c00000000ffffffefffffffffffffffebfffffffffffffff4ffffffff",
            INIT_79 => X"00000000000000000000000e00000000ffffffe5ffffffff0000000100000000",
            INIT_7A => X"0000000300000000ffffffd0ffffffff00000001000000000000000f00000000",
            INIT_7B => X"0000001a000000000000000300000000fffffffeffffffff0000001200000000",
            INIT_7C => X"0000001700000000ffffffffffffffff0000001100000000ffffffd8ffffffff",
            INIT_7D => X"ffffffeefffffffffffffff5ffffffffffffffdaffffffffffffffe2ffffffff",
            INIT_7E => X"00000059000000000000000c000000000000001700000000ffffffd6ffffffff",
            INIT_7F => X"ffffffc4ffffffff0000000d0000000000000009000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE3;


    MEM_IWGHT_LAYER3_INSTANCE4 : if BRAM_NAME = "iwght_layer3_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffdbffffffffffffffe9fffffffffffffff1ffffffff0000001b00000000",
            INIT_01 => X"ffffffd6ffffffff00000033000000000000000200000000ffffffeeffffffff",
            INIT_02 => X"ffffffdbfffffffffffffff3ffffffff0000000300000000ffffffeaffffffff",
            INIT_03 => X"ffffffd6ffffffff000000040000000000000005000000000000000a00000000",
            INIT_04 => X"00000013000000000000000b0000000000000011000000000000001f00000000",
            INIT_05 => X"ffffffeaffffffffffffffefffffffff00000017000000000000000b00000000",
            INIT_06 => X"0000001d0000000000000010000000000000000500000000fffffff2ffffffff",
            INIT_07 => X"ffffffceffffffff00000012000000000000000e00000000fffffffaffffffff",
            INIT_08 => X"00000010000000000000000000000000ffffffedffffffffffffffefffffffff",
            INIT_09 => X"fffffffbffffffff0000001200000000fffffff5ffffffff0000003300000000",
            INIT_0A => X"0000001500000000ffffffe2ffffffffffffffd2ffffffff0000000900000000",
            INIT_0B => X"fffffffffffffffffffffff8ffffffff0000001f000000000000001b00000000",
            INIT_0C => X"fffffff4ffffffff000000100000000000000003000000000000000900000000",
            INIT_0D => X"000000020000000000000009000000000000000000000000ffffffdcffffffff",
            INIT_0E => X"00000013000000000000001f000000000000000000000000ffffffdeffffffff",
            INIT_0F => X"ffffffd2ffffffff0000001300000000fffffff0ffffffff0000001500000000",
            INIT_10 => X"ffffffd5ffffffffffffffe6ffffffff0000000000000000fffffff0ffffffff",
            INIT_11 => X"00000007000000000000000000000000ffffffe8fffffffffffffff7ffffffff",
            INIT_12 => X"ffffffffffffffffffffffecfffffffffffffffbffffffffffffffebffffffff",
            INIT_13 => X"0000000900000000fffffff0fffffffffffffff3ffffffff0000000e00000000",
            INIT_14 => X"fffffffbffffffff00000001000000000000000a00000000fffffff2ffffffff",
            INIT_15 => X"0000000300000000ffffffe2fffffffffffffffdffffffff0000000f00000000",
            INIT_16 => X"ffffffe5ffffffff00000000000000000000000b000000000000000100000000",
            INIT_17 => X"fffffff5ffffffff0000003600000000ffffffc8fffffffffffffff1ffffffff",
            INIT_18 => X"ffffffedffffffff0000000e00000000fffffffcffffffff0000000200000000",
            INIT_19 => X"ffffffe5fffffffffffffff0ffffffffffffffe9ffffffff0000002700000000",
            INIT_1A => X"00000015000000000000000c000000000000000600000000fffffff7ffffffff",
            INIT_1B => X"fffffffbffffffff0000000d000000000000001b00000000ffffffd5ffffffff",
            INIT_1C => X"000000280000000000000000000000000000001e00000000fffffffaffffffff",
            INIT_1D => X"0000000100000000fffffff6ffffffffffffffd1ffffffff0000001800000000",
            INIT_1E => X"0000001000000000fffffff9ffffffff0000002b00000000fffffff9ffffffff",
            INIT_1F => X"ffffffefffffffff0000000a0000000000000004000000000000000800000000",
            INIT_20 => X"ffffffdcfffffffffffffffbffffffff0000000a000000000000000000000000",
            INIT_21 => X"ffffffecffffffffffffffd4ffffffffffffffeffffffffffffffff4ffffffff",
            INIT_22 => X"ffffffc8ffffffffffffffe9ffffffff00000009000000000000000800000000",
            INIT_23 => X"ffffffdfffffffffffffffedffffffffffffffecfffffffffffffff6ffffffff",
            INIT_24 => X"fffffff0fffffffffffffff2fffffffffffffff9fffffffffffffff1ffffffff",
            INIT_25 => X"000000000000000000000006000000000000000000000000fffffffcffffffff",
            INIT_26 => X"00000011000000000000001a00000000ffffffe5ffffffffffffffe9ffffffff",
            INIT_27 => X"ffffffe7ffffffff0000000a000000000000001900000000ffffffedffffffff",
            INIT_28 => X"00000012000000000000001600000000fffffff1fffffffffffffffeffffffff",
            INIT_29 => X"0000000c00000000fffffffaffffffff0000000500000000fffffffcffffffff",
            INIT_2A => X"fffffff5ffffffffffffffd8ffffffffffffffe9fffffffffffffff0ffffffff",
            INIT_2B => X"0000002d00000000fffffff2ffffffff0000000d00000000fffffff2ffffffff",
            INIT_2C => X"000000310000000000000021000000000000000800000000fffffffbffffffff",
            INIT_2D => X"0000000a000000000000001600000000ffffffebffffffff0000002400000000",
            INIT_2E => X"ffffffd5ffffffffffffffaeffffffffffffffe7ffffffffffffffffffffffff",
            INIT_2F => X"0000002c00000000ffffffe1ffffffff0000001100000000fffffffaffffffff",
            INIT_30 => X"ffffffd5ffffffffffffffdaffffffffffffffefffffffffffffffdeffffffff",
            INIT_31 => X"fffffff9ffffffffffffffedffffffffffffffcdffffffff0000000100000000",
            INIT_32 => X"ffffffc9fffffffffffffffefffffffffffffffaffffffff0000001900000000",
            INIT_33 => X"0000001000000000ffffffecfffffffffffffff5ffffffff0000001e00000000",
            INIT_34 => X"0000001d000000000000000600000000fffffff1ffffffff0000000600000000",
            INIT_35 => X"ffffffffffffffff000000080000000000000006000000000000001300000000",
            INIT_36 => X"ffffffeaffffffff0000004900000000ffffffefffffffffffffffedffffffff",
            INIT_37 => X"ffffffe7ffffffff0000002300000000fffffff5ffffffffffffffddffffffff",
            INIT_38 => X"fffffff3ffffffffffffffedffffffff0000001100000000fffffff0ffffffff",
            INIT_39 => X"000000090000000000000003000000000000000e000000000000000e00000000",
            INIT_3A => X"fffffffaffffffffffffffdcffffffffffffffcdffffffff0000000900000000",
            INIT_3B => X"fffffffefffffffffffffff8ffffffff0000001f000000000000001b00000000",
            INIT_3C => X"00000007000000000000001e000000000000001500000000fffffff3ffffffff",
            INIT_3D => X"0000000900000000fffffff4ffffffffffffffe2ffffffff0000001600000000",
            INIT_3E => X"00000001000000000000002300000000fffffff8ffffffffffffffe8ffffffff",
            INIT_3F => X"0000001000000000fffffffeffffffffffffffffffffffff0000000400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe8fffffffffffffff1ffffffffffffffeeffffffffffffffdbffffffff",
            INIT_41 => X"fffffff3fffffffffffffff0ffffffffffffffc3ffffffff0000000a00000000",
            INIT_42 => X"fffffff0ffffffffffffffd3ffffffffffffffe4ffffffff0000001a00000000",
            INIT_43 => X"ffffffe0ffffffff0000003000000000ffffffefffffffffffffffe9ffffffff",
            INIT_44 => X"fffffffaffffffff0000002b000000000000000300000000fffffff4ffffffff",
            INIT_45 => X"ffffffdcffffffffffffffefffffffff0000001300000000fffffffeffffffff",
            INIT_46 => X"0000000d000000000000000d0000000000000011000000000000002000000000",
            INIT_47 => X"00000013000000000000000e000000000000000100000000ffffffefffffffff",
            INIT_48 => X"fffffff5ffffffff00000000000000000000001a00000000ffffffdcffffffff",
            INIT_49 => X"ffffffebffffffff0000000100000000fffffff7ffffffffffffffe4ffffffff",
            INIT_4A => X"fffffffbffffffffffffffe8ffffffffffffffc6fffffffffffffff4ffffffff",
            INIT_4B => X"0000003d000000000000001f00000000fffffff8ffffffff0000000000000000",
            INIT_4C => X"ffffffcbffffffffffffffc7ffffffffffffffddffffffffffffffa2ffffffff",
            INIT_4D => X"0000000e00000000ffffffe3ffffffffffffffe4ffffffff0000001d00000000",
            INIT_4E => X"0000000700000000fffffff4ffffffff00000010000000000000001100000000",
            INIT_4F => X"00000016000000000000000000000000fffffff9ffffffffffffffeeffffffff",
            INIT_50 => X"00000018000000000000002a00000000ffffffe8ffffffff0000002200000000",
            INIT_51 => X"fffffff9ffffffff0000001000000000fffffff9ffffffffffffffd8ffffffff",
            INIT_52 => X"0000000200000000ffffffd6fffffffffffffff7fffffffffffffff8ffffffff",
            INIT_53 => X"00000014000000000000001800000000fffffff4ffffffffffffffc8ffffffff",
            INIT_54 => X"ffffffe5fffffffffffffffbfffffffffffffff8ffffffff0000002300000000",
            INIT_55 => X"ffffffdaffffffff00000003000000000000002f000000000000003400000000",
            INIT_56 => X"0000003100000000ffffffd1ffffffff0000001300000000ffffffe9ffffffff",
            INIT_57 => X"ffffffbfffffffffffffffbfffffffffffffffecffffffffffffffd3ffffffff",
            INIT_58 => X"fffffffdffffffff0000001900000000ffffffdeffffffffffffffdfffffffff",
            INIT_59 => X"0000001200000000ffffffe7ffffffffffffffeffffffffffffffff4ffffffff",
            INIT_5A => X"fffffff2ffffffffffffffc8fffffffffffffffcfffffffffffffff8ffffffff",
            INIT_5B => X"fffffffeffffffff0000000b0000000000000027000000000000000800000000",
            INIT_5C => X"ffffffd3ffffffffffffffc2ffffffffffffffb7ffffffffffffffb9ffffffff",
            INIT_5D => X"0000000300000000ffffffeaffffffffffffffd7ffffffff0000000500000000",
            INIT_5E => X"0000001500000000ffffffd5fffffffffffffff2fffffffffffffffaffffffff",
            INIT_5F => X"fffffff9ffffffff0000000d00000000fffffff8ffffffffffffffd3ffffffff",
            INIT_60 => X"0000000b000000000000003900000000ffffffc8fffffffffffffffbffffffff",
            INIT_61 => X"ffffffd8ffffffff00000023000000000000003e00000000ffffffdbffffffff",
            INIT_62 => X"00000007000000000000001300000000fffffff5ffffffffffffffeaffffffff",
            INIT_63 => X"fffffffdffffffff0000000d000000000000000000000000ffffffb3ffffffff",
            INIT_64 => X"0000001400000000ffffffc5fffffffffffffff5ffffffffffffffe9ffffffff",
            INIT_65 => X"ffffffdaffffffff00000002000000000000002a00000000fffffff4ffffffff",
            INIT_66 => X"0000001400000000ffffffffffffffffffffffeeffffffffffffffd7ffffffff",
            INIT_67 => X"ffffffc0ffffffffffffffe4ffffffff00000016000000000000000400000000",
            INIT_68 => X"0000001700000000ffffffedfffffffffffffff4ffffffffffffffc5ffffffff",
            INIT_69 => X"ffffffe8ffffffff00000006000000000000000b000000000000001600000000",
            INIT_6A => X"0000000500000000fffffff5ffffffff00000025000000000000000000000000",
            INIT_6B => X"00000004000000000000000100000000ffffffddffffffff0000001400000000",
            INIT_6C => X"0000000d00000000ffffffdeffffffffffffffddffffffffffffffadffffffff",
            INIT_6D => X"0000001600000000fffffff5ffffffffffffffccffffffff0000002e00000000",
            INIT_6E => X"00000040000000000000002600000000ffffffecfffffffffffffffdffffffff",
            INIT_6F => X"0000000300000000ffffffe5ffffffff0000000500000000ffffffb3ffffffff",
            INIT_70 => X"fffffffbffffffff0000000300000000ffffffcbfffffffffffffff9ffffffff",
            INIT_71 => X"ffffff83ffffffff000000210000000000000015000000000000000b00000000",
            INIT_72 => X"0000000500000000fffffff3ffffffff0000000400000000ffffffe6ffffffff",
            INIT_73 => X"0000002e000000000000000a00000000ffffffebffffffffffffffccffffffff",
            INIT_74 => X"ffffffb6ffffffff000000180000000000000019000000000000000500000000",
            INIT_75 => X"0000000000000000ffffffedffffffff0000000d000000000000001300000000",
            INIT_76 => X"fffffff3ffffffffffffffe7ffffffff0000001400000000ffffffd3ffffffff",
            INIT_77 => X"00000011000000000000001c00000000ffffffdfffffffff0000001000000000",
            INIT_78 => X"fffffffdffffffff00000017000000000000002f000000000000000c00000000",
            INIT_79 => X"ffffffe4ffffffff000000120000000000000005000000000000002700000000",
            INIT_7A => X"0000000c00000000ffffffdefffffffffffffff6ffffffffffffffeaffffffff",
            INIT_7B => X"0000000e00000000ffffffe0ffffffff0000001f00000000fffffffeffffffff",
            INIT_7C => X"0000001200000000ffffffd9fffffffffffffffdffffffffffffffd5ffffffff",
            INIT_7D => X"00000009000000000000001700000000ffffffeeffffffff0000000300000000",
            INIT_7E => X"ffffffe8ffffffffffffffb6ffffffffffffffe6ffffffff0000001100000000",
            INIT_7F => X"0000002d00000000fffffff4fffffffffffffffbffffffff0000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE4;


    MEM_IWGHT_LAYER3_INSTANCE5 : if BRAM_NAME = "iwght_layer3_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001b0000000000000041000000000000000600000000ffffffceffffffff",
            INIT_01 => X"0000002400000000ffffffe9fffffffffffffff2ffffffff0000001000000000",
            INIT_02 => X"0000000b000000000000001b00000000ffffffbeffffffff0000000700000000",
            INIT_03 => X"0000000a00000000ffffffb0ffffffff00000007000000000000003800000000",
            INIT_04 => X"0000002d00000000ffffffa6fffffffffffffffcffffffff0000001300000000",
            INIT_05 => X"ffffffd8ffffffff0000002000000000fffffffcfffffffffffffff6ffffffff",
            INIT_06 => X"0000000000000000ffffffe9ffffffffffffffddffffffff0000000900000000",
            INIT_07 => X"ffffffe6ffffffff0000001300000000ffffffdaffffffff0000003c00000000",
            INIT_08 => X"000000170000000000000018000000000000003f000000000000001600000000",
            INIT_09 => X"0000000600000000fffffff0ffffffffffffffedffffffff0000000400000000",
            INIT_0A => X"0000000a00000000000000010000000000000008000000000000000000000000",
            INIT_0B => X"ffffffecffffffff0000000800000000ffffffd8ffffffffffffffd2ffffffff",
            INIT_0C => X"ffffffe3ffffffffffffffecffffffffffffffddffffffffffffffd9ffffffff",
            INIT_0D => X"0000001800000000fffffff2ffffffff0000000700000000ffffffeaffffffff",
            INIT_0E => X"ffffffe4ffffffffffffffd5ffffffffffffffedffffffffffffffdbffffffff",
            INIT_0F => X"ffffffeaffffffff0000001800000000fffffff0fffffffffffffff4ffffffff",
            INIT_10 => X"fffffff1ffffffffffffffd8ffffffff00000028000000000000000b00000000",
            INIT_11 => X"0000001200000000fffffff0fffffffffffffff6ffffffff0000000b00000000",
            INIT_12 => X"0000001200000000fffffff7ffffffffffffffc8ffffffffffffffd9ffffffff",
            INIT_13 => X"00000020000000000000000000000000fffffff4ffffffff0000002c00000000",
            INIT_14 => X"0000001700000000ffffffc8ffffffff00000013000000000000002000000000",
            INIT_15 => X"fffffffeffffffff0000001100000000ffffffe7ffffffffffffffd8ffffffff",
            INIT_16 => X"00000006000000000000001900000000ffffffebffffffff0000002500000000",
            INIT_17 => X"ffffffebfffffffffffffff6fffffffffffffff1ffffffff0000001100000000",
            INIT_18 => X"0000000d00000000fffffff3ffffffff0000005400000000ffffffc7ffffffff",
            INIT_19 => X"0000001d000000000000000d0000000000000013000000000000000900000000",
            INIT_1A => X"0000001f000000000000003300000000ffffffd7ffffffff0000001000000000",
            INIT_1B => X"ffffffdaffffffffffffffebffffffffffffffffffffffffffffffefffffffff",
            INIT_1C => X"ffffffefffffffffffffffeeffffffffffffffcffffffffffffffff1ffffffff",
            INIT_1D => X"fffffffeffffffff0000000000000000ffffffffffffffffffffffe8ffffffff",
            INIT_1E => X"ffffffd5ffffffffffffffe8ffffffffffffffe4ffffffff0000001400000000",
            INIT_1F => X"0000003100000000ffffffd5ffffffff00000015000000000000000800000000",
            INIT_20 => X"0000001b000000000000000c000000000000000d000000000000002300000000",
            INIT_21 => X"ffffffc8ffffffff0000001f00000000fffffff9ffffffff0000001c00000000",
            INIT_22 => X"fffffffeffffffff000000280000000000000003000000000000001c00000000",
            INIT_23 => X"000000240000000000000025000000000000001300000000ffffffd3ffffffff",
            INIT_24 => X"fffffff0ffffffffffffffe4ffffffff00000011000000000000001300000000",
            INIT_25 => X"0000003100000000ffffffe7ffffffff00000021000000000000001200000000",
            INIT_26 => X"000000170000000000000000000000000000000e00000000fffffff6ffffffff",
            INIT_27 => X"00000015000000000000001c00000000ffffffefffffffff0000000f00000000",
            INIT_28 => X"0000000900000000fffffff6ffffffff0000002200000000ffffffd6ffffffff",
            INIT_29 => X"0000002700000000ffffffffffffffff00000004000000000000001600000000",
            INIT_2A => X"ffffffe8ffffffff0000001800000000ffffffe0fffffffffffffff3ffffffff",
            INIT_2B => X"0000001a000000000000001c000000000000000f00000000ffffffc0ffffffff",
            INIT_2C => X"0000001900000000ffffffd3ffffffff0000000500000000fffffffeffffffff",
            INIT_2D => X"ffffffffffffffff0000000900000000ffffffa7ffffffff0000000700000000",
            INIT_2E => X"0000001700000000ffffffdbffffffffffffffe5ffffffff0000002e00000000",
            INIT_2F => X"fffffff5fffffffffffffff1ffffffff0000000a000000000000001500000000",
            INIT_30 => X"0000002100000000ffffffd1ffffffffffffffd4fffffffffffffff9ffffffff",
            INIT_31 => X"ffffffbfffffffff0000002e000000000000000300000000ffffffd9ffffffff",
            INIT_32 => X"00000017000000000000003100000000ffffffe4ffffffff0000000f00000000",
            INIT_33 => X"fffffff1ffffffffffffffbffffffffffffffff4ffffffff0000000e00000000",
            INIT_34 => X"ffffffe8ffffffffffffffeeffffffff00000015000000000000002800000000",
            INIT_35 => X"000000130000000000000016000000000000002f000000000000001700000000",
            INIT_36 => X"0000003400000000ffffffe2ffffffffffffffdbffffffff0000001e00000000",
            INIT_37 => X"fffffff6fffffffffffffff9ffffffffffffffc3ffffffffffffffcaffffffff",
            INIT_38 => X"0000001500000000ffffffedffffffff0000001c000000000000000200000000",
            INIT_39 => X"fffffffcffffffff0000000a000000000000000b000000000000000300000000",
            INIT_3A => X"0000002800000000ffffffeeffffffffffffffbdffffffff0000001b00000000",
            INIT_3B => X"ffffffe7ffffffff0000000d000000000000000c00000000ffffffdbffffffff",
            INIT_3C => X"0000001800000000fffffffcffffffff0000002500000000fffffffdffffffff",
            INIT_3D => X"ffffffe1ffffffff0000003e00000000ffffffafffffffffffffffd1ffffffff",
            INIT_3E => X"ffffffe1ffffffffffffffe6ffffffff00000021000000000000003c00000000",
            INIT_3F => X"fffffff3ffffffff00000014000000000000000900000000fffffff1ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffb3ffffffffffffffe8ffffffffffffffd8fffffffffffffff6ffffffff",
            INIT_41 => X"fffffffcffffffff0000001d00000000fffffff8fffffffffffffff4ffffffff",
            INIT_42 => X"ffffffbcffffffff0000001a00000000ffffffebffffffff0000001000000000",
            INIT_43 => X"0000000a000000000000000500000000fffffff0ffffffffffffffefffffffff",
            INIT_44 => X"ffffffcefffffffffffffffbffffffffffffffeeffffffff0000000500000000",
            INIT_45 => X"0000001800000000ffffffdcffffffff0000002d000000000000000e00000000",
            INIT_46 => X"0000001a00000000000000160000000000000016000000000000001a00000000",
            INIT_47 => X"ffffffcefffffffffffffff2ffffffffffffffe8ffffffff0000002000000000",
            INIT_48 => X"0000001600000000ffffffeeffffffff00000037000000000000000e00000000",
            INIT_49 => X"00000026000000000000000900000000fffffff3ffffffffffffffdfffffffff",
            INIT_4A => X"0000003000000000fffffff8ffffffffffffff9affffffff0000001500000000",
            INIT_4B => X"ffffffebffffffffffffffe5ffffffffffffffedffffffffffffffe1ffffffff",
            INIT_4C => X"0000000200000000ffffffeeffffffff00000029000000000000000200000000",
            INIT_4D => X"fffffffafffffffffffffffbffffffffffffffcaffffffffffffffd8ffffffff",
            INIT_4E => X"ffffffd2ffffffff0000002800000000fffffff6ffffffff0000003a00000000",
            INIT_4F => X"00000011000000000000000e00000000fffffff8ffffffff0000000300000000",
            INIT_50 => X"ffffffeeffffffff0000000c00000000ffffffecffffffff0000003e00000000",
            INIT_51 => X"fffffff4ffffffff00000003000000000000001a000000000000000500000000",
            INIT_52 => X"00000011000000000000001a00000000ffffffe7ffffffff0000001300000000",
            INIT_53 => X"0000001b00000000ffffffdafffffffffffffffdffffffff0000001800000000",
            INIT_54 => X"0000000200000000ffffffdfffffffff0000000600000000ffffffe1ffffffff",
            INIT_55 => X"fffffff4ffffffffffffffedffffffffffffffeefffffffffffffffeffffffff",
            INIT_56 => X"fffffff2ffffffff0000000c00000000ffffffccffffffffffffffdeffffffff",
            INIT_57 => X"ffffffebffffffffffffffedffffffffffffffcdffffffff0000000400000000",
            INIT_58 => X"00000016000000000000001000000000fffffff6ffffffff0000000900000000",
            INIT_59 => X"ffffffbbffffffff00000000000000000000000600000000ffffffc6ffffffff",
            INIT_5A => X"ffffffdaffffffff0000001c000000000000000b00000000fffffff3ffffffff",
            INIT_5B => X"ffffffebffffffffffffffeaffffffffffffffddffffffff0000002200000000",
            INIT_5C => X"00000019000000000000001900000000fffffff7ffffffff0000003a00000000",
            INIT_5D => X"fffffff1ffffffff00000000000000000000001300000000ffffffefffffffff",
            INIT_5E => X"ffffffbbffffffffffffffbcffffffff0000002900000000fffffff3ffffffff",
            INIT_5F => X"ffffffdbffffffff000000110000000000000009000000000000000000000000",
            INIT_60 => X"fffffff8ffffffffffffffe9ffffffffffffffedffffffff0000003e00000000",
            INIT_61 => X"0000002a0000000000000012000000000000000a000000000000003800000000",
            INIT_62 => X"0000002d000000000000001f00000000ffffffdaffffffff0000001000000000",
            INIT_63 => X"0000001900000000fffffffbffffffff0000000a000000000000002400000000",
            INIT_64 => X"0000002400000000fffffffaffffffff0000000400000000ffffffffffffffff",
            INIT_65 => X"0000000000000000ffffffddffffffffffffffcaffffffffffffffe5ffffffff",
            INIT_66 => X"ffffffd8ffffffff0000000400000000ffffffcdffffffff0000000600000000",
            INIT_67 => X"0000000800000000ffffffefffffffffffffffc5ffffffff0000000500000000",
            INIT_68 => X"0000000f00000000fffffff0ffffffff0000003d000000000000001700000000",
            INIT_69 => X"fffffffeffffffff0000001600000000ffffffeaffffffffffffffefffffffff",
            INIT_6A => X"ffffffd0ffffffff0000002400000000ffffffd9ffffffff0000000d00000000",
            INIT_6B => X"0000000c0000000000000001000000000000000c000000000000003900000000",
            INIT_6C => X"ffffffe8ffffffff000000250000000000000001000000000000000e00000000",
            INIT_6D => X"00000007000000000000000900000000fffffff5ffffffff0000000200000000",
            INIT_6E => X"fffffff8ffffffff0000003d000000000000000b00000000ffffffbeffffffff",
            INIT_6F => X"fffffffaffffffff0000001b00000000fffffffdffffffffffffffdcffffffff",
            INIT_70 => X"00000012000000000000000000000000ffffffe8ffffffff0000002800000000",
            INIT_71 => X"0000002100000000fffffff5ffffffff0000000b000000000000001000000000",
            INIT_72 => X"00000013000000000000000000000000ffffffc7ffffffff0000001700000000",
            INIT_73 => X"ffffffebffffffff0000003b0000000000000004000000000000001d00000000",
            INIT_74 => X"0000001d000000000000000000000000fffffff9ffffffffffffffdcffffffff",
            INIT_75 => X"fffffffeffffffff0000001c00000000ffffffd3ffffffff0000001700000000",
            INIT_76 => X"fffffff4ffffffff0000002000000000ffffffc9fffffffffffffffdffffffff",
            INIT_77 => X"0000002200000000fffffffffffffffffffffff5ffffffff0000000100000000",
            INIT_78 => X"00000004000000000000000b000000000000003f00000000ffffffe7ffffffff",
            INIT_79 => X"0000001500000000fffffff3ffffffff00000000000000000000000200000000",
            INIT_7A => X"fffffff5ffffffff0000000c00000000ffffffdffffffffffffffff1ffffffff",
            INIT_7B => X"0000001400000000ffffffe2ffffffff0000001600000000ffffffd1ffffffff",
            INIT_7C => X"ffffffefffffffff000000050000000000000024000000000000000c00000000",
            INIT_7D => X"fffffffbffffffff0000001100000000fffffffdffffffffffffffe6ffffffff",
            INIT_7E => X"00000036000000000000000800000000ffffffffffffffffffffffe6ffffffff",
            INIT_7F => X"ffffffecffffffff0000000700000000ffffffeeffffffff0000000300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE5;


    MEM_IWGHT_LAYER3_INSTANCE6 : if BRAM_NAME = "iwght_layer3_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffcffffffffffffffeafffffffffffffffdffffffff0000001600000000",
            INIT_01 => X"0000003f000000000000000600000000ffffffd1ffffffff0000000100000000",
            INIT_02 => X"0000000a000000000000000000000000fffffff6ffffffffffffffbfffffffff",
            INIT_03 => X"0000000600000000fffffff9ffffffff0000001300000000ffffffd8ffffffff",
            INIT_04 => X"ffffffe9ffffffffffffffe2ffffffff0000000800000000fffffffcffffffff",
            INIT_05 => X"0000000400000000fffffffeffffffff0000000b00000000fffffff8ffffffff",
            INIT_06 => X"0000000c00000000ffffffd8fffffffffffffff0fffffffffffffffdffffffff",
            INIT_07 => X"ffffffcafffffffffffffffaffffffffffffffb6ffffffffffffffe8ffffffff",
            INIT_08 => X"0000000e00000000ffffffe8ffffffffffffffe1ffffffffffffffedffffffff",
            INIT_09 => X"fffffff5ffffffff0000001700000000ffffffefffffffffffffffffffffffff",
            INIT_0A => X"0000002000000000fffffff2fffffffffffffffafffffffffffffff9ffffffff",
            INIT_0B => X"ffffffe9ffffffffffffffdffffffffffffffff4fffffffffffffff4ffffffff",
            INIT_0C => X"0000001a000000000000001700000000ffffffdeffffffff0000001400000000",
            INIT_0D => X"ffffffe6ffffffff00000020000000000000000700000000ffffffd7ffffffff",
            INIT_0E => X"fffffffeffffffffffffffc5ffffffff0000003a000000000000001800000000",
            INIT_0F => X"ffffffcbffffffff0000000c00000000ffffffe8ffffffff0000002100000000",
            INIT_10 => X"ffffffb1ffffffffffffffd9ffffffffffffffe5fffffffffffffff7ffffffff",
            INIT_11 => X"fffffff5fffffffffffffff3ffffffffffffffe4ffffffff0000000800000000",
            INIT_12 => X"fffffff7fffffffffffffffeffffffffffffffacffffffff0000002600000000",
            INIT_13 => X"ffffffb9ffffffffffffffebffffffff0000000600000000ffffffe3ffffffff",
            INIT_14 => X"000000200000000000000001000000000000000f00000000ffffffe9ffffffff",
            INIT_15 => X"ffffffd6ffffffff00000015000000000000001900000000fffffff3ffffffff",
            INIT_16 => X"fffffff2ffffffffffffffd9ffffffffffffffd2ffffffff0000003400000000",
            INIT_17 => X"ffffffebffffffff0000000a00000000ffffffdcffffffff0000000200000000",
            INIT_18 => X"0000002f00000000ffffffeffffffffffffffffbffffffff0000003700000000",
            INIT_19 => X"0000002c0000000000000011000000000000000d000000000000002000000000",
            INIT_1A => X"0000000500000000ffffffb7fffffffffffffff2ffffffffffffffe6ffffffff",
            INIT_1B => X"0000001800000000000000070000000000000006000000000000001000000000",
            INIT_1C => X"0000001d00000000ffffffe1fffffffffffffffbfffffffffffffff9ffffffff",
            INIT_1D => X"fffffffcffffffff00000010000000000000002700000000fffffff5ffffffff",
            INIT_1E => X"0000002b000000000000000f00000000ffffffecffffffffffffffb1ffffffff",
            INIT_1F => X"0000002800000000fffffff3ffffffffffffffe9ffffffffffffffdfffffffff",
            INIT_20 => X"ffffffbeffffffffffffffb5fffffffffffffff0fffffffffffffff2ffffffff",
            INIT_21 => X"0000000f000000000000000000000000ffffffdcfffffffffffffffcffffffff",
            INIT_22 => X"fffffff9ffffffffffffffe9fffffffffffffff1fffffffffffffffaffffffff",
            INIT_23 => X"ffffffd2fffffffffffffffdffffffff00000007000000000000001200000000",
            INIT_24 => X"ffffffeffffffffffffffffcfffffffffffffff3fffffffffffffffeffffffff",
            INIT_25 => X"ffffffe9ffffffff0000000d000000000000001d000000000000001800000000",
            INIT_26 => X"fffffff5fffffffffffffff7ffffffffffffffe8ffffffff0000002c00000000",
            INIT_27 => X"fffffffdffffffff0000001800000000ffffffdbfffffffffffffff4ffffffff",
            INIT_28 => X"0000001d00000000ffffffeefffffffffffffff4ffffffffffffffd6ffffffff",
            INIT_29 => X"00000016000000000000001000000000fffffffeffffffff0000002100000000",
            INIT_2A => X"0000002200000000ffffffbaffffffffffffffa0ffffffff0000000600000000",
            INIT_2B => X"ffffffebffffffff00000022000000000000001a00000000fffffff8ffffffff",
            INIT_2C => X"fffffffcffffffffffffffdfffffffffffffffebffffffff0000001900000000",
            INIT_2D => X"ffffffe2ffffffff00000006000000000000001100000000ffffffc5ffffffff",
            INIT_2E => X"fffffffeffffffff00000025000000000000001300000000ffffffedffffffff",
            INIT_2F => X"ffffffeeffffffff00000024000000000000001300000000fffffff3ffffffff",
            INIT_30 => X"fffffffdffffffffffffffdeffffffff0000000d00000000fffffff3ffffffff",
            INIT_31 => X"0000002b000000000000000b00000000ffffffc3ffffffffffffffbeffffffff",
            INIT_32 => X"ffffffc7ffffffff0000000300000000ffffffedffffffffffffffeeffffffff",
            INIT_33 => X"fffffff5fffffffffffffff4fffffffffffffffaffffffff0000000b00000000",
            INIT_34 => X"fffffff6fffffffffffffff3ffffffff00000005000000000000000800000000",
            INIT_35 => X"fffffffaffffffffffffffe9fffffffffffffffaffffffff0000001b00000000",
            INIT_36 => X"0000000600000000fffffff4ffffffffffffffe4ffffffff0000001a00000000",
            INIT_37 => X"fffffff2ffffffff0000001300000000ffffffe2fffffffffffffff2ffffffff",
            INIT_38 => X"fffffffaffffffffffffffeaffffffffffffffe0ffffffffffffffd7ffffffff",
            INIT_39 => X"ffffffd4ffffffff0000000d000000000000001200000000ffffffd8ffffffff",
            INIT_3A => X"fffffffdffffffff0000001200000000ffffffeeffffffff0000000900000000",
            INIT_3B => X"fffffff5ffffffffffffffe4ffffffff0000000c00000000ffffffdfffffffff",
            INIT_3C => X"00000023000000000000000d0000000000000010000000000000002600000000",
            INIT_3D => X"00000000000000000000000800000000ffffffe9ffffffff0000002d00000000",
            INIT_3E => X"fffffffaffffffffffffffcdffffffff00000024000000000000002700000000",
            INIT_3F => X"ffffffecfffffffffffffff4fffffffffffffff0ffffffff0000001300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffc8fffffffffffffffdffffffff0000002200000000ffffffc1ffffffff",
            INIT_41 => X"fffffff7fffffffffffffff1fffffffffffffff1ffffffff0000000600000000",
            INIT_42 => X"fffffff8fffffffffffffff7ffffffffffffffcdffffffff0000000300000000",
            INIT_43 => X"ffffffefffffffff0000000c000000000000001500000000ffffffebffffffff",
            INIT_44 => X"0000000900000000ffffffe1fffffffffffffffbffffffff0000000700000000",
            INIT_45 => X"0000001b00000000000000170000000000000020000000000000000500000000",
            INIT_46 => X"0000000b00000000ffffffe3ffffffff00000009000000000000000d00000000",
            INIT_47 => X"ffffffe6fffffffffffffff8ffffffffffffffbcffffffffffffffefffffffff",
            INIT_48 => X"000000060000000000000010000000000000000800000000ffffffddffffffff",
            INIT_49 => X"0000000200000000ffffffeeffffffff00000007000000000000001900000000",
            INIT_4A => X"fffffff5ffffffffffffffd8fffffffffffffff3ffffffffffffffedffffffff",
            INIT_4B => X"fffffffafffffffffffffff5ffffffffffffffefffffffffffffffbfffffffff",
            INIT_4C => X"ffffffddffffffff00000032000000000000001b000000000000000300000000",
            INIT_4D => X"ffffffe7ffffffff0000000800000000ffffffe8fffffffffffffffaffffffff",
            INIT_4E => X"ffffffdcffffffff0000000400000000ffffffffffffffff0000000500000000",
            INIT_4F => X"fffffff3ffffffffffffffecffffffff00000001000000000000000c00000000",
            INIT_50 => X"ffffffc2ffffffffffffffcffffffffffffffff6ffffffff0000000c00000000",
            INIT_51 => X"fffffffaffffffff0000000200000000ffffffb2ffffffffffffffe4ffffffff",
            INIT_52 => X"ffffff9efffffffffffffff2ffffffffffffffdaffffffff0000000500000000",
            INIT_53 => X"0000000000000000000000040000000000000008000000000000001000000000",
            INIT_54 => X"0000002700000000ffffffedffffffff00000005000000000000001600000000",
            INIT_55 => X"00000003000000000000000200000000ffffffffffffffff0000000500000000",
            INIT_56 => X"00000003000000000000001100000000ffffffe5ffffffff0000001400000000",
            INIT_57 => X"ffffffd6ffffffff0000001000000000ffffffd5ffffffffffffffe1ffffffff",
            INIT_58 => X"ffffffeffffffffffffffffdffffffffffffffe0ffffffffffffffd5ffffffff",
            INIT_59 => X"00000027000000000000000000000000fffffff8ffffffff0000002800000000",
            INIT_5A => X"fffffff9fffffffffffffffeffffffffffffffc0fffffffffffffffeffffffff",
            INIT_5B => X"0000000f00000000ffffffffffffffff0000002900000000ffffffe3ffffffff",
            INIT_5C => X"fffffff3ffffffff0000001d0000000000000018000000000000000b00000000",
            INIT_5D => X"ffffffdfffffffff0000000100000000fffffff3ffffffff0000000100000000",
            INIT_5E => X"ffffffd4ffffffffffffffedffffffffffffffffffffffff0000000d00000000",
            INIT_5F => X"ffffffbcffffffff0000000900000000fffffff8ffffffff0000000c00000000",
            INIT_60 => X"ffffffebffffffffffffffd1ffffffff0000000800000000ffffffe7ffffffff",
            INIT_61 => X"fffffffaffffffffffffffebffffffffffffffe3fffffffffffffff2ffffffff",
            INIT_62 => X"ffffffeeffffffff0000000000000000fffffff0ffffffff0000000e00000000",
            INIT_63 => X"00000010000000000000002e00000000ffffffedffffffffffffffb9ffffffff",
            INIT_64 => X"fffffffbffffffffffffffffffffffff0000000000000000ffffffddffffffff",
            INIT_65 => X"ffffffe5ffffffff00000007000000000000000c00000000fffffffcffffffff",
            INIT_66 => X"ffffffedffffffffffffffeaffffffffffffffd1fffffffffffffff6ffffffff",
            INIT_67 => X"0000000800000000ffffffe6ffffffffffffffb1ffffffffffffffe4ffffffff",
            INIT_68 => X"0000001000000000fffffffbffffffffffffffa3ffffffff0000002700000000",
            INIT_69 => X"fffffff6ffffffffffffffe6ffffffff0000001100000000ffffffd5ffffffff",
            INIT_6A => X"000000170000000000000013000000000000000a00000000ffffffe8ffffffff",
            INIT_6B => X"00000018000000000000002800000000fffffffcffffffffffffffe6ffffffff",
            INIT_6C => X"00000022000000000000000600000000ffffffffffffffffffffffe8ffffffff",
            INIT_6D => X"fffffffeffffffff0000000200000000ffffffe4ffffffffffffffb6ffffffff",
            INIT_6E => X"0000003400000000ffffffbaffffffffffffffd3ffffffffffffffe7ffffffff",
            INIT_6F => X"fffffff4ffffffff00000017000000000000001400000000ffffff84ffffffff",
            INIT_70 => X"ffffffeaffffffff0000002d00000000fffffff2ffffffff0000000000000000",
            INIT_71 => X"ffffffc8ffffffff000000280000000000000016000000000000000c00000000",
            INIT_72 => X"ffffffffffffffffffffffd1fffffffffffffffbffffffffffffffc4ffffffff",
            INIT_73 => X"ffffffffffffffff00000060000000000000000000000000ffffffb9ffffffff",
            INIT_74 => X"ffffffc1ffffffffffffffdffffffffffffffffbffffffff0000001200000000",
            INIT_75 => X"ffffffdcffffffff00000017000000000000002000000000ffffffecffffffff",
            INIT_76 => X"0000002d0000000000000039000000000000001700000000ffffffccffffffff",
            INIT_77 => X"ffffffffffffffff00000012000000000000002a000000000000000400000000",
            INIT_78 => X"00000012000000000000000900000000ffffffecffffffffffffffefffffffff",
            INIT_79 => X"0000000600000000fffffff2fffffffffffffffaffffffffffffffe2ffffffff",
            INIT_7A => X"0000000500000000ffffffe5ffffffff0000002c00000000fffffff8ffffffff",
            INIT_7B => X"fffffff2ffffffff0000002800000000fffffffcffffffffffffffd2ffffffff",
            INIT_7C => X"fffffffdffffffffffffffe8ffffffff0000000b00000000ffffffabffffffff",
            INIT_7D => X"0000000a00000000ffffffd9ffffffff0000003400000000ffffff9bffffffff",
            INIT_7E => X"ffffffd8ffffffffffffffcdffffffffffffffddffffffff0000003600000000",
            INIT_7F => X"fffffffafffffffffffffff8ffffffff0000000c000000000000001a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE6;


    MEM_IWGHT_LAYER3_INSTANCE7 : if BRAM_NAME = "iwght_layer3_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffffffffffffffffffffffbfffffffffffffffeffffffffffffffeeffffffff",
            INIT_01 => X"ffffffdcffffffff0000001500000000fffffffdfffffffffffffffcffffffff",
            INIT_02 => X"fffffff5ffffffffffffffe7fffffffffffffff8ffffffffffffffdbffffffff",
            INIT_03 => X"fffffff2ffffffff0000000000000000ffffffeafffffffffffffffaffffffff",
            INIT_04 => X"0000001e00000000ffffffdaffffffff00000013000000000000000200000000",
            INIT_05 => X"0000000700000000ffffffe5ffffffff0000001e000000000000001c00000000",
            INIT_06 => X"fffffffeffffffff0000002400000000ffffffc5ffffffffffffffbdffffffff",
            INIT_07 => X"fffffff1ffffffffffffffddffffffffffffffcdffffffff0000001800000000",
            INIT_08 => X"fffffffbffffffffffffffefffffffff00000000000000000000002600000000",
            INIT_09 => X"0000000f000000000000001400000000fffffff1ffffffffffffffcfffffffff",
            INIT_0A => X"0000000700000000ffffffdfffffffffffffffefffffffff0000001b00000000",
            INIT_0B => X"0000000a00000000fffffffdffffffff00000013000000000000001c00000000",
            INIT_0C => X"ffffffafffffffffffffffe7ffffffffffffffe0fffffffffffffff4ffffffff",
            INIT_0D => X"0000000c00000000ffffffedffffffffffffffe6ffffffffffffffa6ffffffff",
            INIT_0E => X"00000000000000000000002800000000ffffffdbffffffff0000002700000000",
            INIT_0F => X"fffffff2ffffffff0000000800000000ffffffe8ffffffff0000004b00000000",
            INIT_10 => X"ffffffe6ffffffff000000030000000000000002000000000000001400000000",
            INIT_11 => X"0000001b000000000000001b00000000fffffff7ffffffffffffffc4ffffffff",
            INIT_12 => X"ffffffb3ffffffffffffffcfffffffffffffffd7ffffffffffffffe1ffffffff",
            INIT_13 => X"0000000300000000ffffffedffffffff00000006000000000000002500000000",
            INIT_14 => X"0000003100000000fffffffaffffffffffffffecffffffffffffffd4ffffffff",
            INIT_15 => X"fffffff8ffffffff0000001000000000ffffffe2fffffffffffffff1ffffffff",
            INIT_16 => X"fffffff9ffffffffffffffe3ffffffff00000014000000000000001900000000",
            INIT_17 => X"0000000800000000ffffffadffffffffffffffb8ffffffffffffffc7ffffffff",
            INIT_18 => X"fffffffeffffffff0000001a00000000ffffff9fffffffff0000001100000000",
            INIT_19 => X"0000002a00000000ffffffe7fffffffffffffff6ffffffffffffffedffffffff",
            INIT_1A => X"0000000e00000000fffffff8fffffffffffffffbfffffffffffffffaffffffff",
            INIT_1B => X"0000001700000000000000080000000000000012000000000000002600000000",
            INIT_1C => X"0000001000000000ffffffccffffffff00000021000000000000001800000000",
            INIT_1D => X"fffffff5ffffffffffffffd7ffffffffffffffe9fffffffffffffff2ffffffff",
            INIT_1E => X"000000220000000000000054000000000000000b00000000ffffffe8ffffffff",
            INIT_1F => X"ffffffd8ffffffff0000002900000000fffffff3ffffffffffffffd7ffffffff",
            INIT_20 => X"fffffffdffffffff0000001000000000fffffff1ffffffff0000002800000000",
            INIT_21 => X"0000001e00000000000000290000000000000007000000000000003f00000000",
            INIT_22 => X"0000000c00000000ffffffd5ffffffff0000001500000000ffffffcbffffffff",
            INIT_23 => X"0000006200000000ffffffe0ffffffff0000000b000000000000000200000000",
            INIT_24 => X"ffffffeaffffffffffffffccffffffff00000011000000000000000200000000",
            INIT_25 => X"ffffffd3ffffffffffffffa5ffffffff00000034000000000000002700000000",
            INIT_26 => X"0000004b0000000000000072000000000000003200000000ffffffa8ffffffff",
            INIT_27 => X"fffffff2ffffffffffffffffffffffffffffffe1ffffffffffffffe9ffffffff",
            INIT_28 => X"0000003500000000ffffffe6ffffffffffffffb7ffffffffffffffebffffffff",
            INIT_29 => X"00000000000000000000000c000000000000000400000000ffffffafffffffff",
            INIT_2A => X"0000003400000000ffffffdcffffffffffffffeeffffffff0000000600000000",
            INIT_2B => X"0000000900000000ffffffbfffffffff00000033000000000000004c00000000",
            INIT_2C => X"fffffff4ffffffff00000006000000000000000300000000ffffffe2ffffffff",
            INIT_2D => X"ffffffeaffffffffffffff7fffffffffffffffd6ffffffffffffffd6ffffffff",
            INIT_2E => X"fffffffffffffffffffffff1ffffffff00000017000000000000001500000000",
            INIT_2F => X"ffffffd0ffffffff0000001a00000000ffffffedffffffffffffffdeffffffff",
            INIT_30 => X"0000002500000000fffffffdffffffff0000001a00000000ffffffe3ffffffff",
            INIT_31 => X"ffffffb9ffffffff0000003f000000000000003b00000000ffffffe5ffffffff",
            INIT_32 => X"ffffffc2ffffffff00000000000000000000000100000000fffffff4ffffffff",
            INIT_33 => X"ffffffd4fffffffffffffff4ffffffffffffffe7ffffffff0000000f00000000",
            INIT_34 => X"0000002c00000000ffffffc8ffffffffffffffe8fffffffffffffff4ffffffff",
            INIT_35 => X"ffffffd7ffffffff000000000000000000000007000000000000000800000000",
            INIT_36 => X"ffffffe5ffffffff0000001a00000000fffffff2fffffffffffffff2ffffffff",
            INIT_37 => X"ffffffcdffffffffffffffe0ffffffffffffffddfffffffffffffff3ffffffff",
            INIT_38 => X"0000001600000000fffffff4ffffffffffffffbfffffffff0000002000000000",
            INIT_39 => X"fffffffafffffffffffffff4ffffffff0000001900000000ffffffcaffffffff",
            INIT_3A => X"0000001000000000ffffffe7ffffffff00000047000000000000000000000000",
            INIT_3B => X"00000001000000000000000800000000fffffffaffffffff0000001f00000000",
            INIT_3C => X"0000000a00000000fffffff5ffffffff00000018000000000000001b00000000",
            INIT_3D => X"ffffffeeffffffffffffffe3fffffffffffffff7ffffffffffffffe5ffffffff",
            INIT_3E => X"ffffffcfffffffffffffffd8ffffffffffffffecffffffff0000001b00000000",
            INIT_3F => X"ffffffbafffffffffffffff7ffffffff00000009000000000000005500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffc6ffffffff000000340000000000000012000000000000001a00000000",
            INIT_41 => X"0000001300000000000000140000000000000010000000000000000500000000",
            INIT_42 => X"ffffffccfffffffffffffffcffffffff00000000000000000000001900000000",
            INIT_43 => X"0000000100000000ffffffcfffffffff0000000b00000000ffffffe3ffffffff",
            INIT_44 => X"0000000600000000ffffffffffffffff0000001200000000ffffffceffffffff",
            INIT_45 => X"ffffffc4ffffffff00000003000000000000000b00000000ffffffe3ffffffff",
            INIT_46 => X"0000001f00000000ffffffc3ffffffff0000000700000000ffffffdcffffffff",
            INIT_47 => X"ffffffe6ffffffffffffffe2ffffffffffffffc8ffffffffffffffd0ffffffff",
            INIT_48 => X"0000001300000000fffffff3ffffffffffffff84ffffffff0000000400000000",
            INIT_49 => X"0000000400000000ffffffe8fffffffffffffff1ffffffffffffffd2ffffffff",
            INIT_4A => X"0000000900000000ffffffcfffffffffffffffa4ffffffffffffffedffffffff",
            INIT_4B => X"fffffff5ffffffff0000000a000000000000002e000000000000004100000000",
            INIT_4C => X"fffffffffffffffffffffff5ffffffff0000001e00000000fffffffbffffffff",
            INIT_4D => X"0000001700000000fffffff8ffffffff0000000100000000ffffffcaffffffff",
            INIT_4E => X"ffffffe6ffffffff0000003000000000fffffff8ffffffff0000000300000000",
            INIT_4F => X"0000000b000000000000002b000000000000001200000000ffffffe6ffffffff",
            INIT_50 => X"ffffffe0ffffffff0000002900000000ffffffffffffffff0000001400000000",
            INIT_51 => X"0000001300000000ffffffe8fffffffffffffff1fffffffffffffff8ffffffff",
            INIT_52 => X"00000000000000000000000100000000ffffffdbffffffff0000001300000000",
            INIT_53 => X"0000000000000000ffffffdeffffffffffffffebffffffff0000000300000000",
            INIT_54 => X"0000001c00000000ffffffa6ffffffffffffffeaffffffffffffffbfffffffff",
            INIT_55 => X"ffffffe2ffffffff0000000b00000000ffffffd6ffffffff0000002800000000",
            INIT_56 => X"ffffffd3ffffffffffffffebffffffff00000020000000000000001600000000",
            INIT_57 => X"ffffffe3ffffffffffffffcbffffffffffffffd0ffffffff0000000300000000",
            INIT_58 => X"0000000300000000fffffff0ffffffffffffffb0ffffffff0000003600000000",
            INIT_59 => X"ffffffe3ffffffffffffffffffffffff0000000e00000000ffffffdcffffffff",
            INIT_5A => X"ffffffceffffffffffffffdeffffffffffffffd8ffffffff0000000e00000000",
            INIT_5B => X"0000001700000000fffffff9fffffffffffffffbfffffffffffffff8ffffffff",
            INIT_5C => X"000000340000000000000021000000000000001200000000ffffffd5ffffffff",
            INIT_5D => X"fffffffbffffffff0000000c00000000fffffff6ffffffffffffffdbffffffff",
            INIT_5E => X"00000022000000000000001400000000ffffffddffffffffffffffdaffffffff",
            INIT_5F => X"ffffffd4ffffffff0000001500000000ffffffebffffffff0000000400000000",
            INIT_60 => X"ffffffdcffffffff0000001b00000000ffffffeeffffffff0000002200000000",
            INIT_61 => X"0000001900000000fffffff2ffffffff0000000f000000000000000800000000",
            INIT_62 => X"0000000d000000000000001800000000ffffffceffffffff0000000100000000",
            INIT_63 => X"ffffffdffffffffffffffff0ffffffffffffffe6ffffffffffffffe7ffffffff",
            INIT_64 => X"0000001f00000000ffffffc4ffffffff0000001600000000ffffffd5ffffffff",
            INIT_65 => X"ffffffbeffffffff0000002800000000ffffffd9ffffffff0000000900000000",
            INIT_66 => X"0000001100000000ffffffd4ffffffffffffffd3ffffffffffffffe9ffffffff",
            INIT_67 => X"fffffff5ffffffffffffffe0ffffffffffffffd7fffffffffffffffdffffffff",
            INIT_68 => X"0000001b00000000ffffffeaffffffffffffffa8ffffffffffffffffffffffff",
            INIT_69 => X"fffffff7fffffffffffffff1ffffffffffffffedffffffffffffffebffffffff",
            INIT_6A => X"00000003000000000000000d00000000ffffffeeffffffff0000000800000000",
            INIT_6B => X"00000026000000000000001e0000000000000005000000000000001300000000",
            INIT_6C => X"00000032000000000000000a000000000000001200000000ffffffccffffffff",
            INIT_6D => X"00000008000000000000000600000000fffffff7ffffffffffffffe9ffffffff",
            INIT_6E => X"0000001000000000ffffffc9ffffffffffffffdaffffffff0000000e00000000",
            INIT_6F => X"ffffffedffffffffffffffeeffffffffffffffe8ffffffff0000001200000000",
            INIT_70 => X"ffffffceffffffff0000003800000000ffffffdefffffffffffffff3ffffffff",
            INIT_71 => X"ffffffe9ffffffff0000001a0000000000000004000000000000001600000000",
            INIT_72 => X"fffffffefffffffffffffffbffffffffffffffcafffffffffffffffcffffffff",
            INIT_73 => X"fffffffdffffffff000000030000000000000010000000000000000c00000000",
            INIT_74 => X"fffffffeffffffff0000000000000000fffffff9ffffffffffffffe5ffffffff",
            INIT_75 => X"0000003a000000000000001e000000000000000e00000000ffffffc2ffffffff",
            INIT_76 => X"ffffffa9fffffffffffffffdffffffff0000000c000000000000000600000000",
            INIT_77 => X"ffffffeeffffffff000000250000000000000010000000000000002500000000",
            INIT_78 => X"fffffffdfffffffffffffffeffffffff00000026000000000000000600000000",
            INIT_79 => X"0000000900000000fffffffdffffffff00000011000000000000002100000000",
            INIT_7A => X"ffffffedffffffff0000000200000000ffffffc1ffffffff0000000900000000",
            INIT_7B => X"0000001100000000ffffffc3ffffffffffffffc7ffffffff0000000f00000000",
            INIT_7C => X"fffffff9ffffffffffffffebffffffff0000003300000000ffffffc0ffffffff",
            INIT_7D => X"0000000b000000000000000500000000fffffff9ffffffff0000000d00000000",
            INIT_7E => X"0000000f000000000000005700000000ffffffb4ffffffff0000001900000000",
            INIT_7F => X"0000000800000000fffffff2ffffffffffffffe8ffffffff0000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE7;


    MEM_IWGHT_LAYER3_INSTANCE8 : if BRAM_NAME = "iwght_layer3_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002c00000000fffffffaffffffff0000001500000000ffffffeaffffffff",
            INIT_01 => X"ffffffe3ffffffffffffffebfffffffffffffff9ffffffff0000000000000000",
            INIT_02 => X"ffffffeeffffffff0000001e00000000fffffff6fffffffffffffffbffffffff",
            INIT_03 => X"fffffffbfffffffffffffff6ffffffff00000010000000000000002c00000000",
            INIT_04 => X"0000001300000000ffffffb9ffffffff0000000000000000ffffffd9ffffffff",
            INIT_05 => X"fffffff4ffffffff0000003f000000000000000000000000ffffffd4ffffffff",
            INIT_06 => X"ffffffcbfffffffffffffff1ffffffff0000002700000000fffffff2ffffffff",
            INIT_07 => X"ffffffdcffffffff0000002300000000fffffffafffffffffffffffbffffffff",
            INIT_08 => X"ffffffffffffffffffffffe9fffffffffffffff9ffffffff0000000200000000",
            INIT_09 => X"ffffffdeffffffff0000000f0000000000000017000000000000000500000000",
            INIT_0A => X"fffffffeffffffffffffffd5ffffffffffffffd1ffffffff0000000800000000",
            INIT_0B => X"0000000200000000fffffffcffffffffffffffe0fffffffffffffff7ffffffff",
            INIT_0C => X"0000002200000000fffffffbffffffffffffffe0ffffffffffffffe8ffffffff",
            INIT_0D => X"ffffffe9ffffffff0000002500000000ffffffe9ffffffff0000003500000000",
            INIT_0E => X"fffffff9ffffffffffffffc8fffffffffffffffeffffffffffffff81ffffffff",
            INIT_0F => X"ffffffd6ffffffff0000002200000000fffffff8ffffffffffffffbaffffffff",
            INIT_10 => X"ffffffe5ffffffffffffffe7ffffffff0000001f000000000000002200000000",
            INIT_11 => X"0000003c00000000ffffffcdffffffffffffffd2ffffffffffffffe5ffffffff",
            INIT_12 => X"0000000000000000ffffffddffffffffffffffe4fffffffffffffff4ffffffff",
            INIT_13 => X"00000015000000000000000800000000ffffffe6ffffffff0000000100000000",
            INIT_14 => X"fffffff3ffffffff0000002300000000fffffffcffffffff0000001500000000",
            INIT_15 => X"0000001100000000fffffff8ffffffffffffffd1ffffffffffffffc8ffffffff",
            INIT_16 => X"ffffffd3ffffffff00000008000000000000003c000000000000001300000000",
            INIT_17 => X"ffffffd4ffffffff0000002900000000fffffff0ffffffff0000004600000000",
            INIT_18 => X"fffffffdffffffff0000000c000000000000003000000000fffffff4ffffffff",
            INIT_19 => X"fffffffcffffffff000000020000000000000000000000000000001b00000000",
            INIT_1A => X"ffffffffffffffff00000023000000000000000b00000000ffffffd5ffffffff",
            INIT_1B => X"ffffffdafffffffffffffff2ffffffffffffffe8ffffffffffffffc8ffffffff",
            INIT_1C => X"fffffff4ffffffffffffffe7ffffffff00000004000000000000001500000000",
            INIT_1D => X"ffffffe9ffffffff00000004000000000000000600000000ffffffecffffffff",
            INIT_1E => X"0000000500000000ffffffd2ffffffffffffffe4ffffffffffffffc5ffffffff",
            INIT_1F => X"0000000d00000000ffffffe9ffffffff0000000700000000ffffffc8ffffffff",
            INIT_20 => X"0000001d000000000000001c00000000fffffffbffffffff0000003e00000000",
            INIT_21 => X"00000034000000000000000800000000ffffffe4ffffffff0000003c00000000",
            INIT_22 => X"0000001a00000000fffffff7ffffffffffffffdeffffffffffffffebffffffff",
            INIT_23 => X"ffffffcfffffffffffffffbcffffffff0000001a00000000fffffff7ffffffff",
            INIT_24 => X"00000031000000000000000d00000000fffffff5ffffffff0000001f00000000",
            INIT_25 => X"0000001a00000000fffffffbffffffff00000018000000000000003800000000",
            INIT_26 => X"0000001300000000fffffff0ffffffffffffffe5ffffffff0000003000000000",
            INIT_27 => X"0000000b000000000000000c00000000ffffffe5ffffffff0000000700000000",
            INIT_28 => X"00000016000000000000000e000000000000005200000000ffffffd4ffffffff",
            INIT_29 => X"ffffffccffffffff00000007000000000000000f000000000000001a00000000",
            INIT_2A => X"fffffffcfffffffffffffffaffffffff0000000f00000000ffffffebffffffff",
            INIT_2B => X"0000003a00000000fffffff4ffffffffffffffeeffffffffffffffdaffffffff",
            INIT_2C => X"00000013000000000000001100000000fffffff0ffffffff0000000d00000000",
            INIT_2D => X"00000010000000000000003300000000ffffffd7ffffffffffffffe9ffffffff",
            INIT_2E => X"00000016000000000000002800000000fffffffeffffffff0000004600000000",
            INIT_2F => X"ffffffbeffffffff0000001f00000000fffffffcffffffff0000000400000000",
            INIT_30 => X"fffffff1ffffffff00000001000000000000001c000000000000000f00000000",
            INIT_31 => X"fffffff9ffffffff0000000a0000000000000019000000000000000300000000",
            INIT_32 => X"00000024000000000000002e00000000ffffffa2fffffffffffffff7ffffffff",
            INIT_33 => X"ffffffafffffffffffffffeaffffffff00000006000000000000000400000000",
            INIT_34 => X"ffffffd2ffffffffffffffb7ffffffff0000000c00000000fffffff5ffffffff",
            INIT_35 => X"0000001200000000ffffffdeffffffffffffffa8ffffffffffffffdfffffffff",
            INIT_36 => X"ffffffabffffffffffffff9dfffffffffffffff0ffffffff0000002800000000",
            INIT_37 => X"ffffffeeffffffff0000000800000000fffffffcffffffffffffffcaffffffff",
            INIT_38 => X"fffffffaffffffff0000000e00000000fffffffbffffffff0000001300000000",
            INIT_39 => X"ffffffeeffffffffffffffefffffffffffffffe6ffffffff0000000400000000",
            INIT_3A => X"ffffffb6ffffffffffffffc2ffffffffffffffc4ffffffffffffffdcffffffff",
            INIT_3B => X"ffffffc0ffffffff0000003100000000fffffff6ffffffffffffff81ffffffff",
            INIT_3C => X"ffffffc5ffffffff0000002c00000000ffffffe4ffffffff0000001a00000000",
            INIT_3D => X"ffffffe7ffffffff0000003900000000ffffffecffffffff0000000e00000000",
            INIT_3E => X"ffffffecffffffffffffffdefffffffffffffffaffffffff0000002d00000000",
            INIT_3F => X"00000012000000000000000c00000000ffffffefffffffff0000001e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"fffffff3ffffffffffffffdfffffffffffffffa5ffffffff0000003b00000000",
            INIT_41 => X"ffffffe9ffffffffffffffc1ffffffffffffffe1ffffffff0000000600000000",
            INIT_42 => X"fffffff5ffffffff0000000e00000000ffffffbaffffffff0000001500000000",
            INIT_43 => X"ffffffdcffffffffffffffd0ffffffffffffffeaffffffff0000001100000000",
            INIT_44 => X"ffffffeeffffffffffffffd7fffffffffffffff2ffffffff0000003500000000",
            INIT_45 => X"000000000000000000000014000000000000000000000000ffffffd4ffffffff",
            INIT_46 => X"0000002400000000ffffffe2ffffffffffffffd5fffffffffffffff4ffffffff",
            INIT_47 => X"ffffff84fffffffffffffff8fffffffffffffff8ffffffff0000002500000000",
            INIT_48 => X"fffffff7ffffffff00000001000000000000001e00000000fffffff4ffffffff",
            INIT_49 => X"fffffff3ffffffff0000000c000000000000000e000000000000000e00000000",
            INIT_4A => X"ffffffe5ffffffffffffffddffffffffffffff89fffffffffffffff1ffffffff",
            INIT_4B => X"fffffff2ffffffff0000000900000000fffffff3ffffffffffffffdaffffffff",
            INIT_4C => X"ffffffc7ffffffff0000001100000000ffffffffffffffff0000000700000000",
            INIT_4D => X"fffffff2ffffffff000000270000000000000000000000000000001800000000",
            INIT_4E => X"ffffffe4fffffffffffffff8ffffffff00000022000000000000001400000000",
            INIT_4F => X"ffffffedfffffffffffffff8ffffffff0000001500000000ffffffe2ffffffff",
            INIT_50 => X"0000000300000000fffffffeffffffffffffffc9ffffffff0000001700000000",
            INIT_51 => X"fffffffdffffffff00000000000000000000000300000000ffffffe6ffffffff",
            INIT_52 => X"00000027000000000000001b00000000ffffffd7ffffffffffffffd9ffffffff",
            INIT_53 => X"00000001000000000000000200000000ffffffebffffffffffffffaeffffffff",
            INIT_54 => X"0000003f00000000ffffffb5ffffffff00000000000000000000003400000000",
            INIT_55 => X"fffffff5ffffffff0000000b0000000000000004000000000000002200000000",
            INIT_56 => X"fffffff1ffffffffffffffcafffffffffffffff7ffffffff0000003700000000",
            INIT_57 => X"0000000500000000fffffff1ffffffff00000000000000000000000600000000",
            INIT_58 => X"000000300000000000000001000000000000002700000000ffffffd6ffffffff",
            INIT_59 => X"0000001500000000fffffff6fffffffffffffffaffffffff0000001e00000000",
            INIT_5A => X"000000020000000000000001000000000000002100000000fffffff0ffffffff",
            INIT_5B => X"000000090000000000000007000000000000002200000000ffffffb4ffffffff",
            INIT_5C => X"0000001700000000ffffffe9ffffffffffffffd2ffffffff0000000e00000000",
            INIT_5D => X"0000001400000000fffffff9ffffffffffffffbdffffffff0000001200000000",
            INIT_5E => X"fffffff4ffffffffffffffd4ffffffff0000002f000000000000001000000000",
            INIT_5F => X"0000002100000000ffffffd8ffffffffffffffedffffffffffffffb3ffffffff",
            INIT_60 => X"00000019000000000000000300000000ffffff81ffffffff0000000800000000",
            INIT_61 => X"ffffffa8ffffffff00000041000000000000000700000000ffffffefffffffff",
            INIT_62 => X"ffffffd0ffffffff00000026000000000000001900000000ffffffefffffffff",
            INIT_63 => X"0000000800000000ffffffd3ffffffff0000000000000000ffffffd6ffffffff",
            INIT_64 => X"000000160000000000000010000000000000000c000000000000003a00000000",
            INIT_65 => X"0000000f00000000fffffff2ffffffff0000002c000000000000001600000000",
            INIT_66 => X"0000002400000000fffffff3ffffffff0000003200000000ffffffb9ffffffff",
            INIT_67 => X"ffffffe2ffffffff0000000e0000000000000027000000000000001c00000000",
            INIT_68 => X"00000025000000000000001700000000fffffff9fffffffffffffff7ffffffff",
            INIT_69 => X"0000001700000000fffffff6fffffffffffffff1ffffffff0000000700000000",
            INIT_6A => X"ffffffeaffffffff0000000600000000ffffffe2ffffffff0000000800000000",
            INIT_6B => X"0000001400000000fffffff4ffffffff0000000000000000ffffffe6ffffffff",
            INIT_6C => X"ffffffecffffffffffffffccffffffff0000000a000000000000002c00000000",
            INIT_6D => X"00000017000000000000000500000000ffffff99ffffffff0000000b00000000",
            INIT_6E => X"ffffffe8fffffffffffffff0ffffffff00000031000000000000003200000000",
            INIT_6F => X"ffffffd8fffffffffffffffcffffffff0000000600000000ffffffefffffffff",
            INIT_70 => X"0000004c00000000fffffff0ffffffff00000003000000000000000600000000",
            INIT_71 => X"ffffffc5ffffffff00000038000000000000003900000000ffffffc2ffffffff",
            INIT_72 => X"fffffffeffffffff0000003300000000ffffffe7ffffffffffffffc5ffffffff",
            INIT_73 => X"fffffff5ffffffff0000000c00000000ffffffe8ffffffff0000000300000000",
            INIT_74 => X"ffffffd5ffffffff000000020000000000000008000000000000001e00000000",
            INIT_75 => X"0000003f00000000ffffffe8ffffffff0000000f000000000000001d00000000",
            INIT_76 => X"0000001700000000ffffffa6ffffffff0000000c00000000fffffff5ffffffff",
            INIT_77 => X"ffffffbaffffffff0000001a000000000000000500000000fffffff5ffffffff",
            INIT_78 => X"ffffffffffffffffffffffeeffffffff0000001d000000000000000d00000000",
            INIT_79 => X"0000001000000000fffffff0ffffffffffffffedffffffff0000000100000000",
            INIT_7A => X"0000000500000000ffffffafffffffffffffffa8ffffffffffffffe1ffffffff",
            INIT_7B => X"000000080000000000000002000000000000000700000000ffffffe7ffffffff",
            INIT_7C => X"ffffffaeffffffff0000001100000000fffffff4ffffffffffffffd2ffffffff",
            INIT_7D => X"fffffff5ffffffff0000000400000000ffffffc2ffffffffffffffe4ffffffff",
            INIT_7E => X"ffffffabffffffff000000370000000000000039000000000000004100000000",
            INIT_7F => X"0000001b000000000000001e000000000000000d00000000fffffff9ffffffff",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE8;


    MEM_IWGHT_LAYER3_INSTANCE9 : if BRAM_NAME = "iwght_layer3_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000ffffffe3ffffffffffffffefffffffff0000001100000000",
            INIT_01 => X"00000002000000000000001e000000000000001900000000ffffffa6ffffffff",
            INIT_02 => X"0000001300000000ffffffdcffffffffffffffd4ffffffffffffffc7ffffffff",
            INIT_03 => X"fffffffeffffffffffffffe1ffffffff0000000200000000ffffffd3ffffffff",
            INIT_04 => X"ffffffe0fffffffffffffff7fffffffffffffff1ffffffff0000002c00000000",
            INIT_05 => X"0000000c00000000ffffffbffffffffffffffffaffffffff0000000500000000",
            INIT_06 => X"ffffffe1ffffffffffffffe4ffffffff0000000c000000000000000000000000",
            INIT_07 => X"000000010000000000000017000000000000002c000000000000001f00000000",
            INIT_08 => X"ffffffcdffffffffffffffedfffffffffffffff8ffffffffffffffd5ffffffff",
            INIT_09 => X"ffffffe7fffffffffffffffeffffffff00000000000000000000002500000000",
            INIT_0A => X"0000002100000000ffffffeaffffffff00000011000000000000000d00000000",
            INIT_0B => X"ffffffebffffffffffffffedffffffff00000004000000000000000000000000",
            INIT_0C => X"00000012000000000000000000000000fffffff2ffffffffffffffbaffffffff",
            INIT_0D => X"fffffffbfffffffffffffffbffffffff0000000e000000000000000a00000000",
            INIT_0E => X"fffffff1ffffffffffffffceffffffffffffffcbffffffff0000000300000000",
            INIT_0F => X"0000002400000000ffffffe6ffffffff00000003000000000000001500000000",
            INIT_10 => X"ffffffe6fffffffffffffff3ffffffffffffffecfffffffffffffff4ffffffff",
            INIT_11 => X"fffffff4ffffffff0000000000000000ffffffcdffffffffffffffbaffffffff",
            INIT_12 => X"ffffffdeffffffff000000000000000000000009000000000000002900000000",
            INIT_13 => X"fffffff2ffffffffffffffe7ffffffff0000000500000000ffffffd4ffffffff",
            INIT_14 => X"ffffffefffffffff0000001400000000fffffffcffffffff0000002500000000",
            INIT_15 => X"fffffffbfffffffffffffff5ffffffff00000002000000000000001300000000",
            INIT_16 => X"0000000300000000ffffffd9ffffffff00000010000000000000000000000000",
            INIT_17 => X"ffffffd8ffffffff00000004000000000000000500000000ffffffffffffffff",
            INIT_18 => X"fffffffefffffffffffffffefffffffffffffff6ffffffff0000002200000000",
            INIT_19 => X"0000001a000000000000000900000000fffffff7fffffffffffffffbffffffff",
            INIT_1A => X"0000001d00000000ffffffd1fffffffffffffffbffffffff0000000f00000000",
            INIT_1B => X"0000000700000000ffffffedffffffff0000001600000000ffffffd4ffffffff",
            INIT_1C => X"0000000c00000000fffffff5ffffffff0000000e00000000ffffffdfffffffff",
            INIT_1D => X"0000001400000000ffffffdaffffffff00000005000000000000000700000000",
            INIT_1E => X"ffffffd6ffffffff000000130000000000000025000000000000001300000000",
            INIT_1F => X"0000001600000000fffffff0fffffffffffffffeffffffffffffffe6ffffffff",
            INIT_20 => X"fffffff9ffffffffffffffedfffffffffffffffdffffffffffffffe5ffffffff",
            INIT_21 => X"ffffffcdfffffffffffffffdffffffffffffffd2ffffffffffffffb9ffffffff",
            INIT_22 => X"fffffff3ffffffff00000011000000000000001300000000fffffffeffffffff",
            INIT_23 => X"0000001d00000000ffffffecfffffffffffffff8ffffffffffffffc5ffffffff",
            INIT_24 => X"ffffffe0ffffffffffffffdcffffffff00000009000000000000001100000000",
            INIT_25 => X"0000001c00000000ffffffbeffffffff0000002400000000ffffffcfffffffff",
            INIT_26 => X"ffffffe4ffffffffffffffffffffffff0000000b000000000000001500000000",
            INIT_27 => X"ffffffe4ffffffffffffffeaffffffff0000000b000000000000001600000000",
            INIT_28 => X"fffffff6fffffffffffffff4ffffffffffffffdeffffffffffffffedffffffff",
            INIT_29 => X"0000003500000000fffffff9ffffffff00000011000000000000001300000000",
            INIT_2A => X"000000060000000000000003000000000000002500000000ffffffe4ffffffff",
            INIT_2B => X"ffffffeeffffffffffffffe6fffffffffffffff9fffffffffffffff6ffffffff",
            INIT_2C => X"00000004000000000000002600000000ffffffddffffffff0000000700000000",
            INIT_2D => X"0000001400000000ffffffe2ffffffff0000000c00000000ffffffd5ffffffff",
            INIT_2E => X"ffffffd4ffffffffffffffefffffffff00000005000000000000003300000000",
            INIT_2F => X"0000003600000000ffffffeeffffffff00000009000000000000001800000000",
            INIT_30 => X"00000021000000000000000000000000ffffffe3ffffffffffffffdbffffffff",
            INIT_31 => X"ffffffe0fffffffffffffff7ffffffffffffffe6ffffffffffffffe2ffffffff",
            INIT_32 => X"00000018000000000000001b0000000000000024000000000000000c00000000",
            INIT_33 => X"00000000000000000000001700000000fffffff5ffffffffffffffc3ffffffff",
            INIT_34 => X"ffffffdaffffffff0000000a0000000000000003000000000000000900000000",
            INIT_35 => X"0000000a00000000ffffffb9ffffffffffffffd6ffffffff0000002b00000000",
            INIT_36 => X"ffffffe3ffffffff0000004b00000000fffffffbffffffff0000000600000000",
            INIT_37 => X"0000001f000000000000002b00000000ffffffe9ffffffff0000000700000000",
            INIT_38 => X"fffffff7fffffffffffffffeffffffff0000000400000000fffffffbffffffff",
            INIT_39 => X"fffffff0ffffffffffffffe6fffffffffffffffeffffffff0000000000000000",
            INIT_3A => X"0000000200000000000000170000000000000014000000000000000700000000",
            INIT_3B => X"0000000b00000000ffffffbffffffffffffffff0fffffffffffffff5ffffffff",
            INIT_3C => X"0000001100000000ffffffd9fffffffffffffff9ffffffffffffffc6ffffffff",
            INIT_3D => X"0000001300000000ffffffe4ffffffff0000000f00000000fffffff4ffffffff",
            INIT_3E => X"ffffffefffffffff0000000000000000ffffffeeffffffffffffffefffffffff",
            INIT_3F => X"0000000f0000000000000027000000000000000300000000fffffff9ffffffff",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000a000000000000000500000000ffffffc8ffffffff",
            INIT_41 => X"ffffffadffffffffffffffecffffffffffffff9fffffffffffffffe5ffffffff",
            INIT_42 => X"ffffffedffffffff000000350000000000000010000000000000000c00000000",
            INIT_43 => X"ffffffe6ffffffff00000001000000000000000400000000ffffffd2ffffffff",
            INIT_44 => X"000000170000000000000009000000000000000c000000000000002500000000",
            INIT_45 => X"0000001100000000ffffffe0ffffffff0000000d000000000000002200000000",
            INIT_46 => X"ffffffe8ffffffff00000027000000000000001e00000000ffffffd8ffffffff",
            INIT_47 => X"0000004000000000fffffff8ffffffff0000002900000000fffffff9ffffffff",
            INIT_48 => X"00000000000000000000000a00000000ffffffd3ffffffffffffffefffffffff",
            INIT_49 => X"00000005000000000000000500000000fffffff9ffffffffffffffeeffffffff",
            INIT_4A => X"0000001300000000ffffffc8ffffffff00000064000000000000000b00000000",
            INIT_4B => X"0000003000000000ffffffacfffffffffffffffaffffffffffffffaeffffffff",
            INIT_4C => X"0000000a00000000ffffffc9ffffffffffffffe1fffffffffffffffaffffffff",
            INIT_4D => X"fffffff0ffffffff00000008000000000000001c000000000000003400000000",
            INIT_4E => X"ffffffcefffffffffffffffbffffffff0000000f000000000000000d00000000",
            INIT_4F => X"0000002c0000000000000005000000000000000200000000ffffffeeffffffff",
            INIT_50 => X"000000250000000000000005000000000000000f00000000fffffff8ffffffff",
            INIT_51 => X"ffffffdaffffffff0000000600000000ffffffcbfffffffffffffff7ffffffff",
            INIT_52 => X"fffffff9ffffffffffffffedffffffff0000003400000000fffffff1ffffffff",
            INIT_53 => X"0000001d00000000ffffffbbffffffffffffffe9ffffffff0000000800000000",
            INIT_54 => X"0000000e000000000000000100000000fffffffeffffffff0000004900000000",
            INIT_55 => X"0000000100000000ffffffadffffffff0000004c00000000ffffffbbffffffff",
            INIT_56 => X"ffffffceffffffff000000330000000000000034000000000000000000000000",
            INIT_57 => X"000000170000000000000000000000000000002000000000ffffffc9ffffffff",
            INIT_58 => X"ffffffc6ffffffff00000012000000000000001d000000000000001700000000",
            INIT_59 => X"0000000600000000000000130000000000000009000000000000000c00000000",
            INIT_5A => X"0000001400000000ffffffebffffffff0000004200000000ffffffe0ffffffff",
            INIT_5B => X"ffffffffffffffffffffffcaffffffff0000000700000000ffffffe6ffffffff",
            INIT_5C => X"ffffffcbffffffff0000001c000000000000000b00000000ffffffe0ffffffff",
            INIT_5D => X"000000030000000000000008000000000000000d00000000fffffffeffffffff",
            INIT_5E => X"0000000000000000ffffffe7ffffffffffffffe4ffffffff0000001f00000000",
            INIT_5F => X"0000001d00000000ffffffeaffffffff0000000e00000000ffffffe4ffffffff",
            INIT_60 => X"fffffffaffffffffffffffdaffffffff00000001000000000000000900000000",
            INIT_61 => X"ffffffe7fffffffffffffff0ffffffffffffffb3ffffffffffffffd4ffffffff",
            INIT_62 => X"fffffff9fffffffffffffffdffffffff0000002700000000ffffffe0ffffffff",
            INIT_63 => X"0000001b000000000000000000000000fffffff8ffffffff0000002200000000",
            INIT_64 => X"ffffffe8ffffffff0000002d00000000fffffff2ffffffffffffffedffffffff",
            INIT_65 => X"fffffff7ffffffffffffffebfffffffffffffff8ffffffffffffffefffffffff",
            INIT_66 => X"ffffffc2ffffffff0000004600000000fffffff6ffffffffffffffbbffffffff",
            INIT_67 => X"00000022000000000000000f00000000ffffffe7ffffffffffffffdfffffffff",
            INIT_68 => X"ffffffc8ffffffff0000000100000000fffffff9ffffffff0000002100000000",
            INIT_69 => X"fffffff4ffffffff0000000b000000000000001500000000fffffff2ffffffff",
            INIT_6A => X"fffffffdffffffff0000004200000000fffffff2fffffffffffffffeffffffff",
            INIT_6B => X"0000000000000000ffffffe3ffffffffffffffd6ffffffffffffffc9ffffffff",
            INIT_6C => X"fffffff0ffffffffffffffd4ffffffff0000002e00000000ffffffd9ffffffff",
            INIT_6D => X"fffffffbffffffffffffffceffffffffffffffe9ffffffff0000001200000000",
            INIT_6E => X"0000000700000000ffffffe7ffffffff0000002700000000ffffffb5ffffffff",
            INIT_6F => X"ffffffccffffffff00000004000000000000000c000000000000000900000000",
            INIT_70 => X"000000370000000000000037000000000000007a00000000ffffffc1ffffffff",
            INIT_71 => X"0000000d00000000ffffffa6ffffffffffffff98ffffffff0000002600000000",
            INIT_72 => X"fffffff3ffffffffffffffb1ffffffffffffffebffffffff0000001900000000",
            INIT_73 => X"00000031000000000000000c00000000ffffffffffffffff0000000f00000000",
            INIT_74 => X"ffffffd5ffffffff00000044000000000000000700000000fffffff8ffffffff",
            INIT_75 => X"ffffffdaffffffffffffffe2ffffffffffffffe9ffffffffffffffdfffffffff",
            INIT_76 => X"000000050000000000000053000000000000000e00000000ffffff9fffffffff",
            INIT_77 => X"0000003f00000000ffffffefffffffff0000004200000000ffffffe7ffffffff",
            INIT_78 => X"ffffffbffffffffffffffff7ffffffff0000000700000000ffffffffffffffff",
            INIT_79 => X"0000000000000000fffffffefffffffffffffff4ffffffffffffffd2ffffffff",
            INIT_7A => X"ffffffecffffffff0000001b0000000000000036000000000000001200000000",
            INIT_7B => X"ffffffb1ffffffffffffffe8ffffffffffffffedffffffff0000001f00000000",
            INIT_7C => X"0000000b00000000ffffffeaffffffff0000000000000000ffffffcfffffffff",
            INIT_7D => X"0000000200000000ffffffb7ffffffffffffffc2fffffffffffffff5ffffffff",
            INIT_7E => X"fffffff9ffffffff0000001100000000ffffffd8ffffffff0000000000000000",
            INIT_7F => X"0000000c00000000ffffffeeffffffffffffffe4ffffffff0000005500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE9;


    MEM_IWGHT_LAYER3_INSTANCE10 : if BRAM_NAME = "iwght_layer3_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000090000000000000000000000000000003500000000ffffffbcffffffff",
            INIT_01 => X"ffffffe9ffffffff000000050000000000000010000000000000003700000000",
            INIT_02 => X"fffffff6ffffffffffffffc5ffffffff00000026000000000000005000000000",
            INIT_03 => X"ffffffccffffffffffffffd6fffffffffffffffcffffffff0000003e00000000",
            INIT_04 => X"0000002200000000000000070000000000000012000000000000001e00000000",
            INIT_05 => X"ffffffaaffffffff0000000400000000ffffffeeffffffffffffffd7ffffffff",
            INIT_06 => X"ffffffe2ffffffff0000005500000000fffffff6ffffffffffffffdfffffffff",
            INIT_07 => X"0000000e00000000fffffff3ffffffff0000004000000000ffffffb1ffffffff",
            INIT_08 => X"ffffffb8fffffffffffffff3ffffffff0000002200000000fffffff7ffffffff",
            INIT_09 => X"ffffffc7ffffffff000000150000000000000001000000000000000e00000000",
            INIT_0A => X"ffffffc2ffffffff0000002e0000000000000017000000000000001a00000000",
            INIT_0B => X"ffffffd2ffffffffffffffe2ffffffffffffffc0ffffffff0000002100000000",
            INIT_0C => X"00000005000000000000000100000000ffffffe0ffffffff0000001a00000000",
            INIT_0D => X"fffffff1ffffffffffffffeeffffffff0000000c000000000000003500000000",
            INIT_0E => X"ffffffd1fffffffffffffff9ffffffff0000001500000000ffffffebffffffff",
            INIT_0F => X"ffffffd7ffffffffffffffe9ffffffff0000000b00000000fffffffeffffffff",
            INIT_10 => X"ffffffd5ffffffffffffffe0ffffffff0000002200000000ffffffe6ffffffff",
            INIT_11 => X"fffffff5ffffffffffffffc1ffffffffffffff93ffffffff0000001e00000000",
            INIT_12 => X"00000009000000000000000f0000000000000036000000000000002500000000",
            INIT_13 => X"0000000b00000000ffffffcaffffffffffffffedffffffff0000000600000000",
            INIT_14 => X"ffffffe9ffffffff0000000a00000000fffffffeffffffff0000002800000000",
            INIT_15 => X"ffffffe9fffffffffffffffaffffffffffffffdaffffffffffffffd0ffffffff",
            INIT_16 => X"ffffffe7ffffffffffffffe3fffffffffffffff1ffffffff0000001c00000000",
            INIT_17 => X"fffffffeffffffff000000170000000000000004000000000000002c00000000",
            INIT_18 => X"ffffffe2ffffffffffffffe8ffffffff0000001400000000fffffffbffffffff",
            INIT_19 => X"0000000c00000000fffffff2ffffffff00000010000000000000002200000000",
            INIT_1A => X"fffffff0ffffffffffffff9efffffffffffffffcffffffffffffffe1ffffffff",
            INIT_1B => X"ffffffefffffffffffffff94fffffffffffffff1ffffffff0000001900000000",
            INIT_1C => X"0000001100000000000000040000000000000020000000000000003d00000000",
            INIT_1D => X"fffffffbffffffffffffffe3ffffffff00000009000000000000004600000000",
            INIT_1E => X"ffffffefffffffffffffffdcfffffffffffffff4ffffffff0000001200000000",
            INIT_1F => X"0000000000000000fffffffeffffffff00000002000000000000000700000000",
            INIT_20 => X"0000001b00000000ffffffedffffffff0000002500000000ffffffe1ffffffff",
            INIT_21 => X"00000014000000000000000300000000ffffffa6ffffffff0000001900000000",
            INIT_22 => X"fffffff3ffffffff0000001e00000000fffffff5ffffffff0000000900000000",
            INIT_23 => X"fffffffeffffffff0000000a00000000fffffff0ffffffff0000001200000000",
            INIT_24 => X"ffffffedffffffff0000004b00000000fffffff9fffffffffffffff1ffffffff",
            INIT_25 => X"0000000a00000000ffffffe5ffffffffffffffc4fffffffffffffff8ffffffff",
            INIT_26 => X"ffffffd4ffffffff00000002000000000000000b000000000000001d00000000",
            INIT_27 => X"0000001300000000ffffffe0ffffffff0000001d00000000ffffffe4ffffffff",
            INIT_28 => X"000000130000000000000012000000000000001600000000ffffffefffffffff",
            INIT_29 => X"0000000f000000000000001900000000ffffffe5ffffffff0000002200000000",
            INIT_2A => X"ffffffdfffffffffffffffe4ffffffffffffffe8fffffffffffffff3ffffffff",
            INIT_2B => X"0000001300000000fffffff5ffffffffffffffd1fffffffffffffffeffffffff",
            INIT_2C => X"fffffff0fffffffffffffffcffffffff00000029000000000000003b00000000",
            INIT_2D => X"0000000900000000ffffffecffffffffffffffecfffffffffffffffbffffffff",
            INIT_2E => X"ffffffadfffffffffffffff0ffffffff00000007000000000000002200000000",
            INIT_2F => X"ffffffdcffffffffffffffc5ffffffff0000000600000000fffffff1ffffffff",
            INIT_30 => X"000000140000000000000010000000000000000d000000000000002c00000000",
            INIT_31 => X"fffffff3ffffffff0000000600000000ffffffddffffffff0000001600000000",
            INIT_32 => X"ffffffdcfffffffffffffff3ffffffff0000002300000000fffffff5ffffffff",
            INIT_33 => X"fffffff1ffffffffffffffd5ffffffff00000006000000000000003100000000",
            INIT_34 => X"ffffffedffffffffffffffefffffffff00000012000000000000001700000000",
            INIT_35 => X"0000000a000000000000000a00000000ffffffd8ffffffff0000000d00000000",
            INIT_36 => X"fffffffbffffffffffffffe7ffffffff0000002b000000000000002300000000",
            INIT_37 => X"00000006000000000000001700000000fffffff6ffffffffffffffebffffffff",
            INIT_38 => X"ffffffd4ffffffffffffffefffffffff00000014000000000000000a00000000",
            INIT_39 => X"0000001100000000ffffffedffffffff00000017000000000000002d00000000",
            INIT_3A => X"ffffffceffffffff0000000000000000ffffffefffffffffffffffdfffffffff",
            INIT_3B => X"ffffffefffffffffffffffceffffffffffffffefffffffff0000000400000000",
            INIT_3C => X"fffffff3fffffffffffffff9ffffffff0000002f000000000000002600000000",
            INIT_3D => X"0000001400000000fffffffaffffffff00000014000000000000000d00000000",
            INIT_3E => X"ffffffadffffffff0000000a000000000000002300000000fffffff5ffffffff",
            INIT_3F => X"ffffffedffffffffffffffe7ffffffff0000000e000000000000002800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"ffffffe9ffffffff000000040000000000000016000000000000002b00000000",
            INIT_41 => X"fffffff1ffffffffffffffd8ffffffffffffffc4ffffffff0000001800000000",
            INIT_42 => X"0000002100000000000000190000000000000018000000000000001900000000",
            INIT_43 => X"ffffffe7ffffffff0000000000000000fffffff8ffffffff0000002d00000000",
            INIT_44 => X"ffffffefffffffffffffffd0fffffffffffffff6ffffffff0000000100000000",
            INIT_45 => X"0000001c00000000fffffff6ffffffffffffffbfffffffff0000000500000000",
            INIT_46 => X"ffffffe6fffffffffffffff6ffffffff0000000900000000fffffff9ffffffff",
            INIT_47 => X"0000002b00000000ffffffcefffffffffffffffeffffffff0000001500000000",
            INIT_48 => X"ffffffd0ffffffff00000006000000000000000000000000ffffffedffffffff",
            INIT_49 => X"0000000c00000000fffffffbffffffff0000000600000000ffffffcaffffffff",
            INIT_4A => X"ffffffbefffffffffffffffbffffffffffffffe1ffffffff0000001500000000",
            INIT_4B => X"0000002b00000000000000160000000000000000000000000000000600000000",
            INIT_4C => X"ffffffe9ffffffffffffffe6ffffffffffffffe5ffffffff0000000d00000000",
            INIT_4D => X"0000000200000000ffffffb0ffffffff00000012000000000000002b00000000",
            INIT_4E => X"ffffffffffffffffffffffedffffffffffffffddffffffff0000000f00000000",
            INIT_4F => X"00000005000000000000000200000000fffffff7fffffffffffffff8ffffffff",
            INIT_50 => X"0000002e000000000000001a00000000fffffffdffffffff0000000500000000",
            INIT_51 => X"ffffffb1ffffffffffffffe6ffffffff0000000900000000fffffff3ffffffff",
            INIT_52 => X"00000005000000000000002a000000000000001900000000fffffffeffffffff",
            INIT_53 => X"0000000a000000000000001b000000000000000d000000000000000200000000",
            INIT_54 => X"fffffffdffffffffffffffc6ffffffff0000000300000000ffffffe4ffffffff",
            INIT_55 => X"0000000000000000ffffffedffffffff00000004000000000000004900000000",
            INIT_56 => X"0000000700000000ffffffd7ffffffff0000000700000000ffffffddffffffff",
            INIT_57 => X"0000001b00000000ffffffc5ffffffffffffffdafffffffffffffff4ffffffff",
            INIT_58 => X"ffffffbefffffffffffffff2ffffffffffffffd7ffffffffffffffedffffffff",
            INIT_59 => X"0000000b00000000000000140000000000000000000000000000000500000000",
            INIT_5A => X"ffffffeefffffffffffffffffffffffffffffff3ffffffffffffffefffffffff",
            INIT_5B => X"fffffff0ffffffff0000001b000000000000000f000000000000001900000000",
            INIT_5C => X"000000130000000000000021000000000000001a000000000000003e00000000",
            INIT_5D => X"fffffffeffffffffffffffe5ffffffff0000000c000000000000001e00000000",
            INIT_5E => X"ffffffa3ffffffff00000000000000000000002d000000000000000f00000000",
            INIT_5F => X"00000015000000000000000f000000000000001200000000ffffffe9ffffffff",
            INIT_60 => X"0000001f00000000000000270000000000000022000000000000001100000000",
            INIT_61 => X"0000000400000000fffffff3ffffffff0000003400000000ffffffddffffffff",
            INIT_62 => X"00000020000000000000000a000000000000000200000000fffffffcffffffff",
            INIT_63 => X"0000002e000000000000001100000000fffffff8ffffffffffffffc3ffffffff",
            INIT_64 => X"ffffffefffffffff00000001000000000000000700000000ffffffd7ffffffff",
            INIT_65 => X"0000001b00000000ffffffdaffffffff0000001e000000000000000000000000",
            INIT_66 => X"ffffffe9ffffffffffffffc3ffffffff0000002500000000fffffff8ffffffff",
            INIT_67 => X"0000004700000000ffffffbcffffffff0000001c00000000ffffffd9ffffffff",
            INIT_68 => X"ffffffbeffffffff0000000800000000fffffff1ffffffff0000001900000000",
            INIT_69 => X"ffffffe6ffffffff0000001600000000fffffff3ffffffff0000001500000000",
            INIT_6A => X"0000001e00000000fffffff9ffffffff00000014000000000000000200000000",
            INIT_6B => X"ffffffecffffffff0000001500000000ffffffedffffffff0000000400000000",
            INIT_6C => X"fffffff8ffffffffffffffe7ffffffff0000001b00000000fffffff5ffffffff",
            INIT_6D => X"0000001200000000fffffff2ffffffff0000001a000000000000001600000000",
            INIT_6E => X"ffffffa1fffffffffffffffcffffffff0000001100000000ffffffdeffffffff",
            INIT_6F => X"0000000e00000000fffffffdffffffffffffffebffffffffffffffc4ffffffff",
            INIT_70 => X"0000000c00000000fffffff1ffffffffffffffdefffffffffffffff8ffffffff",
            INIT_71 => X"0000000600000000fffffff7ffffffff0000001c00000000ffffffeeffffffff",
            INIT_72 => X"0000003a0000000000000019000000000000000400000000fffffff4ffffffff",
            INIT_73 => X"ffffffc7ffffffff0000000d00000000ffffffecffffffffffffffd9ffffffff",
            INIT_74 => X"0000000a00000000ffffffa9ffffffff0000000700000000ffffffd1ffffffff",
            INIT_75 => X"0000002a000000000000002a00000000ffffffd7ffffffffffffffccffffffff",
            INIT_76 => X"ffffffbffffffffffffffff9ffffffff00000021000000000000000700000000",
            INIT_77 => X"ffffffdeffffffffffffffadffffffff0000001c000000000000001f00000000",
            INIT_78 => X"00000005000000000000000800000000fffffff6ffffffff0000001300000000",
            INIT_79 => X"ffffffdcfffffffffffffff4ffffffff0000000c00000000ffffffc8ffffffff",
            INIT_7A => X"ffffffedffffffffffffffe6ffffffff0000000e00000000fffffff3ffffffff",
            INIT_7B => X"0000000000000000ffffffb3ffffffffffffffdaffffffff0000002a00000000",
            INIT_7C => X"ffffffbfffffffffffffffe1ffffffffffffff97fffffffffffffff5ffffffff",
            INIT_7D => X"fffffff2ffffffff00000007000000000000007600000000ffffffcaffffffff",
            INIT_7E => X"ffffffe7ffffffffffffffd7ffffffffffffffaafffffffffffffffaffffffff",
            INIT_7F => X"00000005000000000000002200000000fffffff4ffffffff0000002b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE10;


    MEM_IWGHT_LAYER3_INSTANCE11 : if BRAM_NAME = "iwght_layer3_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"ffffffceffffffffffffffa9ffffffff0000000a000000000000001900000000",
            INIT_01 => X"fffffffaffffffffffffffdeffffffffffffffebffffffffffffffd6ffffffff",
            INIT_02 => X"0000002900000000ffffffdcffffffff0000000b00000000ffffffbdffffffff",
            INIT_03 => X"ffffffebffffffffffffffe9fffffffffffffffdffffffffffffffdbffffffff",
            INIT_04 => X"ffffffe4fffffffffffffff6fffffffffffffff1ffffffffffffffebffffffff",
            INIT_05 => X"0000000c00000000fffffff6fffffffffffffff9fffffffffffffffcffffffff",
            INIT_06 => X"00000008000000000000000200000000fffffff0ffffffff0000002800000000",
            INIT_07 => X"0000000f00000000ffffffdfffffffff00000009000000000000003200000000",
            INIT_08 => X"fffffff4fffffffffffffffbffffffff00000006000000000000001300000000",
            INIT_09 => X"0000000000000000ffffffe7ffffffff0000001500000000fffffff7ffffffff",
            INIT_0A => X"000000110000000000000012000000000000001700000000fffffff5ffffffff",
            INIT_0B => X"fffffff8ffffffffffffffbeffffffffffffffd0ffffffff0000001e00000000",
            INIT_0C => X"fffffff6fffffffffffffff4ffffffffffffffd6ffffffffffffffdfffffffff",
            INIT_0D => X"fffffff6ffffffffffffffffffffffff00000039000000000000000800000000",
            INIT_0E => X"ffffffeaffffffff0000000c00000000ffffffb4ffffffffffffffeeffffffff",
            INIT_0F => X"00000033000000000000001f0000000000000012000000000000000000000000",
            INIT_10 => X"ffffffcaffffffff0000001a0000000000000001000000000000001100000000",
            INIT_11 => X"fffffff2ffffffff00000000000000000000000000000000ffffffcaffffffff",
            INIT_12 => X"0000005600000000fffffffbffffffff0000002300000000ffffffdfffffffff",
            INIT_13 => X"fffffff3ffffffff0000000b00000000ffffffe6ffffffffffffffe4ffffffff",
            INIT_14 => X"ffffffcaffffffffffffffffffffffff0000000f00000000ffffffbcffffffff",
            INIT_15 => X"00000005000000000000001000000000ffffffedffffffffffffffc6ffffffff",
            INIT_16 => X"0000001f00000000ffffffd8ffffffff00000002000000000000001500000000",
            INIT_17 => X"0000002d00000000ffffffc3ffffffff00000006000000000000003800000000",
            INIT_18 => X"0000000c00000000fffffff0ffffffffffffffefffffffff0000003c00000000",
            INIT_19 => X"ffffffbefffffffffffffff1fffffffffffffffbffffffff0000000e00000000",
            INIT_1A => X"00000011000000000000000d0000000000000033000000000000000900000000",
            INIT_1B => X"ffffffd6ffffffffffffffe0ffffffffffffffa1ffffffff0000000600000000",
            INIT_1C => X"ffffffe4ffffffffffffffc0ffffffffffffffdeffffffffffffffc5ffffffff",
            INIT_1D => X"0000001400000000000000000000000000000052000000000000002700000000",
            INIT_1E => X"fffffff7ffffffffffffffd9ffffffffffffffc0ffffffffffffffceffffffff",
            INIT_1F => X"00000032000000000000000500000000fffffff2ffffffffffffffc6ffffffff",
            INIT_20 => X"ffffffdfffffffffffffffcfffffffff0000000f000000000000000200000000",
            INIT_21 => X"00000014000000000000000000000000fffffffeffffffffffffffdfffffffff",
            INIT_22 => X"fffffff9ffffffffffffffe2ffffffff",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER3_INSTANCE11;


    MEM_IFMAP_LAYER0_INSTANCE0 : if BRAM_NAME = "ifmap_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE0;


    MEM_IFMAP_LAYER0_INSTANCE1 : if BRAM_NAME = "ifmap_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE1;


    MEM_IFMAP_LAYER0_INSTANCE2 : if BRAM_NAME = "ifmap_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE2;


    MEM_IFMAP_LAYER0_INSTANCE3 : if BRAM_NAME = "ifmap_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE3;


    MEM_IFMAP_LAYER0_INSTANCE4 : if BRAM_NAME = "ifmap_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE4;


    MEM_IFMAP_LAYER0_INSTANCE5 : if BRAM_NAME = "ifmap_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE0 : if BRAM_NAME = "ifmap_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000014000000000000000f0000000000000012000000000000001200000000",
            INIT_01 => X"0000001d000000000000000f000000000000000d000000000000001700000000",
            INIT_02 => X"000000010000000000000000000000000000000a000000000000001d00000000",
            INIT_03 => X"000000160000000000000015000000000000000c000000000000000600000000",
            INIT_04 => X"000000130000000000000013000000000000000f000000000000001200000000",
            INIT_05 => X"0000000000000000000000030000000000000008000000000000000400000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_07 => X"0000000b0000000000000000000000000000000b000000000000000500000000",
            INIT_08 => X"0000001b0000000000000012000000000000001b000000000000001300000000",
            INIT_09 => X"000000000000000000000000000000000000001e000000000000002000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000c00000000000000000000000000000001000000000000000100000000",
            INIT_0C => X"000000000000000000000011000000000000000b000000000000001900000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000300000000000000030000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000001c000000000000000400000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_20 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000007000000000000000400000000",
            INIT_5A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000a000000000000003f000000000000000f000000000000001a00000000",
            INIT_62 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000002000000000000000250000000000000038000000000000003a00000000",
            INIT_64 => X"0000002700000000000000250000000000000029000000000000002200000000",
            INIT_65 => X"00000000000000000000003a000000000000002c000000000000002000000000",
            INIT_66 => X"0000001d000000000000001d000000000000001e000000000000000000000000",
            INIT_67 => X"00000024000000000000001f0000000000000020000000000000002000000000",
            INIT_68 => X"0000002100000000000000280000000000000022000000000000001e00000000",
            INIT_69 => X"0000000e000000000000002f000000000000002f000000000000003000000000",
            INIT_6A => X"0000001d00000000000000190000000000000021000000000000000f00000000",
            INIT_6B => X"00000033000000000000002f0000000000000023000000000000002200000000",
            INIT_6C => X"00000029000000000000003a0000000000000028000000000000003400000000",
            INIT_6D => X"0000002a00000000000000410000000000000031000000000000003300000000",
            INIT_6E => X"00000017000000000000001f000000000000002a000000000000003000000000",
            INIT_6F => X"0000001a000000000000002d0000000000000021000000000000001c00000000",
            INIT_70 => X"0000000000000000000000000000000000000029000000000000001c00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000006000000000000000e0000000000000018000000000000000300000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_7D => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_7E => X"0000000000000000000000060000000000000000000000000000001b00000000",
            INIT_7F => X"0000001e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE0;


    MEM_IFMAP_LAYER1_INSTANCE1 : if BRAM_NAME = "ifmap_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001400000000000000110000000000000000000000000000000000000000",
            INIT_01 => X"0000001d00000000000000000000000000000003000000000000000500000000",
            INIT_02 => X"0000000000000000000000080000000000000000000000000000001000000000",
            INIT_03 => X"000000000000000000000017000000000000000f000000000000000300000000",
            INIT_04 => X"00000006000000000000000a000000000000001a000000000000000000000000",
            INIT_05 => X"0000000300000000000000440000000000000000000000000000000400000000",
            INIT_06 => X"000000020000000000000000000000000000000b000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000000b000000000000001700000000",
            INIT_08 => X"00000000000000000000000b000000000000001e000000000000000c00000000",
            INIT_09 => X"0000000400000000000000000000000000000037000000000000000000000000",
            INIT_0A => X"0000002000000000000000020000000000000011000000000000000a00000000",
            INIT_0B => X"0000000600000000000000000000000000000006000000000000001400000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_0D => X"0000001100000000000000000000000000000000000000000000002000000000",
            INIT_0E => X"00000028000000000000001d0000000000000000000000000000000800000000",
            INIT_0F => X"0000000000000000000000080000000000000011000000000000000400000000",
            INIT_10 => X"00000000000000000000000b000000000000000b000000000000000000000000",
            INIT_11 => X"0000000000000000000000060000000000000000000000000000001000000000",
            INIT_12 => X"0000000000000000000000240000000000000018000000000000000000000000",
            INIT_13 => X"000000120000000000000009000000000000000e000000000000002700000000",
            INIT_14 => X"0000000000000000000000000000000000000015000000000000001200000000",
            INIT_15 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_16 => X"0000005800000000000000000000000000000023000000000000002b00000000",
            INIT_17 => X"00000011000000000000002d0000000000000028000000000000000d00000000",
            INIT_18 => X"00000022000000000000001b0000000000000000000000000000000000000000",
            INIT_19 => X"000000360000000000000000000000000000000b000000000000001f00000000",
            INIT_1A => X"0000000000000000000000450000000000000012000000000000002300000000",
            INIT_1B => X"0000001a0000000000000021000000000000001f000000000000000700000000",
            INIT_1C => X"0000002e00000000000000280000000000000022000000000000001e00000000",
            INIT_1D => X"00000038000000000000002a000000000000002f000000000000002f00000000",
            INIT_1E => X"0000002700000000000000000000000000000025000000000000003300000000",
            INIT_1F => X"0000002a00000000000000240000000000000024000000000000002500000000",
            INIT_20 => X"0000002e000000000000002f0000000000000036000000000000002f00000000",
            INIT_21 => X"00000052000000000000002e000000000000002c000000000000003a00000000",
            INIT_22 => X"00000026000000000000002b0000000000000013000000000000000000000000",
            INIT_23 => X"0000002e000000000000002f000000000000002a000000000000002a00000000",
            INIT_24 => X"000000280000000000000045000000000000002a000000000000002f00000000",
            INIT_25 => X"00000019000000000000002c0000000000000033000000000000002b00000000",
            INIT_26 => X"0000002400000000000000230000000000000028000000000000001900000000",
            INIT_27 => X"0000002e000000000000002d0000000000000031000000000000002e00000000",
            INIT_28 => X"00000000000000000000001f000000000000003a000000000000004300000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000000000000000000000a000000000000000200000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000170000000000000008000000000000001000000000",
            INIT_2F => X"000000000000000000000003000000000000001c000000000000001f00000000",
            INIT_30 => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_31 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000004200000000000000000000000000000000000000000000001100000000",
            INIT_33 => X"000000000000000000000000000000000000003f000000000000002d00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_35 => X"0000002c00000000000000280000000000000000000000000000000e00000000",
            INIT_36 => X"00000026000000000000005a0000000000000000000000000000002500000000",
            INIT_37 => X"0000006c0000000000000000000000000000002a000000000000003b00000000",
            INIT_38 => X"0000003400000000000000000000000000000023000000000000000500000000",
            INIT_39 => X"0000003c0000000000000048000000000000005d000000000000002400000000",
            INIT_3A => X"0000001e0000000000000052000000000000002f000000000000000000000000",
            INIT_3B => X"0000003100000000000000590000000000000000000000000000003e00000000",
            INIT_3C => X"0000002c00000000000000000000000000000000000000000000003700000000",
            INIT_3D => X"000000000000000000000060000000000000003e000000000000006100000000",
            INIT_3E => X"000000310000000000000012000000000000005c000000000000007300000000",
            INIT_3F => X"0000001500000000000000730000000000000048000000000000002500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005a00000000000000000000000000000000000000000000003800000000",
            INIT_41 => X"000000750000000000000000000000000000006a000000000000004a00000000",
            INIT_42 => X"00000037000000000000000c0000000000000012000000000000004700000000",
            INIT_43 => X"0000003100000000000000280000000000000065000000000000004d00000000",
            INIT_44 => X"00000038000000000000008b0000000000000006000000000000000000000000",
            INIT_45 => X"00000050000000000000004f0000000000000000000000000000004600000000",
            INIT_46 => X"0000006800000000000000130000000000000025000000000000000600000000",
            INIT_47 => X"0000002a000000000000000b0000000000000084000000000000004200000000",
            INIT_48 => X"00000000000000000000002c000000000000002e000000000000001300000000",
            INIT_49 => X"00000004000000000000005b0000000000000016000000000000002900000000",
            INIT_4A => X"0000003a000000000000004a0000000000000000000000000000000000000000",
            INIT_4B => X"0000001800000000000000640000000000000000000000000000009f00000000",
            INIT_4C => X"0000003b0000000000000030000000000000004d000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000017000000000000005a00000000",
            INIT_4E => X"00000094000000000000003c000000000000000f000000000000000c00000000",
            INIT_4F => X"00000020000000000000004c0000000000000093000000000000000000000000",
            INIT_50 => X"0000001a00000000000000410000000000000083000000000000007100000000",
            INIT_51 => X"0000003100000000000000200000000000000023000000000000001d00000000",
            INIT_52 => X"00000000000000000000004e000000000000002b000000000000001d00000000",
            INIT_53 => X"0000003c000000000000003a000000000000007300000000000000d800000000",
            INIT_54 => X"0000003c000000000000003d0000000000000038000000000000004700000000",
            INIT_55 => X"0000005f000000000000004f0000000000000040000000000000003e00000000",
            INIT_56 => X"000000af00000000000000820000000000000000000000000000001200000000",
            INIT_57 => X"0000003e000000000000003f0000000000000049000000000000004200000000",
            INIT_58 => X"0000005000000000000000400000000000000038000000000000003900000000",
            INIT_59 => X"00000045000000000000006a000000000000003d000000000000004800000000",
            INIT_5A => X"00000039000000000000005a00000000000000cb000000000000000000000000",
            INIT_5B => X"00000041000000000000003c0000000000000042000000000000004d00000000",
            INIT_5C => X"00000038000000000000004e000000000000004d000000000000004800000000",
            INIT_5D => X"0000003e000000000000004b0000000000000076000000000000007b00000000",
            INIT_5E => X"0000004300000000000000350000000000000048000000000000005400000000",
            INIT_5F => X"0000005500000000000000440000000000000038000000000000004400000000",
            INIT_60 => X"00000080000000000000006f000000000000001a000000000000003a00000000",
            INIT_61 => X"0000000800000000000000080000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000050000000000000003000000000000000600000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_64 => X"0000000700000000000000050000000000000006000000000000000000000000",
            INIT_65 => X"0000000a0000000000000007000000000000000c000000000000000a00000000",
            INIT_66 => X"000000000000000000000000000000000000001a000000000000004900000000",
            INIT_67 => X"0000000000000000000000060000000000000024000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_69 => X"0000000000000000000000070000000000000004000000000000000400000000",
            INIT_6A => X"0000001a000000000000000d0000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000170000000000000007000000000000001500000000",
            INIT_6C => X"0000000900000000000000250000000000000028000000000000000000000000",
            INIT_6D => X"000000370000000000000000000000000000000d000000000000000500000000",
            INIT_6E => X"0000000000000000000000000000000000000005000000000000001b00000000",
            INIT_6F => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_70 => X"0000000b0000000000000013000000000000005a000000000000002600000000",
            INIT_71 => X"0000000e00000000000000060000000000000056000000000000008000000000",
            INIT_72 => X"0000002500000000000000250000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000018000000000000000f00000000",
            INIT_74 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_75 => X"0000001f000000000000001a000000000000002a000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_77 => X"0000000700000000000000060000000000000027000000000000000900000000",
            INIT_78 => X"0000002100000000000000000000000000000004000000000000000000000000",
            INIT_79 => X"000000110000000000000009000000000000000a000000000000000000000000",
            INIT_7A => X"000000170000000000000000000000000000000b000000000000000000000000",
            INIT_7B => X"0000001c00000000000000070000000000000015000000000000001d00000000",
            INIT_7C => X"0000000000000000000000160000000000000019000000000000001000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000004000000000000000b0000000000000004000000000000001000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE1;


    MEM_IFMAP_LAYER1_INSTANCE2 : if BRAM_NAME = "ifmap_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001a00000000000000000000000000000000000000000000001c00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_02 => X"00000000000000000000002f0000000000000003000000000000000000000000",
            INIT_03 => X"0000001100000000000000040000000000000009000000000000000000000000",
            INIT_04 => X"0000000c000000000000004a0000000000000000000000000000000000000000",
            INIT_05 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_07 => X"00000085000000000000009c0000000000000046000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_09 => X"00000000000000000000001b0000000000000041000000000000002000000000",
            INIT_0A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000001200000000000000070000000000000004000000000000000000000000",
            INIT_11 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000001300000000000000140000000000000000000000000000000000000000",
            INIT_18 => X"0000002200000000000000280000000000000000000000000000000400000000",
            INIT_19 => X"000000a200000000000000a3000000000000009d000000000000000000000000",
            INIT_1A => X"000000ac000000000000009d00000000000000a400000000000000a500000000",
            INIT_1B => X"0000007c000000000000009400000000000000ad00000000000000b700000000",
            INIT_1C => X"0000009200000000000000920000000000000084000000000000007c00000000",
            INIT_1D => X"000000ac00000000000000a800000000000000ad00000000000000a200000000",
            INIT_1E => X"000000a000000000000000a9000000000000008c00000000000000a000000000",
            INIT_1F => X"0000003e000000000000002e000000000000003a000000000000007a00000000",
            INIT_20 => X"00000089000000000000008b000000000000006e000000000000004e00000000",
            INIT_21 => X"000000af00000000000000b000000000000000ac000000000000006a00000000",
            INIT_22 => X"0000002d00000000000000480000000000000073000000000000008e00000000",
            INIT_23 => X"00000027000000000000000a000000000000001e000000000000000700000000",
            INIT_24 => X"0000002b000000000000004d0000000000000067000000000000003a00000000",
            INIT_25 => X"0000005900000000000000a200000000000000aa00000000000000a400000000",
            INIT_26 => X"0000000c00000000000000150000000000000027000000000000004d00000000",
            INIT_27 => X"00000025000000000000001b000000000000002d000000000000003300000000",
            INIT_28 => X"00000094000000000000001f0000000000000017000000000000003a00000000",
            INIT_29 => X"000000430000000000000047000000000000004e000000000000006000000000",
            INIT_2A => X"000000310000000000000000000000000000001f000000000000002f00000000",
            INIT_2B => X"0000002f000000000000001c0000000000000017000000000000003900000000",
            INIT_2C => X"00000099000000000000008e0000000000000012000000000000001600000000",
            INIT_2D => X"000000310000000000000045000000000000003b000000000000002500000000",
            INIT_2E => X"0000002a000000000000003e0000000000000000000000000000002d00000000",
            INIT_2F => X"0000000e00000000000000170000000000000012000000000000001000000000",
            INIT_30 => X"0000002f000000000000009f0000000000000062000000000000002a00000000",
            INIT_31 => X"0000002f000000000000002d000000000000003e000000000000003200000000",
            INIT_32 => X"0000001000000000000000280000000000000032000000000000000000000000",
            INIT_33 => X"0000000a000000000000001c0000000000000026000000000000000e00000000",
            INIT_34 => X"0000002600000000000000370000000000000062000000000000002c00000000",
            INIT_35 => X"0000001e00000000000000290000000000000027000000000000002e00000000",
            INIT_36 => X"000000220000000000000009000000000000002d000000000000002f00000000",
            INIT_37 => X"0000002b00000000000000000000000000000014000000000000004100000000",
            INIT_38 => X"0000003600000000000000220000000000000055000000000000000e00000000",
            INIT_39 => X"000000420000000000000054000000000000000d000000000000003000000000",
            INIT_3A => X"00000079000000000000002d000000000000000f000000000000002600000000",
            INIT_3B => X"0000000000000000000000240000000000000005000000000000001000000000",
            INIT_3C => X"0000002800000000000000080000000000000020000000000000003500000000",
            INIT_3D => X"00000006000000000000001d0000000000000034000000000000002d00000000",
            INIT_3E => X"00000000000000000000008a0000000000000062000000000000000900000000",
            INIT_3F => X"0000001700000000000000000000000000000023000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000600000000000000000000000000000000000000000000001a00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"00000000000000000000003a0000000000000006000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000002300000000000000220000000000000000000000000000000000000000",
            INIT_52 => X"00000027000000000000001e0000000000000020000000000000002500000000",
            INIT_53 => X"00000017000000000000001d0000000000000024000000000000002600000000",
            INIT_54 => X"0000001e00000000000000240000000000000026000000000000001a00000000",
            INIT_55 => X"0000002a000000000000002c0000000000000023000000000000001800000000",
            INIT_56 => X"0000000f00000000000000200000000000000028000000000000001f00000000",
            INIT_57 => X"00000000000000000000001d000000000000000e000000000000001d00000000",
            INIT_58 => X"0000001c000000000000002b0000000000000020000000000000000900000000",
            INIT_59 => X"0000002100000000000000280000000000000039000000000000000600000000",
            INIT_5A => X"000000060000000000000000000000000000001a000000000000002700000000",
            INIT_5B => X"000000000000000000000000000000000000002e000000000000002100000000",
            INIT_5C => X"00000000000000000000002c0000000000000025000000000000000000000000",
            INIT_5D => X"0000000f00000000000000290000000000000021000000000000004c00000000",
            INIT_5E => X"0000000000000000000000000000000000000004000000000000002400000000",
            INIT_5F => X"0000000000000000000000090000000000000000000000000000004800000000",
            INIT_60 => X"000000260000000000000000000000000000004a000000000000000000000000",
            INIT_61 => X"0000000b00000000000000090000000000000056000000000000000200000000",
            INIT_62 => X"0000005900000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_64 => X"00000000000000000000000a0000000000000000000000000000002b00000000",
            INIT_65 => X"000000000000000000000013000000000000003e000000000000001a00000000",
            INIT_66 => X"00000000000000000000008e0000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_68 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000036000000000000003f00000000",
            INIT_6A => X"0000000000000000000000000000000000000066000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000015000000000000000a00000000",
            INIT_6C => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_6E => X"0000001d00000000000000000000000000000000000000000000004200000000",
            INIT_6F => X"0000000200000000000000000000000000000008000000000000000f00000000",
            INIT_70 => X"0000001100000000000000040000000000000021000000000000000000000000",
            INIT_71 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_72 => X"00000021000000000000001e0000000000000000000000000000002500000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_74 => X"00000027000000000000000f0000000000000000000000000000002c00000000",
            INIT_75 => X"0000000000000000000000050000000000000002000000000000000000000000",
            INIT_76 => X"0000001400000000000000340000000000000030000000000000000c00000000",
            INIT_77 => X"0000007800000000000000000000000000000004000000000000002a00000000",
            INIT_78 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_79 => X"0000000900000000000000080000000000000000000000000000000000000000",
            INIT_7A => X"0000002000000000000000000000000000000000000000000000000100000000",
            INIT_7B => X"0000000000000000000000400000000000000000000000000000001400000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE2;


    MEM_IFMAP_LAYER1_INSTANCE3 : if BRAM_NAME = "ifmap_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000005d00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000002b00000000000000000000000000000000000000000000000400000000",
            INIT_0A => X"0000002f000000000000002c000000000000002d000000000000003000000000",
            INIT_0B => X"00000037000000000000003a0000000000000030000000000000002900000000",
            INIT_0C => X"0000002700000000000000260000000000000025000000000000002a00000000",
            INIT_0D => X"00000035000000000000002c0000000000000031000000000000002a00000000",
            INIT_0E => X"00000000000000000000002d000000000000002e000000000000003000000000",
            INIT_0F => X"0000000c000000000000003b0000000000000029000000000000001f00000000",
            INIT_10 => X"0000001f000000000000000e0000000000000000000000000000000000000000",
            INIT_11 => X"0000002e0000000000000029000000000000001c000000000000002500000000",
            INIT_12 => X"0000002d000000000000003b0000000000000032000000000000003500000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_14 => X"0000001a00000000000000040000000000000000000000000000000000000000",
            INIT_15 => X"0000003200000000000000230000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000019000000000000002500000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000110000000000000000000000000000000600000000",
            INIT_19 => X"0000000000000000000000180000000000000012000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_1D => X"0000000300000000000000030000000000000038000000000000000b00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000007000000000000003a00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000005000000000000001a00000000",
            INIT_2A => X"0000000400000000000000180000000000000003000000000000000f00000000",
            INIT_2B => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000000000a000000000000001100000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000800000000000000080000000000000011000000000000000a00000000",
            INIT_43 => X"0000000b000000000000000c000000000000000c000000000000000400000000",
            INIT_44 => X"00000023000000000000002d0000000000000021000000000000000b00000000",
            INIT_45 => X"0000000000000000000000060000000000000008000000000000001100000000",
            INIT_46 => X"00000008000000000000000c000000000000000a000000000000000a00000000",
            INIT_47 => X"0000004200000000000000230000000000000005000000000000000000000000",
            INIT_48 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"000000330000000000000035000000000000000a000000000000001700000000",
            INIT_4A => X"0000003700000000000000050000000000000008000000000000000500000000",
            INIT_4B => X"0000000000000000000000000000000000000009000000000000001600000000",
            INIT_4C => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000500000000000000000000000000000000000000000000000c00000000",
            INIT_4E => X"0000000000000000000000000000000000000008000000000000000800000000",
            INIT_4F => X"00000004000000000000001a0000000000000000000000000000000200000000",
            INIT_50 => X"0000000e00000000000000000000000000000006000000000000001000000000",
            INIT_51 => X"0000000e00000000000000020000000000000000000000000000000100000000",
            INIT_52 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_54 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000003e00000000000000030000000000000006000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_57 => X"0000000700000000000000150000000000000014000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000120000000000000018000000000000001c00000000",
            INIT_5A => X"0000000000000000000000110000000000000000000000000000003100000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000003500000000000000350000000000000002000000000000000000000000",
            INIT_5E => X"000000090000000000000000000000000000000e000000000000002100000000",
            INIT_5F => X"00000000000000000000000e0000000000000005000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000026000000000000000000000000",
            INIT_62 => X"0000003000000000000000260000000000000000000000000000000000000000",
            INIT_63 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000002300000000000000000000000000000004000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_66 => X"0000000000000000000000110000000000000036000000000000004e00000000",
            INIT_67 => X"0000000000000000000000030000000000000018000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_69 => X"0000000000000000000000370000000000000051000000000000001e00000000",
            INIT_6A => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000c00000000000000210000000000000035000000000000000a00000000",
            INIT_6C => X"0000000400000000000000280000000000000056000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000003000000000000000500000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001800000000000000000000000000000016000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000b000000000000004f0000000000000018000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_77 => X"0000000300000000000000000000000000000022000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000a0000000000000013000000000000000d000000000000000000000000",
            INIT_7B => X"0000000800000000000000150000000000000009000000000000000e00000000",
            INIT_7C => X"00000022000000000000001c000000000000000c000000000000000600000000",
            INIT_7D => X"0000000200000000000000060000000000000013000000000000001b00000000",
            INIT_7E => X"0000000d0000000000000009000000000000000b000000000000000800000000",
            INIT_7F => X"0000001a000000000000000f0000000000000036000000000000000f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE3;


    MEM_IFMAP_LAYER1_INSTANCE4 : if BRAM_NAME = "ifmap_layer1_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002400000000000000350000000000000034000000000000001f00000000",
            INIT_01 => X"00000026000000000000000a000000000000001a000000000000002100000000",
            INIT_02 => X"00000008000000000000000a000000000000000b000000000000002400000000",
            INIT_03 => X"0000002000000000000000280000000000000033000000000000005100000000",
            INIT_04 => X"0000002b000000000000004b000000000000005e000000000000005300000000",
            INIT_05 => X"000000140000000000000033000000000000001a000000000000001900000000",
            INIT_06 => X"0000002e00000000000000190000000000000012000000000000000e00000000",
            INIT_07 => X"0000005b0000000000000036000000000000002f000000000000004500000000",
            INIT_08 => X"00000015000000000000003b0000000000000042000000000000005d00000000",
            INIT_09 => X"00000015000000000000005e0000000000000071000000000000001b00000000",
            INIT_0A => X"000000640000000000000044000000000000007e000000000000003500000000",
            INIT_0B => X"00000067000000000000003b0000000000000033000000000000003b00000000",
            INIT_0C => X"0000000100000000000000250000000000000039000000000000003800000000",
            INIT_0D => X"000000130000000000000028000000000000009e000000000000007f00000000",
            INIT_0E => X"0000004b000000000000007d000000000000007e00000000000000bd00000000",
            INIT_0F => X"00000050000000000000007f000000000000005b000000000000002e00000000",
            INIT_10 => X"0000007a0000000000000015000000000000003c000000000000004700000000",
            INIT_11 => X"0000005a00000000000000170000000000000043000000000000009400000000",
            INIT_12 => X"0000004e000000000000006500000000000000a8000000000000007500000000",
            INIT_13 => X"0000003b00000000000000460000000000000081000000000000007800000000",
            INIT_14 => X"000000a5000000000000008e0000000000000033000000000000004c00000000",
            INIT_15 => X"000000a500000000000000390000000000000039000000000000004000000000",
            INIT_16 => X"0000005f0000000000000050000000000000006a000000000000008500000000",
            INIT_17 => X"0000004b0000000000000048000000000000004c000000000000007800000000",
            INIT_18 => X"0000006600000000000000b800000000000000b0000000000000002600000000",
            INIT_19 => X"0000005900000000000000660000000000000038000000000000007300000000",
            INIT_1A => X"0000006500000000000000330000000000000051000000000000004e00000000",
            INIT_1B => X"0000000e000000000000002b000000000000002c000000000000004100000000",
            INIT_1C => X"00000075000000000000008600000000000000b300000000000000c000000000",
            INIT_1D => X"00000079000000000000005f0000000000000033000000000000006f00000000",
            INIT_1E => X"000000250000000000000040000000000000005a000000000000004200000000",
            INIT_1F => X"000000c700000000000000270000000000000027000000000000002f00000000",
            INIT_20 => X"0000009e00000000000000a2000000000000008b00000000000000ab00000000",
            INIT_21 => X"0000007900000000000000b90000000000000091000000000000006500000000",
            INIT_22 => X"0000005a00000000000000470000000000000040000000000000003c00000000",
            INIT_23 => X"000000cb00000000000000c10000000000000068000000000000007100000000",
            INIT_24 => X"000000a500000000000000e700000000000000c9000000000000009d00000000",
            INIT_25 => X"0000006f000000000000007c0000000000000085000000000000008a00000000",
            INIT_26 => X"0000008a00000000000000880000000000000080000000000000007800000000",
            INIT_27 => X"000000b100000000000000a1000000000000008c000000000000008e00000000",
            INIT_28 => X"00000075000000000000007a00000000000000af00000000000000e500000000",
            INIT_29 => X"0000008400000000000000760000000000000071000000000000007000000000",
            INIT_2A => X"000000a3000000000000009a0000000000000095000000000000008c00000000",
            INIT_2B => X"000000ef00000000000000a60000000000000085000000000000009d00000000",
            INIT_2C => X"0000007300000000000000790000000000000080000000000000008800000000",
            INIT_2D => X"0000009b000000000000008c0000000000000082000000000000007700000000",
            INIT_2E => X"0000009700000000000000ab00000000000000a3000000000000009300000000",
            INIT_2F => X"0000007400000000000000a7000000000000007f000000000000008f00000000",
            INIT_30 => X"0000007c000000000000007e0000000000000089000000000000007f00000000",
            INIT_31 => X"0000009a00000000000000850000000000000086000000000000008800000000",
            INIT_32 => X"000000000000000000000000000000000000008d00000000000000af00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000000b000000000000001c00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000033000000000000001400000000",
            INIT_39 => X"000000000000000000000000000000000000001e000000000000001400000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_3B => X"00000028000000000000001c000000000000003e000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000190000000000000000000000000000001e000000000000000700000000",
            INIT_3E => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000006000000000000001a0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_43 => X"00000000000000000000001d0000000000000004000000000000000f00000000",
            INIT_44 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_45 => X"000000020000000000000000000000000000002f000000000000002500000000",
            INIT_46 => X"0000000000000000000000000000000000000003000000000000004f00000000",
            INIT_47 => X"0000002600000000000000000000000000000006000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_49 => X"0000000d000000000000000d0000000000000018000000000000000000000000",
            INIT_4A => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_4B => X"0000000800000000000000180000000000000000000000000000000900000000",
            INIT_4C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_4E => X"00000000000000000000001e000000000000003d000000000000000000000000",
            INIT_4F => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_51 => X"0000003200000000000000220000000000000000000000000000002e00000000",
            INIT_52 => X"0000003600000000000000000000000000000000000000000000000300000000",
            INIT_53 => X"00000000000000000000000d000000000000003a000000000000002600000000",
            INIT_54 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000150000000000000012000000000000000000000000",
            INIT_56 => X"00000031000000000000001f000000000000002e000000000000000000000000",
            INIT_57 => X"0000000800000000000000000000000000000000000000000000000100000000",
            INIT_58 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_59 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000000000000000000000000000000000000d000000000000000f00000000",
            INIT_5B => X"0000004100000000000000210000000000000016000000000000000000000000",
            INIT_5C => X"000000a200000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000c0000000000000037000000000000003f000000000000005200000000",
            INIT_5E => X"0000000000000000000000020000000000000000000000000000000600000000",
            INIT_5F => X"00000036000000000000000d0000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000560000000000000041000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_62 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_63 => X"0000002500000000000000000000000000000002000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000006000000000000003e00000000",
            INIT_65 => X"0000000700000000000000000000000000000000000000000000000100000000",
            INIT_66 => X"0000004200000000000000000000000000000000000000000000000a00000000",
            INIT_67 => X"0000003600000000000000180000000000000000000000000000000c00000000",
            INIT_68 => X"0000000000000000000000090000000000000013000000000000002400000000",
            INIT_69 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000000000000000000001f0000000000000004000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"000000070000000000000000000000000000002d000000000000000500000000",
            INIT_79 => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_7B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000300000000000000000000000000000000000000000000003b00000000",
            INIT_7D => X"0000000600000000000000010000000000000010000000000000000000000000",
            INIT_7E => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_7F => X"0000005d00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE4;


    MEM_IFMAP_LAYER1_INSTANCE5 : if BRAM_NAME = "ifmap_layer1_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000000000000000000000f000000000000001c000000000000000000000000",
            INIT_03 => X"0000000000000000000000520000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000130000000000000012000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_06 => X"0000000500000000000000000000000000000017000000000000000c00000000",
            INIT_07 => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000003000000000000001d00000000",
            INIT_09 => X"0000000000000000000000110000000000000000000000000000001600000000",
            INIT_0A => X"0000000800000000000000000000000000000000000000000000001200000000",
            INIT_0B => X"0000001b00000000000000000000000000000011000000000000000000000000",
            INIT_0C => X"0000001900000000000000090000000000000000000000000000000000000000",
            INIT_0D => X"000000030000000000000000000000000000003b000000000000000000000000",
            INIT_0E => X"0000000000000000000000050000000000000000000000000000001000000000",
            INIT_0F => X"0000000000000000000000120000000000000012000000000000000000000000",
            INIT_10 => X"00000000000000000000000d0000000000000033000000000000000000000000",
            INIT_11 => X"0000002d00000000000000000000000000000000000000000000005800000000",
            INIT_12 => X"0000002800000000000000020000000000000000000000000000000400000000",
            INIT_13 => X"0000001d000000000000002c000000000000003e000000000000003300000000",
            INIT_14 => X"0000003b00000000000000000000000000000036000000000000007000000000",
            INIT_15 => X"0000004e000000000000004e000000000000002e000000000000000000000000",
            INIT_16 => X"00000056000000000000004f0000000000000049000000000000004400000000",
            INIT_17 => X"0000005a0000000000000053000000000000005a000000000000005800000000",
            INIT_18 => X"0000000000000000000000080000000000000048000000000000006f00000000",
            INIT_19 => X"0000004c000000000000004a0000000000000048000000000000004900000000",
            INIT_1A => X"00000057000000000000005b000000000000005b000000000000005400000000",
            INIT_1B => X"00000060000000000000005a000000000000005e000000000000005d00000000",
            INIT_1C => X"0000005000000000000000310000000000000000000000000000008a00000000",
            INIT_1D => X"000000570000000000000053000000000000004d000000000000004500000000",
            INIT_1E => X"0000007400000000000000610000000000000064000000000000006100000000",
            INIT_1F => X"0000006700000000000000670000000000000050000000000000005e00000000",
            INIT_20 => X"00000055000000000000005f0000000000000049000000000000004100000000",
            INIT_21 => X"0000005200000000000000520000000000000052000000000000004900000000",
            INIT_22 => X"000000450000000000000053000000000000006b000000000000005e00000000",
            INIT_23 => X"0000002e0000000000000033000000000000002e000000000000002f00000000",
            INIT_24 => X"0000002f0000000000000031000000000000002f000000000000002f00000000",
            INIT_25 => X"00000027000000000000001c0000000000000023000000000000002b00000000",
            INIT_26 => X"0000003200000000000000240000000000000027000000000000002600000000",
            INIT_27 => X"00000034000000000000002d0000000000000035000000000000003200000000",
            INIT_28 => X"0000000400000000000000250000000000000013000000000000005500000000",
            INIT_29 => X"0000002400000000000000150000000000000013000000000000002100000000",
            INIT_2A => X"0000003b000000000000001a0000000000000028000000000000002d00000000",
            INIT_2B => X"0000002c0000000000000038000000000000002e000000000000003400000000",
            INIT_2C => X"0000004f000000000000001a0000000000000000000000000000000000000000",
            INIT_2D => X"000000270000000000000004000000000000000b000000000000000a00000000",
            INIT_2E => X"0000002c00000000000000790000000000000000000000000000003900000000",
            INIT_2F => X"0000001a00000000000000230000000000000025000000000000003600000000",
            INIT_30 => X"0000000000000000000000530000000000000018000000000000000800000000",
            INIT_31 => X"00000053000000000000000e0000000000000000000000000000001200000000",
            INIT_32 => X"00000049000000000000000a0000000000000063000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000001a000000000000002c00000000",
            INIT_34 => X"00000000000000000000000b000000000000005f000000000000000800000000",
            INIT_35 => X"0000000000000000000000390000000000000000000000000000001e00000000",
            INIT_36 => X"00000049000000000000002e0000000000000000000000000000003800000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000230000000000000000000000000000000000000000000000bf00000000",
            INIT_39 => X"000000150000000000000000000000000000000d000000000000000400000000",
            INIT_3A => X"0000005000000000000000610000000000000000000000000000000c00000000",
            INIT_3B => X"000000a400000000000000000000000000000000000000000000000a00000000",
            INIT_3C => X"00000027000000000000001e0000000000000000000000000000000000000000",
            INIT_3D => X"0000000100000000000000000000000000000000000000000000000d00000000",
            INIT_3E => X"0000000000000000000000680000000000000045000000000000000000000000",
            INIT_3F => X"00000000000000000000007c0000000000000000000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000120000000000000022000000000000002a000000000000000000000000",
            INIT_41 => X"0000003c00000000000000000000000000000017000000000000000000000000",
            INIT_42 => X"0000001c00000000000000000000000000000003000000000000001100000000",
            INIT_43 => X"0000000000000000000000220000000000000006000000000000003100000000",
            INIT_44 => X"0000000a0000000000000044000000000000003a000000000000002600000000",
            INIT_45 => X"00000000000000000000004a0000000000000000000000000000001800000000",
            INIT_46 => X"00000017000000000000000e000000000000002a000000000000001900000000",
            INIT_47 => X"0000004800000000000000050000000000000000000000000000000a00000000",
            INIT_48 => X"000000110000000000000051000000000000001c000000000000005600000000",
            INIT_49 => X"0000000b000000000000000000000000000000a3000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000005600000000",
            INIT_4B => X"0000001e000000000000002d0000000000000028000000000000001400000000",
            INIT_4C => X"0000000000000000000000280000000000000040000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000009800000000",
            INIT_4E => X"0000001000000000000000090000000000000000000000000000000000000000",
            INIT_4F => X"000000000000000000000011000000000000000e000000000000001000000000",
            INIT_50 => X"0000001f00000000000000480000000000000041000000000000000300000000",
            INIT_51 => X"0000000a00000000000000050000000000000009000000000000000000000000",
            INIT_52 => X"0000001700000000000000140000000000000010000000000000000800000000",
            INIT_53 => X"0000000000000000000000170000000000000008000000000000001000000000",
            INIT_54 => X"0000000000000000000000000000000000000074000000000000001000000000",
            INIT_55 => X"0000000d00000000000000090000000000000000000000000000001100000000",
            INIT_56 => X"000000000000000000000009000000000000000d000000000000001000000000",
            INIT_57 => X"0000000d00000000000000000000000000000000000000000000002600000000",
            INIT_58 => X"0000001600000000000000000000000000000000000000000000001900000000",
            INIT_59 => X"0000001000000000000000180000000000000009000000000000000c00000000",
            INIT_5A => X"000000030000000000000031000000000000000b000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_61 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000001200000000000000040000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000270000000000000001000000000000000000000000",
            INIT_6B => X"0000000000000000000000080000000000000038000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_71 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE5;


    MEM_IFMAP_LAYER1_INSTANCE6 : if BRAM_NAME = "ifmap_layer1_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_01 => X"00000030000000000000001e0000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_03 => X"000000010000000000000024000000000000001c000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000036000000000000002f0000000000000000000000000000000000000000",
            INIT_14 => X"0000003000000000000000350000000000000035000000000000003300000000",
            INIT_15 => X"0000002b0000000000000036000000000000003b000000000000003900000000",
            INIT_16 => X"0000002800000000000000250000000000000020000000000000002000000000",
            INIT_17 => X"0000003600000000000000380000000000000030000000000000002700000000",
            INIT_18 => X"0000003b00000000000000420000000000000033000000000000003900000000",
            INIT_19 => X"0000000200000000000000020000000000000023000000000000003900000000",
            INIT_1A => X"0000002700000000000000110000000000000006000000000000000600000000",
            INIT_1B => X"0000003900000000000000360000000000000013000000000000003000000000",
            INIT_1C => X"00000000000000000000001e000000000000003d000000000000003700000000",
            INIT_1D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_1E => X"0000001500000000000000170000000000000000000000000000000100000000",
            INIT_1F => X"0000004000000000000000370000000000000032000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000001e000000000000001200000000",
            INIT_21 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_22 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000003300000000000000440000000000000010000000000000003400000000",
            INIT_24 => X"0000000000000000000000000000000000000006000000000000002500000000",
            INIT_25 => X"0000000000000000000000000000000000000009000000000000001000000000",
            INIT_26 => X"00000031000000000000000f0000000000000000000000000000000000000000",
            INIT_27 => X"0000002b000000000000000d000000000000000b000000000000003800000000",
            INIT_28 => X"0000002a0000000000000000000000000000000b000000000000000800000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000003d0000000000000007000000000000002c000000000000000000000000",
            INIT_2B => X"00000017000000000000002e0000000000000011000000000000000e00000000",
            INIT_2C => X"0000000000000000000000130000000000000003000000000000000800000000",
            INIT_2D => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000250000000000000000000000000000001900000000",
            INIT_2F => X"00000000000000000000000a000000000000002e000000000000002200000000",
            INIT_30 => X"000000000000000000000000000000000000000f000000000000001300000000",
            INIT_31 => X"0000001100000000000000150000000000000000000000000000000200000000",
            INIT_32 => X"00000000000000000000001c0000000000000000000000000000000900000000",
            INIT_33 => X"0000002c0000000000000000000000000000000c000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"00000014000000000000000e0000000000000016000000000000002100000000",
            INIT_36 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_37 => X"0000000000000000000000050000000000000006000000000000001f00000000",
            INIT_38 => X"00000028000000000000001e0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000150000000000000014000000000000000500000000",
            INIT_3A => X"0000001700000000000000110000000000000006000000000000002c00000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000003c00000000000000320000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000002c00000000000000290000000000000023000000000000002200000000",
            INIT_4D => X"0000002f000000000000002b0000000000000028000000000000002000000000",
            INIT_4E => X"0000001e000000000000001d0000000000000029000000000000003200000000",
            INIT_4F => X"000000240000000000000028000000000000002e000000000000002900000000",
            INIT_50 => X"0000000e0000000000000021000000000000002c000000000000002400000000",
            INIT_51 => X"00000005000000000000002e0000000000000030000000000000004300000000",
            INIT_52 => X"0000001500000000000000190000000000000029000000000000002100000000",
            INIT_53 => X"000000280000000000000002000000000000003f000000000000002c00000000",
            INIT_54 => X"000000280000000000000020000000000000002a000000000000002900000000",
            INIT_55 => X"0000001c00000000000000000000000000000010000000000000002400000000",
            INIT_56 => X"0000000b000000000000001a0000000000000032000000000000000c00000000",
            INIT_57 => X"00000024000000000000002e0000000000000000000000000000005c00000000",
            INIT_58 => X"000000250000000000000027000000000000000c000000000000003800000000",
            INIT_59 => X"0000001800000000000000230000000000000000000000000000001900000000",
            INIT_5A => X"0000002c00000000000000000000000000000026000000000000001a00000000",
            INIT_5B => X"0000001300000000000000000000000000000041000000000000000500000000",
            INIT_5C => X"000000250000000000000024000000000000002a000000000000002700000000",
            INIT_5D => X"0000001200000000000000380000000000000014000000000000000000000000",
            INIT_5E => X"000000000000000000000024000000000000001a000000000000002b00000000",
            INIT_5F => X"000000000000000000000000000000000000002f000000000000003700000000",
            INIT_60 => X"0000000000000000000000430000000000000025000000000000001600000000",
            INIT_61 => X"0000001d0000000000000007000000000000002a000000000000003400000000",
            INIT_62 => X"0000000e00000000000000240000000000000011000000000000002000000000",
            INIT_63 => X"0000001500000000000000000000000000000000000000000000004600000000",
            INIT_64 => X"0000002b00000000000000000000000000000039000000000000001c00000000",
            INIT_65 => X"000000250000000000000000000000000000000d000000000000002800000000",
            INIT_66 => X"0000003400000000000000290000000000000006000000000000000b00000000",
            INIT_67 => X"0000000b00000000000000350000000000000000000000000000000200000000",
            INIT_68 => X"0000002c00000000000000110000000000000000000000000000001800000000",
            INIT_69 => X"0000000d000000000000000d0000000000000011000000000000000000000000",
            INIT_6A => X"000000340000000000000000000000000000003f000000000000000000000000",
            INIT_6B => X"00000000000000000000001b000000000000000e000000000000000000000000",
            INIT_6C => X"00000000000000000000002b0000000000000005000000000000003f00000000",
            INIT_6D => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_6E => X"00000014000000000000002a0000000000000000000000000000003900000000",
            INIT_6F => X"0000000f000000000000002c000000000000001d000000000000000000000000",
            INIT_70 => X"000000100000000000000000000000000000000f000000000000002f00000000",
            INIT_71 => X"0000003800000000000000000000000000000000000000000000002f00000000",
            INIT_72 => X"0000000000000000000000320000000000000029000000000000000000000000",
            INIT_73 => X"0000000f000000000000002b0000000000000027000000000000000500000000",
            INIT_74 => X"0000002100000000000000110000000000000008000000000000000800000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000005000000000000005200000000",
            INIT_77 => X"0000000000000000000000030000000000000007000000000000000000000000",
            INIT_78 => X"0000001400000000000000030000000000000000000000000000000000000000",
            INIT_79 => X"0000002e00000000000000220000000000000000000000000000000000000000",
            INIT_7A => X"0000000500000000000000020000000000000006000000000000000000000000",
            INIT_7B => X"0000000200000000000000000000000000000000000000000000000100000000",
            INIT_7C => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000000d0000000000000022000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000006000000000000000900000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE6;


    MEM_IFMAP_LAYER1_INSTANCE7 : if BRAM_NAME = "ifmap_layer1_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000013000000000000001500000000",
            INIT_01 => X"0000000000000000000000000000000000000014000000000000000400000000",
            INIT_02 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000001a00000000000000120000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER1_INSTANCE7;


    MEM_IFMAP_LAYER2_INSTANCE0 : if BRAM_NAME = "ifmap_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000210000000000000037000000000000006c000000000000006000000000",
            INIT_0E => X"00000000000000000000004c000000000000000c000000000000003800000000",
            INIT_0F => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000000000002a000000000000000f00000000",
            INIT_11 => X"0000002b00000000000000000000000000000007000000000000001500000000",
            INIT_12 => X"0000001300000000000000110000000000000061000000000000005f00000000",
            INIT_13 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"000000000000000000000073000000000000005d000000000000000000000000",
            INIT_15 => X"0000005a00000000000000b80000000000000046000000000000004300000000",
            INIT_16 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000002300000000000000d600000000",
            INIT_18 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_19 => X"0000001f000000000000003a000000000000001c000000000000000000000000",
            INIT_1A => X"00000000000000000000000e000000000000013a000000000000002700000000",
            INIT_1B => X"00000038000000000000002400000000000000c2000000000000001d00000000",
            INIT_1C => X"000000170000000000000000000000000000006f000000000000008000000000",
            INIT_1D => X"000000000000000000000000000000000000002200000000000001cf00000000",
            INIT_1E => X"000000f200000000000000600000000000000000000000000000001600000000",
            INIT_1F => X"0000017a00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000a00000000000000000000000000000000000000000000009200000000",
            INIT_21 => X"000000ce000000000000009d0000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_23 => X"0000000c000000000000007c0000000000000000000000000000007b00000000",
            INIT_24 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000036000000000000000000000000",
            INIT_2A => X"0000000000000000000000380000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000004b0000000000000000000000000000000000000000",
            INIT_2D => X"0000009d00000000000000000000000000000077000000000000000000000000",
            INIT_2E => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_30 => X"0000002100000000000000000000000000000013000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_34 => X"0000006e00000000000000000000000000000079000000000000000000000000",
            INIT_35 => X"0000006a00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000cb0000000000000000000000000000000000000000",
            INIT_38 => X"00000039000000000000003c0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000037000000000000001b00000000",
            INIT_3A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000b600000000000000320000000000000000000000000000000000000000",
            INIT_3C => X"0000000a00000000000000000000000000000008000000000000000000000000",
            INIT_3D => X"0000000000000000000000670000000000000039000000000000000000000000",
            INIT_3E => X"0000002e00000000000000110000000000000020000000000000000c00000000",
            INIT_3F => X"000000150000000000000000000000000000002a000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000170000000000000009000000000000003600000000",
            INIT_41 => X"0000000b00000000000000090000000000000000000000000000000000000000",
            INIT_42 => X"0000001700000000000000000000000000000006000000000000001900000000",
            INIT_43 => X"000000090000000000000029000000000000000d000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"00000009000000000000000d0000000000000000000000000000001700000000",
            INIT_48 => X"0000001a00000000000000260000000000000016000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000200000000000000010000000000000000000000000000000500000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000e0000000000000000000000000000001b000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000100000000000000000000000000000002000000000000003b00000000",
            INIT_55 => X"0000000000000000000000150000000000000018000000000000000600000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000050000000000000000000000000000000b00000000",
            INIT_58 => X"0000001c00000000000000060000000000000011000000000000000000000000",
            INIT_59 => X"0000001f00000000000000000000000000000001000000000000004000000000",
            INIT_5A => X"0000002d00000000000000170000000000000005000000000000000c00000000",
            INIT_5B => X"0000000800000000000000120000000000000021000000000000000800000000",
            INIT_5C => X"0000000000000000000000300000000000000022000000000000001300000000",
            INIT_5D => X"0000000000000000000000310000000000000038000000000000000000000000",
            INIT_5E => X"000000080000000000000000000000000000001a000000000000002e00000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000004a00000000000000000000000000000000000000000000002200000000",
            INIT_63 => X"000000000000000000000032000000000000002a000000000000004a00000000",
            INIT_64 => X"00000000000000000000000a0000000000000009000000000000000900000000",
            INIT_65 => X"0000000000000000000000000000000000000032000000000000001100000000",
            INIT_66 => X"0000003e00000000000000000000000000000005000000000000000000000000",
            INIT_67 => X"00000000000000000000001f0000000000000019000000000000000400000000",
            INIT_68 => X"00000000000000000000004e0000000000000000000000000000005b00000000",
            INIT_69 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_6A => X"0000000d0000000000000000000000000000005b000000000000005d00000000",
            INIT_6B => X"00000000000000000000005f0000000000000083000000000000000000000000",
            INIT_6C => X"0000005b00000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_72 => X"00000000000000000000003c0000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000360000000000000000000000000000001700000000",
            INIT_74 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_75 => X"000000080000000000000000000000000000001f000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000000e000000000000001700000000",
            INIT_77 => X"0000003b00000000000000aa0000000000000000000000000000000000000000",
            INIT_78 => X"00000000000000000000002f0000000000000027000000000000005600000000",
            INIT_79 => X"0000004d00000000000000560000000000000087000000000000002700000000",
            INIT_7A => X"0000006100000000000000680000000000000072000000000000004c00000000",
            INIT_7B => X"00000000000000000000002d0000000000000094000000000000005100000000",
            INIT_7C => X"0000002500000000000000380000000000000000000000000000004d00000000",
            INIT_7D => X"0000000a000000000000000c0000000000000018000000000000000000000000",
            INIT_7E => X"00000000000000000000002d000000000000009b000000000000000000000000",
            INIT_7F => X"000000000000000000000000000000000000001c000000000000000e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE0;


    MEM_IFMAP_LAYER2_INSTANCE1 : if BRAM_NAME = "ifmap_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003900000000000000390000000000000074000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000001b000000000000003600000000",
            INIT_02 => X"0000001d000000000000004b0000000000000000000000000000001300000000",
            INIT_03 => X"000000920000000000000050000000000000004d000000000000000200000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_05 => X"000000000000000000000000000000000000009e000000000000002400000000",
            INIT_06 => X"0000003200000000000000150000000000000012000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000001c000000000000004b00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_0A => X"0000002c00000000000000370000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_0C => X"0000000000000000000000640000000000000000000000000000000000000000",
            INIT_0D => X"0000001300000000000000110000000000000000000000000000003f00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000002000000000000005f0000000000000000000000000000000000000000",
            INIT_10 => X"0000001400000000000000000000000000000007000000000000000000000000",
            INIT_11 => X"0000000400000000000000530000000000000004000000000000000b00000000",
            INIT_12 => X"00000017000000000000002e0000000000000032000000000000001800000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_19 => X"0000000e00000000000000000000000000000016000000000000000000000000",
            INIT_1A => X"0000000600000000000000000000000000000000000000000000001e00000000",
            INIT_1B => X"0000002100000000000000010000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"000000000000000000000000000000000000001b000000000000001200000000",
            INIT_1E => X"0000004100000000000000380000000000000039000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000007c00000000000000170000000000000000000000000000002300000000",
            INIT_27 => X"00000000000000000000001a0000000000000000000000000000000300000000",
            INIT_28 => X"000000150000000000000000000000000000001a000000000000000000000000",
            INIT_29 => X"0000000000000000000000170000000000000018000000000000000600000000",
            INIT_2A => X"00000024000000000000001e000000000000000c000000000000000000000000",
            INIT_2B => X"0000009200000000000000810000000000000040000000000000003500000000",
            INIT_2C => X"000000000000000000000019000000000000006c000000000000002700000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000003300000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000070000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_31 => X"00000038000000000000004f000000000000001c000000000000000000000000",
            INIT_32 => X"0000000000000000000000360000000000000000000000000000003800000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000650000000000000042000000000000001c000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000066000000000000002600000000",
            INIT_3C => X"000000560000000000000059000000000000004e000000000000006200000000",
            INIT_3D => X"0000004d00000000000000000000000000000019000000000000007700000000",
            INIT_3E => X"000000b700000000000000470000000000000035000000000000006000000000",
            INIT_3F => X"000000250000000000000028000000000000000c000000000000007400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007800000000000000850000000000000039000000000000001800000000",
            INIT_41 => X"00000084000000000000006e0000000000000050000000000000003900000000",
            INIT_42 => X"000000a9000000000000008b000000000000009a000000000000008a00000000",
            INIT_43 => X"000000bb00000000000000ab000000000000009c000000000000009200000000",
            INIT_44 => X"000000a6000000000000000a0000000000000000000000000000000000000000",
            INIT_45 => X"00000050000000000000006700000000000000a900000000000000b500000000",
            INIT_46 => X"00000000000000000000004d0000000000000097000000000000004600000000",
            INIT_47 => X"00000011000000000000002d000000000000001c000000000000000000000000",
            INIT_48 => X"0000002100000000000000000000000000000000000000000000001c00000000",
            INIT_49 => X"0000001d0000000000000068000000000000001d000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000002f000000000000002b0000000000000000000000000000000000000000",
            INIT_4C => X"00000040000000000000006a0000000000000034000000000000003700000000",
            INIT_4D => X"00000056000000000000006700000000000000d1000000000000002400000000",
            INIT_4E => X"0000006100000000000000170000000000000042000000000000007300000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_59 => X"0000009b00000000000000b30000000000000000000000000000006800000000",
            INIT_5A => X"000000c1000000000000007c000000000000009c000000000000007d00000000",
            INIT_5B => X"000000a9000000000000009800000000000000a0000000000000007d00000000",
            INIT_5C => X"0000001c000000000000000600000000000000b000000000000000c200000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000006200000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000500000000000000051000000000000004b000000000000006100000000",
            INIT_6A => X"0000008800000000000000610000000000000041000000000000004900000000",
            INIT_6B => X"0000005a000000000000005e000000000000005b000000000000005300000000",
            INIT_6C => X"00000060000000000000005a0000000000000068000000000000002a00000000",
            INIT_6D => X"0000003c0000000000000073000000000000005f000000000000007600000000",
            INIT_6E => X"0000007b000000000000004e000000000000006d000000000000007600000000",
            INIT_6F => X"0000005c000000000000005d0000000000000041000000000000004600000000",
            INIT_70 => X"0000004f000000000000003b0000000000000046000000000000009700000000",
            INIT_71 => X"0000002e00000000000000230000000000000015000000000000001000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_73 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000057000000000000007b0000000000000073000000000000006300000000",
            INIT_76 => X"000000450000000000000048000000000000004b000000000000005600000000",
            INIT_77 => X"0000000500000000000000400000000000000043000000000000007000000000",
            INIT_78 => X"00000032000000000000002b0000000000000044000000000000001200000000",
            INIT_79 => X"000000240000000000000000000000000000001e000000000000002200000000",
            INIT_7A => X"00000000000000000000005d0000000000000007000000000000003c00000000",
            INIT_7B => X"0000002100000000000000210000000000000000000000000000000900000000",
            INIT_7C => X"0000001500000000000000000000000000000006000000000000000000000000",
            INIT_7D => X"00000000000000000000002b0000000000000017000000000000001900000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE1;


    MEM_IFMAP_LAYER2_INSTANCE2 : if BRAM_NAME = "ifmap_layer2_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000004a000000000000005e000000000000005a000000000000000000000000",
            INIT_02 => X"0000004700000000000000310000000000000026000000000000002c00000000",
            INIT_03 => X"0000002600000000000000000000000000000036000000000000003c00000000",
            INIT_04 => X"00000050000000000000003e000000000000003a000000000000002600000000",
            INIT_05 => X"0000003100000000000000460000000000000002000000000000000e00000000",
            INIT_06 => X"00000035000000000000003f000000000000002d000000000000002e00000000",
            INIT_07 => X"000000350000000000000044000000000000005a000000000000002600000000",
            INIT_08 => X"00000000000000000000001c0000000000000044000000000000004900000000",
            INIT_09 => X"0000001d0000000000000000000000000000002c000000000000000800000000",
            INIT_0A => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_11 => X"0000001100000000000000320000000000000000000000000000000a00000000",
            INIT_12 => X"0000004c00000000000000000000000000000011000000000000000000000000",
            INIT_13 => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_14 => X"0000001c00000000000000760000000000000000000000000000000200000000",
            INIT_15 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_16 => X"0000007b0000000000000012000000000000006e000000000000000000000000",
            INIT_17 => X"0000003e0000000000000018000000000000001a000000000000008600000000",
            INIT_18 => X"00000033000000000000003d00000000000000af000000000000000000000000",
            INIT_19 => X"00000116000000000000004c0000000000000048000000000000003500000000",
            INIT_1A => X"0000007400000000000000d100000000000000be000000000000010a00000000",
            INIT_1B => X"000000f000000000000000be00000000000000c1000000000000006c00000000",
            INIT_1C => X"0000000300000000000000350000000000000015000000000000009600000000",
            INIT_1D => X"0000007b000000000000003e0000000000000055000000000000002b00000000",
            INIT_1E => X"0000001000000000000000000000000000000034000000000000001c00000000",
            INIT_1F => X"0000001100000000000000570000000000000064000000000000004000000000",
            INIT_20 => X"0000001f00000000000000400000000000000000000000000000000a00000000",
            INIT_21 => X"0000002f00000000000000270000000000000030000000000000004000000000",
            INIT_22 => X"0000000000000000000000370000000000000076000000000000001700000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000090000000000000000000000000000006c000000000000000000000000",
            INIT_28 => X"0000000000000000000000970000000000000000000000000000000000000000",
            INIT_29 => X"00000000000000000000006f0000000000000084000000000000006500000000",
            INIT_2A => X"000000b0000000000000000000000000000000ed000000000000000000000000",
            INIT_2B => X"00000000000000000000007900000000000000c4000000000000006200000000",
            INIT_2C => X"0000000000000000000000920000000000000000000000000000005300000000",
            INIT_2D => X"0000007600000000000000250000000000000000000000000000004600000000",
            INIT_2E => X"000000000000000000000000000000000000001f000000000000005300000000",
            INIT_2F => X"00000024000000000000000000000000000000a2000000000000000000000000",
            INIT_30 => X"0000001100000000000000060000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_32 => X"0000001e00000000000000000000000000000006000000000000000000000000",
            INIT_33 => X"000000240000000000000032000000000000005c000000000000001100000000",
            INIT_34 => X"00000034000000000000008a0000000000000050000000000000009e00000000",
            INIT_35 => X"000000420000000000000026000000000000002c000000000000004600000000",
            INIT_36 => X"00000097000000000000002e0000000000000059000000000000003600000000",
            INIT_37 => X"0000002a00000000000000220000000000000036000000000000002200000000",
            INIT_38 => X"0000000000000000000000270000000000000035000000000000003100000000",
            INIT_39 => X"000000a600000000000000af0000000000000017000000000000001f00000000",
            INIT_3A => X"0000002100000000000000660000000000000037000000000000002b00000000",
            INIT_3B => X"0000002800000000000000bd000000000000009a000000000000001c00000000",
            INIT_3C => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000001f000000000000000b0000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001800000000000000300000000000000000000000000000000000000000",
            INIT_46 => X"000000190000000000000020000000000000002a000000000000000500000000",
            INIT_47 => X"00000086000000000000007e0000000000000047000000000000000000000000",
            INIT_48 => X"000000b000000000000000b300000000000000a7000000000000008a00000000",
            INIT_49 => X"000000a300000000000000ae000000000000007d00000000000000d000000000",
            INIT_4A => X"0000000000000000000000e100000000000000bf00000000000000ac00000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_4C => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000004e0000000000000000000000000000002a000000000000002f00000000",
            INIT_4E => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_4F => X"00000000000000000000003a0000000000000000000000000000005300000000",
            INIT_50 => X"0000005000000000000000000000000000000005000000000000001100000000",
            INIT_51 => X"0000001c00000000000000000000000000000025000000000000000000000000",
            INIT_52 => X"000000000000000000000000000000000000008b000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_55 => X"0000001200000000000000000000000000000000000000000000000400000000",
            INIT_56 => X"0000000a0000000000000024000000000000000d000000000000001800000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000005000000000000000040000000000000000000000000000004d00000000",
            INIT_59 => X"0000003300000000000000000000000000000000000000000000001200000000",
            INIT_5A => X"0000003f0000000000000000000000000000001e000000000000000000000000",
            INIT_5B => X"0000000000000000000000910000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000250000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"00000000000000000000000a0000000000000044000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000077000000000000000000000000",
            INIT_60 => X"0000006700000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000a60000000000000005000000000000004200000000",
            INIT_62 => X"0000003800000000000000410000000000000030000000000000006100000000",
            INIT_63 => X"0000000000000000000000030000000000000000000000000000000b00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"00000023000000000000004e0000000000000029000000000000000000000000",
            INIT_66 => X"0000002300000000000000000000000000000022000000000000000000000000",
            INIT_67 => X"00000000000000000000006f000000000000002d000000000000000000000000",
            INIT_68 => X"00000000000000000000005c000000000000002e000000000000000500000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000002e0000000000000003000000000000002b000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000000000000000000053000000000000005e000000000000005e00000000",
            INIT_6E => X"0000003600000000000000300000000000000000000000000000000000000000",
            INIT_6F => X"000000b000000000000000900000000000000039000000000000003000000000",
            INIT_70 => X"0000004a0000000000000067000000000000006700000000000000a200000000",
            INIT_71 => X"0000007900000000000000b4000000000000006a000000000000006800000000",
            INIT_72 => X"000000430000000000000014000000000000003b000000000000002500000000",
            INIT_73 => X"000000000000000000000042000000000000006a000000000000003400000000",
            INIT_74 => X"0000000000000000000000240000000000000000000000000000003400000000",
            INIT_75 => X"000000270000000000000000000000000000002c000000000000002200000000",
            INIT_76 => X"000000330000000000000000000000000000003c000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000008000000000000001700000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_7E => X"0000000a00000000000000160000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000001000000000000002d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE2;


    MEM_IFMAP_LAYER2_INSTANCE3 : if BRAM_NAME = "ifmap_layer2_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002f00000000000000120000000000000017000000000000000300000000",
            INIT_01 => X"000000080000000000000000000000000000001e000000000000004500000000",
            INIT_02 => X"0000006000000000000000000000000000000002000000000000001500000000",
            INIT_03 => X"0000003a00000000000000270000000000000039000000000000004200000000",
            INIT_04 => X"0000000700000000000000690000000000000026000000000000003a00000000",
            INIT_05 => X"00000088000000000000007e000000000000007e000000000000004800000000",
            INIT_06 => X"00000092000000000000006600000000000000bb000000000000009600000000",
            INIT_07 => X"000000ab00000000000000a9000000000000009e000000000000009600000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER2_INSTANCE3;


    MEM_IFMAP_LAYER3_INSTANCE0 : if BRAM_NAME = "ifmap_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000001040000000000000040000000000000001200000000000000a000000000",
            INIT_01 => X"00000000000000000000010100000000000000bc000000000000005100000000",
            INIT_02 => X"0000001c00000000000000000000000000000047000000000000000000000000",
            INIT_03 => X"0000000000000000000000ba0000000000000000000000000000000000000000",
            INIT_04 => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000920000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000200000000000000000000000000000000000000000000010400000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000038000000000000000000000000000000a8000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000370000000000000053000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000134000000000000017a00000000000000a8000000000000000000000000",
            INIT_15 => X"000000b700000000000000820000000000000113000000000000003700000000",
            INIT_16 => X"0000002d00000000000000000000000000000000000000000000003500000000",
            INIT_17 => X"00000062000000000000014d0000000000000000000000000000007900000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000350000000000000010000000000000007e000000000000000000000000",
            INIT_1A => X"000000d10000000000000000000000000000006a000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000a0000000000000000000000000000000b000000000000000b000000000",
            INIT_1D => X"0000008100000000000000d20000000000000077000000000000003300000000",
            INIT_1E => X"000000080000000000000000000000000000000000000000000000c600000000",
            INIT_1F => X"000000650000000000000000000000000000005700000000000000a900000000",
            INIT_20 => X"0000003c00000000000000a1000000000000000000000000000000c800000000",
            INIT_21 => X"00000000000000000000007a0000000000000058000000000000000000000000",
            INIT_22 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000005c00000000",
            INIT_24 => X"0000000000000000000000e6000000000000002c000000000000000000000000",
            INIT_25 => X"000000ff00000000000000000000000000000048000000000000007700000000",
            INIT_26 => X"0000001900000000000000000000000000000000000000000000002400000000",
            INIT_27 => X"0000000000000000000000000000000000000036000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000004d000000000000005d0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000aa000000000000006c00000000000000b500000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000030000000000000001b0000000000000000000000000000003f00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_31 => X"00000012000000000000000000000000000000b3000000000000011900000000",
            INIT_32 => X"000000bd000000000000000000000000000000aa000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000002600000000000000b600000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"00000144000000000000012400000000000000c0000000000000000000000000",
            INIT_39 => X"00000017000000000000006800000000000000d0000000000000014f00000000",
            INIT_3A => X"0000000000000000000000000000000000000040000000000000000000000000",
            INIT_3B => X"0000000000000000000000160000000000000057000000000000000900000000",
            INIT_3C => X"000000000000000000000000000000000000005d00000000000000cf00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000b8000000000000000100000000000000a8000000000000000000000000",
            INIT_42 => X"0000009000000000000000960000000000000028000000000000001e00000000",
            INIT_43 => X"0000000000000000000000000000000000000063000000000000001500000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000009e000000000000011b0000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000006c0000000000000000000000000000000000000000",
            INIT_49 => X"0000007900000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000ff0000000000000004000000000000004300000000000000f800000000",
            INIT_4B => X"0000000000000000000000110000000000000012000000000000006700000000",
            INIT_4C => X"000000690000000000000000000000000000001c000000000000000000000000",
            INIT_4D => X"0000004e00000000000000860000000000000000000000000000004100000000",
            INIT_4E => X"0000009100000000000000000000000000000000000000000000003100000000",
            INIT_4F => X"0000002600000000000000170000000000000051000000000000006c00000000",
            INIT_50 => X"000000fd00000000000000b00000000000000000000000000000004600000000",
            INIT_51 => X"000000000000000000000078000000000000000000000000000000e000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_53 => X"000000ab00000000000000590000000000000000000000000000000000000000",
            INIT_54 => X"0000006a00000000000000ef00000000000000fb00000000000000c100000000",
            INIT_55 => X"00000053000000000000003b00000000000000db000000000000008f00000000",
            INIT_56 => X"0000000000000000000000000000000000000010000000000000001400000000",
            INIT_57 => X"0000006200000000000000ab0000000000000046000000000000007b00000000",
            INIT_58 => X"0000006d00000000000000a2000000000000013c000000000000005a00000000",
            INIT_59 => X"000000510000000000000123000000000000007a000000000000008c00000000",
            INIT_5A => X"00000000000000000000000000000000000000a1000000000000009700000000",
            INIT_5B => X"00000000000000000000003c0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_5D => X"0000010400000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000012f00000000000000a2000000000000004f000000000000001e00000000",
            INIT_60 => X"0000015b00000000000000000000000000000000000000000000008c00000000",
            INIT_61 => X"000000a100000000000000830000000000000161000000000000013a00000000",
            INIT_62 => X"0000000000000000000000120000000000000138000000000000007200000000",
            INIT_63 => X"000000dc00000000000000700000000000000088000000000000000000000000",
            INIT_64 => X"000000cd000000000000013e00000000000000ad00000000000000e000000000",
            INIT_65 => X"000000000000000000000000000000000000000000000000000000ae00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000001f00000000000000c80000000000000000000000000000000000000000",
            INIT_68 => X"0000004e000000000000004b000000000000004600000000000000bf00000000",
            INIT_69 => X"0000001e00000000000000000000000000000026000000000000001b00000000",
            INIT_6A => X"00000036000000000000009f000000000000013b000000000000007300000000",
            INIT_6B => X"000000a500000000000000aa0000000000000006000000000000001e00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000010100000000000000760000000000000043000000000000006a00000000",
            INIT_76 => X"000000000000000000000000000000000000007c000000000000006600000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000005900000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000310000000000000000000000000000006900000000",
            INIT_7B => X"0000003d00000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000003100000000000000100000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000000000000000000000ed000000000000007200000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000012c00000000000000700000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER3_INSTANCE0;


    MEM_IFMAP_LAYER3_INSTANCE1 : if BRAM_NAME = "ifmap_layer3_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000000000000d0000000000000017f00000000",
            INIT_01 => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_02 => X"0000002100000000000000390000000000000008000000000000006700000000",
            INIT_03 => X"000000760000000000000044000000000000006d00000000000000de00000000",
            INIT_04 => X"0000000000000000000000eb0000000000000141000000000000008400000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000003f000000000000006e000000000000007800000000000000b200000000",
            INIT_08 => X"0000000000000000000000000000000000000092000000000000007f00000000",
            INIT_09 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000034000000000000001e0000000000000000000000000000019100000000",
            INIT_0B => X"0000000000000000000000000000000000000148000000000000008700000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000004a00000000000000580000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_0F => X"000000c500000000000000d700000000000000f3000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER3_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE0 : if BRAM_NAME = "gold_layer0_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000014000000000000000f0000000000000012000000000000001200000000",
            INIT_01 => X"0000001d000000000000000f000000000000000d000000000000001700000000",
            INIT_02 => X"000000010000000000000000000000000000000a000000000000001d00000000",
            INIT_03 => X"000000160000000000000015000000000000000c000000000000000600000000",
            INIT_04 => X"000000130000000000000013000000000000000f000000000000001200000000",
            INIT_05 => X"0000000000000000000000030000000000000008000000000000000400000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_07 => X"0000000b0000000000000000000000000000000b000000000000000500000000",
            INIT_08 => X"0000001b0000000000000012000000000000001b000000000000001300000000",
            INIT_09 => X"000000000000000000000000000000000000001e000000000000002000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000c00000000000000000000000000000001000000000000000100000000",
            INIT_0C => X"000000000000000000000011000000000000000b000000000000001900000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000300000000000000030000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000001c000000000000000400000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_20 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000007000000000000000400000000",
            INIT_5A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000a000000000000003f000000000000000f000000000000001a00000000",
            INIT_62 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000002000000000000000250000000000000038000000000000003a00000000",
            INIT_64 => X"0000002700000000000000250000000000000029000000000000002200000000",
            INIT_65 => X"00000000000000000000003a000000000000002c000000000000002000000000",
            INIT_66 => X"0000001d000000000000001d000000000000001e000000000000000000000000",
            INIT_67 => X"00000024000000000000001f0000000000000020000000000000002000000000",
            INIT_68 => X"0000002100000000000000280000000000000022000000000000001e00000000",
            INIT_69 => X"0000000e000000000000002f000000000000002f000000000000003000000000",
            INIT_6A => X"0000001d00000000000000190000000000000021000000000000000f00000000",
            INIT_6B => X"00000033000000000000002f0000000000000023000000000000002200000000",
            INIT_6C => X"00000029000000000000003a0000000000000028000000000000003400000000",
            INIT_6D => X"0000002a00000000000000410000000000000031000000000000003300000000",
            INIT_6E => X"00000017000000000000001f000000000000002a000000000000003000000000",
            INIT_6F => X"0000001a000000000000002d0000000000000021000000000000001c00000000",
            INIT_70 => X"0000000000000000000000000000000000000029000000000000001c00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000006000000000000000e0000000000000018000000000000000300000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_7D => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_7E => X"0000000000000000000000060000000000000000000000000000001b00000000",
            INIT_7F => X"0000001e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE0;


    MEM_GOLD_LAYER0_INSTANCE1 : if BRAM_NAME = "gold_layer0_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001400000000000000110000000000000000000000000000000000000000",
            INIT_01 => X"0000001d00000000000000000000000000000003000000000000000500000000",
            INIT_02 => X"0000000000000000000000080000000000000000000000000000001000000000",
            INIT_03 => X"000000000000000000000017000000000000000f000000000000000300000000",
            INIT_04 => X"00000006000000000000000a000000000000001a000000000000000000000000",
            INIT_05 => X"0000000300000000000000440000000000000000000000000000000400000000",
            INIT_06 => X"000000020000000000000000000000000000000b000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000000b000000000000001700000000",
            INIT_08 => X"00000000000000000000000b000000000000001e000000000000000c00000000",
            INIT_09 => X"0000000400000000000000000000000000000037000000000000000000000000",
            INIT_0A => X"0000002000000000000000020000000000000011000000000000000a00000000",
            INIT_0B => X"0000000600000000000000000000000000000006000000000000001400000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_0D => X"0000001100000000000000000000000000000000000000000000002000000000",
            INIT_0E => X"00000028000000000000001d0000000000000000000000000000000800000000",
            INIT_0F => X"0000000000000000000000080000000000000011000000000000000400000000",
            INIT_10 => X"00000000000000000000000b000000000000000b000000000000000000000000",
            INIT_11 => X"0000000000000000000000060000000000000000000000000000001000000000",
            INIT_12 => X"0000000000000000000000240000000000000018000000000000000000000000",
            INIT_13 => X"000000120000000000000009000000000000000e000000000000002700000000",
            INIT_14 => X"0000000000000000000000000000000000000015000000000000001200000000",
            INIT_15 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_16 => X"0000005800000000000000000000000000000023000000000000002b00000000",
            INIT_17 => X"00000011000000000000002d0000000000000028000000000000000d00000000",
            INIT_18 => X"00000022000000000000001b0000000000000000000000000000000000000000",
            INIT_19 => X"000000360000000000000000000000000000000b000000000000001f00000000",
            INIT_1A => X"0000000000000000000000450000000000000012000000000000002300000000",
            INIT_1B => X"0000001a0000000000000021000000000000001f000000000000000700000000",
            INIT_1C => X"0000002e00000000000000280000000000000022000000000000001e00000000",
            INIT_1D => X"00000038000000000000002a000000000000002f000000000000002f00000000",
            INIT_1E => X"0000002700000000000000000000000000000025000000000000003300000000",
            INIT_1F => X"0000002a00000000000000240000000000000024000000000000002500000000",
            INIT_20 => X"0000002e000000000000002f0000000000000036000000000000002f00000000",
            INIT_21 => X"00000052000000000000002e000000000000002c000000000000003a00000000",
            INIT_22 => X"00000026000000000000002b0000000000000013000000000000000000000000",
            INIT_23 => X"0000002e000000000000002f000000000000002a000000000000002a00000000",
            INIT_24 => X"000000280000000000000045000000000000002a000000000000002f00000000",
            INIT_25 => X"00000019000000000000002c0000000000000033000000000000002b00000000",
            INIT_26 => X"0000002400000000000000230000000000000028000000000000001900000000",
            INIT_27 => X"0000002e000000000000002d0000000000000031000000000000002e00000000",
            INIT_28 => X"00000000000000000000001f000000000000003a000000000000004300000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000000000000000000000a000000000000000200000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000170000000000000008000000000000001000000000",
            INIT_2F => X"000000000000000000000003000000000000001c000000000000001f00000000",
            INIT_30 => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_31 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000004200000000000000000000000000000000000000000000001100000000",
            INIT_33 => X"000000000000000000000000000000000000003f000000000000002d00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_35 => X"0000002c00000000000000280000000000000000000000000000000e00000000",
            INIT_36 => X"00000026000000000000005a0000000000000000000000000000002500000000",
            INIT_37 => X"0000006c0000000000000000000000000000002a000000000000003b00000000",
            INIT_38 => X"0000003400000000000000000000000000000023000000000000000500000000",
            INIT_39 => X"0000003c0000000000000048000000000000005d000000000000002400000000",
            INIT_3A => X"0000001e0000000000000052000000000000002f000000000000000000000000",
            INIT_3B => X"0000003100000000000000590000000000000000000000000000003e00000000",
            INIT_3C => X"0000002c00000000000000000000000000000000000000000000003700000000",
            INIT_3D => X"000000000000000000000060000000000000003e000000000000006100000000",
            INIT_3E => X"000000310000000000000012000000000000005c000000000000007300000000",
            INIT_3F => X"0000001500000000000000730000000000000048000000000000002500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005a00000000000000000000000000000000000000000000003800000000",
            INIT_41 => X"000000750000000000000000000000000000006a000000000000004a00000000",
            INIT_42 => X"00000037000000000000000c0000000000000012000000000000004700000000",
            INIT_43 => X"0000003100000000000000280000000000000065000000000000004d00000000",
            INIT_44 => X"00000038000000000000008b0000000000000006000000000000000000000000",
            INIT_45 => X"00000050000000000000004f0000000000000000000000000000004600000000",
            INIT_46 => X"0000006800000000000000130000000000000025000000000000000600000000",
            INIT_47 => X"0000002a000000000000000b0000000000000084000000000000004200000000",
            INIT_48 => X"00000000000000000000002c000000000000002e000000000000001300000000",
            INIT_49 => X"00000004000000000000005b0000000000000016000000000000002900000000",
            INIT_4A => X"0000003a000000000000004a0000000000000000000000000000000000000000",
            INIT_4B => X"0000001800000000000000640000000000000000000000000000009f00000000",
            INIT_4C => X"0000003b0000000000000030000000000000004d000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000017000000000000005a00000000",
            INIT_4E => X"00000094000000000000003c000000000000000f000000000000000c00000000",
            INIT_4F => X"00000020000000000000004c0000000000000093000000000000000000000000",
            INIT_50 => X"0000001a00000000000000410000000000000083000000000000007100000000",
            INIT_51 => X"0000003100000000000000200000000000000023000000000000001d00000000",
            INIT_52 => X"00000000000000000000004e000000000000002b000000000000001d00000000",
            INIT_53 => X"0000003c000000000000003a000000000000007300000000000000d800000000",
            INIT_54 => X"0000003c000000000000003d0000000000000038000000000000004700000000",
            INIT_55 => X"0000005f000000000000004f0000000000000040000000000000003e00000000",
            INIT_56 => X"000000af00000000000000820000000000000000000000000000001200000000",
            INIT_57 => X"0000003e000000000000003f0000000000000049000000000000004200000000",
            INIT_58 => X"0000005000000000000000400000000000000038000000000000003900000000",
            INIT_59 => X"00000045000000000000006a000000000000003d000000000000004800000000",
            INIT_5A => X"00000039000000000000005a00000000000000cb000000000000000000000000",
            INIT_5B => X"00000041000000000000003c0000000000000042000000000000004d00000000",
            INIT_5C => X"00000038000000000000004e000000000000004d000000000000004800000000",
            INIT_5D => X"0000003e000000000000004b0000000000000076000000000000007b00000000",
            INIT_5E => X"0000004300000000000000350000000000000048000000000000005400000000",
            INIT_5F => X"0000005500000000000000440000000000000038000000000000004400000000",
            INIT_60 => X"00000080000000000000006f000000000000001a000000000000003a00000000",
            INIT_61 => X"0000000800000000000000080000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000050000000000000003000000000000000600000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_64 => X"0000000700000000000000050000000000000006000000000000000000000000",
            INIT_65 => X"0000000a0000000000000007000000000000000c000000000000000a00000000",
            INIT_66 => X"000000000000000000000000000000000000001a000000000000004900000000",
            INIT_67 => X"0000000000000000000000060000000000000024000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_69 => X"0000000000000000000000070000000000000004000000000000000400000000",
            INIT_6A => X"0000001a000000000000000d0000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000170000000000000007000000000000001500000000",
            INIT_6C => X"0000000900000000000000250000000000000028000000000000000000000000",
            INIT_6D => X"000000370000000000000000000000000000000d000000000000000500000000",
            INIT_6E => X"0000000000000000000000000000000000000005000000000000001b00000000",
            INIT_6F => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_70 => X"0000000b0000000000000013000000000000005a000000000000002600000000",
            INIT_71 => X"0000000e00000000000000060000000000000056000000000000008000000000",
            INIT_72 => X"0000002500000000000000250000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000018000000000000000f00000000",
            INIT_74 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_75 => X"0000001f000000000000001a000000000000002a000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_77 => X"0000000700000000000000060000000000000027000000000000000900000000",
            INIT_78 => X"0000002100000000000000000000000000000004000000000000000000000000",
            INIT_79 => X"000000110000000000000009000000000000000a000000000000000000000000",
            INIT_7A => X"000000170000000000000000000000000000000b000000000000000000000000",
            INIT_7B => X"0000001c00000000000000070000000000000015000000000000001d00000000",
            INIT_7C => X"0000000000000000000000160000000000000019000000000000001000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000004000000000000000b0000000000000004000000000000001000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE1;


    MEM_GOLD_LAYER0_INSTANCE2 : if BRAM_NAME = "gold_layer0_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001a00000000000000000000000000000000000000000000001c00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_02 => X"00000000000000000000002f0000000000000003000000000000000000000000",
            INIT_03 => X"0000001100000000000000040000000000000009000000000000000000000000",
            INIT_04 => X"0000000c000000000000004a0000000000000000000000000000000000000000",
            INIT_05 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_07 => X"00000085000000000000009c0000000000000046000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_09 => X"00000000000000000000001b0000000000000041000000000000002000000000",
            INIT_0A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000001200000000000000070000000000000004000000000000000000000000",
            INIT_11 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000001300000000000000140000000000000000000000000000000000000000",
            INIT_18 => X"0000002200000000000000280000000000000000000000000000000400000000",
            INIT_19 => X"000000a200000000000000a3000000000000009d000000000000000000000000",
            INIT_1A => X"000000ac000000000000009d00000000000000a400000000000000a500000000",
            INIT_1B => X"0000007c000000000000009400000000000000ad00000000000000b700000000",
            INIT_1C => X"0000009200000000000000920000000000000084000000000000007c00000000",
            INIT_1D => X"000000ac00000000000000a800000000000000ad00000000000000a200000000",
            INIT_1E => X"000000a000000000000000a9000000000000008c00000000000000a000000000",
            INIT_1F => X"0000003e000000000000002e000000000000003a000000000000007a00000000",
            INIT_20 => X"00000089000000000000008b000000000000006e000000000000004e00000000",
            INIT_21 => X"000000af00000000000000b000000000000000ac000000000000006a00000000",
            INIT_22 => X"0000002d00000000000000480000000000000073000000000000008e00000000",
            INIT_23 => X"00000027000000000000000a000000000000001e000000000000000700000000",
            INIT_24 => X"0000002b000000000000004d0000000000000067000000000000003a00000000",
            INIT_25 => X"0000005900000000000000a200000000000000aa00000000000000a400000000",
            INIT_26 => X"0000000c00000000000000150000000000000027000000000000004d00000000",
            INIT_27 => X"00000025000000000000001b000000000000002d000000000000003300000000",
            INIT_28 => X"00000094000000000000001f0000000000000017000000000000003a00000000",
            INIT_29 => X"000000430000000000000047000000000000004e000000000000006000000000",
            INIT_2A => X"000000310000000000000000000000000000001f000000000000002f00000000",
            INIT_2B => X"0000002f000000000000001c0000000000000017000000000000003900000000",
            INIT_2C => X"00000099000000000000008e0000000000000012000000000000001600000000",
            INIT_2D => X"000000310000000000000045000000000000003b000000000000002500000000",
            INIT_2E => X"0000002a000000000000003e0000000000000000000000000000002d00000000",
            INIT_2F => X"0000000e00000000000000170000000000000012000000000000001000000000",
            INIT_30 => X"0000002f000000000000009f0000000000000062000000000000002a00000000",
            INIT_31 => X"0000002f000000000000002d000000000000003e000000000000003200000000",
            INIT_32 => X"0000001000000000000000280000000000000032000000000000000000000000",
            INIT_33 => X"0000000a000000000000001c0000000000000026000000000000000e00000000",
            INIT_34 => X"0000002600000000000000370000000000000062000000000000002c00000000",
            INIT_35 => X"0000001e00000000000000290000000000000027000000000000002e00000000",
            INIT_36 => X"000000220000000000000009000000000000002d000000000000002f00000000",
            INIT_37 => X"0000002b00000000000000000000000000000014000000000000004100000000",
            INIT_38 => X"0000003600000000000000220000000000000055000000000000000e00000000",
            INIT_39 => X"000000420000000000000054000000000000000d000000000000003000000000",
            INIT_3A => X"00000079000000000000002d000000000000000f000000000000002600000000",
            INIT_3B => X"0000000000000000000000240000000000000005000000000000001000000000",
            INIT_3C => X"0000002800000000000000080000000000000020000000000000003500000000",
            INIT_3D => X"00000006000000000000001d0000000000000034000000000000002d00000000",
            INIT_3E => X"00000000000000000000008a0000000000000062000000000000000900000000",
            INIT_3F => X"0000001700000000000000000000000000000023000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000600000000000000000000000000000000000000000000001a00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"00000000000000000000003a0000000000000006000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000002300000000000000220000000000000000000000000000000000000000",
            INIT_52 => X"00000027000000000000001e0000000000000020000000000000002500000000",
            INIT_53 => X"00000017000000000000001d0000000000000024000000000000002600000000",
            INIT_54 => X"0000001e00000000000000240000000000000026000000000000001a00000000",
            INIT_55 => X"0000002a000000000000002c0000000000000023000000000000001800000000",
            INIT_56 => X"0000000f00000000000000200000000000000028000000000000001f00000000",
            INIT_57 => X"00000000000000000000001d000000000000000e000000000000001d00000000",
            INIT_58 => X"0000001c000000000000002b0000000000000020000000000000000900000000",
            INIT_59 => X"0000002100000000000000280000000000000039000000000000000600000000",
            INIT_5A => X"000000060000000000000000000000000000001a000000000000002700000000",
            INIT_5B => X"000000000000000000000000000000000000002e000000000000002100000000",
            INIT_5C => X"00000000000000000000002c0000000000000025000000000000000000000000",
            INIT_5D => X"0000000f00000000000000290000000000000021000000000000004c00000000",
            INIT_5E => X"0000000000000000000000000000000000000004000000000000002400000000",
            INIT_5F => X"0000000000000000000000090000000000000000000000000000004800000000",
            INIT_60 => X"000000260000000000000000000000000000004a000000000000000000000000",
            INIT_61 => X"0000000b00000000000000090000000000000056000000000000000200000000",
            INIT_62 => X"0000005900000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_64 => X"00000000000000000000000a0000000000000000000000000000002b00000000",
            INIT_65 => X"000000000000000000000013000000000000003e000000000000001a00000000",
            INIT_66 => X"00000000000000000000008e0000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_68 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000036000000000000003f00000000",
            INIT_6A => X"0000000000000000000000000000000000000066000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000015000000000000000a00000000",
            INIT_6C => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_6E => X"0000001d00000000000000000000000000000000000000000000004200000000",
            INIT_6F => X"0000000200000000000000000000000000000008000000000000000f00000000",
            INIT_70 => X"0000001100000000000000040000000000000021000000000000000000000000",
            INIT_71 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_72 => X"00000021000000000000001e0000000000000000000000000000002500000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_74 => X"00000027000000000000000f0000000000000000000000000000002c00000000",
            INIT_75 => X"0000000000000000000000050000000000000002000000000000000000000000",
            INIT_76 => X"0000001400000000000000340000000000000030000000000000000c00000000",
            INIT_77 => X"0000007800000000000000000000000000000004000000000000002a00000000",
            INIT_78 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_79 => X"0000000900000000000000080000000000000000000000000000000000000000",
            INIT_7A => X"0000002000000000000000000000000000000000000000000000000100000000",
            INIT_7B => X"0000000000000000000000400000000000000000000000000000001400000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE2;


    MEM_GOLD_LAYER0_INSTANCE3 : if BRAM_NAME = "gold_layer0_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000005d00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000002b00000000000000000000000000000000000000000000000400000000",
            INIT_0A => X"0000002f000000000000002c000000000000002d000000000000003000000000",
            INIT_0B => X"00000037000000000000003a0000000000000030000000000000002900000000",
            INIT_0C => X"0000002700000000000000260000000000000025000000000000002a00000000",
            INIT_0D => X"00000035000000000000002c0000000000000031000000000000002a00000000",
            INIT_0E => X"00000000000000000000002d000000000000002e000000000000003000000000",
            INIT_0F => X"0000000c000000000000003b0000000000000029000000000000001f00000000",
            INIT_10 => X"0000001f000000000000000e0000000000000000000000000000000000000000",
            INIT_11 => X"0000002e0000000000000029000000000000001c000000000000002500000000",
            INIT_12 => X"0000002d000000000000003b0000000000000032000000000000003500000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_14 => X"0000001a00000000000000040000000000000000000000000000000000000000",
            INIT_15 => X"0000003200000000000000230000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000019000000000000002500000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000110000000000000000000000000000000600000000",
            INIT_19 => X"0000000000000000000000180000000000000012000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_1D => X"0000000300000000000000030000000000000038000000000000000b00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000007000000000000003a00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000005000000000000001a00000000",
            INIT_2A => X"0000000400000000000000180000000000000003000000000000000f00000000",
            INIT_2B => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000000000a000000000000001100000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000800000000000000080000000000000011000000000000000a00000000",
            INIT_43 => X"0000000b000000000000000c000000000000000c000000000000000400000000",
            INIT_44 => X"00000023000000000000002d0000000000000021000000000000000b00000000",
            INIT_45 => X"0000000000000000000000060000000000000008000000000000001100000000",
            INIT_46 => X"00000008000000000000000c000000000000000a000000000000000a00000000",
            INIT_47 => X"0000004200000000000000230000000000000005000000000000000000000000",
            INIT_48 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"000000330000000000000035000000000000000a000000000000001700000000",
            INIT_4A => X"0000003700000000000000050000000000000008000000000000000500000000",
            INIT_4B => X"0000000000000000000000000000000000000009000000000000001600000000",
            INIT_4C => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000500000000000000000000000000000000000000000000000c00000000",
            INIT_4E => X"0000000000000000000000000000000000000008000000000000000800000000",
            INIT_4F => X"00000004000000000000001a0000000000000000000000000000000200000000",
            INIT_50 => X"0000000e00000000000000000000000000000006000000000000001000000000",
            INIT_51 => X"0000000e00000000000000020000000000000000000000000000000100000000",
            INIT_52 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_54 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000003e00000000000000030000000000000006000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_57 => X"0000000700000000000000150000000000000014000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000120000000000000018000000000000001c00000000",
            INIT_5A => X"0000000000000000000000110000000000000000000000000000003100000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000003500000000000000350000000000000002000000000000000000000000",
            INIT_5E => X"000000090000000000000000000000000000000e000000000000002100000000",
            INIT_5F => X"00000000000000000000000e0000000000000005000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000026000000000000000000000000",
            INIT_62 => X"0000003000000000000000260000000000000000000000000000000000000000",
            INIT_63 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000002300000000000000000000000000000004000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_66 => X"0000000000000000000000110000000000000036000000000000004e00000000",
            INIT_67 => X"0000000000000000000000030000000000000018000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_69 => X"0000000000000000000000370000000000000051000000000000001e00000000",
            INIT_6A => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000c00000000000000210000000000000035000000000000000a00000000",
            INIT_6C => X"0000000400000000000000280000000000000056000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000003000000000000000500000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001800000000000000000000000000000016000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000b000000000000004f0000000000000018000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_77 => X"0000000300000000000000000000000000000022000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000a0000000000000013000000000000000d000000000000000000000000",
            INIT_7B => X"0000000800000000000000150000000000000009000000000000000e00000000",
            INIT_7C => X"00000022000000000000001c000000000000000c000000000000000600000000",
            INIT_7D => X"0000000200000000000000060000000000000013000000000000001b00000000",
            INIT_7E => X"0000000d0000000000000009000000000000000b000000000000000800000000",
            INIT_7F => X"0000001a000000000000000f0000000000000036000000000000000f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE3;


    MEM_GOLD_LAYER0_INSTANCE4 : if BRAM_NAME = "gold_layer0_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002400000000000000350000000000000034000000000000001f00000000",
            INIT_01 => X"00000026000000000000000a000000000000001a000000000000002100000000",
            INIT_02 => X"00000008000000000000000a000000000000000b000000000000002400000000",
            INIT_03 => X"0000002000000000000000280000000000000033000000000000005100000000",
            INIT_04 => X"0000002b000000000000004b000000000000005e000000000000005300000000",
            INIT_05 => X"000000140000000000000033000000000000001a000000000000001900000000",
            INIT_06 => X"0000002e00000000000000190000000000000012000000000000000e00000000",
            INIT_07 => X"0000005b0000000000000036000000000000002f000000000000004500000000",
            INIT_08 => X"00000015000000000000003b0000000000000042000000000000005d00000000",
            INIT_09 => X"00000015000000000000005e0000000000000071000000000000001b00000000",
            INIT_0A => X"000000640000000000000044000000000000007e000000000000003500000000",
            INIT_0B => X"00000067000000000000003b0000000000000033000000000000003b00000000",
            INIT_0C => X"0000000100000000000000250000000000000039000000000000003800000000",
            INIT_0D => X"000000130000000000000028000000000000009e000000000000007f00000000",
            INIT_0E => X"0000004b000000000000007d000000000000007e00000000000000bd00000000",
            INIT_0F => X"00000050000000000000007f000000000000005b000000000000002e00000000",
            INIT_10 => X"0000007a0000000000000015000000000000003c000000000000004700000000",
            INIT_11 => X"0000005a00000000000000170000000000000043000000000000009400000000",
            INIT_12 => X"0000004e000000000000006500000000000000a8000000000000007500000000",
            INIT_13 => X"0000003b00000000000000460000000000000081000000000000007800000000",
            INIT_14 => X"000000a5000000000000008e0000000000000033000000000000004c00000000",
            INIT_15 => X"000000a500000000000000390000000000000039000000000000004000000000",
            INIT_16 => X"0000005f0000000000000050000000000000006a000000000000008500000000",
            INIT_17 => X"0000004b0000000000000048000000000000004c000000000000007800000000",
            INIT_18 => X"0000006600000000000000b800000000000000b0000000000000002600000000",
            INIT_19 => X"0000005900000000000000660000000000000038000000000000007300000000",
            INIT_1A => X"0000006500000000000000330000000000000051000000000000004e00000000",
            INIT_1B => X"0000000e000000000000002b000000000000002c000000000000004100000000",
            INIT_1C => X"00000075000000000000008600000000000000b300000000000000c000000000",
            INIT_1D => X"00000079000000000000005f0000000000000033000000000000006f00000000",
            INIT_1E => X"000000250000000000000040000000000000005a000000000000004200000000",
            INIT_1F => X"000000c700000000000000270000000000000027000000000000002f00000000",
            INIT_20 => X"0000009e00000000000000a2000000000000008b00000000000000ab00000000",
            INIT_21 => X"0000007900000000000000b90000000000000091000000000000006500000000",
            INIT_22 => X"0000005a00000000000000470000000000000040000000000000003c00000000",
            INIT_23 => X"000000cb00000000000000c10000000000000068000000000000007100000000",
            INIT_24 => X"000000a500000000000000e700000000000000c9000000000000009d00000000",
            INIT_25 => X"0000006f000000000000007c0000000000000085000000000000008a00000000",
            INIT_26 => X"0000008a00000000000000880000000000000080000000000000007800000000",
            INIT_27 => X"000000b100000000000000a1000000000000008c000000000000008e00000000",
            INIT_28 => X"00000075000000000000007a00000000000000af00000000000000e500000000",
            INIT_29 => X"0000008400000000000000760000000000000071000000000000007000000000",
            INIT_2A => X"000000a3000000000000009a0000000000000095000000000000008c00000000",
            INIT_2B => X"000000ef00000000000000a60000000000000085000000000000009d00000000",
            INIT_2C => X"0000007300000000000000790000000000000080000000000000008800000000",
            INIT_2D => X"0000009b000000000000008c0000000000000082000000000000007700000000",
            INIT_2E => X"0000009700000000000000ab00000000000000a3000000000000009300000000",
            INIT_2F => X"0000007400000000000000a7000000000000007f000000000000008f00000000",
            INIT_30 => X"0000007c000000000000007e0000000000000089000000000000007f00000000",
            INIT_31 => X"0000009a00000000000000850000000000000086000000000000008800000000",
            INIT_32 => X"000000000000000000000000000000000000008d00000000000000af00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000000b000000000000001c00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000033000000000000001400000000",
            INIT_39 => X"000000000000000000000000000000000000001e000000000000001400000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_3B => X"00000028000000000000001c000000000000003e000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000190000000000000000000000000000001e000000000000000700000000",
            INIT_3E => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000006000000000000001a0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_43 => X"00000000000000000000001d0000000000000004000000000000000f00000000",
            INIT_44 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_45 => X"000000020000000000000000000000000000002f000000000000002500000000",
            INIT_46 => X"0000000000000000000000000000000000000003000000000000004f00000000",
            INIT_47 => X"0000002600000000000000000000000000000006000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_49 => X"0000000d000000000000000d0000000000000018000000000000000000000000",
            INIT_4A => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_4B => X"0000000800000000000000180000000000000000000000000000000900000000",
            INIT_4C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_4E => X"00000000000000000000001e000000000000003d000000000000000000000000",
            INIT_4F => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_51 => X"0000003200000000000000220000000000000000000000000000002e00000000",
            INIT_52 => X"0000003600000000000000000000000000000000000000000000000300000000",
            INIT_53 => X"00000000000000000000000d000000000000003a000000000000002600000000",
            INIT_54 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000150000000000000012000000000000000000000000",
            INIT_56 => X"00000031000000000000001f000000000000002e000000000000000000000000",
            INIT_57 => X"0000000800000000000000000000000000000000000000000000000100000000",
            INIT_58 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_59 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000000000000000000000000000000000000d000000000000000f00000000",
            INIT_5B => X"0000004100000000000000210000000000000016000000000000000000000000",
            INIT_5C => X"000000a200000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000c0000000000000037000000000000003f000000000000005200000000",
            INIT_5E => X"0000000000000000000000020000000000000000000000000000000600000000",
            INIT_5F => X"00000036000000000000000d0000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000560000000000000041000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_62 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_63 => X"0000002500000000000000000000000000000002000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000006000000000000003e00000000",
            INIT_65 => X"0000000700000000000000000000000000000000000000000000000100000000",
            INIT_66 => X"0000004200000000000000000000000000000000000000000000000a00000000",
            INIT_67 => X"0000003600000000000000180000000000000000000000000000000c00000000",
            INIT_68 => X"0000000000000000000000090000000000000013000000000000002400000000",
            INIT_69 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000000000000000000001f0000000000000004000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"000000070000000000000000000000000000002d000000000000000500000000",
            INIT_79 => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_7B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000300000000000000000000000000000000000000000000003b00000000",
            INIT_7D => X"0000000600000000000000010000000000000010000000000000000000000000",
            INIT_7E => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_7F => X"0000005d00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE4;


    MEM_GOLD_LAYER0_INSTANCE5 : if BRAM_NAME = "gold_layer0_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000000000000000000000f000000000000001c000000000000000000000000",
            INIT_03 => X"0000000000000000000000520000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000130000000000000012000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_06 => X"0000000500000000000000000000000000000017000000000000000c00000000",
            INIT_07 => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000003000000000000001d00000000",
            INIT_09 => X"0000000000000000000000110000000000000000000000000000001600000000",
            INIT_0A => X"0000000800000000000000000000000000000000000000000000001200000000",
            INIT_0B => X"0000001b00000000000000000000000000000011000000000000000000000000",
            INIT_0C => X"0000001900000000000000090000000000000000000000000000000000000000",
            INIT_0D => X"000000030000000000000000000000000000003b000000000000000000000000",
            INIT_0E => X"0000000000000000000000050000000000000000000000000000001000000000",
            INIT_0F => X"0000000000000000000000120000000000000012000000000000000000000000",
            INIT_10 => X"00000000000000000000000d0000000000000033000000000000000000000000",
            INIT_11 => X"0000002d00000000000000000000000000000000000000000000005800000000",
            INIT_12 => X"0000002800000000000000020000000000000000000000000000000400000000",
            INIT_13 => X"0000001d000000000000002c000000000000003e000000000000003300000000",
            INIT_14 => X"0000003b00000000000000000000000000000036000000000000007000000000",
            INIT_15 => X"0000004e000000000000004e000000000000002e000000000000000000000000",
            INIT_16 => X"00000056000000000000004f0000000000000049000000000000004400000000",
            INIT_17 => X"0000005a0000000000000053000000000000005a000000000000005800000000",
            INIT_18 => X"0000000000000000000000080000000000000048000000000000006f00000000",
            INIT_19 => X"0000004c000000000000004a0000000000000048000000000000004900000000",
            INIT_1A => X"00000057000000000000005b000000000000005b000000000000005400000000",
            INIT_1B => X"00000060000000000000005a000000000000005e000000000000005d00000000",
            INIT_1C => X"0000005000000000000000310000000000000000000000000000008a00000000",
            INIT_1D => X"000000570000000000000053000000000000004d000000000000004500000000",
            INIT_1E => X"0000007400000000000000610000000000000064000000000000006100000000",
            INIT_1F => X"0000006700000000000000670000000000000050000000000000005e00000000",
            INIT_20 => X"00000055000000000000005f0000000000000049000000000000004100000000",
            INIT_21 => X"0000005200000000000000520000000000000052000000000000004900000000",
            INIT_22 => X"000000450000000000000053000000000000006b000000000000005e00000000",
            INIT_23 => X"0000002e0000000000000033000000000000002e000000000000002f00000000",
            INIT_24 => X"0000002f0000000000000031000000000000002f000000000000002f00000000",
            INIT_25 => X"00000027000000000000001c0000000000000023000000000000002b00000000",
            INIT_26 => X"0000003200000000000000240000000000000027000000000000002600000000",
            INIT_27 => X"00000034000000000000002d0000000000000035000000000000003200000000",
            INIT_28 => X"0000000400000000000000250000000000000013000000000000005500000000",
            INIT_29 => X"0000002400000000000000150000000000000013000000000000002100000000",
            INIT_2A => X"0000003b000000000000001a0000000000000028000000000000002d00000000",
            INIT_2B => X"0000002c0000000000000038000000000000002e000000000000003400000000",
            INIT_2C => X"0000004f000000000000001a0000000000000000000000000000000000000000",
            INIT_2D => X"000000270000000000000004000000000000000b000000000000000a00000000",
            INIT_2E => X"0000002c00000000000000790000000000000000000000000000003900000000",
            INIT_2F => X"0000001a00000000000000230000000000000025000000000000003600000000",
            INIT_30 => X"0000000000000000000000530000000000000018000000000000000800000000",
            INIT_31 => X"00000053000000000000000e0000000000000000000000000000001200000000",
            INIT_32 => X"00000049000000000000000a0000000000000063000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000001a000000000000002c00000000",
            INIT_34 => X"00000000000000000000000b000000000000005f000000000000000800000000",
            INIT_35 => X"0000000000000000000000390000000000000000000000000000001e00000000",
            INIT_36 => X"00000049000000000000002e0000000000000000000000000000003800000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000230000000000000000000000000000000000000000000000bf00000000",
            INIT_39 => X"000000150000000000000000000000000000000d000000000000000400000000",
            INIT_3A => X"0000005000000000000000610000000000000000000000000000000c00000000",
            INIT_3B => X"000000a400000000000000000000000000000000000000000000000a00000000",
            INIT_3C => X"00000027000000000000001e0000000000000000000000000000000000000000",
            INIT_3D => X"0000000100000000000000000000000000000000000000000000000d00000000",
            INIT_3E => X"0000000000000000000000680000000000000045000000000000000000000000",
            INIT_3F => X"00000000000000000000007c0000000000000000000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000120000000000000022000000000000002a000000000000000000000000",
            INIT_41 => X"0000003c00000000000000000000000000000017000000000000000000000000",
            INIT_42 => X"0000001c00000000000000000000000000000003000000000000001100000000",
            INIT_43 => X"0000000000000000000000220000000000000006000000000000003100000000",
            INIT_44 => X"0000000a0000000000000044000000000000003a000000000000002600000000",
            INIT_45 => X"00000000000000000000004a0000000000000000000000000000001800000000",
            INIT_46 => X"00000017000000000000000e000000000000002a000000000000001900000000",
            INIT_47 => X"0000004800000000000000050000000000000000000000000000000a00000000",
            INIT_48 => X"000000110000000000000051000000000000001c000000000000005600000000",
            INIT_49 => X"0000000b000000000000000000000000000000a3000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000005600000000",
            INIT_4B => X"0000001e000000000000002d0000000000000028000000000000001400000000",
            INIT_4C => X"0000000000000000000000280000000000000040000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000009800000000",
            INIT_4E => X"0000001000000000000000090000000000000000000000000000000000000000",
            INIT_4F => X"000000000000000000000011000000000000000e000000000000001000000000",
            INIT_50 => X"0000001f00000000000000480000000000000041000000000000000300000000",
            INIT_51 => X"0000000a00000000000000050000000000000009000000000000000000000000",
            INIT_52 => X"0000001700000000000000140000000000000010000000000000000800000000",
            INIT_53 => X"0000000000000000000000170000000000000008000000000000001000000000",
            INIT_54 => X"0000000000000000000000000000000000000074000000000000001000000000",
            INIT_55 => X"0000000d00000000000000090000000000000000000000000000001100000000",
            INIT_56 => X"000000000000000000000009000000000000000d000000000000001000000000",
            INIT_57 => X"0000000d00000000000000000000000000000000000000000000002600000000",
            INIT_58 => X"0000001600000000000000000000000000000000000000000000001900000000",
            INIT_59 => X"0000001000000000000000180000000000000009000000000000000c00000000",
            INIT_5A => X"000000030000000000000031000000000000000b000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_61 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000001200000000000000040000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000270000000000000001000000000000000000000000",
            INIT_6B => X"0000000000000000000000080000000000000038000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_71 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE5;


    MEM_GOLD_LAYER0_INSTANCE6 : if BRAM_NAME = "gold_layer0_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_01 => X"00000030000000000000001e0000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_03 => X"000000010000000000000024000000000000001c000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000036000000000000002f0000000000000000000000000000000000000000",
            INIT_14 => X"0000003000000000000000350000000000000035000000000000003300000000",
            INIT_15 => X"0000002b0000000000000036000000000000003b000000000000003900000000",
            INIT_16 => X"0000002800000000000000250000000000000020000000000000002000000000",
            INIT_17 => X"0000003600000000000000380000000000000030000000000000002700000000",
            INIT_18 => X"0000003b00000000000000420000000000000033000000000000003900000000",
            INIT_19 => X"0000000200000000000000020000000000000023000000000000003900000000",
            INIT_1A => X"0000002700000000000000110000000000000006000000000000000600000000",
            INIT_1B => X"0000003900000000000000360000000000000013000000000000003000000000",
            INIT_1C => X"00000000000000000000001e000000000000003d000000000000003700000000",
            INIT_1D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_1E => X"0000001500000000000000170000000000000000000000000000000100000000",
            INIT_1F => X"0000004000000000000000370000000000000032000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000001e000000000000001200000000",
            INIT_21 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_22 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000003300000000000000440000000000000010000000000000003400000000",
            INIT_24 => X"0000000000000000000000000000000000000006000000000000002500000000",
            INIT_25 => X"0000000000000000000000000000000000000009000000000000001000000000",
            INIT_26 => X"00000031000000000000000f0000000000000000000000000000000000000000",
            INIT_27 => X"0000002b000000000000000d000000000000000b000000000000003800000000",
            INIT_28 => X"0000002a0000000000000000000000000000000b000000000000000800000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000003d0000000000000007000000000000002c000000000000000000000000",
            INIT_2B => X"00000017000000000000002e0000000000000011000000000000000e00000000",
            INIT_2C => X"0000000000000000000000130000000000000003000000000000000800000000",
            INIT_2D => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000250000000000000000000000000000001900000000",
            INIT_2F => X"00000000000000000000000a000000000000002e000000000000002200000000",
            INIT_30 => X"000000000000000000000000000000000000000f000000000000001300000000",
            INIT_31 => X"0000001100000000000000150000000000000000000000000000000200000000",
            INIT_32 => X"00000000000000000000001c0000000000000000000000000000000900000000",
            INIT_33 => X"0000002c0000000000000000000000000000000c000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"00000014000000000000000e0000000000000016000000000000002100000000",
            INIT_36 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_37 => X"0000000000000000000000050000000000000006000000000000001f00000000",
            INIT_38 => X"00000028000000000000001e0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000150000000000000014000000000000000500000000",
            INIT_3A => X"0000001700000000000000110000000000000006000000000000002c00000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000003c00000000000000320000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000002c00000000000000290000000000000023000000000000002200000000",
            INIT_4D => X"0000002f000000000000002b0000000000000028000000000000002000000000",
            INIT_4E => X"0000001e000000000000001d0000000000000029000000000000003200000000",
            INIT_4F => X"000000240000000000000028000000000000002e000000000000002900000000",
            INIT_50 => X"0000000e0000000000000021000000000000002c000000000000002400000000",
            INIT_51 => X"00000005000000000000002e0000000000000030000000000000004300000000",
            INIT_52 => X"0000001500000000000000190000000000000029000000000000002100000000",
            INIT_53 => X"000000280000000000000002000000000000003f000000000000002c00000000",
            INIT_54 => X"000000280000000000000020000000000000002a000000000000002900000000",
            INIT_55 => X"0000001c00000000000000000000000000000010000000000000002400000000",
            INIT_56 => X"0000000b000000000000001a0000000000000032000000000000000c00000000",
            INIT_57 => X"00000024000000000000002e0000000000000000000000000000005c00000000",
            INIT_58 => X"000000250000000000000027000000000000000c000000000000003800000000",
            INIT_59 => X"0000001800000000000000230000000000000000000000000000001900000000",
            INIT_5A => X"0000002c00000000000000000000000000000026000000000000001a00000000",
            INIT_5B => X"0000001300000000000000000000000000000041000000000000000500000000",
            INIT_5C => X"000000250000000000000024000000000000002a000000000000002700000000",
            INIT_5D => X"0000001200000000000000380000000000000014000000000000000000000000",
            INIT_5E => X"000000000000000000000024000000000000001a000000000000002b00000000",
            INIT_5F => X"000000000000000000000000000000000000002f000000000000003700000000",
            INIT_60 => X"0000000000000000000000430000000000000025000000000000001600000000",
            INIT_61 => X"0000001d0000000000000007000000000000002a000000000000003400000000",
            INIT_62 => X"0000000e00000000000000240000000000000011000000000000002000000000",
            INIT_63 => X"0000001500000000000000000000000000000000000000000000004600000000",
            INIT_64 => X"0000002b00000000000000000000000000000039000000000000001c00000000",
            INIT_65 => X"000000250000000000000000000000000000000d000000000000002800000000",
            INIT_66 => X"0000003400000000000000290000000000000006000000000000000b00000000",
            INIT_67 => X"0000000b00000000000000350000000000000000000000000000000200000000",
            INIT_68 => X"0000002c00000000000000110000000000000000000000000000001800000000",
            INIT_69 => X"0000000d000000000000000d0000000000000011000000000000000000000000",
            INIT_6A => X"000000340000000000000000000000000000003f000000000000000000000000",
            INIT_6B => X"00000000000000000000001b000000000000000e000000000000000000000000",
            INIT_6C => X"00000000000000000000002b0000000000000005000000000000003f00000000",
            INIT_6D => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_6E => X"00000014000000000000002a0000000000000000000000000000003900000000",
            INIT_6F => X"0000000f000000000000002c000000000000001d000000000000000000000000",
            INIT_70 => X"000000100000000000000000000000000000000f000000000000002f00000000",
            INIT_71 => X"0000003800000000000000000000000000000000000000000000002f00000000",
            INIT_72 => X"0000000000000000000000320000000000000029000000000000000000000000",
            INIT_73 => X"0000000f000000000000002b0000000000000027000000000000000500000000",
            INIT_74 => X"0000002100000000000000110000000000000008000000000000000800000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000005000000000000005200000000",
            INIT_77 => X"0000000000000000000000030000000000000007000000000000000000000000",
            INIT_78 => X"0000001400000000000000030000000000000000000000000000000000000000",
            INIT_79 => X"0000002e00000000000000220000000000000000000000000000000000000000",
            INIT_7A => X"0000000500000000000000020000000000000006000000000000000000000000",
            INIT_7B => X"0000000200000000000000000000000000000000000000000000000100000000",
            INIT_7C => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000000d0000000000000022000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000006000000000000000900000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE6;


    MEM_GOLD_LAYER0_INSTANCE7 : if BRAM_NAME = "gold_layer0_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000013000000000000001500000000",
            INIT_01 => X"0000000000000000000000000000000000000014000000000000000400000000",
            INIT_02 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000001a00000000000000120000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_INSTANCE7;


    MEM_GOLD_LAYER1_INSTANCE0 : if BRAM_NAME = "gold_layer1_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000210000000000000037000000000000006c000000000000006000000000",
            INIT_0E => X"00000000000000000000004c000000000000000c000000000000003800000000",
            INIT_0F => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000000000002a000000000000000f00000000",
            INIT_11 => X"0000002b00000000000000000000000000000007000000000000001500000000",
            INIT_12 => X"0000001300000000000000110000000000000061000000000000005f00000000",
            INIT_13 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"000000000000000000000073000000000000005d000000000000000000000000",
            INIT_15 => X"0000005a00000000000000b80000000000000046000000000000004300000000",
            INIT_16 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000002300000000000000d600000000",
            INIT_18 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_19 => X"0000001f000000000000003a000000000000001c000000000000000000000000",
            INIT_1A => X"00000000000000000000000e000000000000013a000000000000002700000000",
            INIT_1B => X"00000038000000000000002400000000000000c2000000000000001d00000000",
            INIT_1C => X"000000170000000000000000000000000000006f000000000000008000000000",
            INIT_1D => X"000000000000000000000000000000000000002200000000000001cf00000000",
            INIT_1E => X"000000f200000000000000600000000000000000000000000000001600000000",
            INIT_1F => X"0000017a00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000a00000000000000000000000000000000000000000000009200000000",
            INIT_21 => X"000000ce000000000000009d0000000000000000000000000000000000000000",
            INIT_22 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_23 => X"0000000c000000000000007c0000000000000000000000000000007b00000000",
            INIT_24 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_25 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000036000000000000000000000000",
            INIT_2A => X"0000000000000000000000380000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"00000000000000000000004b0000000000000000000000000000000000000000",
            INIT_2D => X"0000009d00000000000000000000000000000077000000000000000000000000",
            INIT_2E => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_30 => X"0000002100000000000000000000000000000013000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_34 => X"0000006e00000000000000000000000000000079000000000000000000000000",
            INIT_35 => X"0000006a00000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000cb0000000000000000000000000000000000000000",
            INIT_38 => X"00000039000000000000003c0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000037000000000000001b00000000",
            INIT_3A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"000000b600000000000000320000000000000000000000000000000000000000",
            INIT_3C => X"0000000a00000000000000000000000000000008000000000000000000000000",
            INIT_3D => X"0000000000000000000000670000000000000039000000000000000000000000",
            INIT_3E => X"0000002e00000000000000110000000000000020000000000000000c00000000",
            INIT_3F => X"000000150000000000000000000000000000002a000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000170000000000000009000000000000003600000000",
            INIT_41 => X"0000000b00000000000000090000000000000000000000000000000000000000",
            INIT_42 => X"0000001700000000000000000000000000000006000000000000001900000000",
            INIT_43 => X"000000090000000000000029000000000000000d000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"00000009000000000000000d0000000000000000000000000000001700000000",
            INIT_48 => X"0000001a00000000000000260000000000000016000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000200000000000000010000000000000000000000000000000500000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000e0000000000000000000000000000001b000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000100000000000000000000000000000002000000000000003b00000000",
            INIT_55 => X"0000000000000000000000150000000000000018000000000000000600000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000050000000000000000000000000000000b00000000",
            INIT_58 => X"0000001c00000000000000060000000000000011000000000000000000000000",
            INIT_59 => X"0000001f00000000000000000000000000000001000000000000004000000000",
            INIT_5A => X"0000002d00000000000000170000000000000005000000000000000c00000000",
            INIT_5B => X"0000000800000000000000120000000000000021000000000000000800000000",
            INIT_5C => X"0000000000000000000000300000000000000022000000000000001300000000",
            INIT_5D => X"0000000000000000000000310000000000000038000000000000000000000000",
            INIT_5E => X"000000080000000000000000000000000000001a000000000000002e00000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000004a00000000000000000000000000000000000000000000002200000000",
            INIT_63 => X"000000000000000000000032000000000000002a000000000000004a00000000",
            INIT_64 => X"00000000000000000000000a0000000000000009000000000000000900000000",
            INIT_65 => X"0000000000000000000000000000000000000032000000000000001100000000",
            INIT_66 => X"0000003e00000000000000000000000000000005000000000000000000000000",
            INIT_67 => X"00000000000000000000001f0000000000000019000000000000000400000000",
            INIT_68 => X"00000000000000000000004e0000000000000000000000000000005b00000000",
            INIT_69 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_6A => X"0000000d0000000000000000000000000000005b000000000000005d00000000",
            INIT_6B => X"00000000000000000000005f0000000000000083000000000000000000000000",
            INIT_6C => X"0000005b00000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_72 => X"00000000000000000000003c0000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000360000000000000000000000000000001700000000",
            INIT_74 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_75 => X"000000080000000000000000000000000000001f000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000000e000000000000001700000000",
            INIT_77 => X"0000003b00000000000000aa0000000000000000000000000000000000000000",
            INIT_78 => X"00000000000000000000002f0000000000000027000000000000005600000000",
            INIT_79 => X"0000004d00000000000000560000000000000087000000000000002700000000",
            INIT_7A => X"0000006100000000000000680000000000000072000000000000004c00000000",
            INIT_7B => X"00000000000000000000002d0000000000000094000000000000005100000000",
            INIT_7C => X"0000002500000000000000380000000000000000000000000000004d00000000",
            INIT_7D => X"0000000a000000000000000c0000000000000018000000000000000000000000",
            INIT_7E => X"00000000000000000000002d000000000000009b000000000000000000000000",
            INIT_7F => X"000000000000000000000000000000000000001c000000000000000e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE0;


    MEM_GOLD_LAYER1_INSTANCE1 : if BRAM_NAME = "gold_layer1_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003900000000000000390000000000000074000000000000000000000000",
            INIT_01 => X"000000000000000000000000000000000000001b000000000000003600000000",
            INIT_02 => X"0000001d000000000000004b0000000000000000000000000000001300000000",
            INIT_03 => X"000000920000000000000050000000000000004d000000000000000200000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000005000000000",
            INIT_05 => X"000000000000000000000000000000000000009e000000000000002400000000",
            INIT_06 => X"0000003200000000000000150000000000000012000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000001c000000000000004b00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"00000000000000000000004e0000000000000000000000000000000000000000",
            INIT_0A => X"0000002c00000000000000370000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_0C => X"0000000000000000000000640000000000000000000000000000000000000000",
            INIT_0D => X"0000001300000000000000110000000000000000000000000000003f00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000002000000000000005f0000000000000000000000000000000000000000",
            INIT_10 => X"0000001400000000000000000000000000000007000000000000000000000000",
            INIT_11 => X"0000000400000000000000530000000000000004000000000000000b00000000",
            INIT_12 => X"00000017000000000000002e0000000000000032000000000000001800000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_19 => X"0000000e00000000000000000000000000000016000000000000000000000000",
            INIT_1A => X"0000000600000000000000000000000000000000000000000000001e00000000",
            INIT_1B => X"0000002100000000000000010000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"000000000000000000000000000000000000001b000000000000001200000000",
            INIT_1E => X"0000004100000000000000380000000000000039000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000007c00000000000000170000000000000000000000000000002300000000",
            INIT_27 => X"00000000000000000000001a0000000000000000000000000000000300000000",
            INIT_28 => X"000000150000000000000000000000000000001a000000000000000000000000",
            INIT_29 => X"0000000000000000000000170000000000000018000000000000000600000000",
            INIT_2A => X"00000024000000000000001e000000000000000c000000000000000000000000",
            INIT_2B => X"0000009200000000000000810000000000000040000000000000003500000000",
            INIT_2C => X"000000000000000000000019000000000000006c000000000000002700000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000003300000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000070000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_31 => X"00000038000000000000004f000000000000001c000000000000000000000000",
            INIT_32 => X"0000000000000000000000360000000000000000000000000000003800000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000650000000000000042000000000000001c000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000066000000000000002600000000",
            INIT_3C => X"000000560000000000000059000000000000004e000000000000006200000000",
            INIT_3D => X"0000004d00000000000000000000000000000019000000000000007700000000",
            INIT_3E => X"000000b700000000000000470000000000000035000000000000006000000000",
            INIT_3F => X"000000250000000000000028000000000000000c000000000000007400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007800000000000000850000000000000039000000000000001800000000",
            INIT_41 => X"00000084000000000000006e0000000000000050000000000000003900000000",
            INIT_42 => X"000000a9000000000000008b000000000000009a000000000000008a00000000",
            INIT_43 => X"000000bb00000000000000ab000000000000009c000000000000009200000000",
            INIT_44 => X"000000a6000000000000000a0000000000000000000000000000000000000000",
            INIT_45 => X"00000050000000000000006700000000000000a900000000000000b500000000",
            INIT_46 => X"00000000000000000000004d0000000000000097000000000000004600000000",
            INIT_47 => X"00000011000000000000002d000000000000001c000000000000000000000000",
            INIT_48 => X"0000002100000000000000000000000000000000000000000000001c00000000",
            INIT_49 => X"0000001d0000000000000068000000000000001d000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000002f000000000000002b0000000000000000000000000000000000000000",
            INIT_4C => X"00000040000000000000006a0000000000000034000000000000003700000000",
            INIT_4D => X"00000056000000000000006700000000000000d1000000000000002400000000",
            INIT_4E => X"0000006100000000000000170000000000000042000000000000007300000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_59 => X"0000009b00000000000000b30000000000000000000000000000006800000000",
            INIT_5A => X"000000c1000000000000007c000000000000009c000000000000007d00000000",
            INIT_5B => X"000000a9000000000000009800000000000000a0000000000000007d00000000",
            INIT_5C => X"0000001c000000000000000600000000000000b000000000000000c200000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000006200000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000500000000000000051000000000000004b000000000000006100000000",
            INIT_6A => X"0000008800000000000000610000000000000041000000000000004900000000",
            INIT_6B => X"0000005a000000000000005e000000000000005b000000000000005300000000",
            INIT_6C => X"00000060000000000000005a0000000000000068000000000000002a00000000",
            INIT_6D => X"0000003c0000000000000073000000000000005f000000000000007600000000",
            INIT_6E => X"0000007b000000000000004e000000000000006d000000000000007600000000",
            INIT_6F => X"0000005c000000000000005d0000000000000041000000000000004600000000",
            INIT_70 => X"0000004f000000000000003b0000000000000046000000000000009700000000",
            INIT_71 => X"0000002e00000000000000230000000000000015000000000000001000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000002f00000000",
            INIT_73 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000057000000000000007b0000000000000073000000000000006300000000",
            INIT_76 => X"000000450000000000000048000000000000004b000000000000005600000000",
            INIT_77 => X"0000000500000000000000400000000000000043000000000000007000000000",
            INIT_78 => X"00000032000000000000002b0000000000000044000000000000001200000000",
            INIT_79 => X"000000240000000000000000000000000000001e000000000000002200000000",
            INIT_7A => X"00000000000000000000005d0000000000000007000000000000003c00000000",
            INIT_7B => X"0000002100000000000000210000000000000000000000000000000900000000",
            INIT_7C => X"0000001500000000000000000000000000000006000000000000000000000000",
            INIT_7D => X"00000000000000000000002b0000000000000017000000000000001900000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE1;


    MEM_GOLD_LAYER1_INSTANCE2 : if BRAM_NAME = "gold_layer1_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000004a000000000000005e000000000000005a000000000000000000000000",
            INIT_02 => X"0000004700000000000000310000000000000026000000000000002c00000000",
            INIT_03 => X"0000002600000000000000000000000000000036000000000000003c00000000",
            INIT_04 => X"00000050000000000000003e000000000000003a000000000000002600000000",
            INIT_05 => X"0000003100000000000000460000000000000002000000000000000e00000000",
            INIT_06 => X"00000035000000000000003f000000000000002d000000000000002e00000000",
            INIT_07 => X"000000350000000000000044000000000000005a000000000000002600000000",
            INIT_08 => X"00000000000000000000001c0000000000000044000000000000004900000000",
            INIT_09 => X"0000001d0000000000000000000000000000002c000000000000000800000000",
            INIT_0A => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_11 => X"0000001100000000000000320000000000000000000000000000000a00000000",
            INIT_12 => X"0000004c00000000000000000000000000000011000000000000000000000000",
            INIT_13 => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_14 => X"0000001c00000000000000760000000000000000000000000000000200000000",
            INIT_15 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_16 => X"0000007b0000000000000012000000000000006e000000000000000000000000",
            INIT_17 => X"0000003e0000000000000018000000000000001a000000000000008600000000",
            INIT_18 => X"00000033000000000000003d00000000000000af000000000000000000000000",
            INIT_19 => X"00000116000000000000004c0000000000000048000000000000003500000000",
            INIT_1A => X"0000007400000000000000d100000000000000be000000000000010a00000000",
            INIT_1B => X"000000f000000000000000be00000000000000c1000000000000006c00000000",
            INIT_1C => X"0000000300000000000000350000000000000015000000000000009600000000",
            INIT_1D => X"0000007b000000000000003e0000000000000055000000000000002b00000000",
            INIT_1E => X"0000001000000000000000000000000000000034000000000000001c00000000",
            INIT_1F => X"0000001100000000000000570000000000000064000000000000004000000000",
            INIT_20 => X"0000001f00000000000000400000000000000000000000000000000a00000000",
            INIT_21 => X"0000002f00000000000000270000000000000030000000000000004000000000",
            INIT_22 => X"0000000000000000000000370000000000000076000000000000001700000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000090000000000000000000000000000006c000000000000000000000000",
            INIT_28 => X"0000000000000000000000970000000000000000000000000000000000000000",
            INIT_29 => X"00000000000000000000006f0000000000000084000000000000006500000000",
            INIT_2A => X"000000b0000000000000000000000000000000ed000000000000000000000000",
            INIT_2B => X"00000000000000000000007900000000000000c4000000000000006200000000",
            INIT_2C => X"0000000000000000000000920000000000000000000000000000005300000000",
            INIT_2D => X"0000007600000000000000250000000000000000000000000000004600000000",
            INIT_2E => X"000000000000000000000000000000000000001f000000000000005300000000",
            INIT_2F => X"00000024000000000000000000000000000000a2000000000000000000000000",
            INIT_30 => X"0000001100000000000000060000000000000000000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_32 => X"0000001e00000000000000000000000000000006000000000000000000000000",
            INIT_33 => X"000000240000000000000032000000000000005c000000000000001100000000",
            INIT_34 => X"00000034000000000000008a0000000000000050000000000000009e00000000",
            INIT_35 => X"000000420000000000000026000000000000002c000000000000004600000000",
            INIT_36 => X"00000097000000000000002e0000000000000059000000000000003600000000",
            INIT_37 => X"0000002a00000000000000220000000000000036000000000000002200000000",
            INIT_38 => X"0000000000000000000000270000000000000035000000000000003100000000",
            INIT_39 => X"000000a600000000000000af0000000000000017000000000000001f00000000",
            INIT_3A => X"0000002100000000000000660000000000000037000000000000002b00000000",
            INIT_3B => X"0000002800000000000000bd000000000000009a000000000000001c00000000",
            INIT_3C => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000001f000000000000000b0000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001800000000000000300000000000000000000000000000000000000000",
            INIT_46 => X"000000190000000000000020000000000000002a000000000000000500000000",
            INIT_47 => X"00000086000000000000007e0000000000000047000000000000000000000000",
            INIT_48 => X"000000b000000000000000b300000000000000a7000000000000008a00000000",
            INIT_49 => X"000000a300000000000000ae000000000000007d00000000000000d000000000",
            INIT_4A => X"0000000000000000000000e100000000000000bf00000000000000ac00000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_4C => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000004e0000000000000000000000000000002a000000000000002f00000000",
            INIT_4E => X"0000000000000000000000650000000000000000000000000000000000000000",
            INIT_4F => X"00000000000000000000003a0000000000000000000000000000005300000000",
            INIT_50 => X"0000005000000000000000000000000000000005000000000000001100000000",
            INIT_51 => X"0000001c00000000000000000000000000000025000000000000000000000000",
            INIT_52 => X"000000000000000000000000000000000000008b000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_55 => X"0000001200000000000000000000000000000000000000000000000400000000",
            INIT_56 => X"0000000a0000000000000024000000000000000d000000000000001800000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000005000000000000000040000000000000000000000000000004d00000000",
            INIT_59 => X"0000003300000000000000000000000000000000000000000000001200000000",
            INIT_5A => X"0000003f0000000000000000000000000000001e000000000000000000000000",
            INIT_5B => X"0000000000000000000000910000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000250000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"00000000000000000000000a0000000000000044000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000077000000000000000000000000",
            INIT_60 => X"0000006700000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000a60000000000000005000000000000004200000000",
            INIT_62 => X"0000003800000000000000410000000000000030000000000000006100000000",
            INIT_63 => X"0000000000000000000000030000000000000000000000000000000b00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"00000023000000000000004e0000000000000029000000000000000000000000",
            INIT_66 => X"0000002300000000000000000000000000000022000000000000000000000000",
            INIT_67 => X"00000000000000000000006f000000000000002d000000000000000000000000",
            INIT_68 => X"00000000000000000000005c000000000000002e000000000000000500000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000002e0000000000000003000000000000002b000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000000000000000000053000000000000005e000000000000005e00000000",
            INIT_6E => X"0000003600000000000000300000000000000000000000000000000000000000",
            INIT_6F => X"000000b000000000000000900000000000000039000000000000003000000000",
            INIT_70 => X"0000004a0000000000000067000000000000006700000000000000a200000000",
            INIT_71 => X"0000007900000000000000b4000000000000006a000000000000006800000000",
            INIT_72 => X"000000430000000000000014000000000000003b000000000000002500000000",
            INIT_73 => X"000000000000000000000042000000000000006a000000000000003400000000",
            INIT_74 => X"0000000000000000000000240000000000000000000000000000003400000000",
            INIT_75 => X"000000270000000000000000000000000000002c000000000000002200000000",
            INIT_76 => X"000000330000000000000000000000000000003c000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000008000000000000001700000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_7E => X"0000000a00000000000000160000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000001000000000000002d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE2;


    MEM_GOLD_LAYER1_INSTANCE3 : if BRAM_NAME = "gold_layer1_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002f00000000000000120000000000000017000000000000000300000000",
            INIT_01 => X"000000080000000000000000000000000000001e000000000000004500000000",
            INIT_02 => X"0000006000000000000000000000000000000002000000000000001500000000",
            INIT_03 => X"0000003a00000000000000270000000000000039000000000000004200000000",
            INIT_04 => X"0000000700000000000000690000000000000026000000000000003a00000000",
            INIT_05 => X"00000088000000000000007e000000000000007e000000000000004800000000",
            INIT_06 => X"00000092000000000000006600000000000000bb000000000000009600000000",
            INIT_07 => X"000000ab00000000000000a9000000000000009e000000000000009600000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER1_INSTANCE3;


    MEM_GOLD_LAYER2_INSTANCE0 : if BRAM_NAME = "gold_layer2_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000001040000000000000040000000000000001200000000000000a000000000",
            INIT_01 => X"00000000000000000000010100000000000000bc000000000000005100000000",
            INIT_02 => X"0000001c00000000000000000000000000000047000000000000000000000000",
            INIT_03 => X"0000000000000000000000ba0000000000000000000000000000000000000000",
            INIT_04 => X"0000003100000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000920000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000200000000000000000000000000000000000000000000010400000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000038000000000000000000000000000000a8000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000370000000000000053000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000134000000000000017a00000000000000a8000000000000000000000000",
            INIT_15 => X"000000b700000000000000820000000000000113000000000000003700000000",
            INIT_16 => X"0000002d00000000000000000000000000000000000000000000003500000000",
            INIT_17 => X"00000062000000000000014d0000000000000000000000000000007900000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000350000000000000010000000000000007e000000000000000000000000",
            INIT_1A => X"000000d10000000000000000000000000000006a000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"000000a0000000000000000000000000000000b000000000000000b000000000",
            INIT_1D => X"0000008100000000000000d20000000000000077000000000000003300000000",
            INIT_1E => X"000000080000000000000000000000000000000000000000000000c600000000",
            INIT_1F => X"000000650000000000000000000000000000005700000000000000a900000000",
            INIT_20 => X"0000003c00000000000000a1000000000000000000000000000000c800000000",
            INIT_21 => X"00000000000000000000007a0000000000000058000000000000000000000000",
            INIT_22 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000005c00000000",
            INIT_24 => X"0000000000000000000000e6000000000000002c000000000000000000000000",
            INIT_25 => X"000000ff00000000000000000000000000000048000000000000007700000000",
            INIT_26 => X"0000001900000000000000000000000000000000000000000000002400000000",
            INIT_27 => X"0000000000000000000000000000000000000036000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000004d000000000000005d0000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000aa000000000000006c00000000000000b500000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"00000030000000000000001b0000000000000000000000000000003f00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_31 => X"00000012000000000000000000000000000000b3000000000000011900000000",
            INIT_32 => X"000000bd000000000000000000000000000000aa000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000002600000000000000b600000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"00000144000000000000012400000000000000c0000000000000000000000000",
            INIT_39 => X"00000017000000000000006800000000000000d0000000000000014f00000000",
            INIT_3A => X"0000000000000000000000000000000000000040000000000000000000000000",
            INIT_3B => X"0000000000000000000000160000000000000057000000000000000900000000",
            INIT_3C => X"000000000000000000000000000000000000005d00000000000000cf00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000b8000000000000000100000000000000a8000000000000000000000000",
            INIT_42 => X"0000009000000000000000960000000000000028000000000000001e00000000",
            INIT_43 => X"0000000000000000000000000000000000000063000000000000001500000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000009e000000000000011b0000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000006c0000000000000000000000000000000000000000",
            INIT_49 => X"0000007900000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"000000ff0000000000000004000000000000004300000000000000f800000000",
            INIT_4B => X"0000000000000000000000110000000000000012000000000000006700000000",
            INIT_4C => X"000000690000000000000000000000000000001c000000000000000000000000",
            INIT_4D => X"0000004e00000000000000860000000000000000000000000000004100000000",
            INIT_4E => X"0000009100000000000000000000000000000000000000000000003100000000",
            INIT_4F => X"0000002600000000000000170000000000000051000000000000006c00000000",
            INIT_50 => X"000000fd00000000000000b00000000000000000000000000000004600000000",
            INIT_51 => X"000000000000000000000078000000000000000000000000000000e000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_53 => X"000000ab00000000000000590000000000000000000000000000000000000000",
            INIT_54 => X"0000006a00000000000000ef00000000000000fb00000000000000c100000000",
            INIT_55 => X"00000053000000000000003b00000000000000db000000000000008f00000000",
            INIT_56 => X"0000000000000000000000000000000000000010000000000000001400000000",
            INIT_57 => X"0000006200000000000000ab0000000000000046000000000000007b00000000",
            INIT_58 => X"0000006d00000000000000a2000000000000013c000000000000005a00000000",
            INIT_59 => X"000000510000000000000123000000000000007a000000000000008c00000000",
            INIT_5A => X"00000000000000000000000000000000000000a1000000000000009700000000",
            INIT_5B => X"00000000000000000000003c0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_5D => X"0000010400000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000012f00000000000000a2000000000000004f000000000000001e00000000",
            INIT_60 => X"0000015b00000000000000000000000000000000000000000000008c00000000",
            INIT_61 => X"000000a100000000000000830000000000000161000000000000013a00000000",
            INIT_62 => X"0000000000000000000000120000000000000138000000000000007200000000",
            INIT_63 => X"000000dc00000000000000700000000000000088000000000000000000000000",
            INIT_64 => X"000000cd000000000000013e00000000000000ad00000000000000e000000000",
            INIT_65 => X"000000000000000000000000000000000000000000000000000000ae00000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000001f00000000000000c80000000000000000000000000000000000000000",
            INIT_68 => X"0000004e000000000000004b000000000000004600000000000000bf00000000",
            INIT_69 => X"0000001e00000000000000000000000000000026000000000000001b00000000",
            INIT_6A => X"00000036000000000000009f000000000000013b000000000000007300000000",
            INIT_6B => X"000000a500000000000000aa0000000000000006000000000000001e00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000010100000000000000760000000000000043000000000000006a00000000",
            INIT_76 => X"000000000000000000000000000000000000007c000000000000006600000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000005900000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000310000000000000000000000000000006900000000",
            INIT_7B => X"0000003d00000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000003100000000000000100000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000000000000000000000ed000000000000007200000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000012c00000000000000700000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE0;


    MEM_GOLD_LAYER2_INSTANCE1 : if BRAM_NAME = "gold_layer2_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000000000000000000d0000000000000017f00000000",
            INIT_01 => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_02 => X"0000002100000000000000390000000000000008000000000000006700000000",
            INIT_03 => X"000000760000000000000044000000000000006d00000000000000de00000000",
            INIT_04 => X"0000000000000000000000eb0000000000000141000000000000008400000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000003f000000000000006e000000000000007800000000000000b200000000",
            INIT_08 => X"0000000000000000000000000000000000000092000000000000007f00000000",
            INIT_09 => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000034000000000000001e0000000000000000000000000000019100000000",
            INIT_0B => X"0000000000000000000000000000000000000148000000000000008700000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000004a00000000000000580000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_0F => X"000000c500000000000000d700000000000000f3000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER2_INSTANCE1;


    MEM_GOLD_LAYER3_INSTANCE0 : if BRAM_NAME = "gold_layer3_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"fffff5e2fffffffffffef197fffffffffffe4d81fffffffffffdcd4cffffffff",
            INIT_01 => X"fffbdef2fffffffffffebfcffffffffffffe59b4ffffffffffff0ce7ffffffff",
            INIT_02 => X"fffe738afffffffffffd6804ffffffff",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER3_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "sampleifmap_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a600000000000000a5000000000000009f000000000000009e00000000",
            INIT_01 => X"0000009f00000000000000a2000000000000009c00000000000000a000000000",
            INIT_02 => X"000000a000000000000000a1000000000000009f000000000000009e00000000",
            INIT_03 => X"000000aa00000000000000a900000000000000a600000000000000a100000000",
            INIT_04 => X"000000a000000000000000a000000000000000a200000000000000a700000000",
            INIT_05 => X"0000009400000000000000960000000000000095000000000000009c00000000",
            INIT_06 => X"0000008d000000000000008c000000000000008f000000000000009500000000",
            INIT_07 => X"00000074000000000000007e0000000000000089000000000000008f00000000",
            INIT_08 => X"000000a6000000000000009f0000000000000097000000000000009800000000",
            INIT_09 => X"000000a200000000000000a400000000000000a000000000000000a200000000",
            INIT_0A => X"0000009f000000000000009b000000000000009c00000000000000a300000000",
            INIT_0B => X"000000ab00000000000000ab00000000000000aa00000000000000a300000000",
            INIT_0C => X"00000097000000000000009a00000000000000a000000000000000a900000000",
            INIT_0D => X"0000008d000000000000008c000000000000008b000000000000009100000000",
            INIT_0E => X"0000008e00000000000000910000000000000093000000000000009500000000",
            INIT_0F => X"00000077000000000000007d0000000000000088000000000000008f00000000",
            INIT_10 => X"000000a7000000000000009e0000000000000097000000000000009700000000",
            INIT_11 => X"000000a500000000000000a500000000000000a300000000000000a000000000",
            INIT_12 => X"0000009d000000000000009e00000000000000a200000000000000a300000000",
            INIT_13 => X"000000a900000000000000a700000000000000a600000000000000a100000000",
            INIT_14 => X"000000790000000000000091000000000000009f00000000000000aa00000000",
            INIT_15 => X"0000007200000000000000650000000000000062000000000000006e00000000",
            INIT_16 => X"0000008c000000000000008f0000000000000086000000000000007800000000",
            INIT_17 => X"000000780000000000000082000000000000008b000000000000008e00000000",
            INIT_18 => X"000000ae00000000000000a0000000000000009b000000000000009b00000000",
            INIT_19 => X"000000a900000000000000a900000000000000a700000000000000a700000000",
            INIT_1A => X"000000bf00000000000000a700000000000000a500000000000000a500000000",
            INIT_1B => X"000000a400000000000000a2000000000000009d00000000000000b100000000",
            INIT_1C => X"0000006700000000000000680000000000000095000000000000009e00000000",
            INIT_1D => X"0000004a0000000000000050000000000000005c000000000000006200000000",
            INIT_1E => X"0000008400000000000000710000000000000053000000000000005600000000",
            INIT_1F => X"0000007f0000000000000088000000000000008c000000000000008c00000000",
            INIT_20 => X"000000aa00000000000000a1000000000000009c000000000000009b00000000",
            INIT_21 => X"000000a600000000000000a900000000000000a300000000000000a900000000",
            INIT_22 => X"000000f600000000000000ad00000000000000a400000000000000a400000000",
            INIT_23 => X"0000008e0000000000000092000000000000009700000000000000c300000000",
            INIT_24 => X"000000710000000000000055000000000000004e000000000000006f00000000",
            INIT_25 => X"0000005d0000000000000061000000000000006a000000000000007000000000",
            INIT_26 => X"0000006900000000000000550000000000000054000000000000004a00000000",
            INIT_27 => X"000000810000000000000085000000000000008a000000000000008000000000",
            INIT_28 => X"0000009300000000000000820000000000000085000000000000009400000000",
            INIT_29 => X"000000a700000000000000a700000000000000a500000000000000a100000000",
            INIT_2A => X"000000b400000000000000a300000000000000a500000000000000a300000000",
            INIT_2B => X"0000004200000000000000610000000000000080000000000000009d00000000",
            INIT_2C => X"0000007600000000000000590000000000000042000000000000004500000000",
            INIT_2D => X"0000005e00000000000000720000000000000077000000000000007a00000000",
            INIT_2E => X"00000043000000000000003a000000000000005b000000000000006300000000",
            INIT_2F => X"00000086000000000000008a000000000000008c000000000000006c00000000",
            INIT_30 => X"00000058000000000000002f000000000000006d000000000000007f00000000",
            INIT_31 => X"000000aa00000000000000a800000000000000aa000000000000009900000000",
            INIT_32 => X"0000009300000000000000a400000000000000a600000000000000a900000000",
            INIT_33 => X"000000440000000000000064000000000000007f000000000000008100000000",
            INIT_34 => X"0000008400000000000000530000000000000048000000000000004e00000000",
            INIT_35 => X"0000006b0000000000000069000000000000007c000000000000009200000000",
            INIT_36 => X"0000002e000000000000003f0000000000000055000000000000007300000000",
            INIT_37 => X"00000086000000000000008d0000000000000084000000000000004f00000000",
            INIT_38 => X"00000046000000000000002a0000000000000063000000000000008300000000",
            INIT_39 => X"000000a800000000000000a500000000000000a7000000000000008f00000000",
            INIT_3A => X"00000078000000000000008c00000000000000a100000000000000ab00000000",
            INIT_3B => X"0000005800000000000000740000000000000090000000000000008200000000",
            INIT_3C => X"0000007c000000000000004d0000000000000055000000000000005b00000000",
            INIT_3D => X"0000006a0000000000000066000000000000008800000000000000a300000000",
            INIT_3E => X"0000003100000000000000360000000000000055000000000000006400000000",
            INIT_3F => X"00000088000000000000008a000000000000006b000000000000003900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007c0000000000000036000000000000006700000000000000aa00000000",
            INIT_41 => X"000000a600000000000000a300000000000000a1000000000000009900000000",
            INIT_42 => X"0000007d000000000000007100000000000000ae00000000000000a500000000",
            INIT_43 => X"000000560000000000000079000000000000009c000000000000009d00000000",
            INIT_44 => X"0000005100000000000000500000000000000054000000000000005200000000",
            INIT_45 => X"0000005700000000000000710000000000000092000000000000008a00000000",
            INIT_46 => X"0000003800000000000000470000000000000056000000000000005300000000",
            INIT_47 => X"000000890000000000000085000000000000004a000000000000002800000000",
            INIT_48 => X"0000009a000000000000005e000000000000008600000000000000b400000000",
            INIT_49 => X"00000099000000000000009c000000000000009e00000000000000ae00000000",
            INIT_4A => X"0000009c00000000000000cf00000000000000ed00000000000000cf00000000",
            INIT_4B => X"0000005d000000000000007d000000000000009400000000000000ae00000000",
            INIT_4C => X"0000004c000000000000003b000000000000004a000000000000005600000000",
            INIT_4D => X"0000006a0000000000000085000000000000008f000000000000008900000000",
            INIT_4E => X"0000004b00000000000000540000000000000057000000000000005600000000",
            INIT_4F => X"00000084000000000000005f0000000000000028000000000000003200000000",
            INIT_50 => X"000000a5000000000000008e000000000000006c00000000000000b700000000",
            INIT_51 => X"0000007a000000000000009f000000000000009b00000000000000b100000000",
            INIT_52 => X"000000a400000000000000dc00000000000000ed00000000000000d500000000",
            INIT_53 => X"00000078000000000000007d000000000000009c00000000000000b700000000",
            INIT_54 => X"0000005b000000000000002d0000000000000050000000000000004e00000000",
            INIT_55 => X"0000006b000000000000009b000000000000009d00000000000000af00000000",
            INIT_56 => X"0000004e00000000000000580000000000000067000000000000005700000000",
            INIT_57 => X"00000068000000000000003b0000000000000029000000000000003b00000000",
            INIT_58 => X"000000aa0000000000000087000000000000006400000000000000bc00000000",
            INIT_59 => X"0000008600000000000000ad00000000000000a600000000000000bb00000000",
            INIT_5A => X"000000aa00000000000000c700000000000000c2000000000000007500000000",
            INIT_5B => X"00000075000000000000008600000000000000bd00000000000000b900000000",
            INIT_5C => X"0000007d00000000000000260000000000000054000000000000006600000000",
            INIT_5D => X"0000005d000000000000009200000000000000a000000000000000d200000000",
            INIT_5E => X"000000550000000000000068000000000000005e000000000000005300000000",
            INIT_5F => X"0000004c000000000000003e0000000000000037000000000000004900000000",
            INIT_60 => X"000000af000000000000007f000000000000005a00000000000000bd00000000",
            INIT_61 => X"0000009f00000000000000b200000000000000a600000000000000ae00000000",
            INIT_62 => X"0000008900000000000000a800000000000000a8000000000000006100000000",
            INIT_63 => X"0000007b00000000000000a000000000000000d800000000000000ba00000000",
            INIT_64 => X"0000009600000000000000320000000000000073000000000000007800000000",
            INIT_65 => X"0000005b000000000000007b000000000000009b00000000000000c200000000",
            INIT_66 => X"00000056000000000000005f0000000000000054000000000000005400000000",
            INIT_67 => X"00000049000000000000004f0000000000000049000000000000005400000000",
            INIT_68 => X"000000b90000000000000098000000000000005d00000000000000bd00000000",
            INIT_69 => X"000000a700000000000000ad0000000000000088000000000000007700000000",
            INIT_6A => X"000000a700000000000000910000000000000093000000000000006700000000",
            INIT_6B => X"0000008d00000000000000b400000000000000e200000000000000bd00000000",
            INIT_6C => X"0000009a00000000000000470000000000000075000000000000007e00000000",
            INIT_6D => X"000000570000000000000072000000000000009500000000000000ba00000000",
            INIT_6E => X"0000006300000000000000500000000000000048000000000000005000000000",
            INIT_6F => X"0000005e0000000000000061000000000000005a000000000000006400000000",
            INIT_70 => X"000000ba00000000000000a8000000000000006c00000000000000c200000000",
            INIT_71 => X"000000a7000000000000009c0000000000000063000000000000006900000000",
            INIT_72 => X"000000c6000000000000008a0000000000000073000000000000006400000000",
            INIT_73 => X"0000009a000000000000009100000000000000ac00000000000000be00000000",
            INIT_74 => X"0000009800000000000000470000000000000067000000000000009200000000",
            INIT_75 => X"0000006e0000000000000082000000000000008900000000000000b300000000",
            INIT_76 => X"0000006d000000000000005f000000000000005b000000000000005500000000",
            INIT_77 => X"0000007500000000000000610000000000000064000000000000007300000000",
            INIT_78 => X"000000b800000000000000ac000000000000008400000000000000c500000000",
            INIT_79 => X"0000009b000000000000008c000000000000004e000000000000008200000000",
            INIT_7A => X"000000e6000000000000008f0000000000000082000000000000007300000000",
            INIT_7B => X"000000830000000000000087000000000000009100000000000000f200000000",
            INIT_7C => X"00000090000000000000005f000000000000006c000000000000007900000000",
            INIT_7D => X"000000570000000000000070000000000000009800000000000000a800000000",
            INIT_7E => X"0000007000000000000000690000000000000057000000000000004700000000",
            INIT_7F => X"0000008800000000000000790000000000000067000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "sampleifmap_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bf00000000000000a8000000000000009200000000000000cb00000000",
            INIT_01 => X"0000008a000000000000007e000000000000004e00000000000000a800000000",
            INIT_02 => X"000000ad000000000000009a0000000000000060000000000000008a00000000",
            INIT_03 => X"000000710000000000000071000000000000008c00000000000000a200000000",
            INIT_04 => X"000000ab00000000000000700000000000000069000000000000006500000000",
            INIT_05 => X"0000006d00000000000000870000000000000094000000000000009c00000000",
            INIT_06 => X"00000065000000000000005e000000000000004f000000000000004e00000000",
            INIT_07 => X"000000900000000000000097000000000000007d000000000000006b00000000",
            INIT_08 => X"000000b700000000000000a400000000000000a300000000000000d600000000",
            INIT_09 => X"0000009c0000000000000060000000000000005e00000000000000b000000000",
            INIT_0A => X"000000760000000000000081000000000000006a000000000000009400000000",
            INIT_0B => X"0000007300000000000000660000000000000074000000000000007200000000",
            INIT_0C => X"0000007600000000000000900000000000000065000000000000005600000000",
            INIT_0D => X"0000004b00000000000000850000000000000080000000000000004400000000",
            INIT_0E => X"000000660000000000000047000000000000003a000000000000003c00000000",
            INIT_0F => X"0000008c0000000000000096000000000000008f000000000000007400000000",
            INIT_10 => X"000000ad00000000000000a700000000000000b200000000000000d400000000",
            INIT_11 => X"0000008d0000000000000056000000000000007c00000000000000b000000000",
            INIT_12 => X"0000004d00000000000000680000000000000087000000000000009900000000",
            INIT_13 => X"000000930000000000000081000000000000007c000000000000008600000000",
            INIT_14 => X"000000840000000000000096000000000000005c000000000000005500000000",
            INIT_15 => X"00000040000000000000004b000000000000006b000000000000007500000000",
            INIT_16 => X"0000008500000000000000560000000000000041000000000000002c00000000",
            INIT_17 => X"00000097000000000000009a00000000000000a0000000000000009b00000000",
            INIT_18 => X"000000ae00000000000000ab00000000000000bb00000000000000c700000000",
            INIT_19 => X"000000770000000000000056000000000000009000000000000000b100000000",
            INIT_1A => X"0000004600000000000000900000000000000089000000000000007a00000000",
            INIT_1B => X"000000b80000000000000091000000000000006c000000000000008100000000",
            INIT_1C => X"0000008900000000000000830000000000000049000000000000007400000000",
            INIT_1D => X"0000003400000000000000330000000000000059000000000000008600000000",
            INIT_1E => X"000000a30000000000000079000000000000005a000000000000002f00000000",
            INIT_1F => X"00000095000000000000009e00000000000000a400000000000000ab00000000",
            INIT_20 => X"000000b100000000000000b300000000000000c300000000000000a500000000",
            INIT_21 => X"000000830000000000000063000000000000009800000000000000b500000000",
            INIT_22 => X"00000050000000000000005d000000000000006700000000000000ab00000000",
            INIT_23 => X"000000bf00000000000000b2000000000000007a000000000000005d00000000",
            INIT_24 => X"0000005700000000000000590000000000000064000000000000009600000000",
            INIT_25 => X"000000180000000000000026000000000000002e000000000000003c00000000",
            INIT_26 => X"00000090000000000000006c000000000000003c000000000000002e00000000",
            INIT_27 => X"00000078000000000000007f0000000000000080000000000000009000000000",
            INIT_28 => X"000000b200000000000000b100000000000000c3000000000000007500000000",
            INIT_29 => X"000000960000000000000053000000000000008a00000000000000b500000000",
            INIT_2A => X"00000086000000000000008500000000000000db00000000000000f500000000",
            INIT_2B => X"000000c200000000000000be00000000000000b0000000000000009500000000",
            INIT_2C => X"0000003d000000000000006e000000000000007d00000000000000a800000000",
            INIT_2D => X"0000003a00000000000000310000000000000022000000000000002300000000",
            INIT_2E => X"000000480000000000000045000000000000003a000000000000003d00000000",
            INIT_2F => X"00000037000000000000003b0000000000000045000000000000004e00000000",
            INIT_30 => X"000000b000000000000000ae00000000000000af000000000000004f00000000",
            INIT_31 => X"000000d3000000000000006d000000000000008c00000000000000b100000000",
            INIT_32 => X"0000007c00000000000000d000000000000000fc00000000000000fd00000000",
            INIT_33 => X"0000007a0000000000000074000000000000007c000000000000007200000000",
            INIT_34 => X"0000003c00000000000000440000000000000044000000000000006800000000",
            INIT_35 => X"0000003800000000000000330000000000000032000000000000003400000000",
            INIT_36 => X"00000033000000000000002b0000000000000033000000000000003800000000",
            INIT_37 => X"0000002a000000000000002b0000000000000030000000000000003b00000000",
            INIT_38 => X"000000a800000000000000900000000000000060000000000000002900000000",
            INIT_39 => X"000000f600000000000000a500000000000000a500000000000000b200000000",
            INIT_3A => X"0000003c000000000000006e00000000000000e300000000000000fd00000000",
            INIT_3B => X"0000003000000000000000310000000000000031000000000000003500000000",
            INIT_3C => X"0000002a000000000000002e000000000000002a000000000000002d00000000",
            INIT_3D => X"0000002b000000000000002e000000000000002e000000000000002600000000",
            INIT_3E => X"00000032000000000000002e000000000000002e000000000000002a00000000",
            INIT_3F => X"0000002d00000000000000330000000000000035000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000083000000000000003b000000000000001d000000000000001d00000000",
            INIT_41 => X"000000fe00000000000000c2000000000000008400000000000000a600000000",
            INIT_42 => X"00000032000000000000003d000000000000008d00000000000000f100000000",
            INIT_43 => X"0000003200000000000000310000000000000033000000000000003200000000",
            INIT_44 => X"000000220000000000000027000000000000002a000000000000002f00000000",
            INIT_45 => X"0000002a00000000000000260000000000000027000000000000002300000000",
            INIT_46 => X"0000003b000000000000003e0000000000000038000000000000002d00000000",
            INIT_47 => X"00000033000000000000002e0000000000000032000000000000003800000000",
            INIT_48 => X"000000490000000000000022000000000000001e000000000000003000000000",
            INIT_49 => X"0000010000000000000000d70000000000000080000000000000008000000000",
            INIT_4A => X"000000320000000000000036000000000000004200000000000000bb00000000",
            INIT_4B => X"0000002d000000000000002e0000000000000034000000000000003400000000",
            INIT_4C => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_4D => X"0000002e000000000000002b0000000000000028000000000000002800000000",
            INIT_4E => X"0000003b0000000000000040000000000000003e000000000000003b00000000",
            INIT_4F => X"0000005300000000000000460000000000000032000000000000003600000000",
            INIT_50 => X"00000029000000000000001f0000000000000023000000000000003400000000",
            INIT_51 => X"000000f000000000000000e00000000000000080000000000000004200000000",
            INIT_52 => X"000000380000000000000031000000000000003a000000000000007c00000000",
            INIT_53 => X"0000002f000000000000002c000000000000002c000000000000003600000000",
            INIT_54 => X"0000002c000000000000002b000000000000002b000000000000002e00000000",
            INIT_55 => X"0000003a0000000000000036000000000000002d000000000000002c00000000",
            INIT_56 => X"00000024000000000000002b000000000000002e000000000000003600000000",
            INIT_57 => X"0000004c00000000000000550000000000000049000000000000003300000000",
            INIT_58 => X"00000023000000000000001d0000000000000023000000000000003200000000",
            INIT_59 => X"000000d300000000000000ca000000000000004e000000000000002c00000000",
            INIT_5A => X"0000003000000000000000360000000000000041000000000000006100000000",
            INIT_5B => X"0000002d00000000000000280000000000000030000000000000003a00000000",
            INIT_5C => X"0000002e000000000000002f0000000000000030000000000000002f00000000",
            INIT_5D => X"0000003000000000000000270000000000000027000000000000003300000000",
            INIT_5E => X"00000028000000000000001c0000000000000027000000000000002f00000000",
            INIT_5F => X"00000033000000000000002e0000000000000043000000000000004300000000",
            INIT_60 => X"0000002100000000000000200000000000000023000000000000003200000000",
            INIT_61 => X"000000aa0000000000000068000000000000002e000000000000002900000000",
            INIT_62 => X"0000003500000000000000340000000000000036000000000000004000000000",
            INIT_63 => X"0000002d0000000000000036000000000000003a000000000000003d00000000",
            INIT_64 => X"00000031000000000000002e0000000000000029000000000000002a00000000",
            INIT_65 => X"000000270000000000000028000000000000002a000000000000002e00000000",
            INIT_66 => X"0000003f000000000000002c0000000000000028000000000000002500000000",
            INIT_67 => X"00000033000000000000000f000000000000001f000000000000002f00000000",
            INIT_68 => X"00000026000000000000001f000000000000002a000000000000004400000000",
            INIT_69 => X"00000047000000000000002a000000000000002b000000000000002500000000",
            INIT_6A => X"00000026000000000000001b000000000000001f000000000000003100000000",
            INIT_6B => X"00000035000000000000003a0000000000000038000000000000003100000000",
            INIT_6C => X"000000350000000000000039000000000000003c000000000000003800000000",
            INIT_6D => X"000000210000000000000027000000000000002d000000000000003200000000",
            INIT_6E => X"00000049000000000000004f000000000000003e000000000000002a00000000",
            INIT_6F => X"00000028000000000000000d0000000000000026000000000000003800000000",
            INIT_70 => X"0000002b00000000000000230000000000000031000000000000003d00000000",
            INIT_71 => X"00000028000000000000002c000000000000002a000000000000002700000000",
            INIT_72 => X"0000001e0000000000000017000000000000001b000000000000002a00000000",
            INIT_73 => X"0000002f0000000000000024000000000000001d000000000000001b00000000",
            INIT_74 => X"0000004b0000000000000042000000000000003e000000000000003800000000",
            INIT_75 => X"0000002b000000000000002b0000000000000031000000000000004500000000",
            INIT_76 => X"0000005d000000000000006d0000000000000055000000000000003c00000000",
            INIT_77 => X"00000014000000000000001d000000000000001a000000000000003c00000000",
            INIT_78 => X"0000002b000000000000002d0000000000000038000000000000003600000000",
            INIT_79 => X"0000002600000000000000280000000000000028000000000000002800000000",
            INIT_7A => X"0000001d0000000000000016000000000000001a000000000000002400000000",
            INIT_7B => X"000000120000000000000013000000000000001d000000000000001900000000",
            INIT_7C => X"0000004a000000000000003d000000000000002f000000000000002000000000",
            INIT_7D => X"0000002d00000000000000340000000000000035000000000000004200000000",
            INIT_7E => X"0000005900000000000000690000000000000059000000000000004300000000",
            INIT_7F => X"0000001500000000000000220000000000000018000000000000003000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "sampleifmap_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000760000000000000074000000000000006f000000000000007000000000",
            INIT_01 => X"000000710000000000000073000000000000006d000000000000007000000000",
            INIT_02 => X"0000006f00000000000000740000000000000071000000000000006f00000000",
            INIT_03 => X"0000007700000000000000750000000000000075000000000000006f00000000",
            INIT_04 => X"00000070000000000000006f0000000000000071000000000000007500000000",
            INIT_05 => X"0000006a000000000000006b000000000000006b000000000000006d00000000",
            INIT_06 => X"0000006100000000000000620000000000000065000000000000006b00000000",
            INIT_07 => X"00000055000000000000005b000000000000005f000000000000006100000000",
            INIT_08 => X"000000740000000000000072000000000000006e000000000000007000000000",
            INIT_09 => X"0000007200000000000000750000000000000071000000000000007000000000",
            INIT_0A => X"0000006e000000000000006f000000000000006e000000000000007400000000",
            INIT_0B => X"0000007300000000000000750000000000000077000000000000007100000000",
            INIT_0C => X"000000730000000000000070000000000000006f000000000000007300000000",
            INIT_0D => X"0000006400000000000000660000000000000068000000000000006e00000000",
            INIT_0E => X"0000006100000000000000660000000000000066000000000000006900000000",
            INIT_0F => X"00000058000000000000005b000000000000005f000000000000006200000000",
            INIT_10 => X"0000006f000000000000006f000000000000006d000000000000006e00000000",
            INIT_11 => X"0000007500000000000000750000000000000073000000000000006a00000000",
            INIT_12 => X"0000006d00000000000000720000000000000073000000000000007300000000",
            INIT_13 => X"0000007100000000000000720000000000000073000000000000006f00000000",
            INIT_14 => X"00000060000000000000006f0000000000000072000000000000007400000000",
            INIT_15 => X"00000055000000000000004d000000000000004e000000000000005a00000000",
            INIT_16 => X"0000006300000000000000670000000000000060000000000000005600000000",
            INIT_17 => X"00000059000000000000005f0000000000000062000000000000006300000000",
            INIT_18 => X"00000070000000000000006d000000000000006e000000000000006b00000000",
            INIT_19 => X"0000007700000000000000780000000000000075000000000000006e00000000",
            INIT_1A => X"00000092000000000000007b0000000000000075000000000000007300000000",
            INIT_1B => X"000000720000000000000073000000000000006f000000000000008200000000",
            INIT_1C => X"000000570000000000000050000000000000006f000000000000007000000000",
            INIT_1D => X"0000003f000000000000004b000000000000005a000000000000005a00000000",
            INIT_1E => X"000000620000000000000055000000000000003e000000000000004600000000",
            INIT_1F => X"0000005e00000000000000630000000000000065000000000000006600000000",
            INIT_20 => X"0000007200000000000000730000000000000072000000000000006b00000000",
            INIT_21 => X"0000007400000000000000780000000000000071000000000000007200000000",
            INIT_22 => X"000000d600000000000000800000000000000074000000000000007100000000",
            INIT_23 => X"0000006c000000000000006f0000000000000072000000000000009c00000000",
            INIT_24 => X"0000006700000000000000450000000000000035000000000000005000000000",
            INIT_25 => X"0000005e00000000000000660000000000000072000000000000006e00000000",
            INIT_26 => X"000000530000000000000049000000000000004e000000000000004800000000",
            INIT_27 => X"0000005d000000000000005e0000000000000065000000000000006000000000",
            INIT_28 => X"0000007000000000000000640000000000000068000000000000006d00000000",
            INIT_29 => X"0000007300000000000000740000000000000071000000000000007300000000",
            INIT_2A => X"0000008a00000000000000760000000000000074000000000000006f00000000",
            INIT_2B => X"00000032000000000000004b0000000000000066000000000000007a00000000",
            INIT_2C => X"0000007100000000000000530000000000000038000000000000003a00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007900000000",
            INIT_2E => X"0000003a000000000000003a000000000000005b000000000000006400000000",
            INIT_2F => X"0000005f00000000000000620000000000000069000000000000005400000000",
            INIT_30 => X"0000004a0000000000000025000000000000005f000000000000006400000000",
            INIT_31 => X"0000007600000000000000730000000000000076000000000000007500000000",
            INIT_32 => X"0000006b00000000000000780000000000000074000000000000007500000000",
            INIT_33 => X"000000430000000000000057000000000000006c000000000000006200000000",
            INIT_34 => X"000000820000000000000054000000000000004b000000000000005300000000",
            INIT_35 => X"0000006600000000000000630000000000000076000000000000008e00000000",
            INIT_36 => X"0000002f00000000000000470000000000000053000000000000006f00000000",
            INIT_37 => X"0000005d00000000000000630000000000000062000000000000003d00000000",
            INIT_38 => X"00000040000000000000002b0000000000000060000000000000007300000000",
            INIT_39 => X"0000007400000000000000720000000000000075000000000000006f00000000",
            INIT_3A => X"0000005e000000000000006d0000000000000071000000000000007700000000",
            INIT_3B => X"00000057000000000000006a0000000000000083000000000000006e00000000",
            INIT_3C => X"00000076000000000000004d0000000000000058000000000000005f00000000",
            INIT_3D => X"00000062000000000000005d000000000000007c000000000000009900000000",
            INIT_3E => X"00000035000000000000003c0000000000000051000000000000005d00000000",
            INIT_3F => X"0000006100000000000000670000000000000053000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000079000000000000003a000000000000006900000000000000a100000000",
            INIT_41 => X"0000007a00000000000000750000000000000071000000000000007c00000000",
            INIT_42 => X"0000006900000000000000590000000000000087000000000000007900000000",
            INIT_43 => X"00000050000000000000006f000000000000008f000000000000008d00000000",
            INIT_44 => X"00000047000000000000004e0000000000000055000000000000005100000000",
            INIT_45 => X"0000004f00000000000000670000000000000087000000000000007d00000000",
            INIT_46 => X"0000003900000000000000490000000000000052000000000000004d00000000",
            INIT_47 => X"00000067000000000000006a000000000000003b000000000000002300000000",
            INIT_48 => X"0000009a0000000000000064000000000000008b00000000000000b000000000",
            INIT_49 => X"0000007600000000000000740000000000000074000000000000009500000000",
            INIT_4A => X"0000008300000000000000b400000000000000d600000000000000b400000000",
            INIT_4B => X"00000055000000000000006e0000000000000083000000000000009900000000",
            INIT_4C => X"000000440000000000000039000000000000004a000000000000005400000000",
            INIT_4D => X"00000062000000000000007c0000000000000085000000000000007d00000000",
            INIT_4E => X"0000004c00000000000000550000000000000055000000000000005100000000",
            INIT_4F => X"00000067000000000000004b000000000000001e000000000000003100000000",
            INIT_50 => X"000000a90000000000000097000000000000007400000000000000b700000000",
            INIT_51 => X"0000005900000000000000760000000000000070000000000000009c00000000",
            INIT_52 => X"0000008700000000000000bf00000000000000e000000000000000c500000000",
            INIT_53 => X"0000006f000000000000006c0000000000000089000000000000009f00000000",
            INIT_54 => X"00000055000000000000002c0000000000000050000000000000004c00000000",
            INIT_55 => X"000000640000000000000093000000000000009300000000000000a500000000",
            INIT_56 => X"0000004f00000000000000580000000000000066000000000000005300000000",
            INIT_57 => X"00000051000000000000002e0000000000000024000000000000003b00000000",
            INIT_58 => X"000000af0000000000000090000000000000006c00000000000000bf00000000",
            INIT_59 => X"0000005d000000000000007b000000000000007800000000000000a700000000",
            INIT_5A => X"0000008e00000000000000ab00000000000000b6000000000000005f00000000",
            INIT_5B => X"0000006b000000000000007700000000000000ab00000000000000a100000000",
            INIT_5C => X"0000007900000000000000260000000000000054000000000000006200000000",
            INIT_5D => X"00000059000000000000008b000000000000009800000000000000c900000000",
            INIT_5E => X"000000570000000000000068000000000000005d000000000000005000000000",
            INIT_5F => X"0000003800000000000000370000000000000035000000000000004b00000000",
            INIT_60 => X"000000b40000000000000086000000000000006000000000000000c200000000",
            INIT_61 => X"0000006d000000000000007b000000000000007b000000000000009c00000000",
            INIT_62 => X"000000720000000000000090000000000000009a000000000000004400000000",
            INIT_63 => X"00000071000000000000009500000000000000ca00000000000000a600000000",
            INIT_64 => X"0000009300000000000000320000000000000072000000000000007200000000",
            INIT_65 => X"000000580000000000000076000000000000009500000000000000bb00000000",
            INIT_66 => X"00000057000000000000005f0000000000000054000000000000005300000000",
            INIT_67 => X"00000037000000000000004a0000000000000049000000000000005700000000",
            INIT_68 => X"000000bc000000000000009a000000000000005f00000000000000c000000000",
            INIT_69 => X"00000074000000000000007c000000000000006a000000000000006e00000000",
            INIT_6A => X"00000095000000000000007d0000000000000084000000000000004800000000",
            INIT_6B => X"0000008300000000000000ac00000000000000d800000000000000ae00000000",
            INIT_6C => X"0000009800000000000000470000000000000072000000000000007500000000",
            INIT_6D => X"00000055000000000000006e000000000000009000000000000000b500000000",
            INIT_6E => X"0000006400000000000000500000000000000049000000000000005000000000",
            INIT_6F => X"0000004900000000000000590000000000000058000000000000006500000000",
            INIT_70 => X"000000ba00000000000000a7000000000000006b00000000000000c400000000",
            INIT_71 => X"0000007a00000000000000770000000000000059000000000000006d00000000",
            INIT_72 => X"000000b9000000000000007b000000000000006a000000000000004a00000000",
            INIT_73 => X"0000008f000000000000008c00000000000000a500000000000000b400000000",
            INIT_74 => X"0000009800000000000000470000000000000064000000000000008800000000",
            INIT_75 => X"0000006d0000000000000080000000000000008500000000000000af00000000",
            INIT_76 => X"0000006e0000000000000060000000000000005d000000000000005600000000",
            INIT_77 => X"0000005f00000000000000550000000000000060000000000000007400000000",
            INIT_78 => X"000000b200000000000000a7000000000000008100000000000000c500000000",
            INIT_79 => X"0000007d00000000000000780000000000000053000000000000008900000000",
            INIT_7A => X"000000dd00000000000000830000000000000078000000000000005e00000000",
            INIT_7B => X"000000790000000000000082000000000000008a00000000000000ec00000000",
            INIT_7C => X"0000008600000000000000580000000000000068000000000000007000000000",
            INIT_7D => X"00000055000000000000006c0000000000000093000000000000009f00000000",
            INIT_7E => X"0000006d00000000000000680000000000000058000000000000004800000000",
            INIT_7F => X"0000006800000000000000600000000000000056000000000000006e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "sampleifmap_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000a4000000000000009200000000000000cb00000000",
            INIT_01 => X"0000007e000000000000007d000000000000005600000000000000aa00000000",
            INIT_02 => X"000000a3000000000000008f0000000000000050000000000000007900000000",
            INIT_03 => X"0000006a000000000000006a0000000000000084000000000000009800000000",
            INIT_04 => X"0000008f000000000000005a0000000000000065000000000000006500000000",
            INIT_05 => X"000000690000000000000082000000000000008d000000000000008a00000000",
            INIT_06 => X"0000005b000000000000005d000000000000004f000000000000004c00000000",
            INIT_07 => X"00000068000000000000006c0000000000000058000000000000005300000000",
            INIT_08 => X"000000b800000000000000a700000000000000a600000000000000d700000000",
            INIT_09 => X"000000950000000000000060000000000000006600000000000000b600000000",
            INIT_0A => X"000000690000000000000074000000000000005d000000000000008900000000",
            INIT_0B => X"0000006e000000000000005b0000000000000069000000000000006600000000",
            INIT_0C => X"0000006000000000000000800000000000000067000000000000005b00000000",
            INIT_0D => X"00000045000000000000007e0000000000000078000000000000003800000000",
            INIT_0E => X"0000005d00000000000000460000000000000038000000000000003800000000",
            INIT_0F => X"0000006e00000000000000740000000000000070000000000000005e00000000",
            INIT_10 => X"000000b500000000000000af00000000000000b800000000000000d300000000",
            INIT_11 => X"0000008b0000000000000058000000000000008300000000000000b800000000",
            INIT_12 => X"00000040000000000000005a0000000000000080000000000000009400000000",
            INIT_13 => X"0000008f0000000000000075000000000000006f000000000000007900000000",
            INIT_14 => X"00000075000000000000008b0000000000000060000000000000005c00000000",
            INIT_15 => X"0000003b00000000000000440000000000000063000000000000006d00000000",
            INIT_16 => X"000000690000000000000045000000000000003e000000000000002900000000",
            INIT_17 => X"0000006f00000000000000730000000000000078000000000000007700000000",
            INIT_18 => X"000000b300000000000000b000000000000000bd00000000000000c000000000",
            INIT_19 => X"00000079000000000000005a000000000000009500000000000000b600000000",
            INIT_1A => X"0000003b00000000000000860000000000000088000000000000007c00000000",
            INIT_1B => X"000000b000000000000000860000000000000061000000000000007600000000",
            INIT_1C => X"0000007c0000000000000077000000000000004b000000000000007600000000",
            INIT_1D => X"0000003300000000000000310000000000000056000000000000008100000000",
            INIT_1E => X"00000076000000000000005b000000000000005a000000000000003100000000",
            INIT_1F => X"0000006b000000000000006f0000000000000071000000000000007900000000",
            INIT_20 => X"000000ad00000000000000b200000000000000c1000000000000009c00000000",
            INIT_21 => X"000000870000000000000067000000000000009d00000000000000b500000000",
            INIT_22 => X"0000004d000000000000005a000000000000006900000000000000af00000000",
            INIT_23 => X"000000b600000000000000ad0000000000000076000000000000005a00000000",
            INIT_24 => X"0000004d000000000000004e0000000000000064000000000000009400000000",
            INIT_25 => X"00000021000000000000002e0000000000000034000000000000003d00000000",
            INIT_26 => X"0000007d00000000000000640000000000000047000000000000003900000000",
            INIT_27 => X"000000690000000000000071000000000000006d000000000000007b00000000",
            INIT_28 => X"000000a900000000000000b200000000000000c8000000000000007800000000",
            INIT_29 => X"000000990000000000000057000000000000009000000000000000b300000000",
            INIT_2A => X"0000008d000000000000008c00000000000000de00000000000000f700000000",
            INIT_2B => X"000000c000000000000000c400000000000000b6000000000000009c00000000",
            INIT_2C => X"0000003e000000000000006d000000000000008500000000000000ac00000000",
            INIT_2D => X"0000005100000000000000460000000000000036000000000000003100000000",
            INIT_2E => X"0000006500000000000000630000000000000054000000000000005500000000",
            INIT_2F => X"0000005a000000000000005c0000000000000060000000000000006800000000",
            INIT_30 => X"000000ac00000000000000b700000000000000c5000000000000006900000000",
            INIT_31 => X"000000d30000000000000070000000000000009200000000000000b100000000",
            INIT_32 => X"0000008f00000000000000e000000000000000fd00000000000000fc00000000",
            INIT_33 => X"000000850000000000000085000000000000008d000000000000008400000000",
            INIT_34 => X"000000520000000000000057000000000000005d000000000000007c00000000",
            INIT_35 => X"0000005d00000000000000550000000000000054000000000000005400000000",
            INIT_36 => X"000000680000000000000060000000000000005b000000000000005e00000000",
            INIT_37 => X"0000005f00000000000000610000000000000061000000000000006c00000000",
            INIT_38 => X"000000ae00000000000000a80000000000000089000000000000005900000000",
            INIT_39 => X"000000f500000000000000a600000000000000aa00000000000000b600000000",
            INIT_3A => X"00000058000000000000008800000000000000e700000000000000fb00000000",
            INIT_3B => X"00000048000000000000004b000000000000004c000000000000005000000000",
            INIT_3C => X"0000005200000000000000510000000000000051000000000000004f00000000",
            INIT_3D => X"000000570000000000000059000000000000005a000000000000005600000000",
            INIT_3E => X"00000060000000000000005e000000000000005d000000000000005900000000",
            INIT_3F => X"0000005a000000000000005f000000000000005e000000000000006000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009900000000000000660000000000000057000000000000005b00000000",
            INIT_41 => X"000000fa00000000000000bd000000000000008800000000000000b300000000",
            INIT_42 => X"00000054000000000000005e000000000000009f00000000000000f500000000",
            INIT_43 => X"0000005400000000000000530000000000000055000000000000005400000000",
            INIT_44 => X"0000004f00000000000000520000000000000054000000000000005600000000",
            INIT_45 => X"0000005900000000000000550000000000000056000000000000005300000000",
            INIT_46 => X"0000006500000000000000670000000000000067000000000000005c00000000",
            INIT_47 => X"00000067000000000000005e0000000000000063000000000000006600000000",
            INIT_48 => X"0000006a0000000000000055000000000000005e000000000000006f00000000",
            INIT_49 => X"000000fd00000000000000d50000000000000088000000000000009400000000",
            INIT_4A => X"00000058000000000000005b000000000000005d00000000000000c600000000",
            INIT_4B => X"000000520000000000000053000000000000005a000000000000005a00000000",
            INIT_4C => X"0000005300000000000000500000000000000051000000000000005200000000",
            INIT_4D => X"0000005f000000000000005c0000000000000059000000000000005600000000",
            INIT_4E => X"0000006c000000000000006d000000000000006e000000000000006c00000000",
            INIT_4F => X"00000089000000000000007b0000000000000069000000000000006c00000000",
            INIT_50 => X"0000005300000000000000560000000000000063000000000000007200000000",
            INIT_51 => X"000000f500000000000000e50000000000000091000000000000005f00000000",
            INIT_52 => X"0000005e0000000000000057000000000000005c000000000000008f00000000",
            INIT_53 => X"0000005300000000000000520000000000000052000000000000005c00000000",
            INIT_54 => X"0000005800000000000000560000000000000053000000000000005400000000",
            INIT_55 => X"0000006e000000000000006a0000000000000061000000000000005a00000000",
            INIT_56 => X"0000005b000000000000005f0000000000000061000000000000006900000000",
            INIT_57 => X"0000007d000000000000008a0000000000000082000000000000006c00000000",
            INIT_58 => X"0000005600000000000000590000000000000062000000000000006e00000000",
            INIT_59 => X"000000e400000000000000db000000000000006a000000000000005300000000",
            INIT_5A => X"00000057000000000000005e0000000000000068000000000000007e00000000",
            INIT_5B => X"0000005200000000000000500000000000000057000000000000006100000000",
            INIT_5C => X"0000005900000000000000590000000000000057000000000000005400000000",
            INIT_5D => X"00000066000000000000005d000000000000005c000000000000006100000000",
            INIT_5E => X"000000650000000000000055000000000000005d000000000000006500000000",
            INIT_5F => X"000000600000000000000062000000000000007e000000000000008100000000",
            INIT_60 => X"00000058000000000000005c0000000000000061000000000000006c00000000",
            INIT_61 => X"000000c500000000000000850000000000000054000000000000005800000000",
            INIT_62 => X"0000005f000000000000005e0000000000000061000000000000006400000000",
            INIT_63 => X"0000005300000000000000600000000000000064000000000000006700000000",
            INIT_64 => X"0000005c00000000000000580000000000000050000000000000004f00000000",
            INIT_65 => X"0000005c000000000000005d000000000000005f000000000000005c00000000",
            INIT_66 => X"0000007d0000000000000066000000000000005d000000000000005a00000000",
            INIT_67 => X"0000005d000000000000003c000000000000005a000000000000006e00000000",
            INIT_68 => X"0000005b00000000000000580000000000000064000000000000007c00000000",
            INIT_69 => X"0000006b000000000000004f0000000000000059000000000000005700000000",
            INIT_6A => X"000000520000000000000047000000000000004d000000000000005900000000",
            INIT_6B => X"0000005c00000000000000660000000000000064000000000000005d00000000",
            INIT_6C => X"0000006100000000000000630000000000000063000000000000005e00000000",
            INIT_6D => X"000000530000000000000058000000000000005e000000000000005f00000000",
            INIT_6E => X"0000008300000000000000840000000000000070000000000000005b00000000",
            INIT_6F => X"0000005500000000000000400000000000000061000000000000007400000000",
            INIT_70 => X"0000005b00000000000000550000000000000066000000000000007400000000",
            INIT_71 => X"000000510000000000000058000000000000005c000000000000005a00000000",
            INIT_72 => X"0000004a00000000000000430000000000000048000000000000005500000000",
            INIT_73 => X"0000005600000000000000500000000000000049000000000000004700000000",
            INIT_74 => X"00000077000000000000006d0000000000000065000000000000005f00000000",
            INIT_75 => X"000000580000000000000058000000000000005f000000000000007100000000",
            INIT_76 => X"00000091000000000000009c0000000000000082000000000000006900000000",
            INIT_77 => X"0000004000000000000000520000000000000052000000000000007300000000",
            INIT_78 => X"0000005600000000000000590000000000000069000000000000006b00000000",
            INIT_79 => X"000000510000000000000057000000000000005c000000000000005900000000",
            INIT_7A => X"0000004900000000000000420000000000000045000000000000004f00000000",
            INIT_7B => X"0000003a000000000000003f0000000000000049000000000000004500000000",
            INIT_7C => X"0000007700000000000000680000000000000057000000000000004600000000",
            INIT_7D => X"00000057000000000000005f0000000000000060000000000000006f00000000",
            INIT_7E => X"0000008700000000000000920000000000000083000000000000006d00000000",
            INIT_7F => X"000000430000000000000054000000000000004d000000000000006300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "sampleifmap_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000350000000000000033000000000000002f000000000000003100000000",
            INIT_01 => X"0000002d000000000000002f0000000000000029000000000000002e00000000",
            INIT_02 => X"0000003400000000000000290000000000000029000000000000002c00000000",
            INIT_03 => X"0000002c000000000000002d0000000000000029000000000000003100000000",
            INIT_04 => X"0000002b00000000000000270000000000000026000000000000002800000000",
            INIT_05 => X"0000002b000000000000002d000000000000002d000000000000002c00000000",
            INIT_06 => X"00000029000000000000002b0000000000000027000000000000002c00000000",
            INIT_07 => X"0000002100000000000000240000000000000024000000000000002600000000",
            INIT_08 => X"00000038000000000000002d0000000000000028000000000000003300000000",
            INIT_09 => X"0000002d000000000000002f000000000000002b000000000000003100000000",
            INIT_0A => X"0000003600000000000000290000000000000026000000000000002e00000000",
            INIT_0B => X"0000002100000000000000280000000000000029000000000000003400000000",
            INIT_0C => X"0000003200000000000000290000000000000021000000000000001e00000000",
            INIT_0D => X"0000003000000000000000340000000000000037000000000000003500000000",
            INIT_0E => X"00000026000000000000002d000000000000002e000000000000003200000000",
            INIT_0F => X"000000220000000000000020000000000000001f000000000000002200000000",
            INIT_10 => X"0000003000000000000000240000000000000021000000000000002f00000000",
            INIT_11 => X"0000002d000000000000002d000000000000002c000000000000002a00000000",
            INIT_12 => X"000000390000000000000030000000000000002b000000000000002b00000000",
            INIT_13 => X"0000002300000000000000250000000000000026000000000000003300000000",
            INIT_14 => X"000000310000000000000036000000000000002f000000000000002700000000",
            INIT_15 => X"00000032000000000000002f0000000000000032000000000000003400000000",
            INIT_16 => X"0000002700000000000000330000000000000037000000000000003000000000",
            INIT_17 => X"0000002100000000000000220000000000000022000000000000002300000000",
            INIT_18 => X"0000002c000000000000001f0000000000000020000000000000002800000000",
            INIT_19 => X"000000300000000000000030000000000000002e000000000000002b00000000",
            INIT_1A => X"0000005f0000000000000039000000000000002d000000000000002c00000000",
            INIT_1B => X"00000036000000000000002f0000000000000029000000000000004b00000000",
            INIT_1C => X"00000041000000000000002f0000000000000043000000000000003a00000000",
            INIT_1D => X"0000003200000000000000420000000000000054000000000000004c00000000",
            INIT_1E => X"0000002e000000000000002d0000000000000027000000000000003400000000",
            INIT_1F => X"0000002400000000000000270000000000000027000000000000002b00000000",
            INIT_20 => X"0000002f00000000000000310000000000000030000000000000002900000000",
            INIT_21 => X"0000002c000000000000002f0000000000000028000000000000002b00000000",
            INIT_22 => X"000000a4000000000000003b000000000000002a000000000000002900000000",
            INIT_23 => X"00000047000000000000003c0000000000000038000000000000006b00000000",
            INIT_24 => X"000000620000000000000038000000000000001f000000000000003200000000",
            INIT_25 => X"0000005d00000000000000690000000000000076000000000000006f00000000",
            INIT_26 => X"0000002d000000000000002f0000000000000046000000000000004300000000",
            INIT_27 => X"000000240000000000000024000000000000002e000000000000003000000000",
            INIT_28 => X"0000003500000000000000390000000000000040000000000000003600000000",
            INIT_29 => X"0000002900000000000000290000000000000027000000000000002c00000000",
            INIT_2A => X"00000055000000000000002a0000000000000027000000000000002500000000",
            INIT_2B => X"0000001f000000000000002b000000000000003a000000000000004e00000000",
            INIT_2C => X"0000006e000000000000004c000000000000002d000000000000002b00000000",
            INIT_2D => X"000000600000000000000074000000000000007a000000000000007800000000",
            INIT_2E => X"00000025000000000000002f0000000000000056000000000000006100000000",
            INIT_2F => X"00000028000000000000002c000000000000003a000000000000003100000000",
            INIT_30 => X"0000001c00000000000000110000000000000050000000000000003900000000",
            INIT_31 => X"0000002b0000000000000028000000000000002b000000000000003000000000",
            INIT_32 => X"0000003400000000000000270000000000000025000000000000002a00000000",
            INIT_33 => X"000000390000000000000046000000000000004b000000000000003b00000000",
            INIT_34 => X"00000079000000000000004a0000000000000040000000000000004800000000",
            INIT_35 => X"0000005e000000000000005a000000000000006c000000000000008400000000",
            INIT_36 => X"000000270000000000000045000000000000004d000000000000006700000000",
            INIT_37 => X"000000270000000000000030000000000000003a000000000000002400000000",
            INIT_38 => X"000000290000000000000026000000000000005c000000000000005a00000000",
            INIT_39 => X"000000270000000000000024000000000000002a000000000000003800000000",
            INIT_3A => X"0000003100000000000000330000000000000033000000000000003100000000",
            INIT_3B => X"0000004f000000000000005d000000000000006b000000000000004d00000000",
            INIT_3C => X"0000006b00000000000000450000000000000052000000000000005800000000",
            INIT_3D => X"0000005800000000000000510000000000000070000000000000008c00000000",
            INIT_3E => X"00000031000000000000003a000000000000004a000000000000005400000000",
            INIT_3F => X"0000002700000000000000330000000000000032000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000071000000000000003b0000000000000069000000000000009000000000",
            INIT_41 => X"000000320000000000000029000000000000002b000000000000005200000000",
            INIT_42 => X"0000004e000000000000003b000000000000005f000000000000004200000000",
            INIT_43 => X"0000004a00000000000000650000000000000080000000000000007900000000",
            INIT_44 => X"0000003d00000000000000490000000000000052000000000000004d00000000",
            INIT_45 => X"00000046000000000000005d000000000000007b000000000000007000000000",
            INIT_46 => X"000000350000000000000043000000000000004c000000000000004500000000",
            INIT_47 => X"0000002d000000000000003b0000000000000023000000000000001b00000000",
            INIT_48 => X"000000950000000000000069000000000000008f00000000000000a300000000",
            INIT_49 => X"0000003c000000000000002f0000000000000033000000000000007000000000",
            INIT_4A => X"0000007700000000000000a600000000000000c6000000000000009200000000",
            INIT_4B => X"0000004f000000000000006b000000000000007d000000000000009100000000",
            INIT_4C => X"0000003a00000000000000350000000000000047000000000000004f00000000",
            INIT_4D => X"000000590000000000000072000000000000007a000000000000007000000000",
            INIT_4E => X"00000047000000000000004e000000000000004e000000000000004a00000000",
            INIT_4F => X"00000039000000000000002c000000000000000f000000000000002b00000000",
            INIT_50 => X"000000a8000000000000009e000000000000007a00000000000000af00000000",
            INIT_51 => X"0000002f00000000000000330000000000000032000000000000007a00000000",
            INIT_52 => X"0000008300000000000000bc00000000000000e200000000000000b300000000",
            INIT_53 => X"0000006800000000000000680000000000000084000000000000009b00000000",
            INIT_54 => X"0000004d0000000000000028000000000000004d000000000000004500000000",
            INIT_55 => X"0000005c000000000000008a0000000000000089000000000000009a00000000",
            INIT_56 => X"00000049000000000000004f0000000000000060000000000000004d00000000",
            INIT_57 => X"0000002e000000000000001f0000000000000021000000000000003b00000000",
            INIT_58 => X"000000b20000000000000099000000000000007400000000000000bd00000000",
            INIT_59 => X"0000002c0000000000000037000000000000003b000000000000008800000000",
            INIT_5A => X"0000008500000000000000a400000000000000bc000000000000005000000000",
            INIT_5B => X"0000005f000000000000006a000000000000009f000000000000009700000000",
            INIT_5C => X"000000710000000000000022000000000000004f000000000000005900000000",
            INIT_5D => X"000000520000000000000082000000000000008e00000000000000c000000000",
            INIT_5E => X"00000051000000000000005e0000000000000058000000000000004b00000000",
            INIT_5F => X"0000001a00000000000000300000000000000037000000000000004e00000000",
            INIT_60 => X"000000b90000000000000090000000000000006900000000000000c200000000",
            INIT_61 => X"0000002f00000000000000350000000000000044000000000000008500000000",
            INIT_62 => X"0000005e000000000000007e0000000000000098000000000000002c00000000",
            INIT_63 => X"00000062000000000000008100000000000000b7000000000000009400000000",
            INIT_64 => X"0000008c000000000000002f000000000000006d000000000000006900000000",
            INIT_65 => X"00000053000000000000006f000000000000008c00000000000000b200000000",
            INIT_66 => X"0000005100000000000000550000000000000050000000000000004f00000000",
            INIT_67 => X"0000001800000000000000400000000000000049000000000000005900000000",
            INIT_68 => X"000000c000000000000000a3000000000000006700000000000000c100000000",
            INIT_69 => X"00000032000000000000003a0000000000000042000000000000006200000000",
            INIT_6A => X"0000007f00000000000000670000000000000078000000000000002700000000",
            INIT_6B => X"00000075000000000000009d00000000000000c8000000000000009b00000000",
            INIT_6C => X"000000930000000000000044000000000000006d000000000000006b00000000",
            INIT_6D => X"000000500000000000000068000000000000008800000000000000ae00000000",
            INIT_6E => X"0000005e00000000000000480000000000000046000000000000004c00000000",
            INIT_6F => X"0000002200000000000000450000000000000051000000000000006300000000",
            INIT_70 => X"000000bc00000000000000ac000000000000007000000000000000c400000000",
            INIT_71 => X"00000037000000000000003e0000000000000043000000000000006d00000000",
            INIT_72 => X"000000a900000000000000670000000000000058000000000000002200000000",
            INIT_73 => X"00000086000000000000008c000000000000009f00000000000000a900000000",
            INIT_74 => X"000000950000000000000046000000000000005f000000000000007d00000000",
            INIT_75 => X"00000069000000000000007a000000000000007f00000000000000aa00000000",
            INIT_76 => X"00000068000000000000005a000000000000005b000000000000005300000000",
            INIT_77 => X"0000002f00000000000000350000000000000050000000000000006f00000000",
            INIT_78 => X"000000b500000000000000ae000000000000008800000000000000c500000000",
            INIT_79 => X"0000004d0000000000000058000000000000004d000000000000008e00000000",
            INIT_7A => X"000000d30000000000000074000000000000005d000000000000003400000000",
            INIT_7B => X"000000700000000000000082000000000000008900000000000000e600000000",
            INIT_7C => X"00000076000000000000004b000000000000005f000000000000006500000000",
            INIT_7D => X"000000500000000000000065000000000000008a000000000000009200000000",
            INIT_7E => X"0000006300000000000000630000000000000057000000000000004400000000",
            INIT_7F => X"0000003000000000000000300000000000000036000000000000005d00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "sampleifmap_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000bc00000000000000b200000000000000a000000000000000cc00000000",
            INIT_01 => X"00000071000000000000007e000000000000005a00000000000000ac00000000",
            INIT_02 => X"0000009b00000000000000850000000000000025000000000000005200000000",
            INIT_03 => X"0000005a00000000000000580000000000000075000000000000008d00000000",
            INIT_04 => X"00000068000000000000003a0000000000000057000000000000005c00000000",
            INIT_05 => X"000000610000000000000076000000000000007e000000000000006d00000000",
            INIT_06 => X"00000052000000000000005e000000000000004d000000000000004800000000",
            INIT_07 => X"0000002e0000000000000037000000000000002d000000000000003700000000",
            INIT_08 => X"000000c200000000000000b800000000000000b400000000000000d700000000",
            INIT_09 => X"000000910000000000000066000000000000006900000000000000ba00000000",
            INIT_0A => X"0000005f0000000000000069000000000000003d000000000000006f00000000",
            INIT_0B => X"0000006200000000000000490000000000000059000000000000005900000000",
            INIT_0C => X"000000400000000000000066000000000000005f000000000000005800000000",
            INIT_0D => X"0000003d00000000000000730000000000000069000000000000002000000000",
            INIT_0E => X"0000004e00000000000000410000000000000035000000000000003300000000",
            INIT_0F => X"0000003600000000000000400000000000000044000000000000004000000000",
            INIT_10 => X"000000c100000000000000bd00000000000000c000000000000000cd00000000",
            INIT_11 => X"0000008f0000000000000060000000000000008500000000000000bc00000000",
            INIT_12 => X"000000370000000000000050000000000000006f000000000000008d00000000",
            INIT_13 => X"0000008500000000000000640000000000000060000000000000006c00000000",
            INIT_14 => X"0000005d0000000000000078000000000000005d000000000000005d00000000",
            INIT_15 => X"00000034000000000000003a0000000000000056000000000000005c00000000",
            INIT_16 => X"0000003b0000000000000028000000000000003c000000000000002700000000",
            INIT_17 => X"0000002e000000000000002d0000000000000036000000000000003e00000000",
            INIT_18 => X"000000b900000000000000b500000000000000bb00000000000000b400000000",
            INIT_19 => X"000000840000000000000063000000000000009800000000000000b800000000",
            INIT_1A => X"00000033000000000000007e0000000000000087000000000000008200000000",
            INIT_1B => X"000000a8000000000000007b0000000000000056000000000000006c00000000",
            INIT_1C => X"0000006900000000000000670000000000000049000000000000007600000000",
            INIT_1D => X"00000032000000000000002c000000000000004e000000000000007600000000",
            INIT_1E => X"00000044000000000000003c000000000000005d000000000000003400000000",
            INIT_1F => X"0000002e00000000000000320000000000000034000000000000004000000000",
            INIT_20 => X"000000ac00000000000000af00000000000000bb000000000000009200000000",
            INIT_21 => X"00000092000000000000006f00000000000000a000000000000000b400000000",
            INIT_22 => X"000000490000000000000057000000000000006f00000000000000b900000000",
            INIT_23 => X"000000b100000000000000ad0000000000000074000000000000005600000000",
            INIT_24 => X"0000003f00000000000000420000000000000065000000000000009400000000",
            INIT_25 => X"0000002900000000000000330000000000000036000000000000003900000000",
            INIT_26 => X"00000052000000000000004b0000000000000053000000000000004500000000",
            INIT_27 => X"0000003f0000000000000045000000000000003d000000000000004c00000000",
            INIT_28 => X"000000a800000000000000b000000000000000c8000000000000007c00000000",
            INIT_29 => X"0000009f000000000000005b000000000000009300000000000000b300000000",
            INIT_2A => X"00000093000000000000009000000000000000e100000000000000fa00000000",
            INIT_2B => X"000000c500000000000000d000000000000000c000000000000000a400000000",
            INIT_2C => X"0000003e000000000000006d000000000000008f00000000000000b500000000",
            INIT_2D => X"0000006600000000000000570000000000000044000000000000003a00000000",
            INIT_2E => X"00000077000000000000007a000000000000006f000000000000006e00000000",
            INIT_2F => X"0000007300000000000000700000000000000070000000000000007800000000",
            INIT_30 => X"000000b100000000000000c000000000000000d5000000000000008500000000",
            INIT_31 => X"000000d10000000000000071000000000000009600000000000000b600000000",
            INIT_32 => X"0000009d00000000000000e800000000000000fc00000000000000f700000000",
            INIT_33 => X"00000098000000000000009c00000000000000a2000000000000009500000000",
            INIT_34 => X"0000006500000000000000680000000000000077000000000000009400000000",
            INIT_35 => X"0000007d0000000000000073000000000000006e000000000000006f00000000",
            INIT_36 => X"0000008d00000000000000870000000000000082000000000000008300000000",
            INIT_37 => X"0000008400000000000000890000000000000084000000000000008e00000000",
            INIT_38 => X"000000bc00000000000000bc00000000000000a8000000000000008700000000",
            INIT_39 => X"000000ed00000000000000a400000000000000ae00000000000000c000000000",
            INIT_3A => X"0000006f000000000000009900000000000000e400000000000000f100000000",
            INIT_3B => X"00000065000000000000006b0000000000000069000000000000006900000000",
            INIT_3C => X"0000007400000000000000710000000000000078000000000000007300000000",
            INIT_3D => X"00000080000000000000007e000000000000007d000000000000007d00000000",
            INIT_3E => X"000000890000000000000089000000000000008b000000000000008400000000",
            INIT_3F => X"00000085000000000000008b0000000000000086000000000000008700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b000000000000000860000000000000082000000000000008d00000000",
            INIT_41 => X"000000f200000000000000b5000000000000008900000000000000bf00000000",
            INIT_42 => X"00000076000000000000007f00000000000000af00000000000000f500000000",
            INIT_43 => X"0000007400000000000000780000000000000079000000000000007700000000",
            INIT_44 => X"0000007100000000000000730000000000000075000000000000007500000000",
            INIT_45 => X"00000082000000000000007d000000000000007d000000000000007800000000",
            INIT_46 => X"0000008e000000000000008e0000000000000091000000000000008600000000",
            INIT_47 => X"00000095000000000000008c0000000000000090000000000000009200000000",
            INIT_48 => X"00000088000000000000007c000000000000008c00000000000000a200000000",
            INIT_49 => X"000000f900000000000000d1000000000000008f00000000000000a700000000",
            INIT_4A => X"0000007d0000000000000080000000000000007600000000000000cd00000000",
            INIT_4B => X"000000730000000000000079000000000000007f000000000000007f00000000",
            INIT_4C => X"0000007500000000000000710000000000000070000000000000007100000000",
            INIT_4D => X"0000008a00000000000000860000000000000083000000000000007b00000000",
            INIT_4E => X"0000009500000000000000930000000000000098000000000000009600000000",
            INIT_4F => X"000000b600000000000000a70000000000000098000000000000009a00000000",
            INIT_50 => X"0000007a0000000000000082000000000000009300000000000000a500000000",
            INIT_51 => X"000000f700000000000000ea00000000000000a4000000000000007e00000000",
            INIT_52 => X"00000083000000000000007b0000000000000072000000000000009900000000",
            INIT_53 => X"0000007700000000000000770000000000000077000000000000008100000000",
            INIT_54 => X"0000007f000000000000007b0000000000000077000000000000007700000000",
            INIT_55 => X"0000009a0000000000000096000000000000008d000000000000008300000000",
            INIT_56 => X"0000008a000000000000008c000000000000008d000000000000009600000000",
            INIT_57 => X"000000a900000000000000b600000000000000b2000000000000009e00000000",
            INIT_58 => X"00000085000000000000008a000000000000009500000000000000a200000000",
            INIT_59 => X"000000ea00000000000000e9000000000000008a000000000000007e00000000",
            INIT_5A => X"0000007c0000000000000081000000000000007e000000000000008c00000000",
            INIT_5B => X"000000770000000000000074000000000000007b000000000000008500000000",
            INIT_5C => X"000000840000000000000082000000000000007e000000000000007a00000000",
            INIT_5D => X"00000094000000000000008b000000000000008a000000000000008c00000000",
            INIT_5E => X"000000990000000000000085000000000000008b000000000000009300000000",
            INIT_5F => X"0000008b000000000000008e00000000000000b000000000000000b600000000",
            INIT_60 => X"0000008d000000000000008f000000000000009300000000000000a100000000",
            INIT_61 => X"000000d3000000000000009f000000000000007d000000000000008a00000000",
            INIT_62 => X"0000008200000000000000800000000000000079000000000000007700000000",
            INIT_63 => X"0000007800000000000000830000000000000087000000000000008b00000000",
            INIT_64 => X"0000008700000000000000820000000000000078000000000000007600000000",
            INIT_65 => X"00000088000000000000008a000000000000008b000000000000008800000000",
            INIT_66 => X"000000b20000000000000097000000000000008a000000000000008700000000",
            INIT_67 => X"000000880000000000000067000000000000008c00000000000000a400000000",
            INIT_68 => X"000000920000000000000089000000000000009400000000000000b100000000",
            INIT_69 => X"0000008500000000000000710000000000000084000000000000008b00000000",
            INIT_6A => X"0000007500000000000000690000000000000069000000000000007200000000",
            INIT_6B => X"0000008000000000000000890000000000000087000000000000008000000000",
            INIT_6C => X"0000008a000000000000008b0000000000000089000000000000008300000000",
            INIT_6D => X"0000007d00000000000000830000000000000088000000000000008900000000",
            INIT_6E => X"000000b500000000000000b3000000000000009a000000000000008500000000",
            INIT_6F => X"0000007f000000000000006c000000000000009200000000000000a800000000",
            INIT_70 => X"0000008f0000000000000084000000000000009400000000000000a800000000",
            INIT_71 => X"00000070000000000000007d0000000000000086000000000000008b00000000",
            INIT_72 => X"0000006d00000000000000660000000000000068000000000000007300000000",
            INIT_73 => X"000000780000000000000073000000000000006c000000000000006a00000000",
            INIT_74 => X"0000009c00000000000000900000000000000087000000000000008000000000",
            INIT_75 => X"0000007f000000000000007f0000000000000086000000000000009800000000",
            INIT_76 => X"000000be00000000000000c500000000000000aa000000000000009000000000",
            INIT_77 => X"0000006b000000000000007e000000000000008200000000000000a400000000",
            INIT_78 => X"000000860000000000000084000000000000009500000000000000a000000000",
            INIT_79 => X"00000073000000000000007b0000000000000084000000000000008600000000",
            INIT_7A => X"0000006c00000000000000650000000000000069000000000000007200000000",
            INIT_7B => X"000000590000000000000062000000000000006c000000000000006800000000",
            INIT_7C => X"0000009800000000000000890000000000000076000000000000006400000000",
            INIT_7D => X"0000007b00000000000000820000000000000083000000000000009100000000",
            INIT_7E => X"000000af00000000000000b600000000000000a7000000000000009100000000",
            INIT_7F => X"0000006e0000000000000081000000000000007c000000000000009100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "sampleifmap_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e600000000000000e700000000000000e800000000000000e900000000",
            INIT_05 => X"000000e900000000000000e800000000000000e800000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e800000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ec00000000000000ec00000000000000ed00000000",
            INIT_0D => X"000000ec00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ea00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_15 => X"000000ea00000000000000e700000000000000e700000000000000e300000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000df00000000000000e400000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000cf00000000000000d100000000000000ba00000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000ec00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000cb00000000000000db00000000000000e900000000000000ec00000000",
            INIT_25 => X"000000e600000000000000d600000000000000c300000000000000a300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_28 => X"000000ec00000000000000ec00000000000000ec00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_2A => X"000000ed00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e500000000000000eb00000000000000e800000000000000ea00000000",
            INIT_2C => X"000000ae00000000000000b900000000000000c200000000000000d000000000",
            INIT_2D => X"000000e200000000000000cf00000000000000b800000000000000a500000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e700000000000000e800000000000000e400000000000000e400000000",
            INIT_31 => X"000000ec00000000000000ed00000000000000ed00000000000000ea00000000",
            INIT_32 => X"000000ef00000000000000ef00000000000000ed00000000000000ed00000000",
            INIT_33 => X"000000dd00000000000000e900000000000000e000000000000000e100000000",
            INIT_34 => X"0000009a000000000000009f00000000000000a100000000000000b700000000",
            INIT_35 => X"000000c6000000000000009c000000000000008f000000000000009000000000",
            INIT_36 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_37 => X"000000ef00000000000000ed00000000000000ec00000000000000eb00000000",
            INIT_38 => X"000000e300000000000000e600000000000000e000000000000000d400000000",
            INIT_39 => X"000000ee00000000000000ed00000000000000ea00000000000000e500000000",
            INIT_3A => X"000000f000000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_3B => X"000000d600000000000000e900000000000000db00000000000000c900000000",
            INIT_3C => X"000000ad00000000000000b800000000000000b900000000000000c100000000",
            INIT_3D => X"000000ba00000000000000a2000000000000009f00000000000000a500000000",
            INIT_3E => X"000000e900000000000000e900000000000000ea00000000000000e500000000",
            INIT_3F => X"000000ee00000000000000ed00000000000000ec00000000000000ea00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000e100000000000000e100000000000000dd00000000000000d800000000",
            INIT_41 => X"000000ee00000000000000ec00000000000000e700000000000000e300000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_43 => X"000000e600000000000000e900000000000000dc00000000000000c500000000",
            INIT_44 => X"000000d000000000000000db00000000000000d100000000000000d100000000",
            INIT_45 => X"000000da00000000000000d900000000000000d200000000000000d100000000",
            INIT_46 => X"000000e600000000000000e400000000000000e400000000000000e100000000",
            INIT_47 => X"000000ee00000000000000ed00000000000000eb00000000000000e600000000",
            INIT_48 => X"00000088000000000000007c0000000000000077000000000000007600000000",
            INIT_49 => X"000000ed00000000000000eb00000000000000e100000000000000ac00000000",
            INIT_4A => X"000000e900000000000000eb00000000000000eb00000000000000ec00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000e100000000000000e700000000000000e300000000000000e400000000",
            INIT_4D => X"000000b900000000000000c900000000000000d900000000000000e100000000",
            INIT_4E => X"000000ba00000000000000a700000000000000a700000000000000ac00000000",
            INIT_4F => X"000000ee00000000000000ec00000000000000eb00000000000000df00000000",
            INIT_50 => X"0000006f000000000000006c0000000000000067000000000000006d00000000",
            INIT_51 => X"000000e500000000000000e300000000000000de000000000000009200000000",
            INIT_52 => X"000000e600000000000000e700000000000000ea00000000000000ec00000000",
            INIT_53 => X"000000e600000000000000e800000000000000e700000000000000e500000000",
            INIT_54 => X"000000df00000000000000e500000000000000e700000000000000e700000000",
            INIT_55 => X"00000089000000000000009200000000000000a400000000000000bf00000000",
            INIT_56 => X"0000009500000000000000790000000000000080000000000000008600000000",
            INIT_57 => X"000000ed00000000000000eb00000000000000ea00000000000000d800000000",
            INIT_58 => X"000000c800000000000000c700000000000000bc00000000000000c300000000",
            INIT_59 => X"000000d300000000000000d500000000000000df00000000000000d100000000",
            INIT_5A => X"000000d200000000000000db00000000000000dc00000000000000d800000000",
            INIT_5B => X"000000dc00000000000000d800000000000000d300000000000000d100000000",
            INIT_5C => X"000000da00000000000000e100000000000000e200000000000000e100000000",
            INIT_5D => X"000000b200000000000000b500000000000000af00000000000000b700000000",
            INIT_5E => X"000000b9000000000000008e00000000000000aa00000000000000ba00000000",
            INIT_5F => X"000000ec00000000000000ea00000000000000e700000000000000db00000000",
            INIT_60 => X"000000d600000000000000ca00000000000000bf00000000000000c100000000",
            INIT_61 => X"000000ab00000000000000cb00000000000000d600000000000000df00000000",
            INIT_62 => X"0000006200000000000000ae00000000000000cf00000000000000b100000000",
            INIT_63 => X"0000007a000000000000006f0000000000000065000000000000005d00000000",
            INIT_64 => X"000000df00000000000000ca0000000000000099000000000000008900000000",
            INIT_65 => X"000000d900000000000000df00000000000000dc00000000000000da00000000",
            INIT_66 => X"000000de00000000000000c400000000000000d400000000000000dd00000000",
            INIT_67 => X"000000eb00000000000000e800000000000000dd00000000000000db00000000",
            INIT_68 => X"0000007d0000000000000071000000000000006f000000000000007100000000",
            INIT_69 => X"000000be00000000000000bf00000000000000aa000000000000008a00000000",
            INIT_6A => X"00000036000000000000009e00000000000000d800000000000000d000000000",
            INIT_6B => X"0000004200000000000000350000000000000031000000000000002d00000000",
            INIT_6C => X"000000ea00000000000000dd000000000000009f000000000000006600000000",
            INIT_6D => X"000000cf00000000000000df00000000000000e300000000000000e900000000",
            INIT_6E => X"000000c700000000000000d400000000000000d300000000000000ca00000000",
            INIT_6F => X"000000dd00000000000000d300000000000000bc00000000000000b300000000",
            INIT_70 => X"00000044000000000000003f0000000000000045000000000000003d00000000",
            INIT_71 => X"000000c30000000000000097000000000000008b000000000000007b00000000",
            INIT_72 => X"0000006700000000000000a300000000000000ce00000000000000d600000000",
            INIT_73 => X"000000b5000000000000008a0000000000000065000000000000005f00000000",
            INIT_74 => X"000000cd00000000000000db00000000000000dd00000000000000cf00000000",
            INIT_75 => X"000000830000000000000093000000000000009e00000000000000b700000000",
            INIT_76 => X"0000008500000000000000880000000000000082000000000000007d00000000",
            INIT_77 => X"000000c500000000000000b6000000000000008a000000000000008000000000",
            INIT_78 => X"0000007f0000000000000055000000000000003a000000000000002800000000",
            INIT_79 => X"000000a300000000000000770000000000000060000000000000008400000000",
            INIT_7A => X"000000b500000000000000b600000000000000b800000000000000ad00000000",
            INIT_7B => X"000000c800000000000000da00000000000000c600000000000000b700000000",
            INIT_7C => X"000000840000000000000091000000000000009f00000000000000ae00000000",
            INIT_7D => X"00000063000000000000005e0000000000000062000000000000007400000000",
            INIT_7E => X"0000008a000000000000007a000000000000006b000000000000006900000000",
            INIT_7F => X"000000b900000000000000bc000000000000009d000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "sampleifmap_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ce0000000000000086000000000000001a000000000000000d00000000",
            INIT_01 => X"000000ac000000000000008d0000000000000076000000000000008a00000000",
            INIT_02 => X"000000e400000000000000dc00000000000000cf00000000000000b500000000",
            INIT_03 => X"000000b000000000000000e200000000000000e600000000000000e000000000",
            INIT_04 => X"00000091000000000000008e000000000000008a000000000000009000000000",
            INIT_05 => X"0000009a00000000000000950000000000000095000000000000009a00000000",
            INIT_06 => X"000000bb00000000000000ad00000000000000a0000000000000009d00000000",
            INIT_07 => X"0000009d00000000000000a500000000000000b200000000000000be00000000",
            INIT_08 => X"000000e100000000000000c8000000000000003a000000000000000500000000",
            INIT_09 => X"000000e200000000000000d400000000000000c700000000000000c500000000",
            INIT_0A => X"000000e600000000000000e800000000000000e900000000000000e500000000",
            INIT_0B => X"000000d200000000000000dd00000000000000df00000000000000d100000000",
            INIT_0C => X"000000bc00000000000000c100000000000000b400000000000000c600000000",
            INIT_0D => X"000000b800000000000000c000000000000000c200000000000000bd00000000",
            INIT_0E => X"0000009000000000000000a100000000000000ab00000000000000ac00000000",
            INIT_0F => X"0000008a00000000000000800000000000000083000000000000008800000000",
            INIT_10 => X"000000ba00000000000000be0000000000000091000000000000002700000000",
            INIT_11 => X"000000c200000000000000c200000000000000c000000000000000b800000000",
            INIT_12 => X"000000be00000000000000c000000000000000bf00000000000000c200000000",
            INIT_13 => X"00000093000000000000009a00000000000000b400000000000000b100000000",
            INIT_14 => X"000000710000000000000092000000000000009c000000000000009100000000",
            INIT_15 => X"0000006f000000000000007e0000000000000084000000000000007200000000",
            INIT_16 => X"0000005e000000000000005d000000000000005b000000000000005c00000000",
            INIT_17 => X"0000008100000000000000810000000000000079000000000000006900000000",
            INIT_18 => X"00000089000000000000008f00000000000000a2000000000000007a00000000",
            INIT_19 => X"00000082000000000000007f0000000000000080000000000000008300000000",
            INIT_1A => X"00000081000000000000007f0000000000000080000000000000008300000000",
            INIT_1B => X"000000640000000000000068000000000000007c000000000000008100000000",
            INIT_1C => X"0000005e00000000000000700000000000000076000000000000006600000000",
            INIT_1D => X"000000530000000000000057000000000000005e000000000000005e00000000",
            INIT_1E => X"00000065000000000000005d0000000000000053000000000000005000000000",
            INIT_1F => X"0000008200000000000000790000000000000073000000000000006c00000000",
            INIT_20 => X"00000050000000000000004d000000000000004c000000000000004900000000",
            INIT_21 => X"0000005a00000000000000570000000000000057000000000000005400000000",
            INIT_22 => X"00000071000000000000006b0000000000000066000000000000005e00000000",
            INIT_23 => X"0000007800000000000000760000000000000076000000000000007300000000",
            INIT_24 => X"00000064000000000000006a000000000000006e000000000000007300000000",
            INIT_25 => X"00000050000000000000004f0000000000000055000000000000005f00000000",
            INIT_26 => X"000000520000000000000050000000000000004d000000000000005000000000",
            INIT_27 => X"00000088000000000000007d0000000000000071000000000000005c00000000",
            INIT_28 => X"0000001200000000000000090000000000000003000000000000000d00000000",
            INIT_29 => X"0000001600000000000000140000000000000015000000000000001200000000",
            INIT_2A => X"00000030000000000000002a0000000000000022000000000000001a00000000",
            INIT_2B => X"000000460000000000000042000000000000003c000000000000003400000000",
            INIT_2C => X"0000003c00000000000000430000000000000048000000000000004700000000",
            INIT_2D => X"0000003900000000000000350000000000000035000000000000003700000000",
            INIT_2E => X"0000005700000000000000480000000000000039000000000000003900000000",
            INIT_2F => X"0000008900000000000000820000000000000078000000000000006800000000",
            INIT_30 => X"000000200000000000000008000000000000000b000000000000002400000000",
            INIT_31 => X"0000000300000000000000080000000000000016000000000000002400000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_33 => X"0000000300000000000000010000000000000005000000000000000600000000",
            INIT_34 => X"0000001500000000000000150000000000000018000000000000000d00000000",
            INIT_35 => X"00000027000000000000001e0000000000000016000000000000001500000000",
            INIT_36 => X"0000007b00000000000000710000000000000055000000000000003900000000",
            INIT_37 => X"000000990000000000000086000000000000007a000000000000007400000000",
            INIT_38 => X"0000001b000000000000000d000000000000001a000000000000002300000000",
            INIT_39 => X"0000001b00000000000000310000000000000046000000000000004700000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000000a000000000000001f0000000000000039000000000000001100000000",
            INIT_3C => X"0000000e00000000000000070000000000000004000000000000000400000000",
            INIT_3D => X"00000056000000000000003e0000000000000029000000000000001900000000",
            INIT_3E => X"0000007200000000000000840000000000000090000000000000007a00000000",
            INIT_3F => X"000000ac00000000000000920000000000000084000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000030000000000000004000000000000000d000000000000001000000000",
            INIT_41 => X"0000002400000000000000360000000000000041000000000000002d00000000",
            INIT_42 => X"0000000000000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"0000008300000000000000a10000000000000076000000000000000700000000",
            INIT_44 => X"0000006d00000000000000690000000000000069000000000000007000000000",
            INIT_45 => X"00000097000000000000009a000000000000008a000000000000007600000000",
            INIT_46 => X"00000078000000000000006a0000000000000069000000000000007f00000000",
            INIT_47 => X"000000b800000000000000a4000000000000008e000000000000008100000000",
            INIT_48 => X"000000000000000000000000000000000000000c000000000000002800000000",
            INIT_49 => X"000000150000000000000020000000000000001e000000000000000c00000000",
            INIT_4A => X"0000000300000000000000020000000000000002000000000000000700000000",
            INIT_4B => X"000000cd00000000000000b60000000000000044000000000000000000000000",
            INIT_4C => X"000000bb00000000000000c300000000000000c200000000000000c400000000",
            INIT_4D => X"00000067000000000000007b000000000000009600000000000000ac00000000",
            INIT_4E => X"00000081000000000000007a0000000000000068000000000000005f00000000",
            INIT_4F => X"000000b900000000000000ab0000000000000098000000000000008400000000",
            INIT_50 => X"000000010000000000000001000000000000001a000000000000004500000000",
            INIT_51 => X"0000000c0000000000000012000000000000000c000000000000000400000000",
            INIT_52 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_53 => X"000000cb00000000000000990000000000000020000000000000000100000000",
            INIT_54 => X"0000009b00000000000000b300000000000000bf00000000000000c300000000",
            INIT_55 => X"0000005e0000000000000051000000000000005b000000000000007700000000",
            INIT_56 => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_57 => X"000000b800000000000000ad00000000000000a2000000000000009000000000",
            INIT_58 => X"000000020000000000000001000000000000002f000000000000005300000000",
            INIT_59 => X"0000000400000000000000070000000000000005000000000000000200000000",
            INIT_5A => X"0000000300000000000000010000000000000001000000000000000100000000",
            INIT_5B => X"000000cd000000000000008e000000000000001b000000000000000100000000",
            INIT_5C => X"00000055000000000000007900000000000000a900000000000000c600000000",
            INIT_5D => X"0000007900000000000000660000000000000055000000000000004a00000000",
            INIT_5E => X"000000840000000000000079000000000000007a000000000000008000000000",
            INIT_5F => X"000000ba00000000000000b000000000000000a5000000000000009300000000",
            INIT_60 => X"0000000300000000000000060000000000000036000000000000005c00000000",
            INIT_61 => X"0000000100000000000000010000000000000001000000000000000200000000",
            INIT_62 => X"0000000100000000000000010000000000000001000000000000000100000000",
            INIT_63 => X"0000009d0000000000000066000000000000000f000000000000000000000000",
            INIT_64 => X"0000004a0000000000000038000000000000004a000000000000007500000000",
            INIT_65 => X"0000007c000000000000007a0000000000000073000000000000006300000000",
            INIT_66 => X"000000880000000000000080000000000000007d000000000000007b00000000",
            INIT_67 => X"000000bc00000000000000b100000000000000a2000000000000009400000000",
            INIT_68 => X"0000000b0000000000000013000000000000002b000000000000005700000000",
            INIT_69 => X"0000000200000000000000020000000000000005000000000000000800000000",
            INIT_6A => X"0000000200000000000000030000000000000003000000000000000300000000",
            INIT_6B => X"00000047000000000000002a0000000000000004000000000000000000000000",
            INIT_6C => X"0000007100000000000000500000000000000039000000000000003500000000",
            INIT_6D => X"00000074000000000000007b0000000000000086000000000000008400000000",
            INIT_6E => X"0000008f000000000000008b0000000000000083000000000000007800000000",
            INIT_6F => X"000000bc00000000000000b600000000000000a9000000000000009c00000000",
            INIT_70 => X"0000001f0000000000000024000000000000002e000000000000005200000000",
            INIT_71 => X"0000001000000000000000110000000000000016000000000000001b00000000",
            INIT_72 => X"0000001300000000000000140000000000000013000000000000001200000000",
            INIT_73 => X"0000004000000000000000250000000000000017000000000000001300000000",
            INIT_74 => X"0000008000000000000000740000000000000068000000000000005700000000",
            INIT_75 => X"0000007300000000000000750000000000000083000000000000008b00000000",
            INIT_76 => X"00000094000000000000008b0000000000000083000000000000007b00000000",
            INIT_77 => X"000000bb00000000000000b900000000000000ae000000000000009f00000000",
            INIT_78 => X"00000037000000000000003a000000000000003e000000000000005500000000",
            INIT_79 => X"00000030000000000000002e000000000000002f000000000000003300000000",
            INIT_7A => X"0000003700000000000000350000000000000033000000000000003100000000",
            INIT_7B => X"0000006800000000000000510000000000000044000000000000003b00000000",
            INIT_7C => X"0000007f0000000000000085000000000000007f000000000000007400000000",
            INIT_7D => X"0000007a00000000000000720000000000000076000000000000007f00000000",
            INIT_7E => X"00000095000000000000008d0000000000000088000000000000008100000000",
            INIT_7F => X"000000ba00000000000000b400000000000000a8000000000000009e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "sampleifmap_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e900000000000000e900000000000000e700000000000000e700000000",
            INIT_05 => X"000000e900000000000000e800000000000000e700000000000000e800000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e900000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000ea00000000000000ea00000000",
            INIT_0D => X"000000ec00000000000000ec00000000000000ea00000000000000eb00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ec00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000eb00000000000000eb00000000000000ea00000000000000e900000000",
            INIT_15 => X"000000ea00000000000000e900000000000000eb00000000000000e600000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e200000000000000e600000000000000e800000000000000e900000000",
            INIT_1D => X"000000e400000000000000d200000000000000d800000000000000c000000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000d200000000000000e100000000000000ed00000000000000ee00000000",
            INIT_25 => X"000000e500000000000000da00000000000000cd00000000000000ac00000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ef00000000",
            INIT_29 => X"000000eb00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e700000000000000ed00000000000000e900000000000000eb00000000",
            INIT_2C => X"000000bc00000000000000c600000000000000cd00000000000000d800000000",
            INIT_2D => X"000000e400000000000000d700000000000000c400000000000000b300000000",
            INIT_2E => X"000000ec00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e400000000000000e600000000000000e300000000000000e500000000",
            INIT_31 => X"000000ed00000000000000ed00000000000000ec00000000000000e800000000",
            INIT_32 => X"000000ed00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_33 => X"000000e200000000000000ed00000000000000e400000000000000e500000000",
            INIT_34 => X"000000b000000000000000b400000000000000b400000000000000c500000000",
            INIT_35 => X"000000ce00000000000000a9000000000000009f00000000000000a300000000",
            INIT_36 => X"000000eb00000000000000ec00000000000000ed00000000000000ee00000000",
            INIT_37 => X"000000ed00000000000000ed00000000000000ee00000000000000ec00000000",
            INIT_38 => X"000000e800000000000000ea00000000000000e600000000000000dc00000000",
            INIT_39 => X"000000ed00000000000000ee00000000000000ed00000000000000ea00000000",
            INIT_3A => X"000000ee00000000000000ec00000000000000ed00000000000000ed00000000",
            INIT_3B => X"000000da00000000000000ec00000000000000de00000000000000cc00000000",
            INIT_3C => X"000000bf00000000000000c900000000000000c900000000000000cc00000000",
            INIT_3D => X"000000c700000000000000b000000000000000ae00000000000000b600000000",
            INIT_3E => X"000000ee00000000000000ee00000000000000ef00000000000000ef00000000",
            INIT_3F => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ef00000000000000ee00000000000000ec00000000000000ea00000000",
            INIT_41 => X"000000ec00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_43 => X"000000e700000000000000ea00000000000000dd00000000000000c600000000",
            INIT_44 => X"000000da00000000000000e400000000000000d800000000000000d500000000",
            INIT_45 => X"000000eb00000000000000e900000000000000e000000000000000dd00000000",
            INIT_46 => X"000000f000000000000000ef00000000000000ee00000000000000f000000000",
            INIT_47 => X"000000ee00000000000000f000000000000000f000000000000000f000000000",
            INIT_48 => X"0000009b000000000000008e000000000000008a000000000000008c00000000",
            INIT_49 => X"000000ea00000000000000ec00000000000000ea00000000000000bc00000000",
            INIT_4A => X"000000ed00000000000000ed00000000000000eb00000000000000e900000000",
            INIT_4B => X"000000ed00000000000000ea00000000000000e400000000000000d800000000",
            INIT_4C => X"000000e800000000000000ec00000000000000e600000000000000e600000000",
            INIT_4D => X"000000cc00000000000000db00000000000000e900000000000000ed00000000",
            INIT_4E => X"000000c700000000000000b400000000000000b300000000000000bd00000000",
            INIT_4F => X"000000f000000000000000f000000000000000f100000000000000eb00000000",
            INIT_50 => X"0000007f000000000000007d0000000000000079000000000000008200000000",
            INIT_51 => X"000000e200000000000000e400000000000000e5000000000000009f00000000",
            INIT_52 => X"000000ed00000000000000ec00000000000000ea00000000000000e800000000",
            INIT_53 => X"000000eb00000000000000ed00000000000000eb00000000000000ea00000000",
            INIT_54 => X"000000e800000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_55 => X"0000009c00000000000000a500000000000000b800000000000000ce00000000",
            INIT_56 => X"000000a20000000000000085000000000000008c000000000000009500000000",
            INIT_57 => X"000000f000000000000000f000000000000000f100000000000000e400000000",
            INIT_58 => X"000000d300000000000000d300000000000000ca00000000000000d400000000",
            INIT_59 => X"000000d100000000000000d500000000000000e300000000000000d900000000",
            INIT_5A => X"000000dd00000000000000e200000000000000de00000000000000d500000000",
            INIT_5B => X"000000e500000000000000e100000000000000dd00000000000000db00000000",
            INIT_5C => X"000000e700000000000000ed00000000000000ec00000000000000ea00000000",
            INIT_5D => X"000000c200000000000000c800000000000000c600000000000000cc00000000",
            INIT_5E => X"000000c3000000000000009700000000000000b200000000000000c500000000",
            INIT_5F => X"000000f000000000000000f100000000000000f000000000000000e600000000",
            INIT_60 => X"000000d900000000000000d300000000000000ca00000000000000cf00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000db00000000000000e100000000",
            INIT_62 => X"0000007000000000000000b800000000000000d500000000000000b400000000",
            INIT_63 => X"0000008a00000000000000810000000000000079000000000000007200000000",
            INIT_64 => X"000000ec00000000000000d800000000000000a7000000000000009800000000",
            INIT_65 => X"000000e200000000000000ea00000000000000e900000000000000e800000000",
            INIT_66 => X"000000e600000000000000cb00000000000000db00000000000000e400000000",
            INIT_67 => X"000000f100000000000000ef00000000000000e600000000000000e300000000",
            INIT_68 => X"00000083000000000000007d000000000000007d000000000000008200000000",
            INIT_69 => X"000000c700000000000000c900000000000000b6000000000000009100000000",
            INIT_6A => X"0000004700000000000000ac00000000000000e600000000000000db00000000",
            INIT_6B => X"0000005400000000000000490000000000000049000000000000004600000000",
            INIT_6C => X"000000ef00000000000000e300000000000000a8000000000000007200000000",
            INIT_6D => X"000000d300000000000000e400000000000000e700000000000000ed00000000",
            INIT_6E => X"000000ce00000000000000db00000000000000da00000000000000d000000000",
            INIT_6F => X"000000e700000000000000dd00000000000000c500000000000000ba00000000",
            INIT_70 => X"00000055000000000000004f0000000000000056000000000000005100000000",
            INIT_71 => X"000000c8000000000000009d000000000000009b000000000000008d00000000",
            INIT_72 => X"0000007900000000000000b400000000000000df00000000000000e400000000",
            INIT_73 => X"000000c000000000000000970000000000000075000000000000007000000000",
            INIT_74 => X"000000cb00000000000000db00000000000000de00000000000000d400000000",
            INIT_75 => X"0000008a000000000000009a00000000000000a600000000000000ba00000000",
            INIT_76 => X"0000008e0000000000000092000000000000008b000000000000008500000000",
            INIT_77 => X"000000d400000000000000c50000000000000099000000000000008900000000",
            INIT_78 => X"0000009000000000000000620000000000000046000000000000003500000000",
            INIT_79 => X"0000009e0000000000000073000000000000006b000000000000009700000000",
            INIT_7A => X"000000c100000000000000c200000000000000c200000000000000b400000000",
            INIT_7B => X"000000d200000000000000e400000000000000d100000000000000c200000000",
            INIT_7C => X"00000088000000000000009600000000000000a500000000000000b500000000",
            INIT_7D => X"0000006f000000000000006a000000000000006f000000000000007d00000000",
            INIT_7E => X"0000009700000000000000870000000000000079000000000000007600000000",
            INIT_7F => X"000000cb00000000000000ce00000000000000ae00000000000000a400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "sampleifmap_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d8000000000000008c000000000000001d000000000000000f00000000",
            INIT_01 => X"000000a20000000000000085000000000000007b000000000000009600000000",
            INIT_02 => X"000000ea00000000000000e000000000000000d100000000000000b500000000",
            INIT_03 => X"000000bd00000000000000ee00000000000000f100000000000000ea00000000",
            INIT_04 => X"000000a3000000000000009e000000000000009a000000000000009f00000000",
            INIT_05 => X"000000ab00000000000000a500000000000000a500000000000000ab00000000",
            INIT_06 => X"000000cc00000000000000be00000000000000b100000000000000ae00000000",
            INIT_07 => X"000000af00000000000000b700000000000000c400000000000000cf00000000",
            INIT_08 => X"000000e800000000000000cf000000000000003e000000000000000500000000",
            INIT_09 => X"000000e000000000000000d400000000000000cf00000000000000cd00000000",
            INIT_0A => X"000000ee00000000000000ee00000000000000ec00000000000000e600000000",
            INIT_0B => X"000000e400000000000000ee00000000000000ee00000000000000dd00000000",
            INIT_0C => X"000000d500000000000000d800000000000000c800000000000000d900000000",
            INIT_0D => X"000000cc00000000000000d400000000000000d600000000000000d400000000",
            INIT_0E => X"000000a500000000000000b500000000000000bf00000000000000c100000000",
            INIT_0F => X"0000009a000000000000008f0000000000000092000000000000009c00000000",
            INIT_10 => X"000000c400000000000000cc000000000000009b000000000000002d00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000c500000000",
            INIT_12 => X"000000cf00000000000000cf00000000000000cb00000000000000ce00000000",
            INIT_13 => X"000000a900000000000000b000000000000000c600000000000000c100000000",
            INIT_14 => X"0000008500000000000000a300000000000000ab00000000000000a100000000",
            INIT_15 => X"000000870000000000000096000000000000009d000000000000008900000000",
            INIT_16 => X"0000007400000000000000720000000000000070000000000000007300000000",
            INIT_17 => X"0000008e000000000000008d0000000000000085000000000000007d00000000",
            INIT_18 => X"0000009a00000000000000a000000000000000b3000000000000008700000000",
            INIT_19 => X"0000009600000000000000960000000000000098000000000000009800000000",
            INIT_1A => X"0000009500000000000000930000000000000093000000000000009600000000",
            INIT_1B => X"0000007a000000000000007e0000000000000091000000000000009500000000",
            INIT_1C => X"0000006d00000000000000800000000000000086000000000000007800000000",
            INIT_1D => X"0000006700000000000000700000000000000075000000000000007000000000",
            INIT_1E => X"00000075000000000000006f0000000000000067000000000000006100000000",
            INIT_1F => X"000000900000000000000085000000000000007d000000000000007900000000",
            INIT_20 => X"0000005d000000000000005a000000000000005a000000000000005700000000",
            INIT_21 => X"0000006900000000000000660000000000000066000000000000006200000000",
            INIT_22 => X"00000083000000000000007c0000000000000077000000000000006f00000000",
            INIT_23 => X"0000008500000000000000840000000000000088000000000000008900000000",
            INIT_24 => X"00000077000000000000007f0000000000000085000000000000008800000000",
            INIT_25 => X"0000005c00000000000000610000000000000065000000000000006d00000000",
            INIT_26 => X"0000006200000000000000640000000000000064000000000000005e00000000",
            INIT_27 => X"0000009500000000000000870000000000000077000000000000006800000000",
            INIT_28 => X"0000001a0000000000000010000000000000000b000000000000001900000000",
            INIT_29 => X"0000001e00000000000000190000000000000019000000000000001a00000000",
            INIT_2A => X"0000003b0000000000000033000000000000002b000000000000002400000000",
            INIT_2B => X"0000004f000000000000004d000000000000004b000000000000004500000000",
            INIT_2C => X"0000004800000000000000510000000000000058000000000000005700000000",
            INIT_2D => X"0000004500000000000000450000000000000044000000000000004300000000",
            INIT_2E => X"000000640000000000000059000000000000004e000000000000004700000000",
            INIT_2F => X"000000920000000000000088000000000000007c000000000000007100000000",
            INIT_30 => X"0000002c000000000000000d0000000000000010000000000000002e00000000",
            INIT_31 => X"00000008000000000000000b0000000000000019000000000000002d00000000",
            INIT_32 => X"0000000400000000000000020000000000000002000000000000000400000000",
            INIT_33 => X"0000001700000000000000130000000000000012000000000000000d00000000",
            INIT_34 => X"0000001f00000000000000210000000000000026000000000000001d00000000",
            INIT_35 => X"0000003a0000000000000032000000000000002c000000000000002600000000",
            INIT_36 => X"0000007b0000000000000073000000000000005a000000000000004600000000",
            INIT_37 => X"000000a0000000000000008b000000000000007b000000000000007300000000",
            INIT_38 => X"000000290000000000000013000000000000001b000000000000002900000000",
            INIT_39 => X"0000001f00000000000000320000000000000046000000000000005100000000",
            INIT_3A => X"0000000000000000000000020000000000000005000000000000000f00000000",
            INIT_3B => X"0000002400000000000000320000000000000040000000000000001100000000",
            INIT_3C => X"00000023000000000000001e000000000000001e000000000000001e00000000",
            INIT_3D => X"0000006100000000000000470000000000000037000000000000002b00000000",
            INIT_3E => X"0000006900000000000000780000000000000083000000000000007c00000000",
            INIT_3F => X"000000b300000000000000980000000000000086000000000000006f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000000a000000000000000a000000000000000f00000000",
            INIT_41 => X"00000021000000000000002b0000000000000034000000000000002c00000000",
            INIT_42 => X"0000000100000000000000020000000000000004000000000000001200000000",
            INIT_43 => X"00000080000000000000009e0000000000000075000000000000000800000000",
            INIT_44 => X"0000006900000000000000670000000000000069000000000000007000000000",
            INIT_45 => X"0000007e000000000000007e0000000000000073000000000000006b00000000",
            INIT_46 => X"00000074000000000000005e0000000000000056000000000000006a00000000",
            INIT_47 => X"000000c200000000000000ac0000000000000093000000000000008200000000",
            INIT_48 => X"000000040000000000000003000000000000000a000000000000002800000000",
            INIT_49 => X"0000000a000000000000000c000000000000000c000000000000000600000000",
            INIT_4A => X"0000000200000000000000010000000000000001000000000000000600000000",
            INIT_4B => X"000000820000000000000080000000000000003a000000000000000000000000",
            INIT_4C => X"000000710000000000000077000000000000007b000000000000007f00000000",
            INIT_4D => X"00000042000000000000004b0000000000000060000000000000006e00000000",
            INIT_4E => X"000000840000000000000076000000000000005d000000000000004700000000",
            INIT_4F => X"000000c500000000000000b600000000000000a2000000000000008d00000000",
            INIT_50 => X"000000010000000000000001000000000000001d000000000000004d00000000",
            INIT_51 => X"0000000200000000000000030000000000000002000000000000000100000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_53 => X"0000002f000000000000002d000000000000000c000000000000000100000000",
            INIT_54 => X"0000003100000000000000320000000000000030000000000000002e00000000",
            INIT_55 => X"0000004d00000000000000300000000000000026000000000000002a00000000",
            INIT_56 => X"000000870000000000000080000000000000007e000000000000006e00000000",
            INIT_57 => X"000000c600000000000000bb00000000000000b0000000000000009900000000",
            INIT_58 => X"0000000100000000000000010000000000000034000000000000005e00000000",
            INIT_59 => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000002000000000000000190000000000000003000000000000000200000000",
            INIT_5C => X"0000001d00000000000000190000000000000019000000000000001900000000",
            INIT_5D => X"00000071000000000000005c0000000000000042000000000000002900000000",
            INIT_5E => X"0000008b000000000000007f000000000000007e000000000000007c00000000",
            INIT_5F => X"000000c900000000000000bf00000000000000b3000000000000009d00000000",
            INIT_60 => X"000000020000000000000007000000000000003c000000000000006600000000",
            INIT_61 => X"0000000200000000000000030000000000000003000000000000000200000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000001f00000000000000130000000000000001000000000000000300000000",
            INIT_64 => X"0000003a000000000000001b000000000000000d000000000000001100000000",
            INIT_65 => X"0000007c000000000000007e0000000000000073000000000000005a00000000",
            INIT_66 => X"0000009100000000000000870000000000000082000000000000007b00000000",
            INIT_67 => X"000000ca00000000000000c000000000000000b0000000000000009f00000000",
            INIT_68 => X"0000000c00000000000000170000000000000033000000000000006300000000",
            INIT_69 => X"00000007000000000000000a000000000000000b000000000000000a00000000",
            INIT_6A => X"0000000300000000000000040000000000000004000000000000000400000000",
            INIT_6B => X"00000015000000000000000d0000000000000005000000000000000600000000",
            INIT_6C => X"00000062000000000000004d0000000000000032000000000000001b00000000",
            INIT_6D => X"0000007d000000000000007e000000000000007e000000000000007100000000",
            INIT_6E => X"0000009a0000000000000094000000000000008a000000000000008000000000",
            INIT_6F => X"000000ca00000000000000c500000000000000b800000000000000a800000000",
            INIT_70 => X"00000023000000000000002c0000000000000039000000000000006000000000",
            INIT_71 => X"00000017000000000000001a000000000000001c000000000000001e00000000",
            INIT_72 => X"0000001700000000000000160000000000000015000000000000001500000000",
            INIT_73 => X"000000370000000000000028000000000000001f000000000000001b00000000",
            INIT_74 => X"0000007000000000000000660000000000000058000000000000004600000000",
            INIT_75 => X"0000007f000000000000007a000000000000007a000000000000007900000000",
            INIT_76 => X"000000a00000000000000095000000000000008b000000000000008500000000",
            INIT_77 => X"000000ca00000000000000c800000000000000bd00000000000000ac00000000",
            INIT_78 => X"0000003d0000000000000043000000000000004b000000000000006500000000",
            INIT_79 => X"0000003700000000000000350000000000000035000000000000003800000000",
            INIT_7A => X"0000003e000000000000003a0000000000000038000000000000003700000000",
            INIT_7B => X"0000006000000000000000540000000000000047000000000000004300000000",
            INIT_7C => X"000000790000000000000074000000000000006d000000000000006700000000",
            INIT_7D => X"00000083000000000000007d000000000000007c000000000000007f00000000",
            INIT_7E => X"000000a200000000000000980000000000000091000000000000008800000000",
            INIT_7F => X"000000c800000000000000c300000000000000b700000000000000ab00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "sampleifmap_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e800000000000000e800000000000000e700000000000000eb00000000",
            INIT_01 => X"000000e800000000000000e800000000000000e800000000000000e800000000",
            INIT_02 => X"000000e900000000000000e900000000000000e800000000000000e800000000",
            INIT_03 => X"000000e900000000000000e900000000000000e900000000000000e900000000",
            INIT_04 => X"000000e800000000000000e900000000000000e900000000000000e900000000",
            INIT_05 => X"000000e600000000000000e800000000000000ea00000000000000ea00000000",
            INIT_06 => X"000000e800000000000000e800000000000000e900000000000000e700000000",
            INIT_07 => X"000000e800000000000000e900000000000000e900000000000000e800000000",
            INIT_08 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_09 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_0A => X"000000ec00000000000000ec00000000000000eb00000000000000eb00000000",
            INIT_0B => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_0C => X"000000ea00000000000000ea00000000000000e900000000000000e900000000",
            INIT_0D => X"000000eb00000000000000ed00000000000000ee00000000000000ed00000000",
            INIT_0E => X"000000eb00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_0F => X"000000eb00000000000000ec00000000000000ec00000000000000eb00000000",
            INIT_10 => X"000000ea00000000000000ea00000000000000ea00000000000000ed00000000",
            INIT_11 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_12 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_13 => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_14 => X"000000ec00000000000000ea00000000000000e700000000000000e700000000",
            INIT_15 => X"000000ea00000000000000eb00000000000000ee00000000000000e900000000",
            INIT_16 => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_17 => X"000000ea00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_18 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_19 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_1A => X"000000ea00000000000000ea00000000000000ea00000000000000ea00000000",
            INIT_1B => X"000000ea00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_1C => X"000000e700000000000000e800000000000000e700000000000000e600000000",
            INIT_1D => X"000000e600000000000000d500000000000000db00000000000000c500000000",
            INIT_1E => X"000000ea00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_1F => X"000000eb00000000000000eb00000000000000eb00000000000000ea00000000",
            INIT_20 => X"000000eb00000000000000eb00000000000000ea00000000000000ed00000000",
            INIT_21 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_22 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_23 => X"000000eb00000000000000eb00000000000000ea00000000000000ea00000000",
            INIT_24 => X"000000db00000000000000e600000000000000ed00000000000000ec00000000",
            INIT_25 => X"000000e800000000000000dd00000000000000d000000000000000b300000000",
            INIT_26 => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_27 => X"000000ec00000000000000ec00000000000000ec00000000000000ec00000000",
            INIT_28 => X"000000eb00000000000000eb00000000000000eb00000000000000ee00000000",
            INIT_29 => X"000000eb00000000000000eb00000000000000eb00000000000000eb00000000",
            INIT_2A => X"000000ec00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_2B => X"000000e800000000000000ed00000000000000ea00000000000000ec00000000",
            INIT_2C => X"000000c800000000000000cf00000000000000d200000000000000da00000000",
            INIT_2D => X"000000e800000000000000dc00000000000000ca00000000000000bd00000000",
            INIT_2E => X"000000eb00000000000000eb00000000000000eb00000000000000ed00000000",
            INIT_2F => X"000000ed00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_30 => X"000000e600000000000000e700000000000000e400000000000000e500000000",
            INIT_31 => X"000000eb00000000000000eb00000000000000ec00000000000000e900000000",
            INIT_32 => X"000000ee00000000000000ed00000000000000ec00000000000000ec00000000",
            INIT_33 => X"000000e400000000000000ee00000000000000e500000000000000e600000000",
            INIT_34 => X"000000be00000000000000bf00000000000000be00000000000000cc00000000",
            INIT_35 => X"000000d300000000000000b100000000000000ab00000000000000b100000000",
            INIT_36 => X"000000eb00000000000000e900000000000000ea00000000000000ef00000000",
            INIT_37 => X"000000ee00000000000000ed00000000000000ed00000000000000ec00000000",
            INIT_38 => X"000000ea00000000000000ee00000000000000e900000000000000de00000000",
            INIT_39 => X"000000ec00000000000000eb00000000000000ec00000000000000ea00000000",
            INIT_3A => X"000000ef00000000000000ed00000000000000ee00000000000000ee00000000",
            INIT_3B => X"000000da00000000000000eb00000000000000dd00000000000000cb00000000",
            INIT_3C => X"000000cb00000000000000d300000000000000d200000000000000d200000000",
            INIT_3D => X"000000cc00000000000000b900000000000000bb00000000000000c400000000",
            INIT_3E => X"000000ee00000000000000ed00000000000000ee00000000000000f000000000",
            INIT_3F => X"000000ee00000000000000ee00000000000000ee00000000000000ee00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f300000000000000f600000000000000f300000000000000f100000000",
            INIT_41 => X"000000eb00000000000000eb00000000000000ed00000000000000f000000000",
            INIT_42 => X"000000ef00000000000000ed00000000000000ed00000000000000ed00000000",
            INIT_43 => X"000000e500000000000000e700000000000000da00000000000000c400000000",
            INIT_44 => X"000000e300000000000000eb00000000000000de00000000000000d900000000",
            INIT_45 => X"000000f100000000000000f000000000000000eb00000000000000ea00000000",
            INIT_46 => X"000000f000000000000000f000000000000000f000000000000000f300000000",
            INIT_47 => X"000000ee00000000000000ef00000000000000ef00000000000000ef00000000",
            INIT_48 => X"000000a100000000000000990000000000000094000000000000009500000000",
            INIT_49 => X"000000e800000000000000e900000000000000e900000000000000bf00000000",
            INIT_4A => X"000000eb00000000000000ec00000000000000eb00000000000000ea00000000",
            INIT_4B => X"000000ec00000000000000e800000000000000e200000000000000d600000000",
            INIT_4C => X"000000ef00000000000000f100000000000000eb00000000000000e800000000",
            INIT_4D => X"000000d300000000000000e200000000000000f300000000000000f700000000",
            INIT_4E => X"000000c900000000000000b900000000000000ba00000000000000c300000000",
            INIT_4F => X"000000ef00000000000000ef00000000000000ef00000000000000eb00000000",
            INIT_50 => X"0000008900000000000000890000000000000085000000000000008d00000000",
            INIT_51 => X"000000e000000000000000e100000000000000e700000000000000a500000000",
            INIT_52 => X"000000eb00000000000000ea00000000000000ea00000000000000e900000000",
            INIT_53 => X"000000ec00000000000000ee00000000000000ec00000000000000eb00000000",
            INIT_54 => X"000000ee00000000000000f100000000000000f000000000000000ee00000000",
            INIT_55 => X"000000a300000000000000ac00000000000000bf00000000000000d500000000",
            INIT_56 => X"000000a6000000000000008f0000000000000099000000000000009f00000000",
            INIT_57 => X"000000ef00000000000000ee00000000000000ef00000000000000e500000000",
            INIT_58 => X"000000df00000000000000e000000000000000d700000000000000e000000000",
            INIT_59 => X"000000ce00000000000000d300000000000000e700000000000000e300000000",
            INIT_5A => X"000000db00000000000000e100000000000000de00000000000000d600000000",
            INIT_5B => X"000000e900000000000000e600000000000000e100000000000000df00000000",
            INIT_5C => X"000000ed00000000000000f100000000000000ef00000000000000ed00000000",
            INIT_5D => X"000000ca00000000000000cf00000000000000cb00000000000000d000000000",
            INIT_5E => X"000000ca00000000000000a400000000000000c400000000000000d300000000",
            INIT_5F => X"000000ef00000000000000ef00000000000000ee00000000000000e900000000",
            INIT_60 => X"000000ea00000000000000e000000000000000d900000000000000de00000000",
            INIT_61 => X"000000ae00000000000000d000000000000000e300000000000000f100000000",
            INIT_62 => X"0000007900000000000000bc00000000000000d600000000000000b700000000",
            INIT_63 => X"00000093000000000000008b0000000000000084000000000000007e00000000",
            INIT_64 => X"000000ed00000000000000dc00000000000000ae00000000000000a100000000",
            INIT_65 => X"000000e900000000000000f000000000000000ee00000000000000eb00000000",
            INIT_66 => X"000000ed00000000000000d400000000000000e500000000000000ed00000000",
            INIT_67 => X"000000f200000000000000f200000000000000e900000000000000ea00000000",
            INIT_68 => X"00000097000000000000008d0000000000000093000000000000009800000000",
            INIT_69 => X"000000cc00000000000000cd00000000000000c100000000000000a500000000",
            INIT_6A => X"0000005c00000000000000b700000000000000ea00000000000000e200000000",
            INIT_6B => X"00000062000000000000005a000000000000005b000000000000005b00000000",
            INIT_6C => X"000000f100000000000000e900000000000000b3000000000000008100000000",
            INIT_6D => X"000000d900000000000000e900000000000000ed00000000000000f100000000",
            INIT_6E => X"000000d600000000000000df00000000000000dc00000000000000d400000000",
            INIT_6F => X"000000ea00000000000000e300000000000000cd00000000000000c400000000",
            INIT_70 => X"0000006600000000000000640000000000000072000000000000006c00000000",
            INIT_71 => X"000000cf00000000000000a400000000000000a4000000000000009b00000000",
            INIT_72 => X"0000008a00000000000000be00000000000000e400000000000000ea00000000",
            INIT_73 => X"000000cf00000000000000a80000000000000087000000000000008300000000",
            INIT_74 => X"000000d400000000000000e300000000000000e800000000000000df00000000",
            INIT_75 => X"0000009300000000000000a300000000000000ae00000000000000c300000000",
            INIT_76 => X"0000009700000000000000980000000000000090000000000000008c00000000",
            INIT_77 => X"000000d800000000000000cb00000000000000a0000000000000009300000000",
            INIT_78 => X"000000990000000000000074000000000000005e000000000000004d00000000",
            INIT_79 => X"000000a10000000000000076000000000000006e000000000000009c00000000",
            INIT_7A => X"000000c800000000000000c600000000000000c500000000000000b600000000",
            INIT_7B => X"000000d900000000000000ec00000000000000d900000000000000ca00000000",
            INIT_7C => X"00000095000000000000009f00000000000000ac00000000000000ba00000000",
            INIT_7D => X"0000007b0000000000000076000000000000007b000000000000008a00000000",
            INIT_7E => X"000000a100000000000000910000000000000082000000000000008000000000",
            INIT_7F => X"000000d000000000000000d500000000000000b800000000000000ae00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "sampleifmap_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000dc0000000000000097000000000000002f000000000000002300000000",
            INIT_01 => X"000000a20000000000000086000000000000007b000000000000009600000000",
            INIT_02 => X"000000e900000000000000e100000000000000d300000000000000b400000000",
            INIT_03 => X"000000be00000000000000ee00000000000000f000000000000000e800000000",
            INIT_04 => X"000000b100000000000000aa00000000000000a200000000000000a300000000",
            INIT_05 => X"000000bb00000000000000b600000000000000b600000000000000bb00000000",
            INIT_06 => X"000000d900000000000000cc00000000000000bf00000000000000bd00000000",
            INIT_07 => X"000000b700000000000000c100000000000000d000000000000000da00000000",
            INIT_08 => X"000000ef00000000000000d9000000000000004f000000000000001800000000",
            INIT_09 => X"000000e500000000000000da00000000000000d300000000000000d400000000",
            INIT_0A => X"000000ef00000000000000f500000000000000f600000000000000ed00000000",
            INIT_0B => X"000000ea00000000000000f100000000000000ef00000000000000dc00000000",
            INIT_0C => X"000000e500000000000000e600000000000000d600000000000000e400000000",
            INIT_0D => X"000000e000000000000000e800000000000000ea00000000000000e700000000",
            INIT_0E => X"000000b300000000000000c500000000000000d100000000000000d400000000",
            INIT_0F => X"000000a5000000000000009e00000000000000a100000000000000a900000000",
            INIT_10 => X"000000d800000000000000de00000000000000b3000000000000004700000000",
            INIT_11 => X"000000e300000000000000e600000000000000e500000000000000d900000000",
            INIT_12 => X"000000dd00000000000000e400000000000000e400000000000000e300000000",
            INIT_13 => X"000000bc00000000000000c100000000000000d700000000000000cf00000000",
            INIT_14 => X"0000009c00000000000000ba00000000000000c300000000000000b800000000",
            INIT_15 => X"0000009e00000000000000ad00000000000000b400000000000000a100000000",
            INIT_16 => X"0000008300000000000000850000000000000087000000000000008a00000000",
            INIT_17 => X"0000009c000000000000009e0000000000000097000000000000008c00000000",
            INIT_18 => X"000000bd00000000000000c200000000000000cf00000000000000a100000000",
            INIT_19 => X"000000c100000000000000c000000000000000be00000000000000bb00000000",
            INIT_1A => X"000000bd00000000000000bd00000000000000be00000000000000c000000000",
            INIT_1B => X"0000009a00000000000000a300000000000000ba00000000000000bc00000000",
            INIT_1C => X"0000009100000000000000a300000000000000aa000000000000009a00000000",
            INIT_1D => X"0000008800000000000000900000000000000099000000000000009400000000",
            INIT_1E => X"0000008d000000000000008b0000000000000086000000000000008200000000",
            INIT_1F => X"0000009c00000000000000940000000000000092000000000000009000000000",
            INIT_20 => X"0000007f000000000000007a0000000000000071000000000000006d00000000",
            INIT_21 => X"000000960000000000000093000000000000008e000000000000008600000000",
            INIT_22 => X"000000ac00000000000000a500000000000000a0000000000000009800000000",
            INIT_23 => X"000000af00000000000000b400000000000000ba00000000000000b500000000",
            INIT_24 => X"0000009b00000000000000a300000000000000a800000000000000ac00000000",
            INIT_25 => X"0000007f0000000000000084000000000000008b000000000000009400000000",
            INIT_26 => X"0000007a00000000000000810000000000000085000000000000008100000000",
            INIT_27 => X"0000009c0000000000000092000000000000008a000000000000007e00000000",
            INIT_28 => X"0000003000000000000000230000000000000019000000000000002900000000",
            INIT_29 => X"0000003d000000000000003a0000000000000038000000000000003400000000",
            INIT_2A => X"00000057000000000000004d0000000000000046000000000000003e00000000",
            INIT_2B => X"0000007e000000000000007e0000000000000079000000000000006a00000000",
            INIT_2C => X"000000700000000000000078000000000000007e000000000000007f00000000",
            INIT_2D => X"0000006600000000000000670000000000000068000000000000006a00000000",
            INIT_2E => X"000000770000000000000073000000000000006e000000000000006900000000",
            INIT_2F => X"00000095000000000000008d0000000000000088000000000000008000000000",
            INIT_30 => X"0000003500000000000000130000000000000014000000000000003700000000",
            INIT_31 => X"00000018000000000000001e0000000000000029000000000000003a00000000",
            INIT_32 => X"00000014000000000000000f000000000000000f000000000000001100000000",
            INIT_33 => X"0000003e000000000000003c0000000000000038000000000000002a00000000",
            INIT_34 => X"0000004c000000000000004d0000000000000051000000000000004700000000",
            INIT_35 => X"0000005a0000000000000053000000000000004f000000000000004e00000000",
            INIT_36 => X"0000008a000000000000008a0000000000000076000000000000006500000000",
            INIT_37 => X"0000009e00000000000000890000000000000080000000000000007d00000000",
            INIT_38 => X"000000290000000000000012000000000000001a000000000000002d00000000",
            INIT_39 => X"000000250000000000000039000000000000004c000000000000005400000000",
            INIT_3A => X"000000070000000000000007000000000000000b000000000000001500000000",
            INIT_3B => X"0000003e000000000000004e000000000000005b000000000000002300000000",
            INIT_3C => X"00000045000000000000003f000000000000003e000000000000003c00000000",
            INIT_3D => X"0000007b00000000000000630000000000000053000000000000004a00000000",
            INIT_3E => X"0000007200000000000000870000000000000095000000000000009200000000",
            INIT_3F => X"000000af00000000000000920000000000000085000000000000007400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000b00000000000000080000000000000009000000000000001100000000",
            INIT_41 => X"00000023000000000000002f0000000000000039000000000000002e00000000",
            INIT_42 => X"0000000300000000000000040000000000000007000000000000001400000000",
            INIT_43 => X"0000009400000000000000b30000000000000086000000000000000f00000000",
            INIT_44 => X"0000007f000000000000007c000000000000007d000000000000008300000000",
            INIT_45 => X"0000008d00000000000000900000000000000085000000000000007e00000000",
            INIT_46 => X"000000740000000000000061000000000000005b000000000000007400000000",
            INIT_47 => X"000000be00000000000000a50000000000000090000000000000008100000000",
            INIT_48 => X"0000000400000000000000030000000000000007000000000000002300000000",
            INIT_49 => X"0000000c00000000000000110000000000000011000000000000000700000000",
            INIT_4A => X"0000000300000000000000020000000000000003000000000000000700000000",
            INIT_4B => X"0000009400000000000000920000000000000040000000000000000200000000",
            INIT_4C => X"000000810000000000000089000000000000008d000000000000009000000000",
            INIT_4D => X"000000450000000000000053000000000000006a000000000000007a00000000",
            INIT_4E => X"0000007e00000000000000710000000000000058000000000000004600000000",
            INIT_4F => X"000000c200000000000000b0000000000000009e000000000000008700000000",
            INIT_50 => X"0000000200000000000000010000000000000015000000000000004000000000",
            INIT_51 => X"0000000500000000000000090000000000000005000000000000000000000000",
            INIT_52 => X"0000000100000000000000000000000000000000000000000000000200000000",
            INIT_53 => X"00000044000000000000003b000000000000000b000000000000000100000000",
            INIT_54 => X"0000003b00000000000000430000000000000045000000000000004300000000",
            INIT_55 => X"00000047000000000000002e000000000000002a000000000000003100000000",
            INIT_56 => X"0000008000000000000000780000000000000074000000000000006600000000",
            INIT_57 => X"000000c400000000000000b700000000000000ab000000000000009300000000",
            INIT_58 => X"000000020000000000000001000000000000002b000000000000005200000000",
            INIT_59 => X"0000000200000000000000050000000000000002000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000003600000000000000260000000000000002000000000000000000000000",
            INIT_5C => X"000000220000000000000024000000000000002b000000000000002e00000000",
            INIT_5D => X"0000006900000000000000520000000000000038000000000000002700000000",
            INIT_5E => X"0000008300000000000000760000000000000073000000000000007300000000",
            INIT_5F => X"000000c700000000000000bb00000000000000ae000000000000009600000000",
            INIT_60 => X"0000000100000000000000030000000000000032000000000000005d00000000",
            INIT_61 => X"0000000200000000000000030000000000000001000000000000000000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000100000000",
            INIT_63 => X"0000002f000000000000001c0000000000000000000000000000000200000000",
            INIT_64 => X"000000370000000000000016000000000000000c000000000000001700000000",
            INIT_65 => X"00000070000000000000006f0000000000000063000000000000005100000000",
            INIT_66 => X"00000089000000000000007e0000000000000077000000000000007100000000",
            INIT_67 => X"000000c900000000000000bc00000000000000ab000000000000009700000000",
            INIT_68 => X"00000004000000000000000b0000000000000025000000000000005900000000",
            INIT_69 => X"0000000200000000000000040000000000000004000000000000000200000000",
            INIT_6A => X"0000000200000000000000010000000000000001000000000000000100000000",
            INIT_6B => X"00000018000000000000000d0000000000000002000000000000000600000000",
            INIT_6C => X"00000052000000000000003e0000000000000029000000000000001900000000",
            INIT_6D => X"0000006f00000000000000700000000000000071000000000000006500000000",
            INIT_6E => X"000000910000000000000089000000000000007e000000000000007300000000",
            INIT_6F => X"000000c900000000000000c100000000000000b300000000000000a100000000",
            INIT_70 => X"0000001100000000000000160000000000000024000000000000005200000000",
            INIT_71 => X"0000000c000000000000000d000000000000000f000000000000000f00000000",
            INIT_72 => X"0000000f000000000000000e000000000000000d000000000000000c00000000",
            INIT_73 => X"0000002d000000000000001b0000000000000015000000000000001400000000",
            INIT_74 => X"0000005800000000000000550000000000000051000000000000004300000000",
            INIT_75 => X"00000070000000000000006b000000000000006e000000000000006900000000",
            INIT_76 => X"00000097000000000000008a000000000000007f000000000000007700000000",
            INIT_77 => X"000000c800000000000000c400000000000000b700000000000000a400000000",
            INIT_78 => X"0000002500000000000000260000000000000030000000000000005300000000",
            INIT_79 => X"0000002600000000000000220000000000000021000000000000002300000000",
            INIT_7A => X"0000002e000000000000002c0000000000000029000000000000002800000000",
            INIT_7B => X"0000004a000000000000003b0000000000000030000000000000002d00000000",
            INIT_7C => X"000000610000000000000061000000000000005c000000000000005300000000",
            INIT_7D => X"00000075000000000000006c000000000000006a000000000000006b00000000",
            INIT_7E => X"00000099000000000000008d0000000000000085000000000000007b00000000",
            INIT_7F => X"000000c700000000000000bf00000000000000b200000000000000a300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "sampleifmap_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000084000000000000008b000000000000009e000000000000009e00000000",
            INIT_01 => X"000000c100000000000000bb00000000000000b600000000000000a600000000",
            INIT_02 => X"000000ce00000000000000d100000000000000cd00000000000000c700000000",
            INIT_03 => X"000000e600000000000000e300000000000000df00000000000000da00000000",
            INIT_04 => X"000000eb00000000000000e700000000000000e200000000000000d500000000",
            INIT_05 => X"000000ea00000000000000ea00000000000000e800000000000000ec00000000",
            INIT_06 => X"000000ee00000000000000e600000000000000e200000000000000ec00000000",
            INIT_07 => X"000000ee00000000000000ed00000000000000e400000000000000e800000000",
            INIT_08 => X"00000089000000000000009700000000000000ac00000000000000aa00000000",
            INIT_09 => X"000000c700000000000000c500000000000000c100000000000000ae00000000",
            INIT_0A => X"000000d200000000000000d900000000000000d700000000000000ce00000000",
            INIT_0B => X"000000ed00000000000000e900000000000000e700000000000000e100000000",
            INIT_0C => X"000000f200000000000000e800000000000000e400000000000000db00000000",
            INIT_0D => X"000000f200000000000000ec00000000000000ea00000000000000f500000000",
            INIT_0E => X"000000f300000000000000eb00000000000000e400000000000000f100000000",
            INIT_0F => X"000000f600000000000000f600000000000000e800000000000000e900000000",
            INIT_10 => X"0000008e000000000000009d00000000000000b000000000000000ae00000000",
            INIT_11 => X"000000c700000000000000ce00000000000000c900000000000000b500000000",
            INIT_12 => X"000000d400000000000000da00000000000000df00000000000000d100000000",
            INIT_13 => X"000000ef00000000000000e600000000000000e600000000000000e000000000",
            INIT_14 => X"000000ef00000000000000e900000000000000e400000000000000dd00000000",
            INIT_15 => X"000000f300000000000000ec00000000000000d500000000000000e800000000",
            INIT_16 => X"000000f800000000000000ee00000000000000e700000000000000f500000000",
            INIT_17 => X"000000f500000000000000fa00000000000000e600000000000000ed00000000",
            INIT_18 => X"0000009300000000000000a000000000000000b200000000000000b400000000",
            INIT_19 => X"000000cf00000000000000d400000000000000cb00000000000000ba00000000",
            INIT_1A => X"000000d600000000000000dd00000000000000e400000000000000d600000000",
            INIT_1B => X"000000f000000000000000df00000000000000e700000000000000dc00000000",
            INIT_1C => X"000000e400000000000000e900000000000000e400000000000000e000000000",
            INIT_1D => X"000000f300000000000000e600000000000000ac00000000000000b100000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f400000000000000f900000000000000e400000000000000ee00000000",
            INIT_20 => X"0000009300000000000000a500000000000000b900000000000000ba00000000",
            INIT_21 => X"000000cf00000000000000d900000000000000cc00000000000000bd00000000",
            INIT_22 => X"000000d600000000000000de00000000000000e700000000000000d300000000",
            INIT_23 => X"000000eb00000000000000d300000000000000e700000000000000da00000000",
            INIT_24 => X"000000d400000000000000e800000000000000e000000000000000e200000000",
            INIT_25 => X"000000ed00000000000000e000000000000000a8000000000000009f00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f200000000000000f800000000000000ea00000000000000e800000000",
            INIT_28 => X"0000008e00000000000000aa00000000000000be00000000000000c100000000",
            INIT_29 => X"000000d300000000000000db00000000000000cb00000000000000bf00000000",
            INIT_2A => X"000000d600000000000000dd00000000000000ea00000000000000d700000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e400000000000000d600000000",
            INIT_2C => X"000000c100000000000000eb00000000000000ce00000000000000cf00000000",
            INIT_2D => X"000000e600000000000000de000000000000009e000000000000007000000000",
            INIT_2E => X"000000f100000000000000e200000000000000e500000000000000f500000000",
            INIT_2F => X"000000eb00000000000000f300000000000000e700000000000000e400000000",
            INIT_30 => X"0000008500000000000000ac00000000000000bf00000000000000c400000000",
            INIT_31 => X"000000d900000000000000de00000000000000ca00000000000000bf00000000",
            INIT_32 => X"000000d600000000000000da00000000000000eb00000000000000df00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e300000000000000d700000000",
            INIT_34 => X"000000bb00000000000000cd00000000000000ba00000000000000bb00000000",
            INIT_35 => X"000000b700000000000000ac0000000000000089000000000000007800000000",
            INIT_36 => X"000000eb00000000000000d800000000000000df00000000000000db00000000",
            INIT_37 => X"000000eb00000000000000f000000000000000e100000000000000e200000000",
            INIT_38 => X"0000008c00000000000000ae00000000000000c500000000000000cc00000000",
            INIT_39 => X"000000e000000000000000e000000000000000da00000000000000cb00000000",
            INIT_3A => X"000000dc00000000000000dc00000000000000ed00000000000000e800000000",
            INIT_3B => X"000000cd00000000000000c900000000000000dd00000000000000dc00000000",
            INIT_3C => X"000000530000000000000064000000000000008a00000000000000ac00000000",
            INIT_3D => X"0000003c0000000000000041000000000000003e000000000000004700000000",
            INIT_3E => X"000000e400000000000000d100000000000000b6000000000000006800000000",
            INIT_3F => X"000000ec00000000000000ef00000000000000d400000000000000da00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000089000000000000009d00000000000000aa00000000000000af00000000",
            INIT_41 => X"000000c500000000000000af00000000000000ba00000000000000b000000000",
            INIT_42 => X"000000d200000000000000ce00000000000000d400000000000000d100000000",
            INIT_43 => X"000000c100000000000000c100000000000000c900000000000000d400000000",
            INIT_44 => X"0000005b00000000000000590000000000000069000000000000008e00000000",
            INIT_45 => X"00000045000000000000005e0000000000000053000000000000005400000000",
            INIT_46 => X"000000b700000000000000a20000000000000079000000000000004e00000000",
            INIT_47 => X"000000c300000000000000cf00000000000000a300000000000000ae00000000",
            INIT_48 => X"0000006800000000000000710000000000000073000000000000007200000000",
            INIT_49 => X"00000080000000000000006f000000000000006b000000000000006900000000",
            INIT_4A => X"0000009b00000000000000970000000000000092000000000000008b00000000",
            INIT_4B => X"0000009600000000000000970000000000000093000000000000009d00000000",
            INIT_4C => X"0000006300000000000000630000000000000064000000000000007600000000",
            INIT_4D => X"0000005300000000000000560000000000000056000000000000005500000000",
            INIT_4E => X"00000099000000000000009a0000000000000080000000000000008b00000000",
            INIT_4F => X"0000007b0000000000000084000000000000006d000000000000007600000000",
            INIT_50 => X"00000044000000000000004b000000000000004c000000000000004200000000",
            INIT_51 => X"0000005a0000000000000054000000000000005a000000000000005300000000",
            INIT_52 => X"000000670000000000000066000000000000006a000000000000005d00000000",
            INIT_53 => X"0000006c0000000000000072000000000000006b000000000000006a00000000",
            INIT_54 => X"00000055000000000000005b000000000000005a000000000000005a00000000",
            INIT_55 => X"00000072000000000000005f0000000000000042000000000000004800000000",
            INIT_56 => X"000000c70000000000000093000000000000006e000000000000008000000000",
            INIT_57 => X"0000005e000000000000005c0000000000000067000000000000007d00000000",
            INIT_58 => X"0000004d000000000000004b0000000000000041000000000000003500000000",
            INIT_59 => X"000000460000000000000055000000000000006a000000000000006f00000000",
            INIT_5A => X"0000005d000000000000005f0000000000000071000000000000005d00000000",
            INIT_5B => X"00000061000000000000006b0000000000000073000000000000006c00000000",
            INIT_5C => X"000000610000000000000062000000000000005f000000000000006200000000",
            INIT_5D => X"000000bb00000000000000950000000000000055000000000000005a00000000",
            INIT_5E => X"000000cc0000000000000070000000000000009200000000000000b300000000",
            INIT_5F => X"000000550000000000000057000000000000005f000000000000009a00000000",
            INIT_60 => X"0000004a000000000000005e0000000000000056000000000000003a00000000",
            INIT_61 => X"00000055000000000000004d0000000000000064000000000000006400000000",
            INIT_62 => X"0000006c000000000000007f0000000000000085000000000000007800000000",
            INIT_63 => X"000000570000000000000062000000000000006e000000000000006900000000",
            INIT_64 => X"0000005f00000000000000570000000000000051000000000000005100000000",
            INIT_65 => X"000000c300000000000000aa0000000000000070000000000000005f00000000",
            INIT_66 => X"000000ad000000000000007f00000000000000c100000000000000d000000000",
            INIT_67 => X"0000004f0000000000000055000000000000005000000000000000b200000000",
            INIT_68 => X"0000004b00000000000000570000000000000059000000000000004a00000000",
            INIT_69 => X"0000005000000000000000470000000000000044000000000000005200000000",
            INIT_6A => X"0000006f00000000000000760000000000000067000000000000005900000000",
            INIT_6B => X"000000620000000000000069000000000000006a000000000000006500000000",
            INIT_6C => X"0000006d00000000000000620000000000000062000000000000006000000000",
            INIT_6D => X"000000b800000000000000b4000000000000008e000000000000007200000000",
            INIT_6E => X"0000008400000000000000a000000000000000c000000000000000bf00000000",
            INIT_6F => X"00000043000000000000003c000000000000005000000000000000aa00000000",
            INIT_70 => X"0000004e0000000000000052000000000000004f000000000000004d00000000",
            INIT_71 => X"0000005600000000000000460000000000000048000000000000004f00000000",
            INIT_72 => X"0000008500000000000000810000000000000079000000000000006d00000000",
            INIT_73 => X"0000008300000000000000870000000000000088000000000000008900000000",
            INIT_74 => X"0000009600000000000000920000000000000094000000000000009200000000",
            INIT_75 => X"000000b500000000000000b300000000000000a3000000000000009400000000",
            INIT_76 => X"0000006500000000000000aa00000000000000b000000000000000b900000000",
            INIT_77 => X"0000003b00000000000000370000000000000049000000000000005a00000000",
            INIT_78 => X"00000068000000000000006a000000000000005e000000000000006000000000",
            INIT_79 => X"0000008a00000000000000840000000000000083000000000000006d00000000",
            INIT_7A => X"0000009a000000000000009b0000000000000098000000000000009000000000",
            INIT_7B => X"00000094000000000000009e000000000000009b000000000000009b00000000",
            INIT_7C => X"00000092000000000000009c000000000000009d000000000000009600000000",
            INIT_7D => X"000000a900000000000000920000000000000082000000000000007700000000",
            INIT_7E => X"0000006900000000000000a700000000000000a800000000000000b100000000",
            INIT_7F => X"0000004800000000000000560000000000000062000000000000004500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "sampleifmap_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000008300000000000000730000000000000065000000000000006a00000000",
            INIT_01 => X"0000008f00000000000000900000000000000087000000000000008100000000",
            INIT_02 => X"0000009a000000000000009a0000000000000096000000000000009200000000",
            INIT_03 => X"0000009000000000000000970000000000000099000000000000009a00000000",
            INIT_04 => X"0000007f000000000000008b0000000000000086000000000000008200000000",
            INIT_05 => X"0000009f00000000000000920000000000000075000000000000005e00000000",
            INIT_06 => X"0000008400000000000000a200000000000000a300000000000000a700000000",
            INIT_07 => X"00000069000000000000009a00000000000000c0000000000000009000000000",
            INIT_08 => X"0000006d0000000000000076000000000000006c000000000000005f00000000",
            INIT_09 => X"000000910000000000000081000000000000005d000000000000005f00000000",
            INIT_0A => X"0000009000000000000000960000000000000097000000000000009500000000",
            INIT_0B => X"0000007b000000000000007a000000000000007e000000000000008600000000",
            INIT_0C => X"00000094000000000000009b0000000000000085000000000000007a00000000",
            INIT_0D => X"0000009c00000000000000a20000000000000093000000000000008300000000",
            INIT_0E => X"0000009500000000000000990000000000000097000000000000009d00000000",
            INIT_0F => X"00000094000000000000009d00000000000000a4000000000000009f00000000",
            INIT_10 => X"0000004600000000000000490000000000000059000000000000006600000000",
            INIT_11 => X"0000008c000000000000007b000000000000006f000000000000005600000000",
            INIT_12 => X"0000007500000000000000780000000000000081000000000000008f00000000",
            INIT_13 => X"0000008d0000000000000085000000000000007e000000000000007800000000",
            INIT_14 => X"0000009f0000000000000099000000000000008e000000000000009600000000",
            INIT_15 => X"000000a100000000000000a5000000000000009d000000000000009700000000",
            INIT_16 => X"00000090000000000000009a0000000000000098000000000000009900000000",
            INIT_17 => X"00000095000000000000007d0000000000000079000000000000008300000000",
            INIT_18 => X"0000006e0000000000000047000000000000003d000000000000005600000000",
            INIT_19 => X"0000007b0000000000000082000000000000008a000000000000008000000000",
            INIT_1A => X"000000840000000000000076000000000000006c000000000000007600000000",
            INIT_1B => X"00000099000000000000009c0000000000000098000000000000008f00000000",
            INIT_1C => X"0000009a00000000000000910000000000000089000000000000009500000000",
            INIT_1D => X"000000a400000000000000a0000000000000009a000000000000009900000000",
            INIT_1E => X"00000069000000000000007d0000000000000090000000000000009800000000",
            INIT_1F => X"000000840000000000000056000000000000004b000000000000005c00000000",
            INIT_20 => X"00000072000000000000006b0000000000000067000000000000006800000000",
            INIT_21 => X"00000076000000000000007b0000000000000074000000000000007300000000",
            INIT_22 => X"00000090000000000000008d0000000000000086000000000000007400000000",
            INIT_23 => X"000000750000000000000085000000000000008d000000000000008f00000000",
            INIT_24 => X"0000009600000000000000820000000000000059000000000000006200000000",
            INIT_25 => X"000000910000000000000098000000000000009a000000000000009700000000",
            INIT_26 => X"00000050000000000000005a0000000000000060000000000000007500000000",
            INIT_27 => X"0000004100000000000000490000000000000047000000000000004100000000",
            INIT_28 => X"0000006f000000000000006f000000000000006b000000000000006300000000",
            INIT_29 => X"0000007e000000000000007d0000000000000077000000000000007200000000",
            INIT_2A => X"00000081000000000000007d000000000000007d000000000000007500000000",
            INIT_2B => X"0000003d000000000000005b0000000000000082000000000000008300000000",
            INIT_2C => X"0000009400000000000000730000000000000038000000000000003900000000",
            INIT_2D => X"0000005f00000000000000720000000000000082000000000000008b00000000",
            INIT_2E => X"0000003a00000000000000490000000000000053000000000000005600000000",
            INIT_2F => X"0000001b0000000000000033000000000000004b000000000000003c00000000",
            INIT_30 => X"0000007200000000000000740000000000000068000000000000003e00000000",
            INIT_31 => X"0000005b00000000000000660000000000000075000000000000007400000000",
            INIT_32 => X"00000070000000000000004e0000000000000051000000000000005400000000",
            INIT_33 => X"0000004c00000000000000600000000000000082000000000000008500000000",
            INIT_34 => X"0000006c000000000000006b0000000000000056000000000000005300000000",
            INIT_35 => X"0000005100000000000000530000000000000058000000000000006000000000",
            INIT_36 => X"0000002d0000000000000033000000000000003d000000000000004600000000",
            INIT_37 => X"00000018000000000000001e000000000000002e000000000000003400000000",
            INIT_38 => X"00000069000000000000006a0000000000000060000000000000003900000000",
            INIT_39 => X"0000003500000000000000410000000000000068000000000000006b00000000",
            INIT_3A => X"0000006e00000000000000440000000000000040000000000000003b00000000",
            INIT_3B => X"0000006200000000000000730000000000000085000000000000008700000000",
            INIT_3C => X"00000050000000000000004e000000000000004f000000000000005800000000",
            INIT_3D => X"0000003700000000000000460000000000000050000000000000005100000000",
            INIT_3E => X"00000029000000000000002d0000000000000031000000000000002c00000000",
            INIT_3F => X"00000018000000000000001b000000000000001e000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000068000000000000005a000000000000004100000000",
            INIT_41 => X"00000049000000000000004f000000000000006d000000000000006d00000000",
            INIT_42 => X"0000006a00000000000000620000000000000058000000000000005500000000",
            INIT_43 => X"0000004100000000000000440000000000000053000000000000006200000000",
            INIT_44 => X"000000520000000000000051000000000000004a000000000000004600000000",
            INIT_45 => X"0000002c00000000000000290000000000000033000000000000004800000000",
            INIT_46 => X"0000002300000000000000270000000000000037000000000000003d00000000",
            INIT_47 => X"00000019000000000000001b000000000000001e000000000000002000000000",
            INIT_48 => X"0000006700000000000000690000000000000057000000000000004300000000",
            INIT_49 => X"0000005100000000000000580000000000000063000000000000006600000000",
            INIT_4A => X"00000039000000000000003b0000000000000045000000000000004c00000000",
            INIT_4B => X"000000460000000000000042000000000000003f000000000000003a00000000",
            INIT_4C => X"00000036000000000000003e0000000000000044000000000000004800000000",
            INIT_4D => X"0000002c0000000000000031000000000000002f000000000000002e00000000",
            INIT_4E => X"0000001c000000000000001e000000000000002e000000000000003800000000",
            INIT_4F => X"0000001e00000000000000180000000000000019000000000000001d00000000",
            INIT_50 => X"0000003a0000000000000041000000000000003a000000000000003600000000",
            INIT_51 => X"0000002c000000000000002d0000000000000032000000000000003700000000",
            INIT_52 => X"0000003a00000000000000370000000000000033000000000000002e00000000",
            INIT_53 => X"0000003a000000000000003e0000000000000040000000000000003e00000000",
            INIT_54 => X"0000003000000000000000250000000000000026000000000000003300000000",
            INIT_55 => X"00000026000000000000002a0000000000000030000000000000003100000000",
            INIT_56 => X"0000001c000000000000001b0000000000000020000000000000002900000000",
            INIT_57 => X"0000001f000000000000001c0000000000000019000000000000001b00000000",
            INIT_58 => X"0000001b000000000000001a000000000000001d000000000000001e00000000",
            INIT_59 => X"0000002700000000000000210000000000000020000000000000001f00000000",
            INIT_5A => X"0000003300000000000000350000000000000034000000000000003100000000",
            INIT_5B => X"0000002800000000000000260000000000000028000000000000002e00000000",
            INIT_5C => X"000000370000000000000042000000000000002c000000000000002600000000",
            INIT_5D => X"0000002500000000000000240000000000000025000000000000002900000000",
            INIT_5E => X"0000001b000000000000001a000000000000001b000000000000001f00000000",
            INIT_5F => X"000000170000000000000021000000000000001e000000000000001c00000000",
            INIT_60 => X"0000001c000000000000001b000000000000001f000000000000002100000000",
            INIT_61 => X"00000020000000000000001f000000000000001e000000000000001c00000000",
            INIT_62 => X"0000001e000000000000001e0000000000000021000000000000002300000000",
            INIT_63 => X"0000002d00000000000000290000000000000027000000000000002200000000",
            INIT_64 => X"0000003100000000000000490000000000000034000000000000002a00000000",
            INIT_65 => X"0000002000000000000000260000000000000023000000000000001e00000000",
            INIT_66 => X"0000001d000000000000001b000000000000001a000000000000001b00000000",
            INIT_67 => X"0000000d000000000000001a0000000000000026000000000000001e00000000",
            INIT_68 => X"0000001a000000000000001a000000000000001e000000000000001f00000000",
            INIT_69 => X"0000001b000000000000001a0000000000000019000000000000001900000000",
            INIT_6A => X"0000002800000000000000250000000000000020000000000000001d00000000",
            INIT_6B => X"0000002a00000000000000280000000000000029000000000000002a00000000",
            INIT_6C => X"000000260000000000000040000000000000002e000000000000002700000000",
            INIT_6D => X"0000001d000000000000001e0000000000000024000000000000001c00000000",
            INIT_6E => X"0000001c000000000000001b0000000000000019000000000000001a00000000",
            INIT_6F => X"0000000400000000000000090000000000000025000000000000002100000000",
            INIT_70 => X"0000001c0000000000000019000000000000001b000000000000001700000000",
            INIT_71 => X"0000002500000000000000220000000000000020000000000000001e00000000",
            INIT_72 => X"0000002700000000000000280000000000000027000000000000002700000000",
            INIT_73 => X"00000021000000000000001e0000000000000023000000000000002600000000",
            INIT_74 => X"0000002400000000000000390000000000000024000000000000001c00000000",
            INIT_75 => X"0000001d000000000000001d000000000000001d000000000000001e00000000",
            INIT_76 => X"0000001b00000000000000170000000000000018000000000000001800000000",
            INIT_77 => X"0000000500000000000000040000000000000013000000000000002400000000",
            INIT_78 => X"000000220000000000000020000000000000001e000000000000001c00000000",
            INIT_79 => X"0000002500000000000000230000000000000022000000000000002100000000",
            INIT_7A => X"0000002200000000000000240000000000000026000000000000002600000000",
            INIT_7B => X"0000000c000000000000000f0000000000000018000000000000001e00000000",
            INIT_7C => X"00000020000000000000002d0000000000000013000000000000000800000000",
            INIT_7D => X"0000001c000000000000001b000000000000001b000000000000001900000000",
            INIT_7E => X"0000002200000000000000140000000000000015000000000000001800000000",
            INIT_7F => X"0000000700000000000000040000000000000005000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "sampleifmap_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009e00000000000000a600000000000000bb00000000000000be00000000",
            INIT_01 => X"000000d800000000000000d300000000000000d000000000000000c100000000",
            INIT_02 => X"000000da00000000000000de00000000000000dd00000000000000db00000000",
            INIT_03 => X"000000ed00000000000000eb00000000000000e800000000000000e500000000",
            INIT_04 => X"000000ef00000000000000ee00000000000000e900000000000000dc00000000",
            INIT_05 => X"000000f100000000000000f100000000000000ef00000000000000f100000000",
            INIT_06 => X"000000f300000000000000eb00000000000000e700000000000000f200000000",
            INIT_07 => X"000000f100000000000000ef00000000000000e700000000000000ed00000000",
            INIT_08 => X"000000a000000000000000b000000000000000c700000000000000c800000000",
            INIT_09 => X"000000da00000000000000da00000000000000d900000000000000c700000000",
            INIT_0A => X"000000db00000000000000e500000000000000e500000000000000df00000000",
            INIT_0B => X"000000f300000000000000ef00000000000000ee00000000000000e900000000",
            INIT_0C => X"000000f500000000000000ee00000000000000ea00000000000000e100000000",
            INIT_0D => X"000000f500000000000000ef00000000000000ed00000000000000f700000000",
            INIT_0E => X"000000f800000000000000ef00000000000000e900000000000000f500000000",
            INIT_0F => X"000000f700000000000000f600000000000000e800000000000000ec00000000",
            INIT_10 => X"000000a200000000000000b300000000000000c800000000000000c900000000",
            INIT_11 => X"000000d600000000000000df00000000000000dc00000000000000c900000000",
            INIT_12 => X"000000db00000000000000e200000000000000e900000000000000dd00000000",
            INIT_13 => X"000000f400000000000000ea00000000000000ea00000000000000e500000000",
            INIT_14 => X"000000f300000000000000ee00000000000000e900000000000000e200000000",
            INIT_15 => X"000000f100000000000000ea00000000000000d600000000000000eb00000000",
            INIT_16 => X"000000fa00000000000000f000000000000000e900000000000000f700000000",
            INIT_17 => X"000000f400000000000000f900000000000000e500000000000000ee00000000",
            INIT_18 => X"000000a400000000000000b300000000000000c700000000000000cb00000000",
            INIT_19 => X"000000d900000000000000e100000000000000d900000000000000c900000000",
            INIT_1A => X"000000d900000000000000e300000000000000eb00000000000000df00000000",
            INIT_1B => X"000000f400000000000000e200000000000000e800000000000000dd00000000",
            INIT_1C => X"000000eb00000000000000ed00000000000000e700000000000000e400000000",
            INIT_1D => X"000000f100000000000000e400000000000000af00000000000000b800000000",
            INIT_1E => X"000000fa00000000000000ee00000000000000e800000000000000f800000000",
            INIT_1F => X"000000f200000000000000f700000000000000e300000000000000ed00000000",
            INIT_20 => X"000000a100000000000000b500000000000000cc00000000000000cf00000000",
            INIT_21 => X"000000d500000000000000e100000000000000d600000000000000c900000000",
            INIT_22 => X"000000d700000000000000e200000000000000ed00000000000000d700000000",
            INIT_23 => X"000000ec00000000000000d400000000000000e500000000000000d900000000",
            INIT_24 => X"000000e100000000000000ec00000000000000e100000000000000e300000000",
            INIT_25 => X"000000ec00000000000000e000000000000000ae00000000000000aa00000000",
            INIT_26 => X"000000f600000000000000eb00000000000000e700000000000000f700000000",
            INIT_27 => X"000000ef00000000000000f500000000000000e700000000000000e700000000",
            INIT_28 => X"0000009a00000000000000b700000000000000cd00000000000000d000000000",
            INIT_29 => X"000000d700000000000000e200000000000000d400000000000000c900000000",
            INIT_2A => X"000000d700000000000000df00000000000000ee00000000000000da00000000",
            INIT_2B => X"000000cd00000000000000c700000000000000e500000000000000d700000000",
            INIT_2C => X"000000cc00000000000000ef00000000000000d000000000000000d100000000",
            INIT_2D => X"000000e900000000000000e300000000000000a7000000000000007c00000000",
            INIT_2E => X"000000ef00000000000000e100000000000000e500000000000000f600000000",
            INIT_2F => X"000000e800000000000000f100000000000000e600000000000000e200000000",
            INIT_30 => X"0000008b00000000000000b300000000000000c700000000000000cc00000000",
            INIT_31 => X"000000d500000000000000dd00000000000000cb00000000000000c200000000",
            INIT_32 => X"000000d400000000000000d800000000000000e900000000000000db00000000",
            INIT_33 => X"000000b000000000000000bc00000000000000e600000000000000d800000000",
            INIT_34 => X"000000c000000000000000d400000000000000c000000000000000be00000000",
            INIT_35 => X"000000be00000000000000b70000000000000097000000000000008100000000",
            INIT_36 => X"000000e500000000000000d600000000000000e000000000000000e000000000",
            INIT_37 => X"000000e000000000000000eb00000000000000de00000000000000db00000000",
            INIT_38 => X"0000008a00000000000000af00000000000000c600000000000000cd00000000",
            INIT_39 => X"000000cc00000000000000ce00000000000000cb00000000000000c000000000",
            INIT_3A => X"000000d200000000000000d000000000000000df00000000000000d400000000",
            INIT_3B => X"000000ce00000000000000c700000000000000d800000000000000d500000000",
            INIT_3C => X"0000005d0000000000000071000000000000009500000000000000b200000000",
            INIT_3D => X"0000004500000000000000500000000000000050000000000000005500000000",
            INIT_3E => X"000000de00000000000000ce00000000000000b7000000000000006c00000000",
            INIT_3F => X"000000d400000000000000dd00000000000000c500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000085000000000000009a00000000000000a800000000000000ad00000000",
            INIT_41 => X"000000b300000000000000a000000000000000ac00000000000000a500000000",
            INIT_42 => X"000000c300000000000000bd00000000000000c200000000000000be00000000",
            INIT_43 => X"000000c600000000000000c100000000000000bf00000000000000c700000000",
            INIT_44 => X"0000006c000000000000006b0000000000000079000000000000009800000000",
            INIT_45 => X"0000004f000000000000006e0000000000000068000000000000006800000000",
            INIT_46 => X"000000af000000000000009f000000000000007a000000000000005200000000",
            INIT_47 => X"000000af00000000000000be000000000000009500000000000000a300000000",
            INIT_48 => X"0000006900000000000000720000000000000074000000000000007300000000",
            INIT_49 => X"0000007f0000000000000070000000000000006e000000000000006d00000000",
            INIT_4A => X"00000093000000000000008c0000000000000088000000000000008700000000",
            INIT_4B => X"000000a1000000000000009e000000000000008f000000000000009700000000",
            INIT_4C => X"0000007800000000000000780000000000000077000000000000008600000000",
            INIT_4D => X"0000005c0000000000000066000000000000006c000000000000006c00000000",
            INIT_4E => X"0000009100000000000000970000000000000080000000000000008f00000000",
            INIT_4F => X"000000780000000000000082000000000000006a000000000000006e00000000",
            INIT_50 => X"0000005200000000000000560000000000000057000000000000004e00000000",
            INIT_51 => X"0000006400000000000000610000000000000069000000000000006300000000",
            INIT_52 => X"0000006f000000000000006a000000000000006d000000000000006500000000",
            INIT_53 => X"0000007f00000000000000840000000000000076000000000000007200000000",
            INIT_54 => X"0000006b000000000000006e000000000000006d000000000000006d00000000",
            INIT_55 => X"00000077000000000000006c0000000000000057000000000000006000000000",
            INIT_56 => X"000000bf0000000000000090000000000000006f000000000000008400000000",
            INIT_57 => X"000000680000000000000066000000000000006f000000000000007800000000",
            INIT_58 => X"00000062000000000000005f0000000000000055000000000000004a00000000",
            INIT_59 => X"000000510000000000000062000000000000007a000000000000008000000000",
            INIT_5A => X"0000007300000000000000710000000000000081000000000000006800000000",
            INIT_5B => X"0000007b0000000000000086000000000000008b000000000000008400000000",
            INIT_5C => X"0000007700000000000000740000000000000073000000000000007800000000",
            INIT_5D => X"000000bd000000000000009e0000000000000068000000000000007100000000",
            INIT_5E => X"000000c5000000000000006d000000000000009400000000000000b700000000",
            INIT_5F => X"0000006300000000000000630000000000000067000000000000009500000000",
            INIT_60 => X"0000005d0000000000000071000000000000006b000000000000005100000000",
            INIT_61 => X"00000066000000000000005d0000000000000073000000000000007500000000",
            INIT_62 => X"0000008300000000000000950000000000000098000000000000008900000000",
            INIT_63 => X"00000071000000000000007d0000000000000088000000000000008200000000",
            INIT_64 => X"0000007b0000000000000072000000000000006c000000000000006c00000000",
            INIT_65 => X"000000c200000000000000af000000000000007f000000000000007600000000",
            INIT_66 => X"000000a2000000000000007600000000000000bd00000000000000ce00000000",
            INIT_67 => X"000000650000000000000062000000000000005000000000000000a700000000",
            INIT_68 => X"0000005d000000000000006a000000000000006e000000000000006100000000",
            INIT_69 => X"0000006400000000000000590000000000000054000000000000006200000000",
            INIT_6A => X"00000086000000000000008a000000000000007b000000000000006e00000000",
            INIT_6B => X"0000007c00000000000000820000000000000083000000000000007e00000000",
            INIT_6C => X"00000087000000000000007e000000000000007f000000000000007b00000000",
            INIT_6D => X"000000b400000000000000b50000000000000099000000000000008600000000",
            INIT_6E => X"0000007a000000000000009700000000000000b700000000000000b800000000",
            INIT_6F => X"000000590000000000000048000000000000004d00000000000000a000000000",
            INIT_70 => X"0000006100000000000000660000000000000065000000000000006600000000",
            INIT_71 => X"0000006b00000000000000580000000000000058000000000000005f00000000",
            INIT_72 => X"0000009e0000000000000097000000000000008e000000000000008200000000",
            INIT_73 => X"0000009d00000000000000a100000000000000a400000000000000a300000000",
            INIT_74 => X"000000a900000000000000aa00000000000000ad00000000000000ab00000000",
            INIT_75 => X"000000ae00000000000000b100000000000000a900000000000000a200000000",
            INIT_76 => X"0000006200000000000000a400000000000000a800000000000000b000000000",
            INIT_77 => X"0000004b000000000000003f0000000000000046000000000000005700000000",
            INIT_78 => X"0000007c000000000000007f0000000000000076000000000000007b00000000",
            INIT_79 => X"000000a000000000000000980000000000000094000000000000007e00000000",
            INIT_7A => X"000000b400000000000000b300000000000000af00000000000000a700000000",
            INIT_7B => X"000000ae00000000000000b900000000000000b800000000000000b700000000",
            INIT_7C => X"000000a000000000000000af00000000000000b200000000000000ad00000000",
            INIT_7D => X"000000a1000000000000008e0000000000000085000000000000008000000000",
            INIT_7E => X"0000006c00000000000000a600000000000000a200000000000000a900000000",
            INIT_7F => X"000000520000000000000059000000000000005f000000000000004600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "sampleifmap_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000098000000000000008a000000000000007d000000000000008500000000",
            INIT_01 => X"000000a700000000000000a6000000000000009a000000000000009400000000",
            INIT_02 => X"000000b600000000000000b300000000000000ae00000000000000aa00000000",
            INIT_03 => X"000000ab00000000000000b500000000000000b900000000000000b900000000",
            INIT_04 => X"0000008b000000000000009a0000000000000098000000000000009800000000",
            INIT_05 => X"0000009b00000000000000900000000000000078000000000000006600000000",
            INIT_06 => X"0000008800000000000000a300000000000000a200000000000000a500000000",
            INIT_07 => X"0000006c000000000000009900000000000000bb000000000000009100000000",
            INIT_08 => X"00000083000000000000008d0000000000000085000000000000007c00000000",
            INIT_09 => X"000000aa00000000000000980000000000000072000000000000007400000000",
            INIT_0A => X"000000ad00000000000000b000000000000000af00000000000000af00000000",
            INIT_0B => X"00000097000000000000009a00000000000000a000000000000000a700000000",
            INIT_0C => X"000000a000000000000000a80000000000000096000000000000009000000000",
            INIT_0D => X"0000009e00000000000000a50000000000000098000000000000008c00000000",
            INIT_0E => X"00000097000000000000009c000000000000009b00000000000000a300000000",
            INIT_0F => X"000000930000000000000098000000000000009e000000000000009e00000000",
            INIT_10 => X"0000005d00000000000000600000000000000071000000000000008100000000",
            INIT_11 => X"000000a400000000000000940000000000000087000000000000006e00000000",
            INIT_12 => X"000000920000000000000096000000000000009f00000000000000a900000000",
            INIT_13 => X"000000a5000000000000009f0000000000000099000000000000009400000000",
            INIT_14 => X"000000ac00000000000000a800000000000000a000000000000000aa00000000",
            INIT_15 => X"000000a400000000000000a800000000000000a400000000000000a100000000",
            INIT_16 => X"00000092000000000000009e000000000000009e00000000000000a000000000",
            INIT_17 => X"00000096000000000000007d0000000000000079000000000000008400000000",
            INIT_18 => X"0000008700000000000000600000000000000055000000000000007000000000",
            INIT_19 => X"00000093000000000000009c00000000000000a5000000000000009b00000000",
            INIT_1A => X"000000a00000000000000097000000000000008d000000000000008e00000000",
            INIT_1B => X"000000ab00000000000000ae00000000000000ad00000000000000a700000000",
            INIT_1C => X"000000a800000000000000a2000000000000009b00000000000000a700000000",
            INIT_1D => X"000000a600000000000000a300000000000000a100000000000000a300000000",
            INIT_1E => X"0000006f00000000000000820000000000000097000000000000009e00000000",
            INIT_1F => X"0000008a000000000000005c0000000000000052000000000000006200000000",
            INIT_20 => X"0000008f00000000000000870000000000000084000000000000008500000000",
            INIT_21 => X"0000008e0000000000000096000000000000008f000000000000008f00000000",
            INIT_22 => X"000000ab00000000000000a900000000000000a1000000000000008a00000000",
            INIT_23 => X"00000086000000000000009700000000000000a500000000000000a900000000",
            INIT_24 => X"000000a40000000000000094000000000000006b000000000000007400000000",
            INIT_25 => X"00000098000000000000009f00000000000000a300000000000000a300000000",
            INIT_26 => X"0000005b0000000000000066000000000000006c000000000000008000000000",
            INIT_27 => X"000000480000000000000050000000000000004e000000000000004b00000000",
            INIT_28 => X"0000008f0000000000000090000000000000008c000000000000008400000000",
            INIT_29 => X"0000009600000000000000970000000000000093000000000000009000000000",
            INIT_2A => X"0000009a00000000000000940000000000000092000000000000008b00000000",
            INIT_2B => X"0000004e000000000000006e000000000000009c000000000000009f00000000",
            INIT_2C => X"000000a30000000000000084000000000000004a000000000000004b00000000",
            INIT_2D => X"0000006d000000000000007e000000000000008f000000000000009900000000",
            INIT_2E => X"0000004c000000000000005a0000000000000064000000000000006700000000",
            INIT_2F => X"0000002100000000000000390000000000000052000000000000004b00000000",
            INIT_30 => X"0000009200000000000000940000000000000089000000000000005e00000000",
            INIT_31 => X"0000007300000000000000810000000000000091000000000000009200000000",
            INIT_32 => X"0000008700000000000000630000000000000066000000000000006a00000000",
            INIT_33 => X"0000005d0000000000000072000000000000009a000000000000009d00000000",
            INIT_34 => X"0000007c000000000000007d0000000000000068000000000000006500000000",
            INIT_35 => X"000000650000000000000066000000000000006a000000000000007100000000",
            INIT_36 => X"0000003f0000000000000045000000000000004f000000000000005800000000",
            INIT_37 => X"0000001f00000000000000250000000000000035000000000000004300000000",
            INIT_38 => X"000000860000000000000086000000000000007d000000000000005600000000",
            INIT_39 => X"0000004d000000000000005c0000000000000085000000000000008900000000",
            INIT_3A => X"00000083000000000000005c0000000000000059000000000000005200000000",
            INIT_3B => X"0000007300000000000000840000000000000096000000000000009900000000",
            INIT_3C => X"0000006100000000000000600000000000000061000000000000006a00000000",
            INIT_3D => X"0000004f000000000000005f0000000000000065000000000000006300000000",
            INIT_3E => X"00000039000000000000003c0000000000000040000000000000003c00000000",
            INIT_3F => X"0000001f00000000000000220000000000000026000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008300000000000000810000000000000074000000000000005a00000000",
            INIT_41 => X"00000061000000000000006a000000000000008a000000000000008900000000",
            INIT_42 => X"0000007e000000000000007c0000000000000074000000000000006c00000000",
            INIT_43 => X"000000530000000000000054000000000000005f000000000000007100000000",
            INIT_44 => X"000000640000000000000062000000000000005c000000000000005900000000",
            INIT_45 => X"000000450000000000000043000000000000004a000000000000005c00000000",
            INIT_46 => X"0000002e00000000000000330000000000000042000000000000004a00000000",
            INIT_47 => X"0000002000000000000000230000000000000026000000000000002b00000000",
            INIT_48 => X"0000007f00000000000000820000000000000070000000000000005c00000000",
            INIT_49 => X"00000066000000000000006e0000000000000078000000000000007c00000000",
            INIT_4A => X"0000004c0000000000000050000000000000005a000000000000006100000000",
            INIT_4B => X"0000005b00000000000000540000000000000050000000000000004b00000000",
            INIT_4C => X"0000004900000000000000510000000000000059000000000000005f00000000",
            INIT_4D => X"0000003d00000000000000430000000000000041000000000000004100000000",
            INIT_4E => X"00000028000000000000002a000000000000003a000000000000004500000000",
            INIT_4F => X"0000002500000000000000230000000000000028000000000000002a00000000",
            INIT_50 => X"0000004e0000000000000056000000000000004f000000000000004c00000000",
            INIT_51 => X"0000003f00000000000000400000000000000045000000000000004a00000000",
            INIT_52 => X"0000004d000000000000004a0000000000000046000000000000004100000000",
            INIT_53 => X"0000005000000000000000510000000000000052000000000000005100000000",
            INIT_54 => X"000000440000000000000037000000000000003b000000000000004900000000",
            INIT_55 => X"000000320000000000000036000000000000003f000000000000004300000000",
            INIT_56 => X"000000280000000000000028000000000000002d000000000000003600000000",
            INIT_57 => X"0000002500000000000000270000000000000028000000000000002900000000",
            INIT_58 => X"0000002a0000000000000028000000000000002b000000000000002d00000000",
            INIT_59 => X"0000003a00000000000000350000000000000034000000000000003100000000",
            INIT_5A => X"0000004600000000000000480000000000000047000000000000004400000000",
            INIT_5B => X"0000003b000000000000003a000000000000003b000000000000004100000000",
            INIT_5C => X"000000490000000000000055000000000000003f000000000000003800000000",
            INIT_5D => X"0000002f000000000000002f0000000000000033000000000000003900000000",
            INIT_5E => X"0000002800000000000000270000000000000028000000000000002c00000000",
            INIT_5F => X"0000001d000000000000002a000000000000002a000000000000002900000000",
            INIT_60 => X"0000002600000000000000240000000000000028000000000000002b00000000",
            INIT_61 => X"0000003200000000000000310000000000000030000000000000002c00000000",
            INIT_62 => X"0000003100000000000000310000000000000034000000000000003500000000",
            INIT_63 => X"0000003d000000000000003e000000000000003b000000000000003500000000",
            INIT_64 => X"00000042000000000000005e0000000000000045000000000000003700000000",
            INIT_65 => X"00000028000000000000002f000000000000002e000000000000002c00000000",
            INIT_66 => X"0000002a00000000000000280000000000000027000000000000002700000000",
            INIT_67 => X"000000120000000000000020000000000000002e000000000000002900000000",
            INIT_68 => X"0000002400000000000000230000000000000027000000000000002800000000",
            INIT_69 => X"0000002b00000000000000290000000000000029000000000000002700000000",
            INIT_6A => X"0000003a00000000000000380000000000000033000000000000002e00000000",
            INIT_6B => X"00000037000000000000003c000000000000003d000000000000003d00000000",
            INIT_6C => X"000000360000000000000055000000000000003c000000000000002e00000000",
            INIT_6D => X"000000240000000000000025000000000000002e000000000000002800000000",
            INIT_6E => X"0000002a00000000000000280000000000000026000000000000002600000000",
            INIT_6F => X"00000007000000000000000d0000000000000028000000000000002b00000000",
            INIT_70 => X"0000002800000000000000240000000000000026000000000000002200000000",
            INIT_71 => X"000000330000000000000031000000000000002f000000000000002c00000000",
            INIT_72 => X"00000039000000000000003b0000000000000039000000000000003600000000",
            INIT_73 => X"0000002b00000000000000330000000000000037000000000000003900000000",
            INIT_74 => X"00000032000000000000004e0000000000000030000000000000001f00000000",
            INIT_75 => X"0000002300000000000000230000000000000025000000000000002900000000",
            INIT_76 => X"0000002900000000000000240000000000000025000000000000002500000000",
            INIT_77 => X"0000000700000000000000060000000000000014000000000000002d00000000",
            INIT_78 => X"0000002f000000000000002d000000000000002b000000000000002900000000",
            INIT_79 => X"0000003100000000000000300000000000000030000000000000003000000000",
            INIT_7A => X"0000002d00000000000000310000000000000033000000000000003200000000",
            INIT_7B => X"00000011000000000000001a0000000000000022000000000000002800000000",
            INIT_7C => X"0000002c000000000000003f000000000000001b000000000000000800000000",
            INIT_7D => X"0000002300000000000000220000000000000022000000000000002100000000",
            INIT_7E => X"0000002c00000000000000220000000000000022000000000000002300000000",
            INIT_7F => X"0000000800000000000000050000000000000006000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "sampleifmap_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ba00000000000000c200000000000000da00000000000000de00000000",
            INIT_01 => X"000000f100000000000000ee00000000000000ec00000000000000de00000000",
            INIT_02 => X"000000eb00000000000000f400000000000000f500000000000000f300000000",
            INIT_03 => X"000000f500000000000000f200000000000000f100000000000000f000000000",
            INIT_04 => X"000000f800000000000000f500000000000000f000000000000000e300000000",
            INIT_05 => X"000000f300000000000000f300000000000000f300000000000000f900000000",
            INIT_06 => X"000000f700000000000000ef00000000000000eb00000000000000f500000000",
            INIT_07 => X"000000f600000000000000f300000000000000ea00000000000000f100000000",
            INIT_08 => X"000000b800000000000000c900000000000000e200000000000000e500000000",
            INIT_09 => X"000000ee00000000000000f000000000000000f000000000000000df00000000",
            INIT_0A => X"000000e800000000000000f500000000000000f700000000000000f300000000",
            INIT_0B => X"000000f800000000000000f500000000000000f500000000000000f300000000",
            INIT_0C => X"000000fb00000000000000f300000000000000ef00000000000000e600000000",
            INIT_0D => X"000000f400000000000000ee00000000000000ee00000000000000fb00000000",
            INIT_0E => X"000000fc00000000000000f300000000000000ec00000000000000f800000000",
            INIT_0F => X"000000fb00000000000000fa00000000000000ec00000000000000f000000000",
            INIT_10 => X"000000b500000000000000c700000000000000de00000000000000e100000000",
            INIT_11 => X"000000e400000000000000ef00000000000000ee00000000000000db00000000",
            INIT_12 => X"000000e400000000000000ec00000000000000f400000000000000eb00000000",
            INIT_13 => X"000000f700000000000000ee00000000000000ef00000000000000eb00000000",
            INIT_14 => X"000000f600000000000000f100000000000000ec00000000000000e500000000",
            INIT_15 => X"000000ef00000000000000e800000000000000d700000000000000ec00000000",
            INIT_16 => X"000000fc00000000000000f200000000000000eb00000000000000f800000000",
            INIT_17 => X"000000f700000000000000fb00000000000000e800000000000000f100000000",
            INIT_18 => X"000000b300000000000000c200000000000000d800000000000000de00000000",
            INIT_19 => X"000000e100000000000000eb00000000000000e400000000000000d600000000",
            INIT_1A => X"000000dd00000000000000e600000000000000ef00000000000000e500000000",
            INIT_1B => X"000000f700000000000000e600000000000000ec00000000000000e100000000",
            INIT_1C => X"000000ee00000000000000f000000000000000ea00000000000000e600000000",
            INIT_1D => X"000000f100000000000000e500000000000000b000000000000000ba00000000",
            INIT_1E => X"000000fb00000000000000ef00000000000000e900000000000000f800000000",
            INIT_1F => X"000000f300000000000000f800000000000000e400000000000000ee00000000",
            INIT_20 => X"000000ac00000000000000c100000000000000d900000000000000df00000000",
            INIT_21 => X"000000d900000000000000e700000000000000dd00000000000000d200000000",
            INIT_22 => X"000000d700000000000000e100000000000000eb00000000000000da00000000",
            INIT_23 => X"000000ee00000000000000d600000000000000e800000000000000db00000000",
            INIT_24 => X"000000e400000000000000ee00000000000000e300000000000000e500000000",
            INIT_25 => X"000000ef00000000000000e500000000000000b200000000000000b000000000",
            INIT_26 => X"000000f500000000000000ea00000000000000e700000000000000f700000000",
            INIT_27 => X"000000f000000000000000f600000000000000e800000000000000e700000000",
            INIT_28 => X"000000a400000000000000bf00000000000000d500000000000000dc00000000",
            INIT_29 => X"000000d500000000000000e100000000000000d500000000000000ce00000000",
            INIT_2A => X"000000d600000000000000da00000000000000e600000000000000d600000000",
            INIT_2B => X"000000ce00000000000000c800000000000000e300000000000000d600000000",
            INIT_2C => X"000000cf00000000000000ed00000000000000ce00000000000000d000000000",
            INIT_2D => X"000000e900000000000000e600000000000000ad000000000000008200000000",
            INIT_2E => X"000000e800000000000000db00000000000000e100000000000000f400000000",
            INIT_2F => X"000000e600000000000000f200000000000000e700000000000000dd00000000",
            INIT_30 => X"0000009600000000000000b900000000000000ca00000000000000d400000000",
            INIT_31 => X"000000d000000000000000d900000000000000c900000000000000c400000000",
            INIT_32 => X"000000d300000000000000d000000000000000db00000000000000d300000000",
            INIT_33 => X"000000af00000000000000b900000000000000dd00000000000000d400000000",
            INIT_34 => X"000000c500000000000000d200000000000000bd00000000000000bb00000000",
            INIT_35 => X"000000bb00000000000000b8000000000000009d000000000000008900000000",
            INIT_36 => X"000000da00000000000000ce00000000000000dc00000000000000dd00000000",
            INIT_37 => X"000000d800000000000000e700000000000000db00000000000000d100000000",
            INIT_38 => X"0000009300000000000000b300000000000000c900000000000000d300000000",
            INIT_39 => X"000000cb00000000000000ce00000000000000cc00000000000000c500000000",
            INIT_3A => X"000000cd00000000000000c600000000000000d200000000000000d000000000",
            INIT_3B => X"000000cb00000000000000c000000000000000ce00000000000000ce00000000",
            INIT_3C => X"0000006a000000000000007a000000000000009b00000000000000b300000000",
            INIT_3D => X"000000490000000000000058000000000000005e000000000000006400000000",
            INIT_3E => X"000000d700000000000000ca00000000000000b7000000000000006f00000000",
            INIT_3F => X"000000c100000000000000ce00000000000000b900000000000000c600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c00000000000000a000000000000000ad00000000000000b300000000",
            INIT_41 => X"000000b300000000000000a100000000000000af00000000000000aa00000000",
            INIT_42 => X"000000bd00000000000000b400000000000000b800000000000000bb00000000",
            INIT_43 => X"000000c400000000000000ba00000000000000b900000000000000c300000000",
            INIT_44 => X"0000008000000000000000800000000000000089000000000000009f00000000",
            INIT_45 => X"0000005a0000000000000080000000000000007e000000000000007e00000000",
            INIT_46 => X"000000ac000000000000009e000000000000007c000000000000005800000000",
            INIT_47 => X"0000009f00000000000000b00000000000000089000000000000009c00000000",
            INIT_48 => X"00000070000000000000007b000000000000007e000000000000007b00000000",
            INIT_49 => X"0000008000000000000000720000000000000072000000000000007200000000",
            INIT_4A => X"0000009000000000000000890000000000000086000000000000008600000000",
            INIT_4B => X"000000a700000000000000a00000000000000092000000000000009800000000",
            INIT_4C => X"0000008c0000000000000090000000000000008b000000000000009300000000",
            INIT_4D => X"0000006800000000000000780000000000000083000000000000008200000000",
            INIT_4E => X"0000008d00000000000000960000000000000083000000000000009500000000",
            INIT_4F => X"0000007500000000000000800000000000000069000000000000006a00000000",
            INIT_50 => X"0000005800000000000000620000000000000066000000000000005900000000",
            INIT_51 => X"0000006a00000000000000680000000000000073000000000000006b00000000",
            INIT_52 => X"0000007300000000000000710000000000000076000000000000006b00000000",
            INIT_53 => X"0000009200000000000000970000000000000086000000000000007b00000000",
            INIT_54 => X"00000078000000000000007f000000000000007f000000000000008000000000",
            INIT_55 => X"00000080000000000000007a0000000000000068000000000000006f00000000",
            INIT_56 => X"000000b6000000000000008b000000000000006e000000000000008600000000",
            INIT_57 => X"00000070000000000000006d0000000000000075000000000000007200000000",
            INIT_58 => X"0000006a000000000000006e0000000000000068000000000000005800000000",
            INIT_59 => X"0000005e00000000000000710000000000000089000000000000008e00000000",
            INIT_5A => X"0000007d000000000000007f0000000000000092000000000000007400000000",
            INIT_5B => X"0000009700000000000000a500000000000000a5000000000000009400000000",
            INIT_5C => X"0000007f000000000000007f0000000000000082000000000000008e00000000",
            INIT_5D => X"000000bf00000000000000a50000000000000072000000000000007b00000000",
            INIT_5E => X"000000b80000000000000064000000000000008e00000000000000b400000000",
            INIT_5F => X"0000006c000000000000006c000000000000006d000000000000008c00000000",
            INIT_60 => X"0000006800000000000000840000000000000082000000000000006400000000",
            INIT_61 => X"00000076000000000000006d0000000000000082000000000000008100000000",
            INIT_62 => X"0000009700000000000000a800000000000000ab000000000000009a00000000",
            INIT_63 => X"0000008b000000000000009a00000000000000a5000000000000009b00000000",
            INIT_64 => X"0000008c0000000000000081000000000000007d000000000000008200000000",
            INIT_65 => X"000000c100000000000000b30000000000000089000000000000008600000000",
            INIT_66 => X"00000098000000000000007000000000000000b900000000000000cb00000000",
            INIT_67 => X"0000006d0000000000000069000000000000005400000000000000a000000000",
            INIT_68 => X"0000006a000000000000007e0000000000000086000000000000007800000000",
            INIT_69 => X"00000079000000000000006c0000000000000065000000000000007100000000",
            INIT_6A => X"0000009f00000000000000a10000000000000091000000000000008300000000",
            INIT_6B => X"00000095000000000000009e00000000000000a1000000000000009900000000",
            INIT_6C => X"0000009b00000000000000910000000000000093000000000000009200000000",
            INIT_6D => X"000000b100000000000000b600000000000000a1000000000000009600000000",
            INIT_6E => X"00000076000000000000009400000000000000b500000000000000b500000000",
            INIT_6F => X"00000060000000000000004e0000000000000050000000000000009d00000000",
            INIT_70 => X"00000072000000000000007d0000000000000080000000000000007f00000000",
            INIT_71 => X"0000008600000000000000730000000000000071000000000000007400000000",
            INIT_72 => X"000000b800000000000000b000000000000000a8000000000000009f00000000",
            INIT_73 => X"000000b900000000000000be00000000000000bf00000000000000be00000000",
            INIT_74 => X"000000b800000000000000be00000000000000c400000000000000c500000000",
            INIT_75 => X"000000a800000000000000af00000000000000ad00000000000000ac00000000",
            INIT_76 => X"0000006300000000000000a300000000000000a500000000000000ab00000000",
            INIT_77 => X"0000005100000000000000430000000000000047000000000000005700000000",
            INIT_78 => X"00000091000000000000009a0000000000000095000000000000009700000000",
            INIT_79 => X"000000c100000000000000b800000000000000b3000000000000009900000000",
            INIT_7A => X"000000d000000000000000cf00000000000000cd00000000000000c900000000",
            INIT_7B => X"000000c800000000000000d400000000000000d200000000000000d100000000",
            INIT_7C => X"000000ab00000000000000c300000000000000c900000000000000c600000000",
            INIT_7D => X"0000009b000000000000008b0000000000000087000000000000008600000000",
            INIT_7E => X"0000007100000000000000a800000000000000a100000000000000a500000000",
            INIT_7F => X"00000056000000000000005a000000000000005c000000000000004900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "sampleifmap_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b000000000000000a7000000000000009f00000000000000a500000000",
            INIT_01 => X"000000c900000000000000c600000000000000b900000000000000af00000000",
            INIT_02 => X"000000d200000000000000d200000000000000d000000000000000cd00000000",
            INIT_03 => X"000000be00000000000000c900000000000000d000000000000000d200000000",
            INIT_04 => X"0000009400000000000000a900000000000000aa00000000000000aa00000000",
            INIT_05 => X"00000099000000000000008e000000000000007a000000000000006c00000000",
            INIT_06 => X"0000008e00000000000000a700000000000000a500000000000000a700000000",
            INIT_07 => X"0000006f000000000000009800000000000000b5000000000000009300000000",
            INIT_08 => X"0000009d00000000000000ae00000000000000aa000000000000009d00000000",
            INIT_09 => X"000000ca00000000000000b6000000000000008f000000000000008d00000000",
            INIT_0A => X"000000ca00000000000000d100000000000000d300000000000000d000000000",
            INIT_0B => X"000000a200000000000000a700000000000000b500000000000000bf00000000",
            INIT_0C => X"000000a900000000000000b200000000000000a0000000000000009b00000000",
            INIT_0D => X"000000a000000000000000a7000000000000009d000000000000009300000000",
            INIT_0E => X"0000009c00000000000000a100000000000000a200000000000000a900000000",
            INIT_0F => X"0000009400000000000000960000000000000096000000000000009e00000000",
            INIT_10 => X"000000790000000000000080000000000000009400000000000000a200000000",
            INIT_11 => X"000000c200000000000000b100000000000000a4000000000000008a00000000",
            INIT_12 => X"000000ab00000000000000b200000000000000bc00000000000000c700000000",
            INIT_13 => X"000000b000000000000000ac00000000000000ac00000000000000aa00000000",
            INIT_14 => X"000000b500000000000000b000000000000000a800000000000000b400000000",
            INIT_15 => X"000000ac00000000000000af00000000000000ad00000000000000aa00000000",
            INIT_16 => X"0000009600000000000000a300000000000000a500000000000000a800000000",
            INIT_17 => X"00000099000000000000007d0000000000000076000000000000008500000000",
            INIT_18 => X"000000a6000000000000007f0000000000000075000000000000008f00000000",
            INIT_19 => X"000000b000000000000000ba00000000000000c500000000000000bc00000000",
            INIT_1A => X"000000b200000000000000ab00000000000000a300000000000000a900000000",
            INIT_1B => X"000000ba00000000000000bf00000000000000be00000000000000b900000000",
            INIT_1C => X"000000b100000000000000ac00000000000000a500000000000000b400000000",
            INIT_1D => X"000000b200000000000000af00000000000000ac00000000000000ad00000000",
            INIT_1E => X"000000740000000000000088000000000000009c00000000000000a400000000",
            INIT_1F => X"0000009000000000000000620000000000000057000000000000006700000000",
            INIT_20 => X"000000b000000000000000a800000000000000a500000000000000a600000000",
            INIT_21 => X"000000aa00000000000000b300000000000000ae00000000000000b000000000",
            INIT_22 => X"000000bd00000000000000be00000000000000b800000000000000a400000000",
            INIT_23 => X"0000009600000000000000a800000000000000b500000000000000b900000000",
            INIT_24 => X"000000ad000000000000009d0000000000000076000000000000008100000000",
            INIT_25 => X"000000a200000000000000ab00000000000000ad00000000000000ad00000000",
            INIT_26 => X"0000005f000000000000006a0000000000000070000000000000008500000000",
            INIT_27 => X"0000004e00000000000000560000000000000054000000000000005000000000",
            INIT_28 => X"000000af00000000000000b100000000000000ac00000000000000a500000000",
            INIT_29 => X"000000b000000000000000b300000000000000b000000000000000ae00000000",
            INIT_2A => X"000000ad00000000000000ab00000000000000ab00000000000000a400000000",
            INIT_2B => X"0000005e000000000000007e00000000000000ab00000000000000af00000000",
            INIT_2C => X"000000ac000000000000008e0000000000000055000000000000005800000000",
            INIT_2D => X"000000750000000000000088000000000000009800000000000000a200000000",
            INIT_2E => X"00000050000000000000005e0000000000000068000000000000006c00000000",
            INIT_2F => X"00000027000000000000003f0000000000000058000000000000004f00000000",
            INIT_30 => X"000000af00000000000000b200000000000000a6000000000000007c00000000",
            INIT_31 => X"0000008b000000000000009a00000000000000ad00000000000000af00000000",
            INIT_32 => X"0000009a000000000000007a000000000000007e000000000000008200000000",
            INIT_33 => X"0000006c000000000000008300000000000000a900000000000000ae00000000",
            INIT_34 => X"0000008500000000000000860000000000000072000000000000007200000000",
            INIT_35 => X"0000006c000000000000006d0000000000000071000000000000007900000000",
            INIT_36 => X"00000045000000000000004b0000000000000056000000000000005f00000000",
            INIT_37 => X"00000026000000000000002b000000000000003b000000000000004900000000",
            INIT_38 => X"0000009f00000000000000a00000000000000096000000000000006f00000000",
            INIT_39 => X"000000640000000000000074000000000000009e00000000000000a300000000",
            INIT_3A => X"0000009700000000000000730000000000000070000000000000006800000000",
            INIT_3B => X"00000083000000000000009500000000000000a800000000000000ac00000000",
            INIT_3C => X"0000006a000000000000006a000000000000006b000000000000007700000000",
            INIT_3D => X"000000540000000000000064000000000000006c000000000000006a00000000",
            INIT_3E => X"0000004100000000000000440000000000000049000000000000004500000000",
            INIT_3F => X"000000250000000000000028000000000000002c000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009a0000000000000097000000000000008a000000000000007100000000",
            INIT_41 => X"00000077000000000000008000000000000000a200000000000000a100000000",
            INIT_42 => X"0000009200000000000000900000000000000088000000000000008100000000",
            INIT_43 => X"0000006200000000000000650000000000000072000000000000008400000000",
            INIT_44 => X"0000006c000000000000006d0000000000000067000000000000006500000000",
            INIT_45 => X"0000004b00000000000000480000000000000050000000000000006300000000",
            INIT_46 => X"0000003a000000000000003d000000000000004d000000000000005500000000",
            INIT_47 => X"000000270000000000000029000000000000002d000000000000003400000000",
            INIT_48 => X"00000097000000000000009a0000000000000088000000000000007400000000",
            INIT_49 => X"0000007c0000000000000084000000000000008f000000000000009400000000",
            INIT_4A => X"00000057000000000000005b0000000000000067000000000000007600000000",
            INIT_4B => X"000000650000000000000063000000000000005b000000000000005600000000",
            INIT_4C => X"00000052000000000000005e0000000000000063000000000000006500000000",
            INIT_4D => X"00000045000000000000004a0000000000000048000000000000004800000000",
            INIT_4E => X"0000003200000000000000340000000000000044000000000000004e00000000",
            INIT_4F => X"00000030000000000000002f0000000000000030000000000000003300000000",
            INIT_50 => X"00000063000000000000006a0000000000000064000000000000006000000000",
            INIT_51 => X"0000005100000000000000520000000000000056000000000000005c00000000",
            INIT_52 => X"000000540000000000000051000000000000004f000000000000005200000000",
            INIT_53 => X"00000058000000000000005e000000000000005b000000000000005700000000",
            INIT_54 => X"0000004c00000000000000440000000000000044000000000000004d00000000",
            INIT_55 => X"0000003b00000000000000400000000000000048000000000000004a00000000",
            INIT_56 => X"0000003200000000000000310000000000000036000000000000003f00000000",
            INIT_57 => X"0000003000000000000000340000000000000030000000000000003100000000",
            INIT_58 => X"0000003700000000000000360000000000000039000000000000003b00000000",
            INIT_59 => X"00000044000000000000003e000000000000003d000000000000003c00000000",
            INIT_5A => X"0000004d000000000000004f000000000000004f000000000000004e00000000",
            INIT_5B => X"0000004200000000000000450000000000000044000000000000004800000000",
            INIT_5C => X"0000005200000000000000610000000000000047000000000000003d00000000",
            INIT_5D => X"000000390000000000000038000000000000003c000000000000004100000000",
            INIT_5E => X"0000003100000000000000300000000000000031000000000000003500000000",
            INIT_5F => X"0000002300000000000000320000000000000032000000000000003200000000",
            INIT_60 => X"0000002d000000000000002c0000000000000030000000000000003200000000",
            INIT_61 => X"0000003700000000000000350000000000000035000000000000003100000000",
            INIT_62 => X"000000380000000000000038000000000000003b000000000000003a00000000",
            INIT_63 => X"0000004400000000000000470000000000000042000000000000003c00000000",
            INIT_64 => X"0000004b0000000000000068000000000000004b000000000000003b00000000",
            INIT_65 => X"00000033000000000000003a0000000000000038000000000000003500000000",
            INIT_66 => X"0000003300000000000000310000000000000030000000000000003100000000",
            INIT_67 => X"0000001400000000000000250000000000000035000000000000003200000000",
            INIT_68 => X"000000290000000000000028000000000000002c000000000000002d00000000",
            INIT_69 => X"00000030000000000000002e000000000000002e000000000000002c00000000",
            INIT_6A => X"00000041000000000000003f0000000000000039000000000000003300000000",
            INIT_6B => X"0000003d00000000000000440000000000000044000000000000004400000000",
            INIT_6C => X"0000003f000000000000005d0000000000000042000000000000003200000000",
            INIT_6D => X"0000002f00000000000000300000000000000038000000000000003100000000",
            INIT_6E => X"000000330000000000000031000000000000002f000000000000002f00000000",
            INIT_6F => X"00000005000000000000000e000000000000002e000000000000003400000000",
            INIT_70 => X"0000002d0000000000000029000000000000002b000000000000002700000000",
            INIT_71 => X"0000003b00000000000000380000000000000036000000000000003200000000",
            INIT_72 => X"0000004000000000000000420000000000000040000000000000003e00000000",
            INIT_73 => X"00000031000000000000003a000000000000003d000000000000004000000000",
            INIT_74 => X"0000003b00000000000000550000000000000035000000000000002400000000",
            INIT_75 => X"0000002f000000000000002f0000000000000030000000000000003200000000",
            INIT_76 => X"00000032000000000000002d000000000000002e000000000000002e00000000",
            INIT_77 => X"0000000300000000000000030000000000000018000000000000003600000000",
            INIT_78 => X"0000003600000000000000340000000000000032000000000000002f00000000",
            INIT_79 => X"0000003a00000000000000380000000000000038000000000000003800000000",
            INIT_7A => X"0000003200000000000000350000000000000037000000000000003a00000000",
            INIT_7B => X"00000014000000000000001e0000000000000027000000000000002d00000000",
            INIT_7C => X"0000003600000000000000480000000000000021000000000000000b00000000",
            INIT_7D => X"0000002e000000000000002d000000000000002d000000000000002c00000000",
            INIT_7E => X"00000034000000000000002b000000000000002c000000000000002c00000000",
            INIT_7F => X"0000000700000000000000030000000000000008000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "sampleifmap_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000be00000000000000b000000000000000a7000000000000009b00000000",
            INIT_01 => X"000000a600000000000000a800000000000000a600000000000000b100000000",
            INIT_02 => X"000000bb00000000000000bb00000000000000b300000000000000aa00000000",
            INIT_03 => X"000000b800000000000000b800000000000000bb00000000000000bb00000000",
            INIT_04 => X"000000ba00000000000000b800000000000000b400000000000000b600000000",
            INIT_05 => X"000000bd00000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000c000000000000000ca00000000000000c900000000000000c900000000",
            INIT_08 => X"000000bb00000000000000ab00000000000000a3000000000000009900000000",
            INIT_09 => X"0000009f000000000000009a000000000000009b00000000000000b300000000",
            INIT_0A => X"000000af00000000000000ab00000000000000a5000000000000009f00000000",
            INIT_0B => X"000000a500000000000000a200000000000000ab00000000000000a900000000",
            INIT_0C => X"000000a500000000000000a600000000000000a400000000000000aa00000000",
            INIT_0D => X"000000a800000000000000a900000000000000ad00000000000000a700000000",
            INIT_0E => X"000000ca00000000000000be00000000000000ad00000000000000a900000000",
            INIT_0F => X"000000bd00000000000000cb00000000000000ca00000000000000cc00000000",
            INIT_10 => X"000000b800000000000000a800000000000000a0000000000000009b00000000",
            INIT_11 => X"000000bc00000000000000b000000000000000ae00000000000000bb00000000",
            INIT_12 => X"000000be00000000000000b100000000000000b300000000000000b600000000",
            INIT_13 => X"000000b900000000000000bc00000000000000c200000000000000c000000000",
            INIT_14 => X"000000c200000000000000c100000000000000c200000000000000c100000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c500000000000000c300000000",
            INIT_16 => X"000000cf00000000000000ce00000000000000c500000000000000bf00000000",
            INIT_17 => X"000000bd00000000000000cc00000000000000ce00000000000000d000000000",
            INIT_18 => X"000000b100000000000000a6000000000000009d000000000000009700000000",
            INIT_19 => X"000000c500000000000000c700000000000000b900000000000000b400000000",
            INIT_1A => X"000000c600000000000000cd00000000000000cc00000000000000b600000000",
            INIT_1B => X"000000cb00000000000000c400000000000000c500000000000000d200000000",
            INIT_1C => X"000000cb00000000000000d200000000000000cf00000000000000cd00000000",
            INIT_1D => X"000000cc00000000000000c500000000000000d200000000000000cf00000000",
            INIT_1E => X"000000c900000000000000cc00000000000000c600000000000000d000000000",
            INIT_1F => X"000000c000000000000000ce00000000000000cf00000000000000d100000000",
            INIT_20 => X"000000ae00000000000000a8000000000000009e000000000000009700000000",
            INIT_21 => X"000000c400000000000000bf00000000000000b500000000000000b100000000",
            INIT_22 => X"000000b900000000000000bd00000000000000c200000000000000b700000000",
            INIT_23 => X"000000ca00000000000000b900000000000000b900000000000000c400000000",
            INIT_24 => X"000000c000000000000000c800000000000000c700000000000000c700000000",
            INIT_25 => X"000000bc00000000000000be00000000000000c700000000000000c300000000",
            INIT_26 => X"000000c400000000000000c900000000000000c700000000000000c900000000",
            INIT_27 => X"000000c400000000000000cf00000000000000cc00000000000000ce00000000",
            INIT_28 => X"000000ae00000000000000a7000000000000009c000000000000009400000000",
            INIT_29 => X"000000c300000000000000c400000000000000ae00000000000000ab00000000",
            INIT_2A => X"000000b800000000000000bd00000000000000be00000000000000c000000000",
            INIT_2B => X"000000bf00000000000000bd00000000000000bd00000000000000bb00000000",
            INIT_2C => X"000000c600000000000000bb00000000000000c300000000000000be00000000",
            INIT_2D => X"000000c100000000000000c000000000000000bc00000000000000c000000000",
            INIT_2E => X"000000d100000000000000cb00000000000000ce00000000000000cd00000000",
            INIT_2F => X"000000c400000000000000d100000000000000d000000000000000d400000000",
            INIT_30 => X"000000ae00000000000000a50000000000000099000000000000009400000000",
            INIT_31 => X"000000c300000000000000cb00000000000000b000000000000000a800000000",
            INIT_32 => X"000000be00000000000000bb00000000000000bc00000000000000bc00000000",
            INIT_33 => X"000000c300000000000000c500000000000000c200000000000000b600000000",
            INIT_34 => X"000000cd00000000000000c800000000000000c100000000000000c400000000",
            INIT_35 => X"000000c900000000000000c500000000000000c500000000000000c600000000",
            INIT_36 => X"000000c300000000000000c600000000000000c800000000000000c500000000",
            INIT_37 => X"000000c300000000000000cf00000000000000cb00000000000000c500000000",
            INIT_38 => X"000000ac00000000000000a3000000000000009b000000000000009900000000",
            INIT_39 => X"000000d100000000000000c700000000000000bc00000000000000ac00000000",
            INIT_3A => X"000000bf00000000000000bd00000000000000be00000000000000c400000000",
            INIT_3B => X"000000c400000000000000bb00000000000000bc00000000000000c100000000",
            INIT_3C => X"000000ce00000000000000c400000000000000c200000000000000ca00000000",
            INIT_3D => X"000000c800000000000000c400000000000000c900000000000000c200000000",
            INIT_3E => X"000000c900000000000000c800000000000000bb00000000000000b500000000",
            INIT_3F => X"000000bd00000000000000c700000000000000c400000000000000c800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ac00000000000000a3000000000000009f00000000000000a000000000",
            INIT_41 => X"000000be00000000000000b000000000000000b000000000000000ae00000000",
            INIT_42 => X"000000b000000000000000b000000000000000af00000000000000b400000000",
            INIT_43 => X"000000b600000000000000ac00000000000000aa00000000000000b500000000",
            INIT_44 => X"000000bb00000000000000b500000000000000b200000000000000bb00000000",
            INIT_45 => X"000000bb00000000000000b400000000000000bc00000000000000b100000000",
            INIT_46 => X"000000bc00000000000000bc00000000000000c400000000000000c700000000",
            INIT_47 => X"000000b800000000000000c200000000000000c000000000000000c500000000",
            INIT_48 => X"000000ac00000000000000a200000000000000a700000000000000ab00000000",
            INIT_49 => X"000000b000000000000000b400000000000000ab00000000000000aa00000000",
            INIT_4A => X"0000009c0000000000000096000000000000009c000000000000009b00000000",
            INIT_4B => X"0000009e00000000000000990000000000000092000000000000009600000000",
            INIT_4C => X"0000009d00000000000000a400000000000000a600000000000000a600000000",
            INIT_4D => X"000000a6000000000000009c00000000000000a2000000000000009d00000000",
            INIT_4E => X"000000bd00000000000000bc00000000000000c700000000000000c800000000",
            INIT_4F => X"000000b600000000000000c200000000000000c100000000000000c500000000",
            INIT_50 => X"000000b000000000000000a800000000000000b400000000000000af00000000",
            INIT_51 => X"000000ae00000000000000b600000000000000b100000000000000ad00000000",
            INIT_52 => X"0000009a000000000000009f00000000000000a0000000000000009c00000000",
            INIT_53 => X"000000ad00000000000000a800000000000000a3000000000000009f00000000",
            INIT_54 => X"000000a200000000000000a000000000000000a400000000000000aa00000000",
            INIT_55 => X"000000ac00000000000000a700000000000000a800000000000000a000000000",
            INIT_56 => X"000000c400000000000000c400000000000000c300000000000000c200000000",
            INIT_57 => X"000000b700000000000000c100000000000000bf00000000000000c500000000",
            INIT_58 => X"000000bb00000000000000b200000000000000bb00000000000000b500000000",
            INIT_59 => X"000000b600000000000000ae00000000000000aa00000000000000b700000000",
            INIT_5A => X"000000b500000000000000b400000000000000b300000000000000b300000000",
            INIT_5B => X"000000c100000000000000c100000000000000bb00000000000000b800000000",
            INIT_5C => X"000000b900000000000000bc00000000000000c000000000000000c100000000",
            INIT_5D => X"000000c000000000000000c000000000000000ba00000000000000b800000000",
            INIT_5E => X"000000bd00000000000000c000000000000000bc00000000000000bb00000000",
            INIT_5F => X"000000ba00000000000000c400000000000000bf00000000000000be00000000",
            INIT_60 => X"000000ab00000000000000ba00000000000000be00000000000000b900000000",
            INIT_61 => X"000000c100000000000000950000000000000084000000000000009900000000",
            INIT_62 => X"000000bc00000000000000ba00000000000000bf00000000000000c600000000",
            INIT_63 => X"000000c400000000000000c300000000000000c100000000000000bf00000000",
            INIT_64 => X"000000bc00000000000000be00000000000000c000000000000000c300000000",
            INIT_65 => X"000000bf00000000000000c000000000000000be00000000000000bc00000000",
            INIT_66 => X"000000c500000000000000c300000000000000c100000000000000bf00000000",
            INIT_67 => X"000000c100000000000000cc00000000000000ca00000000000000ca00000000",
            INIT_68 => X"0000009e00000000000000bc00000000000000c200000000000000ba00000000",
            INIT_69 => X"0000006d000000000000005e0000000000000074000000000000008400000000",
            INIT_6A => X"000000c200000000000000c200000000000000b1000000000000009100000000",
            INIT_6B => X"000000c700000000000000c400000000000000c100000000000000bf00000000",
            INIT_6C => X"000000c600000000000000c800000000000000c700000000000000c700000000",
            INIT_6D => X"000000c600000000000000c700000000000000c400000000000000c400000000",
            INIT_6E => X"000000c400000000000000c400000000000000c400000000000000c500000000",
            INIT_6F => X"000000b900000000000000c600000000000000c500000000000000c600000000",
            INIT_70 => X"000000c600000000000000c400000000000000c500000000000000ba00000000",
            INIT_71 => X"0000005c000000000000008d00000000000000b800000000000000c200000000",
            INIT_72 => X"000000b3000000000000008e0000000000000068000000000000005400000000",
            INIT_73 => X"000000cc00000000000000cc00000000000000c900000000000000c300000000",
            INIT_74 => X"000000c700000000000000cc00000000000000cc00000000000000cc00000000",
            INIT_75 => X"000000bf00000000000000c200000000000000c200000000000000c200000000",
            INIT_76 => X"000000be00000000000000be00000000000000be00000000000000bd00000000",
            INIT_77 => X"000000b500000000000000c000000000000000be00000000000000bf00000000",
            INIT_78 => X"000000c800000000000000c600000000000000c700000000000000b800000000",
            INIT_79 => X"000000b100000000000000c900000000000000c800000000000000c500000000",
            INIT_7A => X"00000080000000000000005d0000000000000054000000000000007500000000",
            INIT_7B => X"000000cd00000000000000d000000000000000ca00000000000000ad00000000",
            INIT_7C => X"000000c700000000000000c700000000000000c800000000000000ca00000000",
            INIT_7D => X"000000c300000000000000c500000000000000c400000000000000c300000000",
            INIT_7E => X"000000bf00000000000000c200000000000000c300000000000000c100000000",
            INIT_7F => X"000000b200000000000000be00000000000000bd00000000000000bf00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "sampleifmap_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d000000000000000cb00000000000000c900000000000000b900000000",
            INIT_01 => X"000000d600000000000000d000000000000000ce00000000000000cd00000000",
            INIT_02 => X"0000005b000000000000004c000000000000005c00000000000000af00000000",
            INIT_03 => X"000000cb00000000000000b5000000000000008c000000000000006900000000",
            INIT_04 => X"000000c200000000000000c500000000000000ca00000000000000ce00000000",
            INIT_05 => X"000000c200000000000000c200000000000000c200000000000000c100000000",
            INIT_06 => X"000000bf00000000000000c100000000000000c300000000000000c200000000",
            INIT_07 => X"000000b400000000000000be00000000000000be00000000000000c100000000",
            INIT_08 => X"000000d600000000000000cf00000000000000cc00000000000000bb00000000",
            INIT_09 => X"000000d000000000000000d300000000000000d400000000000000d400000000",
            INIT_0A => X"000000570000000000000047000000000000007c00000000000000cb00000000",
            INIT_0B => X"0000008400000000000000630000000000000054000000000000005400000000",
            INIT_0C => X"000000cb00000000000000cb00000000000000be00000000000000a700000000",
            INIT_0D => X"000000c400000000000000c500000000000000c000000000000000c300000000",
            INIT_0E => X"000000bf00000000000000c000000000000000c200000000000000c200000000",
            INIT_0F => X"000000b700000000000000c000000000000000bf00000000000000c100000000",
            INIT_10 => X"000000d600000000000000cf00000000000000cf00000000000000be00000000",
            INIT_11 => X"000000d000000000000000d300000000000000d300000000000000d400000000",
            INIT_12 => X"000000570000000000000048000000000000008900000000000000d300000000",
            INIT_13 => X"0000005300000000000000560000000000000054000000000000005300000000",
            INIT_14 => X"0000009b0000000000000083000000000000006b000000000000005900000000",
            INIT_15 => X"000000cc00000000000000cb00000000000000b600000000000000a300000000",
            INIT_16 => X"000000bf00000000000000c200000000000000c600000000000000ca00000000",
            INIT_17 => X"000000b600000000000000bf00000000000000c000000000000000c100000000",
            INIT_18 => X"000000d700000000000000d100000000000000d200000000000000bf00000000",
            INIT_19 => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1A => X"0000003a000000000000002f000000000000007100000000000000cc00000000",
            INIT_1B => X"0000005d0000000000000057000000000000004c000000000000003f00000000",
            INIT_1C => X"0000003e00000000000000460000000000000050000000000000005a00000000",
            INIT_1D => X"0000009f000000000000007a000000000000004d000000000000003a00000000",
            INIT_1E => X"000000c800000000000000c900000000000000c200000000000000b400000000",
            INIT_1F => X"000000b900000000000000c400000000000000c400000000000000c800000000",
            INIT_20 => X"000000d300000000000000cf00000000000000d000000000000000bf00000000",
            INIT_21 => X"000000d400000000000000d100000000000000d200000000000000d100000000",
            INIT_22 => X"0000002500000000000000410000000000000065000000000000009d00000000",
            INIT_23 => X"00000058000000000000004a0000000000000044000000000000003300000000",
            INIT_24 => X"0000004900000000000000550000000000000056000000000000005b00000000",
            INIT_25 => X"00000048000000000000003e000000000000002e000000000000003700000000",
            INIT_26 => X"0000009e0000000000000085000000000000006b000000000000004e00000000",
            INIT_27 => X"000000ba00000000000000c400000000000000c300000000000000b800000000",
            INIT_28 => X"000000d100000000000000cb00000000000000ca00000000000000ba00000000",
            INIT_29 => X"000000c800000000000000d100000000000000ce00000000000000cf00000000",
            INIT_2A => X"000000640000000000000097000000000000008c000000000000009500000000",
            INIT_2B => X"0000006000000000000000320000000000000035000000000000002d00000000",
            INIT_2C => X"00000048000000000000008000000000000000a0000000000000009c00000000",
            INIT_2D => X"0000004200000000000000590000000000000070000000000000006200000000",
            INIT_2E => X"000000a300000000000000a60000000000000083000000000000004300000000",
            INIT_2F => X"000000b200000000000000bc00000000000000b700000000000000ad00000000",
            INIT_30 => X"000000d200000000000000ca00000000000000c900000000000000b900000000",
            INIT_31 => X"000000d100000000000000d100000000000000d000000000000000d200000000",
            INIT_32 => X"000000bd00000000000000d700000000000000d300000000000000d200000000",
            INIT_33 => X"000000a800000000000000940000000000000092000000000000009000000000",
            INIT_34 => X"0000009a00000000000000c000000000000000ce00000000000000ca00000000",
            INIT_35 => X"0000009f00000000000000b100000000000000b200000000000000a300000000",
            INIT_36 => X"000000c200000000000000bf00000000000000b2000000000000009c00000000",
            INIT_37 => X"000000b000000000000000bc00000000000000c100000000000000c400000000",
            INIT_38 => X"000000c400000000000000c000000000000000bc00000000000000b000000000",
            INIT_39 => X"000000b700000000000000b900000000000000bc00000000000000c000000000",
            INIT_3A => X"000000ad00000000000000b300000000000000b200000000000000b600000000",
            INIT_3B => X"000000ad00000000000000ab00000000000000aa00000000000000aa00000000",
            INIT_3C => X"000000a700000000000000a100000000000000a000000000000000a900000000",
            INIT_3D => X"000000aa00000000000000a500000000000000a100000000000000a500000000",
            INIT_3E => X"00000096000000000000009800000000000000a000000000000000aa00000000",
            INIT_3F => X"0000009c00000000000000a400000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006b000000000000006e0000000000000063000000000000007200000000",
            INIT_41 => X"0000005d000000000000005e0000000000000061000000000000006600000000",
            INIT_42 => X"0000005000000000000000580000000000000055000000000000005800000000",
            INIT_43 => X"000000650000000000000053000000000000004e000000000000004d00000000",
            INIT_44 => X"0000006b000000000000006a000000000000006c000000000000007100000000",
            INIT_45 => X"00000071000000000000006f000000000000006e000000000000006c00000000",
            INIT_46 => X"0000007700000000000000780000000000000077000000000000007500000000",
            INIT_47 => X"0000007c000000000000007a0000000000000079000000000000007800000000",
            INIT_48 => X"000000750000000000000071000000000000006d000000000000007a00000000",
            INIT_49 => X"0000007100000000000000720000000000000070000000000000007300000000",
            INIT_4A => X"0000006d000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006c000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006b00000000000000690000000000000070000000000000007300000000",
            INIT_4D => X"000000680000000000000065000000000000006a000000000000006c00000000",
            INIT_4E => X"0000006d000000000000006d000000000000006b000000000000006a00000000",
            INIT_4F => X"00000065000000000000005e0000000000000066000000000000006700000000",
            INIT_50 => X"00000070000000000000006b0000000000000061000000000000007800000000",
            INIT_51 => X"0000005e00000000000000620000000000000068000000000000006d00000000",
            INIT_52 => X"000000560000000000000058000000000000005d000000000000005e00000000",
            INIT_53 => X"0000004e0000000000000050000000000000004f000000000000005200000000",
            INIT_54 => X"000000450000000000000048000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000042000000000000004300000000",
            INIT_56 => X"0000004000000000000000420000000000000041000000000000004000000000",
            INIT_57 => X"0000004d0000000000000035000000000000003f000000000000004300000000",
            INIT_58 => X"0000004500000000000000410000000000000037000000000000005b00000000",
            INIT_59 => X"0000003d000000000000003f0000000000000042000000000000004200000000",
            INIT_5A => X"00000039000000000000003c0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003a00000000000000400000000000000042000000000000003f00000000",
            INIT_5D => X"0000003c000000000000003b0000000000000039000000000000003800000000",
            INIT_5E => X"0000003900000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000005c000000000000004b0000000000000031000000000000003400000000",
            INIT_60 => X"000000440000000000000042000000000000003c000000000000005d00000000",
            INIT_61 => X"0000004100000000000000400000000000000043000000000000004300000000",
            INIT_62 => X"0000003b000000000000003e0000000000000041000000000000004500000000",
            INIT_63 => X"0000003d000000000000003c000000000000003b000000000000003b00000000",
            INIT_64 => X"00000038000000000000003a000000000000003f000000000000004000000000",
            INIT_65 => X"0000003800000000000000380000000000000037000000000000003700000000",
            INIT_66 => X"000000350000000000000038000000000000003a000000000000003900000000",
            INIT_67 => X"000000510000000000000061000000000000005d000000000000004100000000",
            INIT_68 => X"00000039000000000000003d0000000000000039000000000000005900000000",
            INIT_69 => X"0000003b0000000000000039000000000000003b000000000000003900000000",
            INIT_6A => X"000000360000000000000038000000000000003a000000000000003c00000000",
            INIT_6B => X"0000003d000000000000003b000000000000003d000000000000003c00000000",
            INIT_6C => X"00000039000000000000003a000000000000003d000000000000004100000000",
            INIT_6D => X"0000003d000000000000003d000000000000003c000000000000003c00000000",
            INIT_6E => X"000000460000000000000039000000000000003e000000000000004200000000",
            INIT_6F => X"00000043000000000000003b0000000000000059000000000000006100000000",
            INIT_70 => X"0000003e000000000000003f000000000000003c000000000000005900000000",
            INIT_71 => X"0000003f000000000000003e000000000000003e000000000000003e00000000",
            INIT_72 => X"000000520000000000000041000000000000003d000000000000003e00000000",
            INIT_73 => X"00000051000000000000004e0000000000000051000000000000005400000000",
            INIT_74 => X"0000005300000000000000550000000000000054000000000000005800000000",
            INIT_75 => X"0000004000000000000000420000000000000043000000000000005000000000",
            INIT_76 => X"0000006700000000000000560000000000000038000000000000003400000000",
            INIT_77 => X"0000004b000000000000003d0000000000000039000000000000004c00000000",
            INIT_78 => X"0000003c000000000000003d000000000000003c000000000000005c00000000",
            INIT_79 => X"0000004100000000000000430000000000000042000000000000003f00000000",
            INIT_7A => X"0000004800000000000000410000000000000043000000000000004200000000",
            INIT_7B => X"0000004600000000000000480000000000000049000000000000004900000000",
            INIT_7C => X"0000004b000000000000004b000000000000004a000000000000004900000000",
            INIT_7D => X"0000003e00000000000000400000000000000040000000000000004b00000000",
            INIT_7E => X"0000004000000000000000580000000000000056000000000000004100000000",
            INIT_7F => X"000000490000000000000040000000000000003c000000000000003900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "sampleifmap_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c000000000000000b300000000000000b0000000000000009c00000000",
            INIT_01 => X"000000ad00000000000000ad00000000000000ab00000000000000b900000000",
            INIT_02 => X"000000b800000000000000b600000000000000b300000000000000af00000000",
            INIT_03 => X"000000b500000000000000b600000000000000b800000000000000b900000000",
            INIT_04 => X"000000b900000000000000b700000000000000b300000000000000b300000000",
            INIT_05 => X"000000bd00000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000b700000000000000ca00000000000000c400000000000000c500000000",
            INIT_08 => X"000000c300000000000000b800000000000000b3000000000000009b00000000",
            INIT_09 => X"000000a4000000000000009f00000000000000a200000000000000be00000000",
            INIT_0A => X"000000b000000000000000a900000000000000a500000000000000a300000000",
            INIT_0B => X"000000a700000000000000a400000000000000ae00000000000000ab00000000",
            INIT_0C => X"000000a600000000000000a800000000000000a600000000000000ac00000000",
            INIT_0D => X"000000a900000000000000ab00000000000000af00000000000000a900000000",
            INIT_0E => X"000000cc00000000000000bf00000000000000ae00000000000000aa00000000",
            INIT_0F => X"000000be00000000000000d700000000000000d000000000000000ce00000000",
            INIT_10 => X"000000c400000000000000b900000000000000b2000000000000009a00000000",
            INIT_11 => X"000000a800000000000000b200000000000000c100000000000000cb00000000",
            INIT_12 => X"000000c400000000000000be00000000000000af00000000000000a000000000",
            INIT_13 => X"000000bc00000000000000be00000000000000c500000000000000c300000000",
            INIT_14 => X"000000c300000000000000c200000000000000c300000000000000c400000000",
            INIT_15 => X"000000bf00000000000000c100000000000000c600000000000000c400000000",
            INIT_16 => X"000000cd00000000000000cd00000000000000c400000000000000c000000000",
            INIT_17 => X"000000bf00000000000000d700000000000000d000000000000000ce00000000",
            INIT_18 => X"000000c300000000000000bc00000000000000b2000000000000009a00000000",
            INIT_19 => X"0000008000000000000000bc00000000000000c500000000000000ca00000000",
            INIT_1A => X"0000009b000000000000009a0000000000000098000000000000006c00000000",
            INIT_1B => X"0000009400000000000000950000000000000095000000000000009e00000000",
            INIT_1C => X"000000ad00000000000000a300000000000000a100000000000000a700000000",
            INIT_1D => X"0000009f00000000000000ae00000000000000a300000000000000a800000000",
            INIT_1E => X"000000ce00000000000000cc00000000000000d000000000000000bc00000000",
            INIT_1F => X"000000bc00000000000000d400000000000000cd00000000000000cc00000000",
            INIT_20 => X"000000bf00000000000000bb00000000000000b1000000000000009a00000000",
            INIT_21 => X"0000007e00000000000000bd00000000000000c400000000000000c600000000",
            INIT_22 => X"0000006b000000000000006a000000000000008b000000000000008000000000",
            INIT_23 => X"0000007100000000000000760000000000000078000000000000007300000000",
            INIT_24 => X"0000007e00000000000000720000000000000072000000000000007700000000",
            INIT_25 => X"0000007000000000000000880000000000000070000000000000007600000000",
            INIT_26 => X"000000ce00000000000000c900000000000000cb00000000000000a000000000",
            INIT_27 => X"000000be00000000000000d600000000000000cd00000000000000ce00000000",
            INIT_28 => X"000000bd00000000000000bb00000000000000ae000000000000009700000000",
            INIT_29 => X"0000009300000000000000b700000000000000c800000000000000c500000000",
            INIT_2A => X"000000a5000000000000009100000000000000a800000000000000a900000000",
            INIT_2B => X"0000009d0000000000000095000000000000009200000000000000aa00000000",
            INIT_2C => X"000000bd00000000000000b000000000000000b200000000000000b400000000",
            INIT_2D => X"000000b100000000000000bc00000000000000b300000000000000b000000000",
            INIT_2E => X"000000d000000000000000cf00000000000000d000000000000000c400000000",
            INIT_2F => X"000000be00000000000000d800000000000000d100000000000000d000000000",
            INIT_30 => X"000000bd00000000000000b900000000000000ac000000000000009800000000",
            INIT_31 => X"00000060000000000000009300000000000000c600000000000000c200000000",
            INIT_32 => X"0000009800000000000000900000000000000097000000000000009500000000",
            INIT_33 => X"0000008b00000000000000800000000000000079000000000000009800000000",
            INIT_34 => X"000000a200000000000000aa0000000000000097000000000000009c00000000",
            INIT_35 => X"000000a4000000000000009600000000000000ad000000000000009600000000",
            INIT_36 => X"000000d200000000000000cc00000000000000a6000000000000009c00000000",
            INIT_37 => X"000000bc00000000000000d400000000000000cf00000000000000d300000000",
            INIT_38 => X"000000bb00000000000000b600000000000000ac000000000000009b00000000",
            INIT_39 => X"00000065000000000000007700000000000000b500000000000000c200000000",
            INIT_3A => X"0000007800000000000000830000000000000083000000000000007b00000000",
            INIT_3B => X"0000007f00000000000000870000000000000087000000000000009200000000",
            INIT_3C => X"0000007b0000000000000083000000000000007b000000000000007b00000000",
            INIT_3D => X"0000009f000000000000007b0000000000000084000000000000006d00000000",
            INIT_3E => X"000000c700000000000000bf0000000000000084000000000000007b00000000",
            INIT_3F => X"000000ba00000000000000d000000000000000c900000000000000c900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b900000000000000b400000000000000af00000000000000a100000000",
            INIT_41 => X"000000af00000000000000ab00000000000000ba00000000000000c000000000",
            INIT_42 => X"000000a600000000000000ac00000000000000a500000000000000a200000000",
            INIT_43 => X"000000aa00000000000000ad00000000000000ac00000000000000af00000000",
            INIT_44 => X"000000af00000000000000b200000000000000b200000000000000ac00000000",
            INIT_45 => X"000000be00000000000000b200000000000000ac00000000000000a300000000",
            INIT_46 => X"000000cd00000000000000c800000000000000b000000000000000ac00000000",
            INIT_47 => X"000000b900000000000000d100000000000000c900000000000000c800000000",
            INIT_48 => X"000000ba00000000000000b400000000000000b700000000000000ac00000000",
            INIT_49 => X"000000b700000000000000c200000000000000c000000000000000be00000000",
            INIT_4A => X"000000a300000000000000a200000000000000a500000000000000a000000000",
            INIT_4B => X"000000a200000000000000a4000000000000009e000000000000009f00000000",
            INIT_4C => X"000000a200000000000000ac00000000000000ae00000000000000a700000000",
            INIT_4D => X"000000b600000000000000a500000000000000a300000000000000a000000000",
            INIT_4E => X"000000cd00000000000000ca00000000000000c600000000000000c800000000",
            INIT_4F => X"000000b800000000000000d000000000000000ca00000000000000ca00000000",
            INIT_50 => X"000000be00000000000000ba00000000000000c400000000000000b100000000",
            INIT_51 => X"000000b700000000000000c100000000000000c100000000000000c000000000",
            INIT_52 => X"0000009f00000000000000a500000000000000a700000000000000a300000000",
            INIT_53 => X"000000ac00000000000000aa00000000000000a600000000000000a400000000",
            INIT_54 => X"000000ab00000000000000a600000000000000a600000000000000a800000000",
            INIT_55 => X"000000b200000000000000ab00000000000000ad00000000000000a800000000",
            INIT_56 => X"000000c700000000000000c700000000000000c600000000000000c700000000",
            INIT_57 => X"000000b800000000000000d000000000000000c800000000000000c800000000",
            INIT_58 => X"000000c800000000000000c300000000000000cc00000000000000b700000000",
            INIT_59 => X"000000c600000000000000be00000000000000bb00000000000000c900000000",
            INIT_5A => X"000000c100000000000000c100000000000000c100000000000000c200000000",
            INIT_5B => X"000000c600000000000000c600000000000000c200000000000000c100000000",
            INIT_5C => X"000000c600000000000000c300000000000000c300000000000000c600000000",
            INIT_5D => X"000000c500000000000000c400000000000000c400000000000000c500000000",
            INIT_5E => X"000000c900000000000000c900000000000000cb00000000000000c900000000",
            INIT_5F => X"000000bb00000000000000d100000000000000c800000000000000ca00000000",
            INIT_60 => X"000000b200000000000000c600000000000000cd00000000000000b900000000",
            INIT_61 => X"000000c4000000000000009a000000000000008d00000000000000a600000000",
            INIT_62 => X"000000c500000000000000c700000000000000ca00000000000000ca00000000",
            INIT_63 => X"000000ca00000000000000c900000000000000c700000000000000c500000000",
            INIT_64 => X"000000c400000000000000c600000000000000c700000000000000c900000000",
            INIT_65 => X"000000c600000000000000c700000000000000c600000000000000c400000000",
            INIT_66 => X"000000ce00000000000000cb00000000000000ca00000000000000c700000000",
            INIT_67 => X"000000bd00000000000000d400000000000000ce00000000000000cf00000000",
            INIT_68 => X"000000a500000000000000c800000000000000d000000000000000ba00000000",
            INIT_69 => X"0000006b000000000000005f000000000000007c000000000000009000000000",
            INIT_6A => X"000000c700000000000000c700000000000000b3000000000000008f00000000",
            INIT_6B => X"000000cc00000000000000c900000000000000c600000000000000c500000000",
            INIT_6C => X"000000cc00000000000000ce00000000000000cd00000000000000cc00000000",
            INIT_6D => X"000000cd00000000000000cd00000000000000c900000000000000c900000000",
            INIT_6E => X"000000cb00000000000000cb00000000000000cb00000000000000cc00000000",
            INIT_6F => X"000000b700000000000000cf00000000000000ca00000000000000ca00000000",
            INIT_70 => X"000000cc00000000000000d000000000000000d400000000000000ba00000000",
            INIT_71 => X"0000005b000000000000008f00000000000000c100000000000000ce00000000",
            INIT_72 => X"000000b5000000000000008e0000000000000065000000000000005100000000",
            INIT_73 => X"000000cf00000000000000cf00000000000000cc00000000000000c600000000",
            INIT_74 => X"000000ca00000000000000cf00000000000000cf00000000000000cf00000000",
            INIT_75 => X"000000c500000000000000c600000000000000c500000000000000c500000000",
            INIT_76 => X"000000c500000000000000c500000000000000c500000000000000c500000000",
            INIT_77 => X"000000b500000000000000cc00000000000000c500000000000000c400000000",
            INIT_78 => X"000000ce00000000000000d200000000000000d600000000000000b800000000",
            INIT_79 => X"000000b300000000000000cf00000000000000d400000000000000d100000000",
            INIT_7A => X"00000080000000000000005d0000000000000053000000000000007400000000",
            INIT_7B => X"000000ce00000000000000d200000000000000cb00000000000000ae00000000",
            INIT_7C => X"000000c900000000000000ca00000000000000ca00000000000000cc00000000",
            INIT_7D => X"000000c900000000000000c900000000000000c700000000000000c600000000",
            INIT_7E => X"000000c700000000000000c900000000000000ca00000000000000c800000000",
            INIT_7F => X"000000b400000000000000cb00000000000000c600000000000000c600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "sampleifmap_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d500000000000000d600000000000000d700000000000000ba00000000",
            INIT_01 => X"000000d900000000000000d400000000000000d600000000000000d600000000",
            INIT_02 => X"000000560000000000000049000000000000005b00000000000000af00000000",
            INIT_03 => X"000000cc00000000000000b5000000000000008a000000000000006500000000",
            INIT_04 => X"000000c600000000000000c700000000000000cb00000000000000d000000000",
            INIT_05 => X"000000c800000000000000c900000000000000c900000000000000c700000000",
            INIT_06 => X"000000c900000000000000c900000000000000ca00000000000000c800000000",
            INIT_07 => X"000000b600000000000000cc00000000000000c800000000000000ca00000000",
            INIT_08 => X"000000d900000000000000d800000000000000d800000000000000bb00000000",
            INIT_09 => X"000000d300000000000000d600000000000000d900000000000000db00000000",
            INIT_0A => X"000000520000000000000044000000000000007b00000000000000cc00000000",
            INIT_0B => X"0000008200000000000000610000000000000051000000000000004f00000000",
            INIT_0C => X"000000ca00000000000000c900000000000000bc00000000000000a500000000",
            INIT_0D => X"000000c600000000000000c700000000000000c100000000000000c400000000",
            INIT_0E => X"000000c800000000000000c800000000000000c700000000000000c600000000",
            INIT_0F => X"000000b600000000000000cc00000000000000c700000000000000c900000000",
            INIT_10 => X"000000d600000000000000d500000000000000d900000000000000bc00000000",
            INIT_11 => X"000000d200000000000000d600000000000000d800000000000000d800000000",
            INIT_12 => X"000000530000000000000046000000000000008800000000000000d400000000",
            INIT_13 => X"0000004d00000000000000500000000000000050000000000000004e00000000",
            INIT_14 => X"00000097000000000000007e0000000000000066000000000000005300000000",
            INIT_15 => X"000000cc00000000000000c900000000000000b2000000000000009f00000000",
            INIT_16 => X"000000c600000000000000c800000000000000c900000000000000cb00000000",
            INIT_17 => X"000000b400000000000000c900000000000000c500000000000000c700000000",
            INIT_18 => X"000000d500000000000000d600000000000000da00000000000000bb00000000",
            INIT_19 => X"000000d800000000000000d700000000000000d800000000000000d700000000",
            INIT_1A => X"00000037000000000000002d000000000000007000000000000000cc00000000",
            INIT_1B => X"00000051000000000000004d0000000000000045000000000000003a00000000",
            INIT_1C => X"0000003e0000000000000046000000000000004d000000000000005000000000",
            INIT_1D => X"000000a0000000000000007c000000000000004f000000000000003b00000000",
            INIT_1E => X"000000cd00000000000000cd00000000000000c400000000000000b500000000",
            INIT_1F => X"000000b400000000000000ca00000000000000c800000000000000cb00000000",
            INIT_20 => X"000000d100000000000000d200000000000000d800000000000000bc00000000",
            INIT_21 => X"000000d400000000000000d400000000000000d600000000000000d300000000",
            INIT_22 => X"00000021000000000000003a000000000000005f000000000000009a00000000",
            INIT_23 => X"0000004d0000000000000041000000000000003e000000000000003000000000",
            INIT_24 => X"0000004800000000000000540000000000000054000000000000005200000000",
            INIT_25 => X"00000048000000000000003f000000000000002f000000000000003800000000",
            INIT_26 => X"0000009e0000000000000084000000000000006b000000000000004e00000000",
            INIT_27 => X"000000b600000000000000ca00000000000000c100000000000000b500000000",
            INIT_28 => X"000000cf00000000000000ce00000000000000d200000000000000b800000000",
            INIT_29 => X"000000c800000000000000d400000000000000d300000000000000d100000000",
            INIT_2A => X"00000061000000000000008f0000000000000085000000000000009100000000",
            INIT_2B => X"0000005a000000000000002e0000000000000032000000000000002d00000000",
            INIT_2C => X"00000047000000000000007f000000000000009e000000000000009600000000",
            INIT_2D => X"0000004100000000000000580000000000000070000000000000006100000000",
            INIT_2E => X"000000a200000000000000a50000000000000082000000000000004300000000",
            INIT_2F => X"000000b000000000000000c500000000000000b500000000000000a800000000",
            INIT_30 => X"000000d000000000000000cd00000000000000d200000000000000b700000000",
            INIT_31 => X"000000d200000000000000d500000000000000d400000000000000d300000000",
            INIT_32 => X"000000bf00000000000000d400000000000000d100000000000000d100000000",
            INIT_33 => X"000000a600000000000000930000000000000093000000000000009400000000",
            INIT_34 => X"0000009d00000000000000c300000000000000d000000000000000c800000000",
            INIT_35 => X"000000a200000000000000b400000000000000b500000000000000a600000000",
            INIT_36 => X"000000c500000000000000c100000000000000b4000000000000009f00000000",
            INIT_37 => X"000000b100000000000000c700000000000000c100000000000000c300000000",
            INIT_38 => X"000000c200000000000000c300000000000000c400000000000000ae00000000",
            INIT_39 => X"000000b900000000000000bb00000000000000be00000000000000c200000000",
            INIT_3A => X"000000b500000000000000b700000000000000b500000000000000b800000000",
            INIT_3B => X"000000ad00000000000000ae00000000000000b000000000000000b200000000",
            INIT_3C => X"000000ac00000000000000a600000000000000a400000000000000aa00000000",
            INIT_3D => X"000000b000000000000000aa00000000000000a600000000000000aa00000000",
            INIT_3E => X"0000009b000000000000009d00000000000000a500000000000000af00000000",
            INIT_3F => X"0000009e00000000000000af00000000000000a3000000000000009d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000070000000000000006c000000000000007000000000",
            INIT_41 => X"0000006000000000000000610000000000000064000000000000006700000000",
            INIT_42 => X"00000057000000000000005e000000000000005a000000000000005c00000000",
            INIT_43 => X"0000006700000000000000570000000000000053000000000000005400000000",
            INIT_44 => X"00000070000000000000006f0000000000000070000000000000007300000000",
            INIT_45 => X"0000007600000000000000740000000000000073000000000000007100000000",
            INIT_46 => X"0000007b000000000000007c000000000000007b000000000000007a00000000",
            INIT_47 => X"0000007c0000000000000084000000000000007a000000000000007900000000",
            INIT_48 => X"0000007000000000000000710000000000000073000000000000007500000000",
            INIT_49 => X"000000710000000000000071000000000000006f000000000000007100000000",
            INIT_4A => X"0000006e000000000000006f0000000000000070000000000000006f00000000",
            INIT_4B => X"0000006b000000000000006e000000000000006d000000000000006e00000000",
            INIT_4C => X"0000006e000000000000006c0000000000000073000000000000007300000000",
            INIT_4D => X"0000006b0000000000000068000000000000006d000000000000006f00000000",
            INIT_4E => X"000000700000000000000070000000000000006e000000000000006d00000000",
            INIT_4F => X"000000650000000000000062000000000000005f000000000000006400000000",
            INIT_50 => X"0000006a00000000000000690000000000000066000000000000007100000000",
            INIT_51 => X"0000005d00000000000000610000000000000066000000000000006a00000000",
            INIT_52 => X"000000550000000000000059000000000000005e000000000000005f00000000",
            INIT_53 => X"0000004e000000000000004f000000000000004e000000000000005200000000",
            INIT_54 => X"000000440000000000000047000000000000004f000000000000005000000000",
            INIT_55 => X"0000004100000000000000410000000000000041000000000000004300000000",
            INIT_56 => X"0000004100000000000000420000000000000042000000000000004100000000",
            INIT_57 => X"0000006400000000000000470000000000000037000000000000003c00000000",
            INIT_58 => X"000000400000000000000041000000000000003c000000000000005400000000",
            INIT_59 => X"0000003c000000000000003e0000000000000040000000000000004000000000",
            INIT_5A => X"00000038000000000000003d0000000000000040000000000000004200000000",
            INIT_5B => X"0000003f000000000000003d000000000000003c000000000000003900000000",
            INIT_5C => X"0000003b00000000000000410000000000000043000000000000004000000000",
            INIT_5D => X"0000003c000000000000003b000000000000003a000000000000003800000000",
            INIT_5E => X"0000003800000000000000380000000000000039000000000000003a00000000",
            INIT_5F => X"0000008000000000000000750000000000000048000000000000003800000000",
            INIT_60 => X"0000003e000000000000003f000000000000003b000000000000005300000000",
            INIT_61 => X"0000003f000000000000003d0000000000000041000000000000003f00000000",
            INIT_62 => X"00000039000000000000003c000000000000003e000000000000004300000000",
            INIT_63 => X"0000003d000000000000003c000000000000003a000000000000003a00000000",
            INIT_64 => X"0000003e00000000000000400000000000000044000000000000004100000000",
            INIT_65 => X"0000003d000000000000003e000000000000003c000000000000003d00000000",
            INIT_66 => X"00000041000000000000003d000000000000003a000000000000003a00000000",
            INIT_67 => X"0000006300000000000000890000000000000088000000000000005b00000000",
            INIT_68 => X"00000039000000000000003d0000000000000035000000000000004f00000000",
            INIT_69 => X"0000003c000000000000003a000000000000003b000000000000003700000000",
            INIT_6A => X"000000370000000000000039000000000000003c000000000000003d00000000",
            INIT_6B => X"0000003f000000000000003d000000000000003e000000000000003c00000000",
            INIT_6C => X"0000003b000000000000003c000000000000003f000000000000004300000000",
            INIT_6D => X"0000003f0000000000000040000000000000003e000000000000003e00000000",
            INIT_6E => X"0000006e0000000000000047000000000000003c000000000000003e00000000",
            INIT_6F => X"0000004a000000000000004f0000000000000077000000000000008e00000000",
            INIT_70 => X"000000410000000000000042000000000000003a000000000000005200000000",
            INIT_71 => X"0000003e000000000000003e000000000000003e000000000000003f00000000",
            INIT_72 => X"0000004f0000000000000041000000000000003e000000000000003f00000000",
            INIT_73 => X"0000004d000000000000004a000000000000004c000000000000004f00000000",
            INIT_74 => X"0000004e00000000000000500000000000000050000000000000005400000000",
            INIT_75 => X"00000041000000000000003e000000000000003f000000000000004c00000000",
            INIT_76 => X"0000008d000000000000007c0000000000000056000000000000004200000000",
            INIT_77 => X"0000004500000000000000400000000000000042000000000000006600000000",
            INIT_78 => X"0000003a000000000000003a0000000000000034000000000000004e00000000",
            INIT_79 => X"00000039000000000000003b000000000000003a000000000000003a00000000",
            INIT_7A => X"00000045000000000000003a000000000000003b000000000000003a00000000",
            INIT_7B => X"0000004500000000000000460000000000000047000000000000004700000000",
            INIT_7C => X"0000004a00000000000000490000000000000048000000000000004800000000",
            INIT_7D => X"00000044000000000000003f000000000000003f000000000000004900000000",
            INIT_7E => X"0000005800000000000000800000000000000080000000000000005a00000000",
            INIT_7F => X"000000440000000000000041000000000000003f000000000000004200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "sampleifmap_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000cd00000000000000c100000000000000bb000000000000009500000000",
            INIT_01 => X"000000b400000000000000b500000000000000b700000000000000ca00000000",
            INIT_02 => X"000000c000000000000000c100000000000000bd00000000000000b600000000",
            INIT_03 => X"000000bd00000000000000bd00000000000000c000000000000000c000000000",
            INIT_04 => X"000000c000000000000000bd00000000000000b900000000000000ba00000000",
            INIT_05 => X"000000be00000000000000c000000000000000c100000000000000c100000000",
            INIT_06 => X"000000c300000000000000bc00000000000000bb00000000000000bb00000000",
            INIT_07 => X"000000ab00000000000000d400000000000000d100000000000000ca00000000",
            INIT_08 => X"000000e300000000000000d700000000000000cc000000000000009d00000000",
            INIT_09 => X"000000b300000000000000b300000000000000be00000000000000e000000000",
            INIT_0A => X"000000c300000000000000c300000000000000bb00000000000000b300000000",
            INIT_0B => X"000000b700000000000000b400000000000000be00000000000000bb00000000",
            INIT_0C => X"000000b700000000000000b800000000000000b700000000000000bc00000000",
            INIT_0D => X"000000bc00000000000000bc00000000000000bf00000000000000b900000000",
            INIT_0E => X"000000e000000000000000d300000000000000c200000000000000be00000000",
            INIT_0F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_10 => X"000000db00000000000000d500000000000000c9000000000000009900000000",
            INIT_11 => X"000000b800000000000000c400000000000000d500000000000000df00000000",
            INIT_12 => X"000000d400000000000000d300000000000000c300000000000000b100000000",
            INIT_13 => X"000000ca00000000000000cc00000000000000d200000000000000d000000000",
            INIT_14 => X"000000d100000000000000d000000000000000d100000000000000d100000000",
            INIT_15 => X"000000d000000000000000d000000000000000d400000000000000d200000000",
            INIT_16 => X"000000df00000000000000de00000000000000d500000000000000d000000000",
            INIT_17 => X"000000b800000000000000e000000000000000d700000000000000da00000000",
            INIT_18 => X"000000de00000000000000d300000000000000cf00000000000000a600000000",
            INIT_19 => X"0000008300000000000000c900000000000000dc00000000000000e200000000",
            INIT_1A => X"000000b100000000000000a6000000000000009e000000000000007700000000",
            INIT_1B => X"000000ab00000000000000a600000000000000a700000000000000b200000000",
            INIT_1C => X"000000ba00000000000000b200000000000000b200000000000000b700000000",
            INIT_1D => X"000000a500000000000000b400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000dd00000000000000dc00000000000000e400000000000000cf00000000",
            INIT_1F => X"000000ba00000000000000e600000000000000df00000000000000e000000000",
            INIT_20 => X"000000da00000000000000ca00000000000000cb00000000000000a700000000",
            INIT_21 => X"0000008e00000000000000d600000000000000e100000000000000e000000000",
            INIT_22 => X"0000008100000000000000780000000000000098000000000000009900000000",
            INIT_23 => X"00000083000000000000007c000000000000007e000000000000008100000000",
            INIT_24 => X"0000008a00000000000000820000000000000084000000000000008600000000",
            INIT_25 => X"0000007b000000000000008d0000000000000088000000000000008800000000",
            INIT_26 => X"000000d900000000000000da00000000000000e300000000000000ba00000000",
            INIT_27 => X"000000b900000000000000e300000000000000dc00000000000000de00000000",
            INIT_28 => X"000000d900000000000000cb00000000000000c900000000000000a400000000",
            INIT_29 => X"000000a500000000000000d100000000000000da00000000000000dc00000000",
            INIT_2A => X"000000b4000000000000009c00000000000000b500000000000000c400000000",
            INIT_2B => X"000000ac00000000000000a300000000000000a000000000000000b300000000",
            INIT_2C => X"000000c900000000000000be00000000000000c100000000000000bf00000000",
            INIT_2D => X"000000be00000000000000c600000000000000c000000000000000bf00000000",
            INIT_2E => X"000000e100000000000000e100000000000000e100000000000000d400000000",
            INIT_2F => X"000000bc00000000000000e800000000000000e100000000000000df00000000",
            INIT_30 => X"000000d900000000000000c800000000000000c600000000000000a400000000",
            INIT_31 => X"0000006800000000000000ac00000000000000d600000000000000d900000000",
            INIT_32 => X"000000af00000000000000a600000000000000a5000000000000009e00000000",
            INIT_33 => X"000000a00000000000000097000000000000009000000000000000a500000000",
            INIT_34 => X"000000b600000000000000bd00000000000000ad00000000000000b200000000",
            INIT_35 => X"000000b900000000000000ad00000000000000b700000000000000aa00000000",
            INIT_36 => X"000000e200000000000000dc00000000000000b200000000000000a600000000",
            INIT_37 => X"000000bc00000000000000e700000000000000e000000000000000dd00000000",
            INIT_38 => X"000000d800000000000000c700000000000000c900000000000000a900000000",
            INIT_39 => X"0000006f000000000000009200000000000000cb00000000000000da00000000",
            INIT_3A => X"00000090000000000000009d0000000000000095000000000000008600000000",
            INIT_3B => X"00000090000000000000008f000000000000008f000000000000009b00000000",
            INIT_3C => X"0000008e0000000000000094000000000000008e000000000000009300000000",
            INIT_3D => X"000000b0000000000000008e000000000000008d000000000000007f00000000",
            INIT_3E => X"000000dc00000000000000d10000000000000095000000000000008900000000",
            INIT_3F => X"000000ba00000000000000e400000000000000dc00000000000000d900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d900000000000000c700000000000000ce00000000000000b100000000",
            INIT_41 => X"000000c500000000000000c100000000000000cd00000000000000db00000000",
            INIT_42 => X"000000b800000000000000bb00000000000000b700000000000000b800000000",
            INIT_43 => X"000000bd00000000000000bb00000000000000ba00000000000000c000000000",
            INIT_44 => X"000000bf00000000000000c200000000000000c200000000000000c000000000",
            INIT_45 => X"000000c800000000000000bc00000000000000ba00000000000000b200000000",
            INIT_46 => X"000000db00000000000000d600000000000000c600000000000000c100000000",
            INIT_47 => X"000000b900000000000000e400000000000000dd00000000000000db00000000",
            INIT_48 => X"000000d600000000000000c500000000000000d400000000000000ba00000000",
            INIT_49 => X"000000d200000000000000dc00000000000000d600000000000000d700000000",
            INIT_4A => X"000000ba00000000000000b600000000000000bb00000000000000b900000000",
            INIT_4B => X"000000ba00000000000000b900000000000000b400000000000000b600000000",
            INIT_4C => X"000000b800000000000000c300000000000000c600000000000000c100000000",
            INIT_4D => X"000000c600000000000000b600000000000000b600000000000000b500000000",
            INIT_4E => X"000000df00000000000000dd00000000000000de00000000000000de00000000",
            INIT_4F => X"000000b700000000000000e300000000000000de00000000000000df00000000",
            INIT_50 => X"000000d800000000000000c800000000000000de00000000000000bc00000000",
            INIT_51 => X"000000cc00000000000000d600000000000000d400000000000000d700000000",
            INIT_52 => X"000000b000000000000000b600000000000000b800000000000000b500000000",
            INIT_53 => X"000000bf00000000000000bc00000000000000b800000000000000b500000000",
            INIT_54 => X"000000b900000000000000b800000000000000ba00000000000000bd00000000",
            INIT_55 => X"000000c900000000000000ba00000000000000b800000000000000b600000000",
            INIT_56 => X"000000db00000000000000dc00000000000000dd00000000000000df00000000",
            INIT_57 => X"000000b800000000000000e300000000000000dc00000000000000db00000000",
            INIT_58 => X"000000e000000000000000cf00000000000000e200000000000000bf00000000",
            INIT_59 => X"000000de00000000000000d700000000000000d100000000000000dc00000000",
            INIT_5A => X"000000d700000000000000d600000000000000d700000000000000d900000000",
            INIT_5B => X"000000df00000000000000df00000000000000db00000000000000d900000000",
            INIT_5C => X"000000da00000000000000db00000000000000dd00000000000000df00000000",
            INIT_5D => X"000000db00000000000000d900000000000000d600000000000000d800000000",
            INIT_5E => X"000000d600000000000000d900000000000000db00000000000000db00000000",
            INIT_5F => X"000000ba00000000000000e300000000000000db00000000000000d700000000",
            INIT_60 => X"000000ce00000000000000d400000000000000dc00000000000000bc00000000",
            INIT_61 => X"000000d900000000000000ac000000000000009900000000000000b500000000",
            INIT_62 => X"000000dc00000000000000dd00000000000000e100000000000000e200000000",
            INIT_63 => X"000000e200000000000000e100000000000000df00000000000000de00000000",
            INIT_64 => X"000000da00000000000000dc00000000000000dd00000000000000e100000000",
            INIT_65 => X"000000da00000000000000dc00000000000000db00000000000000d900000000",
            INIT_66 => X"000000e000000000000000de00000000000000dc00000000000000d900000000",
            INIT_67 => X"000000bb00000000000000e600000000000000e000000000000000e000000000",
            INIT_68 => X"000000c100000000000000d600000000000000df00000000000000bd00000000",
            INIT_69 => X"000000730000000000000063000000000000007e000000000000009d00000000",
            INIT_6A => X"000000dd00000000000000dd00000000000000c6000000000000009d00000000",
            INIT_6B => X"000000e200000000000000df00000000000000dc00000000000000da00000000",
            INIT_6C => X"000000df00000000000000e100000000000000e000000000000000e200000000",
            INIT_6D => X"000000e000000000000000e000000000000000dd00000000000000dc00000000",
            INIT_6E => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_6F => X"000000b700000000000000e200000000000000dd00000000000000dd00000000",
            INIT_70 => X"000000e900000000000000de00000000000000e200000000000000bd00000000",
            INIT_71 => X"0000005a000000000000009200000000000000c400000000000000dc00000000",
            INIT_72 => X"000000ca00000000000000a10000000000000071000000000000005400000000",
            INIT_73 => X"000000e400000000000000e300000000000000e000000000000000da00000000",
            INIT_74 => X"000000dc00000000000000e000000000000000e100000000000000e200000000",
            INIT_75 => X"000000d900000000000000d800000000000000d700000000000000d700000000",
            INIT_76 => X"000000d800000000000000d800000000000000d800000000000000d800000000",
            INIT_77 => X"000000b600000000000000e100000000000000da00000000000000d700000000",
            INIT_78 => X"000000ea00000000000000e000000000000000e500000000000000bb00000000",
            INIT_79 => X"000000b300000000000000da00000000000000e100000000000000e100000000",
            INIT_7A => X"00000091000000000000006a0000000000000058000000000000007300000000",
            INIT_7B => X"000000e100000000000000e400000000000000dd00000000000000c000000000",
            INIT_7C => X"000000d900000000000000da00000000000000db00000000000000df00000000",
            INIT_7D => X"000000db00000000000000d900000000000000d600000000000000d600000000",
            INIT_7E => X"000000da00000000000000dc00000000000000dd00000000000000db00000000",
            INIT_7F => X"000000b700000000000000e200000000000000dc00000000000000d900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "sampleifmap_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000e900000000000000de00000000000000e900000000000000be00000000",
            INIT_01 => X"000000e100000000000000e000000000000000e200000000000000e400000000",
            INIT_02 => X"0000005b0000000000000050000000000000006200000000000000b500000000",
            INIT_03 => X"000000d900000000000000c00000000000000092000000000000006a00000000",
            INIT_04 => X"000000da00000000000000dd00000000000000e100000000000000e000000000",
            INIT_05 => X"000000d900000000000000da00000000000000da00000000000000d900000000",
            INIT_06 => X"000000dd00000000000000dd00000000000000dd00000000000000da00000000",
            INIT_07 => X"000000bc00000000000000e300000000000000dc00000000000000dd00000000",
            INIT_08 => X"000000e900000000000000dd00000000000000ea00000000000000bf00000000",
            INIT_09 => X"000000dd00000000000000e200000000000000e300000000000000e700000000",
            INIT_0A => X"0000004f0000000000000049000000000000008200000000000000d500000000",
            INIT_0B => X"0000008800000000000000640000000000000050000000000000004b00000000",
            INIT_0C => X"000000dc00000000000000d700000000000000c800000000000000ad00000000",
            INIT_0D => X"000000de00000000000000df00000000000000d900000000000000d900000000",
            INIT_0E => X"000000db00000000000000db00000000000000dd00000000000000dd00000000",
            INIT_0F => X"000000bd00000000000000e300000000000000db00000000000000da00000000",
            INIT_10 => X"000000e400000000000000d900000000000000e800000000000000bd00000000",
            INIT_11 => X"000000dc00000000000000e200000000000000e100000000000000e300000000",
            INIT_12 => X"00000050000000000000004a000000000000009000000000000000dd00000000",
            INIT_13 => X"0000004c000000000000004e000000000000004c000000000000004a00000000",
            INIT_14 => X"000000a100000000000000810000000000000064000000000000005300000000",
            INIT_15 => X"000000e200000000000000e100000000000000c900000000000000b000000000",
            INIT_16 => X"000000d700000000000000d900000000000000dc00000000000000df00000000",
            INIT_17 => X"000000bb00000000000000e100000000000000d900000000000000d700000000",
            INIT_18 => X"000000e100000000000000d700000000000000e800000000000000bb00000000",
            INIT_19 => X"000000e200000000000000e300000000000000e100000000000000e000000000",
            INIT_1A => X"000000380000000000000032000000000000007700000000000000d500000000",
            INIT_1B => X"00000052000000000000004d0000000000000045000000000000003b00000000",
            INIT_1C => X"0000003f00000000000000420000000000000048000000000000005000000000",
            INIT_1D => X"000000a20000000000000085000000000000005b000000000000004100000000",
            INIT_1E => X"000000df00000000000000da00000000000000cc00000000000000b800000000",
            INIT_1F => X"000000bc00000000000000e300000000000000dd00000000000000dd00000000",
            INIT_20 => X"000000df00000000000000de00000000000000e700000000000000b700000000",
            INIT_21 => X"000000e100000000000000e400000000000000e600000000000000df00000000",
            INIT_22 => X"00000027000000000000003c000000000000006200000000000000a200000000",
            INIT_23 => X"0000004e00000000000000440000000000000043000000000000003500000000",
            INIT_24 => X"0000004800000000000000530000000000000052000000000000005100000000",
            INIT_25 => X"00000043000000000000003f0000000000000031000000000000003900000000",
            INIT_26 => X"000000a8000000000000008b000000000000006d000000000000004b00000000",
            INIT_27 => X"000000c300000000000000df00000000000000d700000000000000c600000000",
            INIT_28 => X"000000de00000000000000e200000000000000e200000000000000b000000000",
            INIT_29 => X"000000d400000000000000e200000000000000e200000000000000de00000000",
            INIT_2A => X"0000006a0000000000000096000000000000008b000000000000009b00000000",
            INIT_2B => X"0000005e00000000000000330000000000000039000000000000003500000000",
            INIT_2C => X"00000049000000000000008200000000000000a1000000000000009a00000000",
            INIT_2D => X"00000043000000000000005a0000000000000072000000000000006300000000",
            INIT_2E => X"000000a900000000000000ab0000000000000086000000000000004500000000",
            INIT_2F => X"000000be00000000000000d000000000000000c500000000000000b700000000",
            INIT_30 => X"000000df00000000000000e100000000000000e100000000000000af00000000",
            INIT_31 => X"000000de00000000000000de00000000000000de00000000000000df00000000",
            INIT_32 => X"000000cc00000000000000e400000000000000e000000000000000de00000000",
            INIT_33 => X"000000b300000000000000a0000000000000009f000000000000009f00000000",
            INIT_34 => X"000000a900000000000000cf00000000000000dc00000000000000d600000000",
            INIT_35 => X"000000ad00000000000000c000000000000000c100000000000000b200000000",
            INIT_36 => X"000000d600000000000000d200000000000000c300000000000000ab00000000",
            INIT_37 => X"000000bd00000000000000d200000000000000d100000000000000d800000000",
            INIT_38 => X"000000d100000000000000d700000000000000d400000000000000a600000000",
            INIT_39 => X"000000c700000000000000c900000000000000cc00000000000000ce00000000",
            INIT_3A => X"000000c200000000000000c500000000000000c300000000000000c700000000",
            INIT_3B => X"000000c400000000000000c200000000000000c100000000000000c000000000",
            INIT_3C => X"000000ca00000000000000c400000000000000c200000000000000c400000000",
            INIT_3D => X"000000cd00000000000000c800000000000000c400000000000000c800000000",
            INIT_3E => X"000000bf00000000000000c000000000000000c500000000000000ce00000000",
            INIT_3F => X"000000b500000000000000c900000000000000c500000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007800000000000000820000000000000078000000000000006500000000",
            INIT_41 => X"0000006a000000000000006b0000000000000070000000000000007600000000",
            INIT_42 => X"0000006300000000000000660000000000000062000000000000006500000000",
            INIT_43 => X"00000080000000000000006c0000000000000065000000000000006200000000",
            INIT_44 => X"0000009300000000000000920000000000000092000000000000009000000000",
            INIT_45 => X"0000009e00000000000000980000000000000096000000000000009400000000",
            INIT_46 => X"000000a800000000000000a800000000000000a600000000000000a400000000",
            INIT_47 => X"0000009200000000000000a700000000000000a500000000000000a800000000",
            INIT_48 => X"0000008600000000000000860000000000000082000000000000006f00000000",
            INIT_49 => X"0000008800000000000000890000000000000088000000000000008a00000000",
            INIT_4A => X"0000007e00000000000000830000000000000086000000000000008400000000",
            INIT_4B => X"0000008300000000000000830000000000000080000000000000007f00000000",
            INIT_4C => X"00000081000000000000007f0000000000000086000000000000008a00000000",
            INIT_4D => X"0000007e000000000000007c0000000000000080000000000000008100000000",
            INIT_4E => X"0000008400000000000000840000000000000082000000000000008100000000",
            INIT_4F => X"0000006000000000000000730000000000000073000000000000007700000000",
            INIT_50 => X"0000007800000000000000780000000000000071000000000000006800000000",
            INIT_51 => X"00000064000000000000006c0000000000000076000000000000007a00000000",
            INIT_52 => X"000000590000000000000055000000000000005b000000000000006000000000",
            INIT_53 => X"0000005600000000000000570000000000000055000000000000005800000000",
            INIT_54 => X"000000430000000000000046000000000000004f000000000000005600000000",
            INIT_55 => X"0000003c000000000000003f0000000000000041000000000000004200000000",
            INIT_56 => X"0000003b000000000000003c000000000000003c000000000000003b00000000",
            INIT_57 => X"0000004b000000000000003f0000000000000032000000000000003600000000",
            INIT_58 => X"00000039000000000000003d0000000000000037000000000000003d00000000",
            INIT_59 => X"00000036000000000000003b000000000000003f000000000000003a00000000",
            INIT_5A => X"0000002f000000000000002f0000000000000033000000000000003800000000",
            INIT_5B => X"0000003200000000000000310000000000000032000000000000003000000000",
            INIT_5C => X"0000002f00000000000000350000000000000037000000000000003300000000",
            INIT_5D => X"000000370000000000000032000000000000002e000000000000002d00000000",
            INIT_5E => X"0000003400000000000000340000000000000034000000000000003600000000",
            INIT_5F => X"000000680000000000000068000000000000003a000000000000003000000000",
            INIT_60 => X"0000003c0000000000000041000000000000003d000000000000004400000000",
            INIT_61 => X"000000390000000000000037000000000000003d000000000000003e00000000",
            INIT_62 => X"0000003a00000000000000370000000000000038000000000000003d00000000",
            INIT_63 => X"0000003600000000000000380000000000000038000000000000003b00000000",
            INIT_64 => X"000000340000000000000037000000000000003b000000000000003900000000",
            INIT_65 => X"0000003400000000000000340000000000000033000000000000003300000000",
            INIT_66 => X"0000003900000000000000370000000000000035000000000000003300000000",
            INIT_67 => X"0000004b00000000000000780000000000000071000000000000004b00000000",
            INIT_68 => X"00000035000000000000003b0000000000000034000000000000003e00000000",
            INIT_69 => X"0000003600000000000000340000000000000039000000000000003900000000",
            INIT_6A => X"0000003200000000000000300000000000000032000000000000003600000000",
            INIT_6B => X"0000003500000000000000340000000000000038000000000000003900000000",
            INIT_6C => X"0000003300000000000000340000000000000036000000000000003900000000",
            INIT_6D => X"0000003000000000000000350000000000000037000000000000003600000000",
            INIT_6E => X"0000005f000000000000003d0000000000000034000000000000003200000000",
            INIT_6F => X"00000032000000000000003e0000000000000065000000000000007c00000000",
            INIT_70 => X"00000037000000000000003a0000000000000035000000000000003e00000000",
            INIT_71 => X"0000003c000000000000003c000000000000003d000000000000003b00000000",
            INIT_72 => X"0000004b000000000000003a0000000000000037000000000000003900000000",
            INIT_73 => X"0000004500000000000000440000000000000048000000000000004c00000000",
            INIT_74 => X"00000049000000000000004b000000000000004a000000000000004b00000000",
            INIT_75 => X"000000350000000000000037000000000000003a000000000000004600000000",
            INIT_76 => X"0000007f000000000000006b0000000000000045000000000000003300000000",
            INIT_77 => X"000000330000000000000036000000000000003a000000000000005b00000000",
            INIT_78 => X"0000002e00000000000000330000000000000033000000000000004000000000",
            INIT_79 => X"0000003500000000000000390000000000000038000000000000003300000000",
            INIT_7A => X"0000003e00000000000000320000000000000033000000000000003400000000",
            INIT_7B => X"00000039000000000000003c000000000000003e000000000000004000000000",
            INIT_7C => X"000000400000000000000040000000000000003e000000000000003c00000000",
            INIT_7D => X"0000003700000000000000340000000000000035000000000000004000000000",
            INIT_7E => X"0000004800000000000000690000000000000067000000000000004600000000",
            INIT_7F => X"0000003200000000000000340000000000000032000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "sampleifmap_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e00000000000000300000000000000046000000000000004100000000",
            INIT_01 => X"0000002d000000000000002c0000000000000028000000000000001700000000",
            INIT_02 => X"0000000f000000000000000a0000000000000028000000000000002d00000000",
            INIT_03 => X"0000003000000000000000330000000000000035000000000000002c00000000",
            INIT_04 => X"0000005b000000000000005d000000000000005a000000000000004100000000",
            INIT_05 => X"00000037000000000000003c0000000000000051000000000000005f00000000",
            INIT_06 => X"000000440000000000000029000000000000006f000000000000007000000000",
            INIT_07 => X"0000004300000000000000360000000000000033000000000000004d00000000",
            INIT_08 => X"0000001e000000000000003c000000000000004f000000000000004500000000",
            INIT_09 => X"0000003100000000000000310000000000000041000000000000002900000000",
            INIT_0A => X"0000001900000000000000070000000000000023000000000000003100000000",
            INIT_0B => X"0000003100000000000000370000000000000045000000000000004100000000",
            INIT_0C => X"0000005000000000000000530000000000000055000000000000004d00000000",
            INIT_0D => X"0000003b00000000000000370000000000000051000000000000005700000000",
            INIT_0E => X"0000002f000000000000001f0000000000000079000000000000008300000000",
            INIT_0F => X"0000003d00000000000000410000000000000036000000000000003800000000",
            INIT_10 => X"0000002900000000000000480000000000000054000000000000004900000000",
            INIT_11 => X"000000360000000000000032000000000000004a000000000000004000000000",
            INIT_12 => X"00000024000000000000000b0000000000000020000000000000003600000000",
            INIT_13 => X"00000027000000000000002f0000000000000043000000000000003c00000000",
            INIT_14 => X"0000003e000000000000003b000000000000004d000000000000004b00000000",
            INIT_15 => X"0000003f00000000000000300000000000000055000000000000005300000000",
            INIT_16 => X"0000002900000000000000170000000000000080000000000000008b00000000",
            INIT_17 => X"000000300000000000000049000000000000004e000000000000004600000000",
            INIT_18 => X"000000360000000000000050000000000000004b000000000000005800000000",
            INIT_19 => X"0000003f00000000000000370000000000000044000000000000005000000000",
            INIT_1A => X"000000250000000000000011000000000000001c000000000000003a00000000",
            INIT_1B => X"0000002700000000000000280000000000000033000000000000002b00000000",
            INIT_1C => X"00000046000000000000004b0000000000000062000000000000005500000000",
            INIT_1D => X"0000004400000000000000320000000000000054000000000000005600000000",
            INIT_1E => X"0000004b000000000000002f0000000000000089000000000000008e00000000",
            INIT_1F => X"000000260000000000000041000000000000005d000000000000006400000000",
            INIT_20 => X"00000042000000000000006f0000000000000059000000000000005f00000000",
            INIT_21 => X"00000044000000000000003d000000000000003d000000000000005100000000",
            INIT_22 => X"00000016000000000000000f0000000000000016000000000000003e00000000",
            INIT_23 => X"0000003f00000000000000330000000000000023000000000000001f00000000",
            INIT_24 => X"000000470000000000000048000000000000004b000000000000004800000000",
            INIT_25 => X"0000004e00000000000000330000000000000053000000000000004d00000000",
            INIT_26 => X"000000570000000000000057000000000000009c000000000000009500000000",
            INIT_27 => X"00000058000000000000004b000000000000005f000000000000006300000000",
            INIT_28 => X"0000004d00000000000000520000000000000053000000000000005200000000",
            INIT_29 => X"000000390000000000000040000000000000003a000000000000004700000000",
            INIT_2A => X"0000001c00000000000000110000000000000014000000000000003b00000000",
            INIT_2B => X"000000470000000000000047000000000000003d000000000000003200000000",
            INIT_2C => X"0000003800000000000000440000000000000043000000000000004500000000",
            INIT_2D => X"0000004e00000000000000460000000000000053000000000000002900000000",
            INIT_2E => X"00000059000000000000006200000000000000ac000000000000009c00000000",
            INIT_2F => X"000000630000000000000070000000000000006f000000000000005e00000000",
            INIT_30 => X"0000003b00000000000000200000000000000040000000000000004500000000",
            INIT_31 => X"000000310000000000000049000000000000004a000000000000004800000000",
            INIT_32 => X"0000003e000000000000001d0000000000000012000000000000003100000000",
            INIT_33 => X"0000003f00000000000000560000000000000055000000000000005200000000",
            INIT_34 => X"0000002b000000000000005f0000000000000034000000000000002200000000",
            INIT_35 => X"0000004e0000000000000055000000000000005e000000000000001900000000",
            INIT_36 => X"0000006b000000000000006d00000000000000b400000000000000a600000000",
            INIT_37 => X"0000002f00000000000000560000000000000083000000000000006c00000000",
            INIT_38 => X"0000004600000000000000190000000000000035000000000000003b00000000",
            INIT_39 => X"0000003d0000000000000050000000000000004e000000000000005100000000",
            INIT_3A => X"0000005e0000000000000035000000000000000a000000000000002800000000",
            INIT_3B => X"00000019000000000000004b0000000000000058000000000000005700000000",
            INIT_3C => X"00000039000000000000005c000000000000002d000000000000000d00000000",
            INIT_3D => X"0000006200000000000000590000000000000065000000000000003200000000",
            INIT_3E => X"0000007c000000000000007800000000000000b3000000000000009000000000",
            INIT_3F => X"0000001800000000000000340000000000000080000000000000007c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000660000000000000031000000000000002f000000000000004400000000",
            INIT_41 => X"0000004f000000000000003f0000000000000059000000000000007700000000",
            INIT_42 => X"0000006000000000000000510000000000000022000000000000004200000000",
            INIT_43 => X"0000000e0000000000000029000000000000005a000000000000005900000000",
            INIT_44 => X"000000470000000000000043000000000000005c000000000000003400000000",
            INIT_45 => X"00000073000000000000006e0000000000000071000000000000006f00000000",
            INIT_46 => X"0000007f0000000000000079000000000000009c000000000000008800000000",
            INIT_47 => X"00000016000000000000001f0000000000000073000000000000007c00000000",
            INIT_48 => X"0000007200000000000000370000000000000035000000000000004d00000000",
            INIT_49 => X"000000370000000000000041000000000000007b000000000000008000000000",
            INIT_4A => X"0000006e000000000000006f0000000000000052000000000000004f00000000",
            INIT_4B => X"0000002500000000000000140000000000000045000000000000006a00000000",
            INIT_4C => X"0000006100000000000000530000000000000069000000000000005c00000000",
            INIT_4D => X"0000005c00000000000000730000000000000078000000000000007600000000",
            INIT_4E => X"0000007f000000000000007d0000000000000093000000000000009000000000",
            INIT_4F => X"00000017000000000000000e000000000000005f000000000000007700000000",
            INIT_50 => X"000000700000000000000036000000000000003a000000000000005500000000",
            INIT_51 => X"0000003100000000000000640000000000000084000000000000008100000000",
            INIT_52 => X"0000006d00000000000000680000000000000054000000000000002700000000",
            INIT_53 => X"00000053000000000000003f000000000000005d000000000000007d00000000",
            INIT_54 => X"0000006e0000000000000068000000000000005e000000000000006100000000",
            INIT_55 => X"000000390000000000000055000000000000007f000000000000006d00000000",
            INIT_56 => X"0000007c000000000000007b0000000000000096000000000000009800000000",
            INIT_57 => X"00000015000000000000000c000000000000005d000000000000007200000000",
            INIT_58 => X"0000006b00000000000000320000000000000035000000000000006c00000000",
            INIT_59 => X"0000004b00000000000000800000000000000083000000000000007e00000000",
            INIT_5A => X"0000006b0000000000000055000000000000005b000000000000003300000000",
            INIT_5B => X"000000930000000000000081000000000000006e000000000000008a00000000",
            INIT_5C => X"0000007700000000000000710000000000000078000000000000008400000000",
            INIT_5D => X"0000005d000000000000005a0000000000000073000000000000007500000000",
            INIT_5E => X"0000007d0000000000000071000000000000008d00000000000000a000000000",
            INIT_5F => X"00000009000000000000000e0000000000000065000000000000007900000000",
            INIT_60 => X"0000005c000000000000002b000000000000002a000000000000006000000000",
            INIT_61 => X"0000007700000000000000820000000000000080000000000000006a00000000",
            INIT_62 => X"000000890000000000000072000000000000007b000000000000007800000000",
            INIT_63 => X"000000840000000000000069000000000000006e000000000000009400000000",
            INIT_64 => X"0000008600000000000000800000000000000087000000000000009200000000",
            INIT_65 => X"00000077000000000000007e0000000000000078000000000000008c00000000",
            INIT_66 => X"0000006a00000000000000630000000000000091000000000000009800000000",
            INIT_67 => X"0000002800000000000000120000000000000063000000000000008200000000",
            INIT_68 => X"00000059000000000000003b0000000000000042000000000000006100000000",
            INIT_69 => X"000000880000000000000085000000000000006f000000000000006400000000",
            INIT_6A => X"000000910000000000000096000000000000008c000000000000009300000000",
            INIT_6B => X"0000007f00000000000000830000000000000088000000000000008e00000000",
            INIT_6C => X"000000930000000000000088000000000000007b000000000000007d00000000",
            INIT_6D => X"00000088000000000000009c000000000000008e000000000000009700000000",
            INIT_6E => X"00000070000000000000006d0000000000000090000000000000009200000000",
            INIT_6F => X"000000530000000000000032000000000000005c000000000000008200000000",
            INIT_70 => X"0000005f000000000000004b0000000000000048000000000000006900000000",
            INIT_71 => X"000000850000000000000085000000000000005e000000000000006800000000",
            INIT_72 => X"0000008500000000000000800000000000000087000000000000008f00000000",
            INIT_73 => X"0000009800000000000000a00000000000000096000000000000009300000000",
            INIT_74 => X"0000008700000000000000840000000000000090000000000000009100000000",
            INIT_75 => X"000000a500000000000000a2000000000000008a000000000000008a00000000",
            INIT_76 => X"00000077000000000000007e000000000000007f00000000000000a300000000",
            INIT_77 => X"0000004d000000000000003b000000000000005f000000000000007600000000",
            INIT_78 => X"0000005b00000000000000440000000000000044000000000000005e00000000",
            INIT_79 => X"00000083000000000000007b0000000000000062000000000000006500000000",
            INIT_7A => X"0000004f000000000000008a00000000000000c1000000000000009300000000",
            INIT_7B => X"000000a200000000000000930000000000000093000000000000007c00000000",
            INIT_7C => X"00000090000000000000009800000000000000ab00000000000000b400000000",
            INIT_7D => X"000000b300000000000000940000000000000079000000000000009000000000",
            INIT_7E => X"0000007b000000000000008000000000000000a000000000000000b400000000",
            INIT_7F => X"00000054000000000000001a000000000000003f000000000000007000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "sampleifmap_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000004a000000000000004f000000000000005800000000",
            INIT_01 => X"0000008100000000000000780000000000000078000000000000006e00000000",
            INIT_02 => X"0000005700000000000000c000000000000000b8000000000000007800000000",
            INIT_03 => X"000000a600000000000000a4000000000000009c000000000000007200000000",
            INIT_04 => X"000000b600000000000000b700000000000000a1000000000000009a00000000",
            INIT_05 => X"0000008f000000000000009400000000000000ad00000000000000bb00000000",
            INIT_06 => X"0000007c000000000000008e00000000000000c300000000000000b500000000",
            INIT_07 => X"000000760000000000000029000000000000002c000000000000006b00000000",
            INIT_08 => X"0000006000000000000000670000000000000059000000000000005b00000000",
            INIT_09 => X"0000006a000000000000006f0000000000000064000000000000007400000000",
            INIT_0A => X"000000a800000000000000bb0000000000000080000000000000007200000000",
            INIT_0B => X"000000ac00000000000000ac0000000000000099000000000000008c00000000",
            INIT_0C => X"000000a3000000000000009d00000000000000a400000000000000a700000000",
            INIT_0D => X"0000009c00000000000000ab00000000000000a500000000000000a100000000",
            INIT_0E => X"0000007200000000000000a7000000000000009100000000000000a100000000",
            INIT_0F => X"0000005e000000000000002a000000000000004a000000000000006a00000000",
            INIT_10 => X"0000007a00000000000000780000000000000061000000000000006500000000",
            INIT_11 => X"0000005b000000000000005f000000000000004e000000000000007200000000",
            INIT_12 => X"000000cc0000000000000081000000000000006e000000000000007300000000",
            INIT_13 => X"0000009900000000000000a0000000000000008900000000000000a700000000",
            INIT_14 => X"000000b200000000000000aa00000000000000ba00000000000000b300000000",
            INIT_15 => X"000000a500000000000000a2000000000000009c00000000000000b300000000",
            INIT_16 => X"000000480000000000000068000000000000008c000000000000009c00000000",
            INIT_17 => X"0000007200000000000000460000000000000059000000000000005400000000",
            INIT_18 => X"00000060000000000000007a000000000000006b000000000000006e00000000",
            INIT_19 => X"000000640000000000000048000000000000004c000000000000005a00000000",
            INIT_1A => X"0000008c0000000000000057000000000000007f000000000000006d00000000",
            INIT_1B => X"000000b400000000000000a6000000000000009f00000000000000bd00000000",
            INIT_1C => X"000000bc00000000000000be00000000000000ad00000000000000ae00000000",
            INIT_1D => X"000000a100000000000000a2000000000000009900000000000000a200000000",
            INIT_1E => X"0000004a000000000000004b0000000000000095000000000000009900000000",
            INIT_1F => X"0000008a0000000000000070000000000000003e000000000000004200000000",
            INIT_20 => X"0000004e0000000000000059000000000000006a000000000000007700000000",
            INIT_21 => X"00000067000000000000003c0000000000000047000000000000005900000000",
            INIT_22 => X"000000420000000000000072000000000000005f000000000000004b00000000",
            INIT_23 => X"000000be00000000000000ae00000000000000b5000000000000007f00000000",
            INIT_24 => X"000000c100000000000000b800000000000000ab00000000000000ba00000000",
            INIT_25 => X"000000a500000000000000ab00000000000000a000000000000000a400000000",
            INIT_26 => X"0000005c0000000000000068000000000000008b000000000000009200000000",
            INIT_27 => X"000000730000000000000070000000000000005e000000000000004d00000000",
            INIT_28 => X"00000067000000000000003a000000000000005e000000000000007e00000000",
            INIT_29 => X"0000005f0000000000000048000000000000004c000000000000006a00000000",
            INIT_2A => X"0000006300000000000000780000000000000041000000000000005e00000000",
            INIT_2B => X"000000bc00000000000000c400000000000000a1000000000000005b00000000",
            INIT_2C => X"000000a700000000000000a700000000000000c100000000000000b600000000",
            INIT_2D => X"000000a1000000000000009a00000000000000a000000000000000aa00000000",
            INIT_2E => X"00000051000000000000006e000000000000008a000000000000009100000000",
            INIT_2F => X"00000064000000000000006d0000000000000088000000000000006900000000",
            INIT_30 => X"0000006800000000000000460000000000000052000000000000006f00000000",
            INIT_31 => X"000000540000000000000045000000000000005e000000000000007100000000",
            INIT_32 => X"0000007d0000000000000055000000000000006d000000000000007400000000",
            INIT_33 => X"000000c800000000000000ba000000000000009b000000000000007f00000000",
            INIT_34 => X"0000009d00000000000000b100000000000000bb00000000000000bb00000000",
            INIT_35 => X"000000a600000000000000a400000000000000a2000000000000009400000000",
            INIT_36 => X"000000610000000000000079000000000000009500000000000000a200000000",
            INIT_37 => X"0000006100000000000000610000000000000073000000000000007800000000",
            INIT_38 => X"000000b4000000000000008c000000000000005c000000000000006500000000",
            INIT_39 => X"0000004c0000000000000055000000000000007b000000000000009700000000",
            INIT_3A => X"00000054000000000000005a000000000000007c000000000000006700000000",
            INIT_3B => X"000000c800000000000000ad00000000000000af000000000000009200000000",
            INIT_3C => X"0000009f00000000000000ad00000000000000ad00000000000000bc00000000",
            INIT_3D => X"000000ad00000000000000a300000000000000ac000000000000009f00000000",
            INIT_3E => X"000000830000000000000083000000000000008b00000000000000a400000000",
            INIT_3F => X"000000600000000000000064000000000000005f000000000000007000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000c00000000000000090000000000000007700000000",
            INIT_41 => X"0000006c000000000000007f000000000000009d00000000000000c200000000",
            INIT_42 => X"0000006f000000000000006a000000000000005e000000000000006a00000000",
            INIT_43 => X"000000c500000000000000b000000000000000af000000000000007c00000000",
            INIT_44 => X"000000a500000000000000b000000000000000aa00000000000000b800000000",
            INIT_45 => X"000000a300000000000000af00000000000000c5000000000000009c00000000",
            INIT_46 => X"00000065000000000000007a0000000000000083000000000000009300000000",
            INIT_47 => X"00000066000000000000006b0000000000000060000000000000006400000000",
            INIT_48 => X"000000a9000000000000008a0000000000000074000000000000006e00000000",
            INIT_49 => X"0000008800000000000000a000000000000000c400000000000000c500000000",
            INIT_4A => X"0000008a000000000000005c0000000000000063000000000000008100000000",
            INIT_4B => X"000000a900000000000000b4000000000000009f000000000000009200000000",
            INIT_4C => X"000000b200000000000000af000000000000008d000000000000008e00000000",
            INIT_4D => X"0000009700000000000000b300000000000000bc00000000000000a600000000",
            INIT_4E => X"0000003a0000000000000070000000000000009a000000000000008f00000000",
            INIT_4F => X"0000004900000000000000660000000000000065000000000000005b00000000",
            INIT_50 => X"0000006b000000000000004a0000000000000057000000000000005b00000000",
            INIT_51 => X"000000a300000000000000bf00000000000000b900000000000000a500000000",
            INIT_52 => X"00000066000000000000006a0000000000000080000000000000008600000000",
            INIT_53 => X"0000007400000000000000920000000000000084000000000000007600000000",
            INIT_54 => X"000000b600000000000000a10000000000000063000000000000004d00000000",
            INIT_55 => X"000000a700000000000000ad000000000000009f00000000000000b700000000",
            INIT_56 => X"0000002b000000000000005e0000000000000087000000000000009c00000000",
            INIT_57 => X"0000004d0000000000000044000000000000005c000000000000005b00000000",
            INIT_58 => X"0000002c0000000000000032000000000000005f000000000000005100000000",
            INIT_59 => X"000000bb00000000000000a60000000000000094000000000000005f00000000",
            INIT_5A => X"00000072000000000000007e000000000000009000000000000000ae00000000",
            INIT_5B => X"0000006b00000000000000770000000000000072000000000000006800000000",
            INIT_5C => X"000000b6000000000000009d0000000000000052000000000000005100000000",
            INIT_5D => X"0000009600000000000000a900000000000000b200000000000000a900000000",
            INIT_5E => X"0000003f000000000000002c000000000000006c000000000000009800000000",
            INIT_5F => X"0000005600000000000000500000000000000045000000000000006100000000",
            INIT_60 => X"000000150000000000000034000000000000005f000000000000005a00000000",
            INIT_61 => X"000000b00000000000000092000000000000006d000000000000001c00000000",
            INIT_62 => X"0000007f000000000000008e00000000000000b500000000000000ca00000000",
            INIT_63 => X"0000008200000000000000720000000000000077000000000000007800000000",
            INIT_64 => X"000000a900000000000000900000000000000076000000000000008100000000",
            INIT_65 => X"0000009800000000000000b400000000000000ad000000000000009f00000000",
            INIT_66 => X"00000055000000000000002c0000000000000044000000000000007700000000",
            INIT_67 => X"0000006a00000000000000a70000000000000072000000000000003300000000",
            INIT_68 => X"000000340000000000000039000000000000005b000000000000005f00000000",
            INIT_69 => X"0000009c00000000000000770000000000000031000000000000001800000000",
            INIT_6A => X"0000009b00000000000000ba00000000000000cb00000000000000bb00000000",
            INIT_6B => X"0000007500000000000000740000000000000085000000000000008d00000000",
            INIT_6C => X"00000099000000000000008b0000000000000077000000000000006d00000000",
            INIT_6D => X"0000007d000000000000009c00000000000000a7000000000000009f00000000",
            INIT_6E => X"0000004000000000000000440000000000000041000000000000006500000000",
            INIT_6F => X"0000007a00000000000000aa0000000000000090000000000000003700000000",
            INIT_70 => X"000000490000000000000020000000000000004b000000000000005e00000000",
            INIT_71 => X"0000007300000000000000360000000000000021000000000000002e00000000",
            INIT_72 => X"000000c200000000000000c300000000000000b0000000000000009600000000",
            INIT_73 => X"000000920000000000000088000000000000009b00000000000000b100000000",
            INIT_74 => X"00000077000000000000005e0000000000000065000000000000008b00000000",
            INIT_75 => X"000000690000000000000060000000000000005f000000000000006500000000",
            INIT_76 => X"0000006d000000000000006b0000000000000076000000000000008300000000",
            INIT_77 => X"0000006a000000000000009a000000000000008f000000000000008000000000",
            INIT_78 => X"0000004c00000000000000180000000000000023000000000000004e00000000",
            INIT_79 => X"0000003b000000000000001b0000000000000028000000000000004100000000",
            INIT_7A => X"000000b000000000000000960000000000000088000000000000007800000000",
            INIT_7B => X"000000ba00000000000000a500000000000000b700000000000000c000000000",
            INIT_7C => X"00000056000000000000006b00000000000000aa00000000000000cf00000000",
            INIT_7D => X"0000008c00000000000000700000000000000055000000000000004200000000",
            INIT_7E => X"000000890000000000000089000000000000009500000000000000a900000000",
            INIT_7F => X"00000080000000000000009a000000000000008f000000000000009600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "sampleifmap_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002e00000000000000400000000000000051000000000000004400000000",
            INIT_01 => X"00000050000000000000004b0000000000000039000000000000002100000000",
            INIT_02 => X"0000002200000000000000140000000000000046000000000000005300000000",
            INIT_03 => X"000000420000000000000046000000000000004b000000000000004700000000",
            INIT_04 => X"00000079000000000000007c0000000000000078000000000000005700000000",
            INIT_05 => X"000000520000000000000054000000000000006c000000000000007e00000000",
            INIT_06 => X"0000005b000000000000003b0000000000000081000000000000008800000000",
            INIT_07 => X"00000057000000000000004c0000000000000043000000000000006000000000",
            INIT_08 => X"0000002f000000000000004a0000000000000066000000000000005000000000",
            INIT_09 => X"000000540000000000000054000000000000005c000000000000003800000000",
            INIT_0A => X"000000300000000000000012000000000000003e000000000000005800000000",
            INIT_0B => X"00000049000000000000004d000000000000005c000000000000005d00000000",
            INIT_0C => X"0000006a000000000000006f0000000000000075000000000000006b00000000",
            INIT_0D => X"00000053000000000000004d000000000000006c000000000000007500000000",
            INIT_0E => X"00000041000000000000002d000000000000008b000000000000009700000000",
            INIT_0F => X"00000051000000000000005a0000000000000042000000000000004700000000",
            INIT_10 => X"000000380000000000000058000000000000006d000000000000005f00000000",
            INIT_11 => X"0000005a00000000000000560000000000000069000000000000005400000000",
            INIT_12 => X"0000003c00000000000000140000000000000035000000000000005c00000000",
            INIT_13 => X"0000003c00000000000000420000000000000058000000000000005900000000",
            INIT_14 => X"00000054000000000000004e0000000000000066000000000000006700000000",
            INIT_15 => X"0000005600000000000000420000000000000072000000000000007200000000",
            INIT_16 => X"000000370000000000000023000000000000008f000000000000009e00000000",
            INIT_17 => X"0000003b00000000000000620000000000000062000000000000005400000000",
            INIT_18 => X"0000004900000000000000640000000000000064000000000000007400000000",
            INIT_19 => X"0000006000000000000000580000000000000066000000000000006d00000000",
            INIT_1A => X"00000038000000000000001a000000000000002d000000000000005e00000000",
            INIT_1B => X"0000003700000000000000360000000000000043000000000000004100000000",
            INIT_1C => X"0000006200000000000000610000000000000075000000000000006a00000000",
            INIT_1D => X"0000005b00000000000000450000000000000072000000000000007600000000",
            INIT_1E => X"0000005d0000000000000040000000000000009600000000000000a000000000",
            INIT_1F => X"00000032000000000000005e000000000000007e000000000000007800000000",
            INIT_20 => X"0000005d00000000000000800000000000000068000000000000007800000000",
            INIT_21 => X"0000005e000000000000005a000000000000005e000000000000007200000000",
            INIT_22 => X"00000024000000000000001a0000000000000027000000000000005d00000000",
            INIT_23 => X"0000005600000000000000490000000000000037000000000000002f00000000",
            INIT_24 => X"00000065000000000000006b0000000000000071000000000000006900000000",
            INIT_25 => X"00000067000000000000004a000000000000006d000000000000006700000000",
            INIT_26 => X"00000074000000000000007000000000000000ac00000000000000a200000000",
            INIT_27 => X"0000006c00000000000000670000000000000084000000000000008100000000",
            INIT_28 => X"0000006200000000000000620000000000000066000000000000006900000000",
            INIT_29 => X"0000004e000000000000005b0000000000000059000000000000005f00000000",
            INIT_2A => X"0000002b000000000000001b0000000000000023000000000000005800000000",
            INIT_2B => X"0000006c000000000000006a000000000000005d000000000000004d00000000",
            INIT_2C => X"0000004e00000000000000640000000000000065000000000000006700000000",
            INIT_2D => X"000000660000000000000062000000000000006e000000000000003900000000",
            INIT_2E => X"0000007f000000000000008200000000000000ba00000000000000a700000000",
            INIT_2F => X"0000007800000000000000840000000000000090000000000000008100000000",
            INIT_30 => X"0000004f00000000000000300000000000000060000000000000005e00000000",
            INIT_31 => X"0000003f000000000000005d0000000000000064000000000000005a00000000",
            INIT_32 => X"0000005a0000000000000026000000000000001d000000000000004a00000000",
            INIT_33 => X"0000006300000000000000820000000000000081000000000000007e00000000",
            INIT_34 => X"0000003900000000000000730000000000000047000000000000003a00000000",
            INIT_35 => X"0000006a0000000000000071000000000000007b000000000000002500000000",
            INIT_36 => X"0000008c000000000000008d00000000000000c100000000000000b700000000",
            INIT_37 => X"0000003b000000000000006500000000000000a0000000000000008900000000",
            INIT_38 => X"00000069000000000000002f0000000000000054000000000000005600000000",
            INIT_39 => X"00000047000000000000005e0000000000000061000000000000006700000000",
            INIT_3A => X"0000008b00000000000000490000000000000014000000000000003800000000",
            INIT_3B => X"000000290000000000000072000000000000008c000000000000008a00000000",
            INIT_3C => X"0000004f00000000000000730000000000000041000000000000001a00000000",
            INIT_3D => X"0000008c0000000000000078000000000000007d000000000000003b00000000",
            INIT_3E => X"00000094000000000000009600000000000000c300000000000000b000000000",
            INIT_3F => X"00000018000000000000003f000000000000009b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008c000000000000004a000000000000004e000000000000006200000000",
            INIT_41 => X"0000005c00000000000000500000000000000072000000000000009500000000",
            INIT_42 => X"000000900000000000000071000000000000002c000000000000004700000000",
            INIT_43 => X"00000017000000000000003f0000000000000086000000000000008800000000",
            INIT_44 => X"00000056000000000000005e000000000000007c000000000000004500000000",
            INIT_45 => X"000000a5000000000000009b000000000000008b000000000000007000000000",
            INIT_46 => X"00000096000000000000009600000000000000b100000000000000aa00000000",
            INIT_47 => X"000000160000000000000029000000000000008e000000000000009200000000",
            INIT_48 => X"00000094000000000000004e0000000000000051000000000000007400000000",
            INIT_49 => X"000000450000000000000054000000000000009b00000000000000a300000000",
            INIT_4A => X"0000008e0000000000000089000000000000005a000000000000005100000000",
            INIT_4B => X"000000380000000000000021000000000000005d000000000000008a00000000",
            INIT_4C => X"000000800000000000000073000000000000008f000000000000007c00000000",
            INIT_4D => X"00000081000000000000009c000000000000009c000000000000009700000000",
            INIT_4E => X"0000009a000000000000009800000000000000ad00000000000000a700000000",
            INIT_4F => X"0000001800000000000000160000000000000079000000000000009400000000",
            INIT_50 => X"000000910000000000000049000000000000004f000000000000007800000000",
            INIT_51 => X"00000041000000000000007f00000000000000a600000000000000a500000000",
            INIT_52 => X"0000007f000000000000008e0000000000000072000000000000003600000000",
            INIT_53 => X"0000006c0000000000000047000000000000005d000000000000007e00000000",
            INIT_54 => X"000000a100000000000000920000000000000085000000000000008700000000",
            INIT_55 => X"00000057000000000000007500000000000000a5000000000000009c00000000",
            INIT_56 => X"0000009c000000000000009700000000000000af00000000000000a900000000",
            INIT_57 => X"0000001700000000000000130000000000000074000000000000009100000000",
            INIT_58 => X"0000008a00000000000000420000000000000045000000000000007b00000000",
            INIT_59 => X"0000005f00000000000000a500000000000000a800000000000000a100000000",
            INIT_5A => X"00000070000000000000008a000000000000008c000000000000004b00000000",
            INIT_5B => X"000000a200000000000000880000000000000066000000000000006d00000000",
            INIT_5C => X"000000870000000000000097000000000000009a000000000000009900000000",
            INIT_5D => X"0000008800000000000000760000000000000085000000000000007c00000000",
            INIT_5E => X"0000009d000000000000009200000000000000aa00000000000000bd00000000",
            INIT_5F => X"0000000b00000000000000140000000000000077000000000000009400000000",
            INIT_60 => X"00000079000000000000003c0000000000000039000000000000006a00000000",
            INIT_61 => X"0000009800000000000000ad00000000000000a4000000000000008700000000",
            INIT_62 => X"00000076000000000000007f0000000000000093000000000000009000000000",
            INIT_63 => X"0000008b0000000000000066000000000000005c000000000000007300000000",
            INIT_64 => X"000000740000000000000085000000000000008a000000000000008d00000000",
            INIT_65 => X"000000880000000000000077000000000000006b000000000000007800000000",
            INIT_66 => X"00000091000000000000008700000000000000ae00000000000000b000000000",
            INIT_67 => X"0000002b000000000000001a000000000000007200000000000000a100000000",
            INIT_68 => X"00000074000000000000004e0000000000000055000000000000007400000000",
            INIT_69 => X"000000ab00000000000000ac000000000000008c000000000000007f00000000",
            INIT_6A => X"000000780000000000000082000000000000007c000000000000009900000000",
            INIT_6B => X"0000006e00000000000000710000000000000076000000000000007700000000",
            INIT_6C => X"0000007d0000000000000077000000000000006c000000000000006900000000",
            INIT_6D => X"000000750000000000000081000000000000007a000000000000008300000000",
            INIT_6E => X"0000009a000000000000008d00000000000000a2000000000000009000000000",
            INIT_6F => X"0000005f0000000000000041000000000000007000000000000000a600000000",
            INIT_70 => X"0000007800000000000000630000000000000060000000000000008400000000",
            INIT_71 => X"000000a800000000000000a50000000000000072000000000000008200000000",
            INIT_72 => X"000000700000000000000068000000000000006b000000000000008b00000000",
            INIT_73 => X"00000084000000000000008e0000000000000081000000000000007c00000000",
            INIT_74 => X"0000006f000000000000006b0000000000000077000000000000007a00000000",
            INIT_75 => X"00000090000000000000008d0000000000000076000000000000007300000000",
            INIT_76 => X"0000009f0000000000000092000000000000007b000000000000008e00000000",
            INIT_77 => X"0000005e00000000000000480000000000000070000000000000009d00000000",
            INIT_78 => X"00000076000000000000005d000000000000005a000000000000007900000000",
            INIT_79 => X"000000a60000000000000097000000000000007c000000000000007f00000000",
            INIT_7A => X"00000045000000000000007900000000000000ab000000000000009900000000",
            INIT_7B => X"0000008b000000000000007b000000000000007c000000000000006b00000000",
            INIT_7C => X"0000007700000000000000800000000000000090000000000000009b00000000",
            INIT_7D => X"000000a700000000000000830000000000000067000000000000007a00000000",
            INIT_7E => X"000000a00000000000000080000000000000008c000000000000009f00000000",
            INIT_7F => X"000000680000000000000022000000000000004b000000000000009500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "sampleifmap_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000007e00000000000000640000000000000064000000000000007000000000",
            INIT_01 => X"000000a300000000000000950000000000000098000000000000008d00000000",
            INIT_02 => X"0000004700000000000000a600000000000000a3000000000000008a00000000",
            INIT_03 => X"0000008d000000000000008b0000000000000085000000000000006400000000",
            INIT_04 => X"0000009e00000000000000a00000000000000088000000000000008100000000",
            INIT_05 => X"0000007e000000000000007d000000000000009700000000000000a300000000",
            INIT_06 => X"0000008f000000000000007a00000000000000b100000000000000a900000000",
            INIT_07 => X"0000008b0000000000000033000000000000003d000000000000008f00000000",
            INIT_08 => X"0000008100000000000000830000000000000070000000000000007000000000",
            INIT_09 => X"000000890000000000000090000000000000007c000000000000009300000000",
            INIT_0A => X"0000009900000000000000a80000000000000079000000000000008f00000000",
            INIT_0B => X"000000930000000000000092000000000000007f000000000000007a00000000",
            INIT_0C => X"0000008a0000000000000084000000000000008b000000000000008d00000000",
            INIT_0D => X"000000860000000000000099000000000000008f000000000000008600000000",
            INIT_0E => X"0000007a00000000000000920000000000000082000000000000009100000000",
            INIT_0F => X"0000006f000000000000003a0000000000000064000000000000008600000000",
            INIT_10 => X"0000008e00000000000000950000000000000076000000000000007900000000",
            INIT_11 => X"00000076000000000000007b0000000000000061000000000000008d00000000",
            INIT_12 => X"000000bb0000000000000079000000000000007e000000000000008f00000000",
            INIT_13 => X"000000820000000000000088000000000000006e000000000000009100000000",
            INIT_14 => X"0000009a000000000000009400000000000000a1000000000000009a00000000",
            INIT_15 => X"0000009100000000000000960000000000000086000000000000009700000000",
            INIT_16 => X"000000570000000000000061000000000000007b000000000000008600000000",
            INIT_17 => X"0000008600000000000000610000000000000077000000000000006700000000",
            INIT_18 => X"0000006f00000000000000970000000000000087000000000000008800000000",
            INIT_19 => X"0000007d000000000000005d0000000000000065000000000000007a00000000",
            INIT_1A => X"0000007d00000000000000600000000000000099000000000000008600000000",
            INIT_1B => X"000000a00000000000000092000000000000008800000000000000a900000000",
            INIT_1C => X"000000a700000000000000a60000000000000094000000000000009600000000",
            INIT_1D => X"0000009100000000000000900000000000000080000000000000008d00000000",
            INIT_1E => X"0000005e000000000000004b0000000000000082000000000000008400000000",
            INIT_1F => X"000000a900000000000000950000000000000057000000000000005300000000",
            INIT_20 => X"0000005e0000000000000070000000000000008c000000000000009400000000",
            INIT_21 => X"0000008200000000000000540000000000000068000000000000007900000000",
            INIT_22 => X"0000004a000000000000008d0000000000000074000000000000006600000000",
            INIT_23 => X"000000aa000000000000009b00000000000000a3000000000000007600000000",
            INIT_24 => X"000000a7000000000000009d000000000000009500000000000000a500000000",
            INIT_25 => X"0000009100000000000000930000000000000089000000000000009200000000",
            INIT_26 => X"00000071000000000000006d000000000000007c000000000000007f00000000",
            INIT_27 => X"000000a1000000000000009c0000000000000077000000000000006000000000",
            INIT_28 => X"0000007d00000000000000480000000000000077000000000000009800000000",
            INIT_29 => X"0000007900000000000000630000000000000065000000000000008100000000",
            INIT_2A => X"0000007d000000000000009a000000000000005b000000000000007800000000",
            INIT_2B => X"000000a900000000000000b50000000000000096000000000000005d00000000",
            INIT_2C => X"0000008f000000000000009100000000000000ad00000000000000a200000000",
            INIT_2D => X"0000008b00000000000000810000000000000087000000000000008f00000000",
            INIT_2E => X"0000006600000000000000750000000000000078000000000000007d00000000",
            INIT_2F => X"00000099000000000000009a00000000000000ab000000000000008100000000",
            INIT_30 => X"0000007b00000000000000520000000000000068000000000000008800000000",
            INIT_31 => X"0000007300000000000000620000000000000076000000000000008800000000",
            INIT_32 => X"000000940000000000000075000000000000008d000000000000009600000000",
            INIT_33 => X"000000b300000000000000ad0000000000000095000000000000008100000000",
            INIT_34 => X"0000008f000000000000009f00000000000000a800000000000000a500000000",
            INIT_35 => X"0000008d000000000000008c000000000000008b000000000000007e00000000",
            INIT_36 => X"0000006d000000000000007a0000000000000085000000000000008800000000",
            INIT_37 => X"00000095000000000000009600000000000000a4000000000000009800000000",
            INIT_38 => X"000000bf0000000000000096000000000000006f000000000000007d00000000",
            INIT_39 => X"0000006f0000000000000079000000000000009e00000000000000ac00000000",
            INIT_3A => X"0000006900000000000000730000000000000099000000000000009100000000",
            INIT_3B => X"000000ac000000000000009a00000000000000a1000000000000009400000000",
            INIT_3C => X"0000008d000000000000009c000000000000009b00000000000000a100000000",
            INIT_3D => X"0000008f00000000000000880000000000000093000000000000008900000000",
            INIT_3E => X"00000086000000000000007b000000000000008c000000000000008900000000",
            INIT_3F => X"00000095000000000000009e0000000000000095000000000000009c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000dc00000000000000c800000000000000a2000000000000009500000000",
            INIT_41 => X"0000009300000000000000aa00000000000000bd00000000000000d100000000",
            INIT_42 => X"00000088000000000000007d000000000000007a000000000000009100000000",
            INIT_43 => X"000000a40000000000000096000000000000009f000000000000008b00000000",
            INIT_44 => X"0000008e000000000000009f000000000000009b000000000000009b00000000",
            INIT_45 => X"00000088000000000000009300000000000000a9000000000000008500000000",
            INIT_46 => X"00000072000000000000006b000000000000007e000000000000007f00000000",
            INIT_47 => X"0000009c00000000000000a0000000000000008f000000000000009a00000000",
            INIT_48 => X"000000be000000000000009d0000000000000089000000000000008b00000000",
            INIT_49 => X"000000b000000000000000bf00000000000000d700000000000000d500000000",
            INIT_4A => X"000000a30000000000000075000000000000008400000000000000a900000000",
            INIT_4B => X"0000008f000000000000009a000000000000009700000000000000ad00000000",
            INIT_4C => X"0000009800000000000000990000000000000081000000000000007c00000000",
            INIT_4D => X"0000007c000000000000009500000000000000a3000000000000009100000000",
            INIT_4E => X"0000004a00000000000000600000000000000083000000000000007700000000",
            INIT_4F => X"0000007800000000000000970000000000000095000000000000009100000000",
            INIT_50 => X"000000860000000000000061000000000000006f000000000000007300000000",
            INIT_51 => X"000000c100000000000000d300000000000000cf00000000000000bf00000000",
            INIT_52 => X"0000007f000000000000009100000000000000ad00000000000000b100000000",
            INIT_53 => X"000000680000000000000086000000000000008f000000000000009000000000",
            INIT_54 => X"0000009b000000000000008b000000000000005c000000000000004900000000",
            INIT_55 => X"0000008e0000000000000094000000000000008a00000000000000a100000000",
            INIT_56 => X"0000003c00000000000000550000000000000075000000000000008300000000",
            INIT_57 => X"0000006d000000000000006f0000000000000091000000000000009200000000",
            INIT_58 => X"0000004000000000000000410000000000000072000000000000006a00000000",
            INIT_59 => X"000000d500000000000000c300000000000000b2000000000000007800000000",
            INIT_5A => X"0000009900000000000000ad00000000000000b900000000000000ca00000000",
            INIT_5B => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_5C => X"0000009a000000000000008e0000000000000060000000000000006c00000000",
            INIT_5D => X"0000007f000000000000009500000000000000a1000000000000009000000000",
            INIT_5E => X"0000006100000000000000310000000000000062000000000000008300000000",
            INIT_5F => X"000000750000000000000076000000000000006c000000000000009300000000",
            INIT_60 => X"00000026000000000000003e0000000000000070000000000000007400000000",
            INIT_61 => X"000000c700000000000000b40000000000000087000000000000002900000000",
            INIT_62 => X"000000b200000000000000b700000000000000cc00000000000000d400000000",
            INIT_63 => X"000000a1000000000000009e00000000000000a400000000000000ab00000000",
            INIT_64 => X"0000008d0000000000000087000000000000008b000000000000009d00000000",
            INIT_65 => X"0000007e000000000000009c0000000000000099000000000000008700000000",
            INIT_66 => X"0000007c000000000000003b0000000000000042000000000000006700000000",
            INIT_67 => X"0000008300000000000000c50000000000000088000000000000005400000000",
            INIT_68 => X"0000004e000000000000004f000000000000007b000000000000007f00000000",
            INIT_69 => X"000000bf00000000000000950000000000000042000000000000002500000000",
            INIT_6A => X"000000c200000000000000d600000000000000db00000000000000d000000000",
            INIT_6B => X"0000009f00000000000000a500000000000000b400000000000000b800000000",
            INIT_6C => X"00000083000000000000007b000000000000007d000000000000008700000000",
            INIT_6D => X"0000007200000000000000870000000000000093000000000000008a00000000",
            INIT_6E => X"0000005b0000000000000055000000000000004f000000000000006c00000000",
            INIT_6F => X"0000008f00000000000000c900000000000000ac000000000000004e00000000",
            INIT_70 => X"0000006b00000000000000340000000000000068000000000000007d00000000",
            INIT_71 => X"00000097000000000000004e0000000000000030000000000000004300000000",
            INIT_72 => X"000000da00000000000000d900000000000000cb00000000000000bd00000000",
            INIT_73 => X"000000b600000000000000b400000000000000c300000000000000cd00000000",
            INIT_74 => X"0000007a000000000000005e000000000000007400000000000000a500000000",
            INIT_75 => X"0000006f00000000000000590000000000000059000000000000006100000000",
            INIT_76 => X"000000860000000000000082000000000000008a000000000000009600000000",
            INIT_77 => X"0000008100000000000000bc00000000000000b5000000000000009f00000000",
            INIT_78 => X"0000007300000000000000280000000000000033000000000000006600000000",
            INIT_79 => X"0000004e0000000000000029000000000000003a000000000000006000000000",
            INIT_7A => X"000000cf00000000000000b900000000000000b500000000000000a000000000",
            INIT_7B => X"000000ce00000000000000c400000000000000d200000000000000da00000000",
            INIT_7C => X"00000071000000000000007c00000000000000b400000000000000d600000000",
            INIT_7D => X"000000a000000000000000840000000000000066000000000000005600000000",
            INIT_7E => X"000000a700000000000000a700000000000000a700000000000000ba00000000",
            INIT_7F => X"0000009c00000000000000b900000000000000b300000000000000b400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "sampleifmap_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000002e0000000000000040000000000000003200000000",
            INIT_01 => X"0000003900000000000000370000000000000024000000000000001600000000",
            INIT_02 => X"00000012000000000000000c0000000000000036000000000000003b00000000",
            INIT_03 => X"000000320000000000000031000000000000002c000000000000002b00000000",
            INIT_04 => X"0000004d0000000000000051000000000000004d000000000000003a00000000",
            INIT_05 => X"000000390000000000000038000000000000004e000000000000005300000000",
            INIT_06 => X"0000003a000000000000001f000000000000005d000000000000006100000000",
            INIT_07 => X"0000004200000000000000350000000000000029000000000000004100000000",
            INIT_08 => X"0000001d00000000000000390000000000000051000000000000003a00000000",
            INIT_09 => X"0000003c000000000000003b000000000000003d000000000000002300000000",
            INIT_0A => X"0000001b0000000000000007000000000000002f000000000000004000000000",
            INIT_0B => X"0000002f000000000000003b000000000000003e000000000000003800000000",
            INIT_0C => X"00000044000000000000004a000000000000004a000000000000004400000000",
            INIT_0D => X"0000003c00000000000000330000000000000051000000000000004e00000000",
            INIT_0E => X"0000002700000000000000150000000000000060000000000000006f00000000",
            INIT_0F => X"000000420000000000000045000000000000002c000000000000002d00000000",
            INIT_10 => X"0000002300000000000000460000000000000057000000000000004800000000",
            INIT_11 => X"00000041000000000000003c0000000000000048000000000000003500000000",
            INIT_12 => X"0000002300000000000000070000000000000026000000000000004500000000",
            INIT_13 => X"0000002100000000000000300000000000000041000000000000003400000000",
            INIT_14 => X"0000003700000000000000320000000000000042000000000000004300000000",
            INIT_15 => X"0000003e000000000000002d0000000000000052000000000000004d00000000",
            INIT_16 => X"0000002600000000000000100000000000000063000000000000007400000000",
            INIT_17 => X"00000033000000000000004d000000000000004b000000000000003f00000000",
            INIT_18 => X"0000002f0000000000000050000000000000004c000000000000005e00000000",
            INIT_19 => X"0000004a00000000000000410000000000000048000000000000004700000000",
            INIT_1A => X"00000022000000000000000c000000000000001e000000000000004800000000",
            INIT_1B => X"0000001e00000000000000230000000000000034000000000000002800000000",
            INIT_1C => X"0000004500000000000000440000000000000057000000000000004b00000000",
            INIT_1D => X"00000043000000000000002e000000000000004d000000000000005100000000",
            INIT_1E => X"00000049000000000000002a000000000000006b000000000000007700000000",
            INIT_1F => X"0000002200000000000000440000000000000060000000000000005f00000000",
            INIT_20 => X"0000003c000000000000006a000000000000004f000000000000006100000000",
            INIT_21 => X"0000004c00000000000000480000000000000044000000000000004b00000000",
            INIT_22 => X"00000011000000000000000c0000000000000018000000000000004900000000",
            INIT_23 => X"0000003b00000000000000330000000000000025000000000000001c00000000",
            INIT_24 => X"00000047000000000000004b000000000000004f000000000000004800000000",
            INIT_25 => X"0000004d000000000000002d0000000000000049000000000000004700000000",
            INIT_26 => X"0000005500000000000000520000000000000081000000000000008000000000",
            INIT_27 => X"0000005000000000000000490000000000000061000000000000005e00000000",
            INIT_28 => X"00000043000000000000004b000000000000004d000000000000005200000000",
            INIT_29 => X"0000003d000000000000004d0000000000000045000000000000003d00000000",
            INIT_2A => X"00000016000000000000000d0000000000000013000000000000004300000000",
            INIT_2B => X"000000490000000000000047000000000000003b000000000000002c00000000",
            INIT_2C => X"0000003500000000000000490000000000000048000000000000004800000000",
            INIT_2D => X"0000004d000000000000003e0000000000000049000000000000002200000000",
            INIT_2E => X"0000005b00000000000000600000000000000093000000000000008800000000",
            INIT_2F => X"0000005c0000000000000068000000000000006e000000000000005c00000000",
            INIT_30 => X"0000003300000000000000190000000000000046000000000000004800000000",
            INIT_31 => X"00000032000000000000004f000000000000004f000000000000003e00000000",
            INIT_32 => X"000000360000000000000018000000000000000f000000000000003800000000",
            INIT_33 => X"0000003e000000000000004d000000000000004b000000000000004900000000",
            INIT_34 => X"0000002a00000000000000600000000000000033000000000000002200000000",
            INIT_35 => X"0000004a00000000000000480000000000000058000000000000001600000000",
            INIT_36 => X"0000006c000000000000006800000000000000a1000000000000009500000000",
            INIT_37 => X"0000002b00000000000000510000000000000083000000000000006b00000000",
            INIT_38 => X"000000460000000000000015000000000000003b000000000000003f00000000",
            INIT_39 => X"0000003a000000000000004b0000000000000048000000000000004d00000000",
            INIT_3A => X"00000051000000000000002f0000000000000008000000000000002900000000",
            INIT_3B => X"00000012000000000000003e000000000000004b000000000000004b00000000",
            INIT_3C => X"0000004000000000000000590000000000000027000000000000000600000000",
            INIT_3D => X"000000530000000000000048000000000000005e000000000000002a00000000",
            INIT_3E => X"00000078000000000000007200000000000000a2000000000000008300000000",
            INIT_3F => X"0000001500000000000000340000000000000085000000000000007600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006800000000000000310000000000000035000000000000004900000000",
            INIT_41 => X"0000004600000000000000390000000000000058000000000000007900000000",
            INIT_42 => X"0000005300000000000000470000000000000017000000000000003300000000",
            INIT_43 => X"000000070000000000000022000000000000004f000000000000004e00000000",
            INIT_44 => X"0000003e000000000000003c0000000000000051000000000000002800000000",
            INIT_45 => X"0000005d000000000000005b0000000000000063000000000000005000000000",
            INIT_46 => X"000000790000000000000078000000000000008d000000000000007300000000",
            INIT_47 => X"000000140000000000000021000000000000007c000000000000007900000000",
            INIT_48 => X"000000760000000000000038000000000000003a000000000000005600000000",
            INIT_49 => X"000000330000000000000040000000000000007f000000000000008300000000",
            INIT_4A => X"0000006300000000000000610000000000000040000000000000003b00000000",
            INIT_4B => X"0000001c000000000000000d000000000000003a000000000000005e00000000",
            INIT_4C => X"000000500000000000000049000000000000005d000000000000005300000000",
            INIT_4D => X"0000004a000000000000005f0000000000000069000000000000006200000000",
            INIT_4E => X"0000007e00000000000000770000000000000084000000000000007400000000",
            INIT_4F => X"00000017000000000000000d0000000000000065000000000000007f00000000",
            INIT_50 => X"000000740000000000000035000000000000003b000000000000005b00000000",
            INIT_51 => X"0000003000000000000000670000000000000087000000000000008400000000",
            INIT_52 => X"000000610000000000000060000000000000004b000000000000002000000000",
            INIT_53 => X"000000490000000000000032000000000000004a000000000000006600000000",
            INIT_54 => X"0000006100000000000000590000000000000052000000000000005a00000000",
            INIT_55 => X"000000310000000000000047000000000000006c000000000000006200000000",
            INIT_56 => X"0000008a0000000000000077000000000000007c000000000000007700000000",
            INIT_57 => X"00000014000000000000000a000000000000005b000000000000007b00000000",
            INIT_58 => X"0000006e000000000000002f0000000000000033000000000000006500000000",
            INIT_59 => X"0000004800000000000000870000000000000087000000000000008100000000",
            INIT_5A => X"0000004f00000000000000520000000000000054000000000000002e00000000",
            INIT_5B => X"0000008700000000000000750000000000000056000000000000005e00000000",
            INIT_5C => X"0000005e000000000000005d0000000000000066000000000000007800000000",
            INIT_5D => X"00000058000000000000004a0000000000000058000000000000005c00000000",
            INIT_5E => X"0000008d00000000000000760000000000000073000000000000008400000000",
            INIT_5F => X"00000007000000000000000b000000000000005b000000000000007700000000",
            INIT_60 => X"0000006000000000000000280000000000000028000000000000005800000000",
            INIT_61 => X"00000077000000000000008b0000000000000083000000000000006b00000000",
            INIT_62 => X"0000005900000000000000570000000000000066000000000000006b00000000",
            INIT_63 => X"0000006c0000000000000051000000000000004a000000000000005f00000000",
            INIT_64 => X"0000005d0000000000000064000000000000006e000000000000007600000000",
            INIT_65 => X"0000005f00000000000000570000000000000055000000000000006600000000",
            INIT_66 => X"0000007100000000000000650000000000000078000000000000007c00000000",
            INIT_67 => X"00000020000000000000000f0000000000000059000000000000007b00000000",
            INIT_68 => X"0000005c0000000000000037000000000000003f000000000000005f00000000",
            INIT_69 => X"00000089000000000000008b000000000000006e000000000000006400000000",
            INIT_6A => X"0000005c00000000000000650000000000000061000000000000007b00000000",
            INIT_6B => X"0000005600000000000000560000000000000058000000000000005a00000000",
            INIT_6C => X"0000006c00000000000000640000000000000058000000000000005500000000",
            INIT_6D => X"0000005f000000000000006e000000000000006c000000000000007200000000",
            INIT_6E => X"00000073000000000000006b0000000000000075000000000000006d00000000",
            INIT_6F => X"0000004c00000000000000310000000000000058000000000000008000000000",
            INIT_70 => X"0000006000000000000000470000000000000045000000000000006a00000000",
            INIT_71 => X"0000008700000000000000860000000000000056000000000000006800000000",
            INIT_72 => X"0000005800000000000000510000000000000057000000000000007400000000",
            INIT_73 => X"0000006a000000000000006e0000000000000060000000000000006000000000",
            INIT_74 => X"0000005c0000000000000057000000000000005f000000000000006200000000",
            INIT_75 => X"00000080000000000000007f000000000000006b000000000000006100000000",
            INIT_76 => X"000000770000000000000074000000000000005e000000000000007a00000000",
            INIT_77 => X"000000460000000000000035000000000000005c000000000000007a00000000",
            INIT_78 => X"0000005c00000000000000400000000000000040000000000000006000000000",
            INIT_79 => X"000000850000000000000079000000000000005f000000000000006700000000",
            INIT_7A => X"0000003300000000000000640000000000000096000000000000008100000000",
            INIT_7B => X"0000007100000000000000620000000000000065000000000000005800000000",
            INIT_7C => X"0000005f00000000000000650000000000000077000000000000008300000000",
            INIT_7D => X"0000009800000000000000710000000000000053000000000000006000000000",
            INIT_7E => X"0000007c00000000000000620000000000000078000000000000009400000000",
            INIT_7F => X"00000048000000000000000d0000000000000039000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "sampleifmap_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005a0000000000000047000000000000004c000000000000005700000000",
            INIT_01 => X"000000820000000000000078000000000000007c000000000000007300000000",
            INIT_02 => X"0000003a0000000000000096000000000000008e000000000000006e00000000",
            INIT_03 => X"0000007800000000000000770000000000000074000000000000005400000000",
            INIT_04 => X"0000008600000000000000850000000000000071000000000000006c00000000",
            INIT_05 => X"0000006e0000000000000067000000000000007e000000000000008900000000",
            INIT_06 => X"00000072000000000000006300000000000000a3000000000000009f00000000",
            INIT_07 => X"0000006b0000000000000021000000000000002a000000000000007500000000",
            INIT_08 => X"0000005d00000000000000640000000000000058000000000000005600000000",
            INIT_09 => X"0000006900000000000000750000000000000063000000000000007500000000",
            INIT_0A => X"0000008b000000000000009b0000000000000066000000000000006e00000000",
            INIT_0B => X"000000810000000000000081000000000000006f000000000000006b00000000",
            INIT_0C => X"00000076000000000000006d0000000000000077000000000000007c00000000",
            INIT_0D => X"00000071000000000000007c0000000000000076000000000000007100000000",
            INIT_0E => X"0000006300000000000000830000000000000075000000000000008300000000",
            INIT_0F => X"0000005700000000000000270000000000000048000000000000006900000000",
            INIT_10 => X"0000007300000000000000780000000000000060000000000000005f00000000",
            INIT_11 => X"0000005600000000000000630000000000000047000000000000006d00000000",
            INIT_12 => X"000000b0000000000000006a0000000000000063000000000000006c00000000",
            INIT_13 => X"00000075000000000000007b000000000000005e000000000000008200000000",
            INIT_14 => X"000000880000000000000081000000000000008d000000000000008900000000",
            INIT_15 => X"000000790000000000000078000000000000006f000000000000008300000000",
            INIT_16 => X"000000430000000000000050000000000000006b000000000000007500000000",
            INIT_17 => X"0000006e00000000000000430000000000000051000000000000004800000000",
            INIT_18 => X"00000057000000000000007d0000000000000070000000000000006d00000000",
            INIT_19 => X"0000005e00000000000000470000000000000048000000000000005800000000",
            INIT_1A => X"0000007300000000000000490000000000000079000000000000006400000000",
            INIT_1B => X"0000009400000000000000870000000000000076000000000000009800000000",
            INIT_1C => X"0000009500000000000000940000000000000082000000000000008500000000",
            INIT_1D => X"0000007a00000000000000790000000000000071000000000000007d00000000",
            INIT_1E => X"0000004e000000000000003a0000000000000071000000000000007200000000",
            INIT_1F => X"0000008a00000000000000730000000000000038000000000000003d00000000",
            INIT_20 => X"0000004300000000000000590000000000000074000000000000007700000000",
            INIT_21 => X"00000066000000000000003c0000000000000048000000000000005800000000",
            INIT_22 => X"00000037000000000000006d0000000000000057000000000000004800000000",
            INIT_23 => X"0000009c000000000000008d0000000000000092000000000000006500000000",
            INIT_24 => X"00000098000000000000008c0000000000000088000000000000009800000000",
            INIT_25 => X"0000007c000000000000007f000000000000007b000000000000008600000000",
            INIT_26 => X"00000062000000000000005d0000000000000069000000000000006d00000000",
            INIT_27 => X"00000077000000000000007a0000000000000062000000000000004d00000000",
            INIT_28 => X"0000005d00000000000000320000000000000061000000000000007e00000000",
            INIT_29 => X"00000060000000000000004b0000000000000046000000000000006000000000",
            INIT_2A => X"000000610000000000000076000000000000003b000000000000005a00000000",
            INIT_2B => X"0000009700000000000000a20000000000000083000000000000004900000000",
            INIT_2C => X"0000007f000000000000008400000000000000a3000000000000009600000000",
            INIT_2D => X"00000075000000000000006e0000000000000076000000000000007d00000000",
            INIT_2E => X"0000004f000000000000005e0000000000000066000000000000006900000000",
            INIT_2F => X"0000006a0000000000000070000000000000008e000000000000006b00000000",
            INIT_30 => X"0000005900000000000000370000000000000051000000000000007000000000",
            INIT_31 => X"000000590000000000000045000000000000004e000000000000005c00000000",
            INIT_32 => X"000000760000000000000053000000000000006b000000000000007700000000",
            INIT_33 => X"0000009c0000000000000097000000000000007d000000000000006b00000000",
            INIT_34 => X"0000007e0000000000000094000000000000009b000000000000009400000000",
            INIT_35 => X"000000750000000000000078000000000000007b000000000000006c00000000",
            INIT_36 => X"0000005600000000000000540000000000000066000000000000007200000000",
            INIT_37 => X"0000006900000000000000630000000000000079000000000000008100000000",
            INIT_38 => X"0000009a00000000000000780000000000000056000000000000006200000000",
            INIT_39 => X"0000004e0000000000000045000000000000005f000000000000007700000000",
            INIT_3A => X"0000004e0000000000000057000000000000007e000000000000007300000000",
            INIT_3B => X"000000960000000000000084000000000000008b000000000000007d00000000",
            INIT_3C => X"0000007e0000000000000092000000000000008e000000000000008d00000000",
            INIT_3D => X"0000007b00000000000000760000000000000084000000000000007900000000",
            INIT_3E => X"0000006f00000000000000520000000000000058000000000000007300000000",
            INIT_3F => X"00000067000000000000006a0000000000000065000000000000007900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a70000000000000088000000000000007400000000",
            INIT_41 => X"0000005c00000000000000600000000000000077000000000000009f00000000",
            INIT_42 => X"0000006f0000000000000066000000000000005a000000000000006600000000",
            INIT_43 => X"0000008f00000000000000830000000000000088000000000000007000000000",
            INIT_44 => X"000000800000000000000096000000000000008e000000000000008600000000",
            INIT_45 => X"000000770000000000000084000000000000009c000000000000007500000000",
            INIT_46 => X"00000053000000000000004e0000000000000059000000000000006600000000",
            INIT_47 => X"0000006c00000000000000710000000000000060000000000000006a00000000",
            INIT_48 => X"000000920000000000000071000000000000006d000000000000006c00000000",
            INIT_49 => X"00000069000000000000007b000000000000009e00000000000000a600000000",
            INIT_4A => X"0000008c00000000000000550000000000000052000000000000006600000000",
            INIT_4B => X"0000007b0000000000000086000000000000007e000000000000009100000000",
            INIT_4C => X"00000089000000000000008a0000000000000073000000000000006800000000",
            INIT_4D => X"0000006a000000000000008a0000000000000096000000000000008300000000",
            INIT_4E => X"0000002d000000000000004a000000000000006f000000000000006100000000",
            INIT_4F => X"0000004b00000000000000690000000000000065000000000000006000000000",
            INIT_50 => X"0000005600000000000000370000000000000055000000000000005800000000",
            INIT_51 => X"0000007e00000000000000970000000000000097000000000000008b00000000",
            INIT_52 => X"0000005700000000000000570000000000000068000000000000006800000000",
            INIT_53 => X"00000052000000000000006e000000000000006e000000000000006f00000000",
            INIT_54 => X"0000008c0000000000000079000000000000004b000000000000003500000000",
            INIT_55 => X"0000007a00000000000000810000000000000078000000000000009100000000",
            INIT_56 => X"00000020000000000000003e0000000000000062000000000000007400000000",
            INIT_57 => X"0000004000000000000000410000000000000062000000000000006100000000",
            INIT_58 => X"000000200000000000000022000000000000005c000000000000005200000000",
            INIT_59 => X"0000009c00000000000000860000000000000075000000000000004b00000000",
            INIT_5A => X"000000570000000000000062000000000000006d000000000000008d00000000",
            INIT_5B => X"0000005f000000000000005b000000000000005a000000000000005200000000",
            INIT_5C => X"0000008b00000000000000790000000000000046000000000000005200000000",
            INIT_5D => X"0000006b0000000000000080000000000000008f000000000000008100000000",
            INIT_5E => X"0000003f000000000000001d000000000000004e000000000000007100000000",
            INIT_5F => X"0000004200000000000000470000000000000047000000000000006300000000",
            INIT_60 => X"0000000d00000000000000230000000000000056000000000000005a00000000",
            INIT_61 => X"000000940000000000000072000000000000004e000000000000000f00000000",
            INIT_62 => X"00000062000000000000006f000000000000008b00000000000000a200000000",
            INIT_63 => X"000000710000000000000056000000000000005b000000000000006100000000",
            INIT_64 => X"0000007e0000000000000073000000000000006a000000000000007800000000",
            INIT_65 => X"0000006a00000000000000870000000000000087000000000000007600000000",
            INIT_66 => X"0000005b0000000000000026000000000000002a000000000000004f00000000",
            INIT_67 => X"0000005300000000000000990000000000000060000000000000002c00000000",
            INIT_68 => X"00000025000000000000002d0000000000000056000000000000005c00000000",
            INIT_69 => X"0000007a0000000000000057000000000000001f000000000000000d00000000",
            INIT_6A => X"0000007a000000000000009e00000000000000ad000000000000009600000000",
            INIT_6B => X"0000005c000000000000005d0000000000000072000000000000007500000000",
            INIT_6C => X"0000007100000000000000670000000000000055000000000000004d00000000",
            INIT_6D => X"0000005b00000000000000730000000000000085000000000000007e00000000",
            INIT_6E => X"0000003c000000000000003b0000000000000032000000000000004e00000000",
            INIT_6F => X"000000620000000000000086000000000000006c000000000000002a00000000",
            INIT_70 => X"0000003800000000000000180000000000000047000000000000005200000000",
            INIT_71 => X"0000005400000000000000230000000000000017000000000000002400000000",
            INIT_72 => X"000000a500000000000000a50000000000000092000000000000007600000000",
            INIT_73 => X"00000079000000000000006f0000000000000082000000000000009600000000",
            INIT_74 => X"00000062000000000000003f0000000000000042000000000000006c00000000",
            INIT_75 => X"0000005600000000000000460000000000000045000000000000004e00000000",
            INIT_76 => X"000000620000000000000060000000000000006c000000000000007500000000",
            INIT_77 => X"00000059000000000000007b0000000000000074000000000000007800000000",
            INIT_78 => X"000000400000000000000011000000000000001b000000000000004100000000",
            INIT_79 => X"00000025000000000000000f000000000000001d000000000000003400000000",
            INIT_7A => X"0000009600000000000000740000000000000064000000000000005900000000",
            INIT_7B => X"0000009c0000000000000088000000000000009800000000000000aa00000000",
            INIT_7C => X"0000004a0000000000000045000000000000007900000000000000a600000000",
            INIT_7D => X"0000007f00000000000000660000000000000047000000000000002f00000000",
            INIT_7E => X"000000820000000000000083000000000000008b000000000000009c00000000",
            INIT_7F => X"0000007500000000000000920000000000000088000000000000009300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "sampleifmap_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000058000000000000004d000000000000008b00000000000000b300000000",
            INIT_01 => X"00000097000000000000009c000000000000009d000000000000008d00000000",
            INIT_02 => X"000000970000000000000090000000000000009e000000000000009c00000000",
            INIT_03 => X"0000007600000000000000790000000000000088000000000000009700000000",
            INIT_04 => X"000000540000000000000054000000000000006c000000000000007e00000000",
            INIT_05 => X"00000053000000000000005e0000000000000062000000000000006200000000",
            INIT_06 => X"0000006000000000000000540000000000000056000000000000005a00000000",
            INIT_07 => X"0000004d000000000000004c0000000000000057000000000000007500000000",
            INIT_08 => X"000000920000000000000080000000000000008500000000000000b800000000",
            INIT_09 => X"000000a7000000000000009e000000000000009f000000000000009f00000000",
            INIT_0A => X"0000009a000000000000009900000000000000a200000000000000a500000000",
            INIT_0B => X"0000007d00000000000000880000000000000096000000000000009600000000",
            INIT_0C => X"00000052000000000000005a000000000000006d000000000000008100000000",
            INIT_0D => X"00000058000000000000005e0000000000000062000000000000005d00000000",
            INIT_0E => X"0000006a000000000000005b000000000000004c000000000000004e00000000",
            INIT_0F => X"0000005a000000000000005b0000000000000062000000000000007600000000",
            INIT_10 => X"000000aa00000000000000b0000000000000009800000000000000b400000000",
            INIT_11 => X"000000a4000000000000009b000000000000009800000000000000a400000000",
            INIT_12 => X"0000009f00000000000000a200000000000000aa00000000000000a200000000",
            INIT_13 => X"0000008c00000000000000920000000000000097000000000000009c00000000",
            INIT_14 => X"000000470000000000000058000000000000007c000000000000009200000000",
            INIT_15 => X"0000006b00000000000000670000000000000062000000000000005500000000",
            INIT_16 => X"0000006f000000000000006f000000000000006d000000000000006500000000",
            INIT_17 => X"0000005f000000000000005d0000000000000065000000000000006f00000000",
            INIT_18 => X"000000b500000000000000b800000000000000ae00000000000000af00000000",
            INIT_19 => X"000000a300000000000000a4000000000000009800000000000000a800000000",
            INIT_1A => X"000000a800000000000000a700000000000000b300000000000000a600000000",
            INIT_1B => X"000000a4000000000000009f00000000000000a200000000000000ae00000000",
            INIT_1C => X"0000003a00000000000000590000000000000089000000000000009700000000",
            INIT_1D => X"0000006b0000000000000063000000000000005a000000000000004800000000",
            INIT_1E => X"00000079000000000000007d0000000000000080000000000000007500000000",
            INIT_1F => X"0000006f000000000000006d0000000000000061000000000000006900000000",
            INIT_20 => X"000000ac00000000000000a700000000000000ae00000000000000af00000000",
            INIT_21 => X"000000af00000000000000b000000000000000a100000000000000a200000000",
            INIT_22 => X"000000b400000000000000b300000000000000b200000000000000b200000000",
            INIT_23 => X"000000a400000000000000a000000000000000a800000000000000b000000000",
            INIT_24 => X"000000450000000000000078000000000000009c00000000000000ad00000000",
            INIT_25 => X"0000005e0000000000000063000000000000005a000000000000004200000000",
            INIT_26 => X"0000007b000000000000007f000000000000007c000000000000006900000000",
            INIT_27 => X"0000007400000000000000710000000000000068000000000000007000000000",
            INIT_28 => X"000000aa000000000000009000000000000000ae00000000000000b500000000",
            INIT_29 => X"000000b300000000000000b000000000000000a600000000000000a900000000",
            INIT_2A => X"000000b500000000000000b400000000000000b400000000000000b400000000",
            INIT_2B => X"00000096000000000000009f00000000000000ae00000000000000b000000000",
            INIT_2C => X"00000074000000000000009b00000000000000af00000000000000b500000000",
            INIT_2D => X"000000700000000000000083000000000000007d000000000000006000000000",
            INIT_2E => X"00000079000000000000007a0000000000000078000000000000007500000000",
            INIT_2F => X"0000007c00000000000000760000000000000078000000000000007900000000",
            INIT_30 => X"000000b2000000000000008a000000000000009c00000000000000c000000000",
            INIT_31 => X"000000af00000000000000b000000000000000ae00000000000000af00000000",
            INIT_32 => X"000000b800000000000000ba00000000000000b400000000000000b800000000",
            INIT_33 => X"0000009900000000000000ad00000000000000bb00000000000000bb00000000",
            INIT_34 => X"000000a700000000000000ad00000000000000ad00000000000000a600000000",
            INIT_35 => X"0000007900000000000000940000000000000095000000000000009600000000",
            INIT_36 => X"0000006f000000000000006d0000000000000075000000000000007300000000",
            INIT_37 => X"00000080000000000000007b000000000000007a000000000000007800000000",
            INIT_38 => X"000000ab000000000000009c000000000000007d00000000000000b900000000",
            INIT_39 => X"000000b800000000000000af00000000000000af00000000000000ad00000000",
            INIT_3A => X"000000c200000000000000c100000000000000b700000000000000bc00000000",
            INIT_3B => X"000000a600000000000000b800000000000000b900000000000000bd00000000",
            INIT_3C => X"000000b000000000000000b100000000000000ac00000000000000a400000000",
            INIT_3D => X"0000007a000000000000008f000000000000008900000000000000aa00000000",
            INIT_3E => X"000000670000000000000060000000000000006e000000000000006b00000000",
            INIT_3F => X"0000007d000000000000007b0000000000000076000000000000007500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a0000000000000009f0000000000000095000000000000009b00000000",
            INIT_41 => X"000000b400000000000000b200000000000000ad00000000000000ac00000000",
            INIT_42 => X"000000bf00000000000000ba00000000000000ba00000000000000bb00000000",
            INIT_43 => X"000000a000000000000000ac00000000000000af00000000000000bb00000000",
            INIT_44 => X"000000b000000000000000a60000000000000097000000000000009a00000000",
            INIT_45 => X"0000008500000000000000a6000000000000009b00000000000000b700000000",
            INIT_46 => X"0000007700000000000000700000000000000068000000000000006800000000",
            INIT_47 => X"0000007d000000000000007a000000000000007a000000000000007600000000",
            INIT_48 => X"000000a900000000000000930000000000000098000000000000009a00000000",
            INIT_49 => X"000000aa00000000000000b700000000000000b200000000000000b200000000",
            INIT_4A => X"000000c100000000000000c600000000000000bc00000000000000b000000000",
            INIT_4B => X"000000a900000000000000a500000000000000a700000000000000ae00000000",
            INIT_4C => X"000000a90000000000000092000000000000008c000000000000009d00000000",
            INIT_4D => X"0000008d00000000000000ab00000000000000a000000000000000b300000000",
            INIT_4E => X"0000007700000000000000750000000000000068000000000000005f00000000",
            INIT_4F => X"0000007d0000000000000076000000000000007b000000000000007400000000",
            INIT_50 => X"000000b1000000000000009f0000000000000070000000000000008600000000",
            INIT_51 => X"000000ba00000000000000b800000000000000b800000000000000ae00000000",
            INIT_52 => X"000000b000000000000000bf00000000000000c200000000000000ba00000000",
            INIT_53 => X"000000bb00000000000000a7000000000000009e000000000000009b00000000",
            INIT_54 => X"000000970000000000000086000000000000009300000000000000ae00000000",
            INIT_55 => X"0000007c000000000000009b000000000000009c00000000000000a000000000",
            INIT_56 => X"0000006600000000000000690000000000000066000000000000004a00000000",
            INIT_57 => X"0000007f000000000000007b0000000000000075000000000000006b00000000",
            INIT_58 => X"0000009d00000000000000ae000000000000005b000000000000004100000000",
            INIT_59 => X"000000be00000000000000bf00000000000000b1000000000000009300000000",
            INIT_5A => X"000000b000000000000000ac00000000000000b000000000000000bc00000000",
            INIT_5B => X"000000a3000000000000009400000000000000ae00000000000000b800000000",
            INIT_5C => X"000000950000000000000085000000000000009a00000000000000b000000000",
            INIT_5D => X"0000005000000000000000830000000000000095000000000000009800000000",
            INIT_5E => X"0000006600000000000000670000000000000061000000000000004200000000",
            INIT_5F => X"0000007d00000000000000780000000000000071000000000000006700000000",
            INIT_60 => X"000000b100000000000000bf000000000000005c000000000000001500000000",
            INIT_61 => X"000000b600000000000000bd00000000000000ca00000000000000bc00000000",
            INIT_62 => X"000000bc00000000000000a5000000000000009c00000000000000b300000000",
            INIT_63 => X"00000072000000000000009800000000000000ae00000000000000c800000000",
            INIT_64 => X"000000890000000000000078000000000000007f000000000000005f00000000",
            INIT_65 => X"0000004e00000000000000720000000000000088000000000000009700000000",
            INIT_66 => X"0000006200000000000000590000000000000049000000000000004000000000",
            INIT_67 => X"0000007600000000000000750000000000000071000000000000006200000000",
            INIT_68 => X"000000ad00000000000000a80000000000000063000000000000002c00000000",
            INIT_69 => X"000000bb00000000000000bc00000000000000c300000000000000c800000000",
            INIT_6A => X"000000c200000000000000b4000000000000009500000000000000a500000000",
            INIT_6B => X"0000009a00000000000000a800000000000000a800000000000000b900000000",
            INIT_6C => X"0000008a00000000000000910000000000000092000000000000006b00000000",
            INIT_6D => X"000000480000000000000064000000000000007f000000000000009c00000000",
            INIT_6E => X"0000006000000000000000530000000000000040000000000000003900000000",
            INIT_6F => X"0000006f000000000000006c000000000000006a000000000000006200000000",
            INIT_70 => X"0000009f00000000000000750000000000000076000000000000006900000000",
            INIT_71 => X"000000bb00000000000000b400000000000000be00000000000000c400000000",
            INIT_72 => X"000000c100000000000000c600000000000000ad00000000000000ad00000000",
            INIT_73 => X"000000bc00000000000000b400000000000000a500000000000000ab00000000",
            INIT_74 => X"000000b300000000000000ad00000000000000bb00000000000000ae00000000",
            INIT_75 => X"000000480000000000000069000000000000008000000000000000a000000000",
            INIT_76 => X"0000006c00000000000000570000000000000045000000000000004300000000",
            INIT_77 => X"0000006600000000000000610000000000000064000000000000006300000000",
            INIT_78 => X"0000009d00000000000000680000000000000071000000000000008a00000000",
            INIT_79 => X"000000a800000000000000b400000000000000c400000000000000c600000000",
            INIT_7A => X"000000cd00000000000000cb00000000000000bf00000000000000b400000000",
            INIT_7B => X"000000c800000000000000c400000000000000bf00000000000000d200000000",
            INIT_7C => X"000000be00000000000000bc00000000000000bb00000000000000c000000000",
            INIT_7D => X"000000500000000000000071000000000000009900000000000000a800000000",
            INIT_7E => X"0000008700000000000000600000000000000040000000000000004600000000",
            INIT_7F => X"00000062000000000000005a000000000000005a000000000000007800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "sampleifmap_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000930000000000000073000000000000008a000000000000009600000000",
            INIT_01 => X"0000009600000000000000b000000000000000bb00000000000000be00000000",
            INIT_02 => X"000000c600000000000000d300000000000000c700000000000000ab00000000",
            INIT_03 => X"000000cb00000000000000be00000000000000c200000000000000d300000000",
            INIT_04 => X"000000bd00000000000000b800000000000000ba00000000000000bf00000000",
            INIT_05 => X"00000046000000000000006400000000000000a600000000000000be00000000",
            INIT_06 => X"0000008f000000000000006a0000000000000038000000000000002f00000000",
            INIT_07 => X"0000005e000000000000004a000000000000005c000000000000009500000000",
            INIT_08 => X"000000a50000000000000092000000000000009b000000000000009b00000000",
            INIT_09 => X"0000009100000000000000bf00000000000000c000000000000000bd00000000",
            INIT_0A => X"0000009500000000000000a900000000000000d2000000000000009c00000000",
            INIT_0B => X"000000a800000000000000b200000000000000c200000000000000c000000000",
            INIT_0C => X"000000a700000000000000aa00000000000000b500000000000000a900000000",
            INIT_0D => X"0000002b00000000000000430000000000000075000000000000009a00000000",
            INIT_0E => X"0000008f00000000000000680000000000000031000000000000002200000000",
            INIT_0F => X"00000050000000000000003f000000000000006a000000000000009c00000000",
            INIT_10 => X"000000a6000000000000008a00000000000000a200000000000000a500000000",
            INIT_11 => X"0000008900000000000000ba00000000000000be00000000000000c400000000",
            INIT_12 => X"000000a9000000000000009d00000000000000c9000000000000007400000000",
            INIT_13 => X"0000008f000000000000008000000000000000b600000000000000d200000000",
            INIT_14 => X"00000061000000000000007f0000000000000093000000000000007c00000000",
            INIT_15 => X"00000033000000000000002f0000000000000038000000000000005200000000",
            INIT_16 => X"0000009d00000000000000690000000000000040000000000000002b00000000",
            INIT_17 => X"000000410000000000000039000000000000007b000000000000009d00000000",
            INIT_18 => X"0000009e0000000000000078000000000000009600000000000000a900000000",
            INIT_19 => X"0000009800000000000000be00000000000000be00000000000000be00000000",
            INIT_1A => X"000000b900000000000000bc0000000000000099000000000000003c00000000",
            INIT_1B => X"000000ce000000000000009000000000000000a500000000000000c300000000",
            INIT_1C => X"0000003d0000000000000065000000000000008900000000000000b100000000",
            INIT_1D => X"0000005000000000000000470000000000000033000000000000003700000000",
            INIT_1E => X"000000a0000000000000006e000000000000004a000000000000003700000000",
            INIT_1F => X"000000320000000000000036000000000000008e00000000000000b000000000",
            INIT_20 => X"000000a6000000000000009600000000000000a000000000000000aa00000000",
            INIT_21 => X"0000009a00000000000000ba00000000000000bc00000000000000ba00000000",
            INIT_22 => X"00000092000000000000007e0000000000000031000000000000002000000000",
            INIT_23 => X"000000c0000000000000008c000000000000008c000000000000009b00000000",
            INIT_24 => X"0000003e0000000000000061000000000000009c00000000000000cc00000000",
            INIT_25 => X"0000005700000000000000520000000000000049000000000000004900000000",
            INIT_26 => X"000000a6000000000000006b000000000000003e000000000000003a00000000",
            INIT_27 => X"00000033000000000000004800000000000000a700000000000000bc00000000",
            INIT_28 => X"0000009c000000000000009700000000000000ab00000000000000b200000000",
            INIT_29 => X"0000007c00000000000000a300000000000000b200000000000000b500000000",
            INIT_2A => X"000000370000000000000028000000000000001d000000000000002400000000",
            INIT_2B => X"0000008200000000000000650000000000000063000000000000004e00000000",
            INIT_2C => X"00000037000000000000005f000000000000007b000000000000009000000000",
            INIT_2D => X"00000055000000000000003c0000000000000033000000000000003400000000",
            INIT_2E => X"000000990000000000000066000000000000004d000000000000004e00000000",
            INIT_2F => X"00000037000000000000005900000000000000b100000000000000bb00000000",
            INIT_30 => X"00000098000000000000009200000000000000ab00000000000000b500000000",
            INIT_31 => X"00000069000000000000009500000000000000a700000000000000a900000000",
            INIT_32 => X"0000002e0000000000000042000000000000005e000000000000004f00000000",
            INIT_33 => X"00000078000000000000005c0000000000000047000000000000002f00000000",
            INIT_34 => X"0000002900000000000000380000000000000037000000000000005a00000000",
            INIT_35 => X"00000037000000000000001e0000000000000022000000000000002300000000",
            INIT_36 => X"0000007700000000000000610000000000000056000000000000005200000000",
            INIT_37 => X"0000003c000000000000006a00000000000000ae00000000000000ad00000000",
            INIT_38 => X"000000a3000000000000009e000000000000009c00000000000000b100000000",
            INIT_39 => X"00000089000000000000009400000000000000a0000000000000009c00000000",
            INIT_3A => X"0000006b00000000000000660000000000000076000000000000008f00000000",
            INIT_3B => X"00000067000000000000007d000000000000006d000000000000006e00000000",
            INIT_3C => X"0000001300000000000000100000000000000011000000000000002f00000000",
            INIT_3D => X"00000013000000000000000e000000000000001c000000000000001800000000",
            INIT_3E => X"0000006300000000000000600000000000000041000000000000002b00000000",
            INIT_3F => X"00000043000000000000008500000000000000ad000000000000008c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b600000000000000a7000000000000008b000000000000009e00000000",
            INIT_41 => X"000000c000000000000000ab000000000000008c000000000000009700000000",
            INIT_42 => X"000000880000000000000085000000000000007400000000000000ac00000000",
            INIT_43 => X"00000065000000000000007f000000000000008d000000000000009200000000",
            INIT_44 => X"0000001900000000000000200000000000000025000000000000004100000000",
            INIT_45 => X"0000000f000000000000000a0000000000000011000000000000001800000000",
            INIT_46 => X"0000004e00000000000000610000000000000042000000000000001400000000",
            INIT_47 => X"00000069000000000000009c0000000000000094000000000000006200000000",
            INIT_48 => X"000000ab00000000000000ae00000000000000a400000000000000a000000000",
            INIT_49 => X"000000b100000000000000940000000000000088000000000000009e00000000",
            INIT_4A => X"0000009700000000000000a9000000000000009300000000000000b800000000",
            INIT_4B => X"0000007d000000000000008e000000000000008b000000000000007f00000000",
            INIT_4C => X"0000002b000000000000003f000000000000004d000000000000006700000000",
            INIT_4D => X"0000001a00000000000000110000000000000018000000000000002100000000",
            INIT_4E => X"000000320000000000000048000000000000003e000000000000001f00000000",
            INIT_4F => X"000000880000000000000078000000000000005a000000000000004800000000",
            INIT_50 => X"000000a700000000000000a700000000000000a300000000000000a000000000",
            INIT_51 => X"00000078000000000000008c00000000000000a800000000000000b100000000",
            INIT_52 => X"000000820000000000000076000000000000008f00000000000000ab00000000",
            INIT_53 => X"0000009100000000000000a6000000000000009c000000000000007b00000000",
            INIT_54 => X"0000004e000000000000005b0000000000000069000000000000007c00000000",
            INIT_55 => X"0000004300000000000000380000000000000042000000000000004c00000000",
            INIT_56 => X"0000004900000000000000410000000000000041000000000000004600000000",
            INIT_57 => X"0000006a0000000000000051000000000000007b000000000000006400000000",
            INIT_58 => X"00000093000000000000008c000000000000009f000000000000009c00000000",
            INIT_59 => X"0000007b000000000000009900000000000000aa00000000000000b400000000",
            INIT_5A => X"0000007e0000000000000073000000000000009c000000000000008b00000000",
            INIT_5B => X"000000a200000000000000a8000000000000009e000000000000008300000000",
            INIT_5C => X"00000078000000000000007b0000000000000077000000000000007f00000000",
            INIT_5D => X"0000007700000000000000690000000000000068000000000000007000000000",
            INIT_5E => X"0000006d00000000000000680000000000000069000000000000007400000000",
            INIT_5F => X"00000068000000000000005c0000000000000086000000000000007a00000000",
            INIT_60 => X"0000008b000000000000007b000000000000009e00000000000000a400000000",
            INIT_61 => X"0000008c000000000000008d000000000000009c00000000000000ad00000000",
            INIT_62 => X"000000a100000000000000820000000000000079000000000000008d00000000",
            INIT_63 => X"000000a800000000000000a6000000000000009d000000000000009700000000",
            INIT_64 => X"00000084000000000000008f000000000000008a000000000000009000000000",
            INIT_65 => X"00000094000000000000008a0000000000000085000000000000008100000000",
            INIT_66 => X"0000008400000000000000860000000000000089000000000000008f00000000",
            INIT_67 => X"0000009300000000000000730000000000000064000000000000007800000000",
            INIT_68 => X"000000a800000000000000900000000000000095000000000000008e00000000",
            INIT_69 => X"0000009e000000000000009e00000000000000a100000000000000a700000000",
            INIT_6A => X"000000a90000000000000097000000000000009000000000000000a500000000",
            INIT_6B => X"000000a2000000000000009e00000000000000a000000000000000a100000000",
            INIT_6C => X"0000007f00000000000000890000000000000091000000000000009900000000",
            INIT_6D => X"0000009e00000000000000960000000000000095000000000000008d00000000",
            INIT_6E => X"0000008f00000000000000940000000000000096000000000000009f00000000",
            INIT_6F => X"0000009f000000000000008b0000000000000077000000000000007b00000000",
            INIT_70 => X"000000b900000000000000b300000000000000a6000000000000009800000000",
            INIT_71 => X"000000a800000000000000aa00000000000000a700000000000000a700000000",
            INIT_72 => X"000000b200000000000000ad00000000000000a400000000000000a700000000",
            INIT_73 => X"000000850000000000000089000000000000009d00000000000000a900000000",
            INIT_74 => X"00000088000000000000008c000000000000008f000000000000009200000000",
            INIT_75 => X"0000009d00000000000000980000000000000097000000000000008c00000000",
            INIT_76 => X"000000900000000000000099000000000000009c00000000000000a600000000",
            INIT_77 => X"0000009900000000000000900000000000000083000000000000008500000000",
            INIT_78 => X"000000ab00000000000000b700000000000000b2000000000000009f00000000",
            INIT_79 => X"0000009f0000000000000091000000000000007d000000000000008b00000000",
            INIT_7A => X"0000009c0000000000000095000000000000008b00000000000000a200000000",
            INIT_7B => X"0000007300000000000000830000000000000098000000000000009e00000000",
            INIT_7C => X"0000008f0000000000000094000000000000008e000000000000008400000000",
            INIT_7D => X"000000a1000000000000009c000000000000009d000000000000009000000000",
            INIT_7E => X"0000009c0000000000000094000000000000009f00000000000000a700000000",
            INIT_7F => X"0000009800000000000000990000000000000096000000000000009c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "sampleifmap_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003b00000000000000310000000000000060000000000000007600000000",
            INIT_01 => X"000000530000000000000054000000000000005f000000000000006000000000",
            INIT_02 => X"0000005a00000000000000530000000000000061000000000000005f00000000",
            INIT_03 => X"0000004f000000000000004b0000000000000052000000000000005c00000000",
            INIT_04 => X"00000032000000000000003b0000000000000050000000000000005b00000000",
            INIT_05 => X"0000003300000000000000380000000000000038000000000000003700000000",
            INIT_06 => X"0000003a00000000000000330000000000000038000000000000003c00000000",
            INIT_07 => X"0000002f000000000000002f0000000000000035000000000000004c00000000",
            INIT_08 => X"0000006900000000000000590000000000000058000000000000008200000000",
            INIT_09 => X"00000068000000000000005d0000000000000060000000000000006c00000000",
            INIT_0A => X"0000005b000000000000005a0000000000000062000000000000006500000000",
            INIT_0B => X"00000048000000000000004f0000000000000057000000000000005400000000",
            INIT_0C => X"00000032000000000000003d0000000000000048000000000000005200000000",
            INIT_0D => X"0000003300000000000000370000000000000038000000000000003700000000",
            INIT_0E => X"0000004100000000000000350000000000000028000000000000002b00000000",
            INIT_0F => X"00000039000000000000003a000000000000003d000000000000004b00000000",
            INIT_10 => X"0000007a00000000000000810000000000000068000000000000008400000000",
            INIT_11 => X"0000006a000000000000005f0000000000000059000000000000006c00000000",
            INIT_12 => X"0000005e00000000000000620000000000000069000000000000006200000000",
            INIT_13 => X"0000004c000000000000004f0000000000000050000000000000005500000000",
            INIT_14 => X"0000002a0000000000000036000000000000004c000000000000005500000000",
            INIT_15 => X"00000042000000000000003f000000000000003a000000000000003300000000",
            INIT_16 => X"0000004200000000000000430000000000000042000000000000003c00000000",
            INIT_17 => X"000000390000000000000038000000000000003e000000000000004300000000",
            INIT_18 => X"000000840000000000000088000000000000007f000000000000008100000000",
            INIT_19 => X"000000690000000000000068000000000000005a000000000000007000000000",
            INIT_1A => X"0000006600000000000000650000000000000071000000000000006500000000",
            INIT_1B => X"0000005d0000000000000057000000000000005a000000000000006700000000",
            INIT_1C => X"0000001f0000000000000033000000000000004e000000000000004f00000000",
            INIT_1D => X"0000003e00000000000000390000000000000033000000000000002a00000000",
            INIT_1E => X"0000004a000000000000004b000000000000004d000000000000004600000000",
            INIT_1F => X"0000004500000000000000430000000000000037000000000000003c00000000",
            INIT_20 => X"0000007f0000000000000079000000000000007f000000000000008000000000",
            INIT_21 => X"0000007200000000000000720000000000000063000000000000006d00000000",
            INIT_22 => X"000000710000000000000070000000000000006f000000000000006f00000000",
            INIT_23 => X"0000005c00000000000000590000000000000063000000000000006c00000000",
            INIT_24 => X"0000002c000000000000004e0000000000000059000000000000005e00000000",
            INIT_25 => X"0000002e00000000000000380000000000000034000000000000002700000000",
            INIT_26 => X"0000004900000000000000470000000000000043000000000000003500000000",
            INIT_27 => X"000000470000000000000045000000000000003b000000000000004200000000",
            INIT_28 => X"0000007f00000000000000680000000000000083000000000000008900000000",
            INIT_29 => X"000000740000000000000071000000000000006a000000000000007600000000",
            INIT_2A => X"0000007100000000000000740000000000000075000000000000007300000000",
            INIT_2B => X"00000054000000000000005a0000000000000069000000000000006d00000000",
            INIT_2C => X"0000004f00000000000000670000000000000068000000000000006a00000000",
            INIT_2D => X"0000003d0000000000000052000000000000004d000000000000003a00000000",
            INIT_2E => X"000000460000000000000043000000000000003f000000000000003e00000000",
            INIT_2F => X"0000004b00000000000000460000000000000048000000000000004900000000",
            INIT_30 => X"0000008700000000000000660000000000000077000000000000009800000000",
            INIT_31 => X"0000006f00000000000000730000000000000075000000000000007a00000000",
            INIT_32 => X"00000070000000000000007c000000000000007b000000000000007900000000",
            INIT_33 => X"0000005c00000000000000660000000000000071000000000000007300000000",
            INIT_34 => X"0000006e000000000000006d0000000000000065000000000000006400000000",
            INIT_35 => X"00000043000000000000005b0000000000000057000000000000005c00000000",
            INIT_36 => X"0000003b00000000000000380000000000000040000000000000003e00000000",
            INIT_37 => X"0000004e000000000000004a0000000000000048000000000000004500000000",
            INIT_38 => X"0000007e00000000000000780000000000000059000000000000009300000000",
            INIT_39 => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_3A => X"00000073000000000000007c000000000000007a000000000000008000000000",
            INIT_3B => X"00000064000000000000006c000000000000006d000000000000007300000000",
            INIT_3C => X"0000006a000000000000006d0000000000000068000000000000006500000000",
            INIT_3D => X"000000480000000000000057000000000000004b000000000000006600000000",
            INIT_3E => X"00000035000000000000002e000000000000003c000000000000003b00000000",
            INIT_3F => X"0000004b00000000000000490000000000000044000000000000004200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000720000000000000078000000000000006f000000000000007600000000",
            INIT_41 => X"0000007700000000000000750000000000000074000000000000007700000000",
            INIT_42 => X"0000006d000000000000006f000000000000007a000000000000008000000000",
            INIT_43 => X"0000005e00000000000000610000000000000067000000000000007300000000",
            INIT_44 => X"0000006400000000000000610000000000000059000000000000005e00000000",
            INIT_45 => X"000000590000000000000072000000000000005f000000000000006d00000000",
            INIT_46 => X"000000470000000000000040000000000000003a000000000000003e00000000",
            INIT_47 => X"0000004b00000000000000480000000000000048000000000000004600000000",
            INIT_48 => X"0000007800000000000000690000000000000071000000000000007700000000",
            INIT_49 => X"0000006f000000000000007b000000000000007a000000000000007c00000000",
            INIT_4A => X"00000079000000000000007d000000000000007b000000000000007600000000",
            INIT_4B => X"0000006f0000000000000065000000000000006d000000000000007600000000",
            INIT_4C => X"0000006000000000000000520000000000000055000000000000006900000000",
            INIT_4D => X"00000067000000000000007a0000000000000064000000000000006a00000000",
            INIT_4E => X"000000490000000000000047000000000000003e000000000000003d00000000",
            INIT_4F => X"0000004b0000000000000044000000000000004b000000000000004700000000",
            INIT_50 => X"0000007e00000000000000720000000000000048000000000000006400000000",
            INIT_51 => X"0000007e000000000000007c000000000000007f000000000000007800000000",
            INIT_52 => X"0000007b00000000000000800000000000000081000000000000007f00000000",
            INIT_53 => X"0000009000000000000000780000000000000077000000000000007900000000",
            INIT_54 => X"00000058000000000000004f0000000000000063000000000000008300000000",
            INIT_55 => X"0000005b000000000000006c0000000000000061000000000000005f00000000",
            INIT_56 => X"0000003b000000000000003d000000000000003e000000000000002e00000000",
            INIT_57 => X"0000004c00000000000000490000000000000046000000000000004000000000",
            INIT_58 => X"00000069000000000000007f0000000000000034000000000000002200000000",
            INIT_59 => X"000000830000000000000084000000000000007a000000000000005d00000000",
            INIT_5A => X"0000008c00000000000000780000000000000073000000000000008100000000",
            INIT_5B => X"000000850000000000000074000000000000009700000000000000a600000000",
            INIT_5C => X"000000610000000000000056000000000000006e000000000000008d00000000",
            INIT_5D => X"000000310000000000000056000000000000005c000000000000006000000000",
            INIT_5E => X"0000003c000000000000003e000000000000003c000000000000002a00000000",
            INIT_5F => X"0000004a00000000000000450000000000000042000000000000003e00000000",
            INIT_60 => X"0000007d000000000000008e0000000000000040000000000000000400000000",
            INIT_61 => X"00000084000000000000008c000000000000009a000000000000008c00000000",
            INIT_62 => X"0000009c000000000000007b000000000000006b000000000000007f00000000",
            INIT_63 => X"000000530000000000000077000000000000009300000000000000b200000000",
            INIT_64 => X"000000640000000000000053000000000000005b000000000000004000000000",
            INIT_65 => X"00000031000000000000004d000000000000005c000000000000006f00000000",
            INIT_66 => X"000000390000000000000037000000000000002f000000000000002900000000",
            INIT_67 => X"0000004400000000000000420000000000000043000000000000003b00000000",
            INIT_68 => X"0000007b000000000000007a0000000000000048000000000000001800000000",
            INIT_69 => X"0000008d000000000000008f0000000000000096000000000000009c00000000",
            INIT_6A => X"000000a0000000000000008f000000000000006a000000000000007700000000",
            INIT_6B => X"0000007700000000000000800000000000000081000000000000009700000000",
            INIT_6C => X"0000006d00000000000000730000000000000074000000000000004d00000000",
            INIT_6D => X"0000002d0000000000000044000000000000005a000000000000007b00000000",
            INIT_6E => X"000000370000000000000033000000000000002b000000000000002300000000",
            INIT_6F => X"0000003e000000000000003a000000000000003e000000000000003b00000000",
            INIT_70 => X"00000070000000000000004a0000000000000052000000000000004500000000",
            INIT_71 => X"0000008f00000000000000860000000000000091000000000000009600000000",
            INIT_72 => X"0000009c00000000000000a10000000000000084000000000000008300000000",
            INIT_73 => X"0000009700000000000000850000000000000072000000000000007d00000000",
            INIT_74 => X"00000098000000000000009200000000000000a0000000000000009100000000",
            INIT_75 => X"0000002f000000000000004b000000000000005d000000000000008100000000",
            INIT_76 => X"0000004400000000000000380000000000000030000000000000002f00000000",
            INIT_77 => X"000000390000000000000036000000000000003c000000000000003c00000000",
            INIT_78 => X"00000070000000000000003b0000000000000041000000000000005700000000",
            INIT_79 => X"0000007d00000000000000860000000000000096000000000000009800000000",
            INIT_7A => X"000000a500000000000000a7000000000000009b000000000000008f00000000",
            INIT_7B => X"000000a0000000000000008f0000000000000084000000000000009b00000000",
            INIT_7C => X"000000a1000000000000009f000000000000009e00000000000000a200000000",
            INIT_7D => X"0000003900000000000000540000000000000078000000000000008900000000",
            INIT_7E => X"0000005f0000000000000040000000000000002b000000000000003300000000",
            INIT_7F => X"0000003900000000000000360000000000000037000000000000005100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "sampleifmap_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000660000000000000040000000000000004e000000000000005800000000",
            INIT_01 => X"0000006c0000000000000081000000000000008d000000000000009000000000",
            INIT_02 => X"0000009d00000000000000af00000000000000a5000000000000008b00000000",
            INIT_03 => X"0000009f00000000000000860000000000000086000000000000009e00000000",
            INIT_04 => X"0000009800000000000000930000000000000094000000000000009a00000000",
            INIT_05 => X"0000003100000000000000490000000000000087000000000000009a00000000",
            INIT_06 => X"00000067000000000000004b0000000000000023000000000000001e00000000",
            INIT_07 => X"00000039000000000000002c000000000000003d000000000000006f00000000",
            INIT_08 => X"0000007400000000000000570000000000000057000000000000005600000000",
            INIT_09 => X"0000006900000000000000910000000000000093000000000000008f00000000",
            INIT_0A => X"0000006c000000000000008500000000000000b3000000000000008000000000",
            INIT_0B => X"00000079000000000000007a000000000000008b000000000000009100000000",
            INIT_0C => X"00000079000000000000007c0000000000000087000000000000007d00000000",
            INIT_0D => X"00000018000000000000002a0000000000000058000000000000007200000000",
            INIT_0E => X"000000660000000000000049000000000000001d000000000000001300000000",
            INIT_0F => X"0000002e00000000000000270000000000000050000000000000007500000000",
            INIT_10 => X"00000076000000000000004d000000000000005c000000000000005c00000000",
            INIT_11 => X"0000006200000000000000910000000000000099000000000000009c00000000",
            INIT_12 => X"0000007a000000000000007400000000000000aa000000000000005c00000000",
            INIT_13 => X"00000062000000000000004b000000000000008300000000000000a500000000",
            INIT_14 => X"0000004000000000000000550000000000000061000000000000004c00000000",
            INIT_15 => X"0000001b0000000000000011000000000000001b000000000000003600000000",
            INIT_16 => X"0000007500000000000000450000000000000028000000000000001a00000000",
            INIT_17 => X"0000002800000000000000240000000000000064000000000000007f00000000",
            INIT_18 => X"0000006e000000000000003c0000000000000054000000000000005e00000000",
            INIT_19 => X"00000073000000000000009b00000000000000a3000000000000009c00000000",
            INIT_1A => X"000000890000000000000094000000000000007c000000000000002700000000",
            INIT_1B => X"0000009c00000000000000570000000000000071000000000000009500000000",
            INIT_1C => X"00000027000000000000003d0000000000000050000000000000007800000000",
            INIT_1D => X"0000002e00000000000000220000000000000018000000000000002700000000",
            INIT_1E => X"000000780000000000000045000000000000002d000000000000001f00000000",
            INIT_1F => X"000000200000000000000022000000000000007b000000000000009900000000",
            INIT_20 => X"000000720000000000000059000000000000005d000000000000006100000000",
            INIT_21 => X"00000075000000000000009800000000000000a2000000000000009600000000",
            INIT_22 => X"000000740000000000000064000000000000001d000000000000000d00000000",
            INIT_23 => X"0000007c00000000000000490000000000000056000000000000007300000000",
            INIT_24 => X"0000001b000000000000002f000000000000005b000000000000008600000000",
            INIT_25 => X"0000003200000000000000310000000000000032000000000000003100000000",
            INIT_26 => X"0000007d0000000000000042000000000000001e000000000000001900000000",
            INIT_27 => X"000000200000000000000038000000000000009600000000000000a200000000",
            INIT_28 => X"0000006300000000000000570000000000000068000000000000006a00000000",
            INIT_29 => X"0000005700000000000000810000000000000096000000000000008d00000000",
            INIT_2A => X"000000250000000000000016000000000000000b000000000000000f00000000",
            INIT_2B => X"0000003e00000000000000290000000000000039000000000000003600000000",
            INIT_2C => X"0000001a00000000000000360000000000000048000000000000005300000000",
            INIT_2D => X"0000003300000000000000220000000000000023000000000000002000000000",
            INIT_2E => X"00000070000000000000003e000000000000002b000000000000002800000000",
            INIT_2F => X"0000001f000000000000004a000000000000009e000000000000009b00000000",
            INIT_30 => X"0000005a000000000000004f0000000000000068000000000000007000000000",
            INIT_31 => X"0000004200000000000000730000000000000089000000000000007b00000000",
            INIT_32 => X"0000001700000000000000280000000000000042000000000000002f00000000",
            INIT_33 => X"00000045000000000000002c0000000000000026000000000000001b00000000",
            INIT_34 => X"0000001d0000000000000026000000000000001f000000000000003600000000",
            INIT_35 => X"0000001f000000000000000f0000000000000016000000000000001900000000",
            INIT_36 => X"0000004e000000000000003a0000000000000033000000000000003100000000",
            INIT_37 => X"0000001f00000000000000570000000000000094000000000000008600000000",
            INIT_38 => X"0000006000000000000000590000000000000058000000000000006d00000000",
            INIT_39 => X"0000005e00000000000000730000000000000081000000000000006900000000",
            INIT_3A => X"0000003c00000000000000360000000000000047000000000000006100000000",
            INIT_3B => X"0000003c000000000000004b000000000000003e000000000000004200000000",
            INIT_3C => X"0000000e0000000000000009000000000000000a000000000000001a00000000",
            INIT_3D => X"0000000c000000000000000b0000000000000013000000000000001100000000",
            INIT_3E => X"0000003b000000000000003a000000000000001f000000000000001700000000",
            INIT_3F => X"0000002300000000000000690000000000000088000000000000005e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007000000000000000600000000000000046000000000000005b00000000",
            INIT_41 => X"0000009300000000000000890000000000000068000000000000006000000000",
            INIT_42 => X"000000430000000000000045000000000000003a000000000000007500000000",
            INIT_43 => X"00000035000000000000003f0000000000000045000000000000004a00000000",
            INIT_44 => X"0000000d00000000000000130000000000000019000000000000002900000000",
            INIT_45 => X"00000012000000000000000d0000000000000009000000000000000c00000000",
            INIT_46 => X"00000027000000000000003e0000000000000024000000000000000c00000000",
            INIT_47 => X"0000004700000000000000790000000000000068000000000000003400000000",
            INIT_48 => X"000000620000000000000062000000000000005c000000000000005b00000000",
            INIT_49 => X"0000008600000000000000690000000000000056000000000000006100000000",
            INIT_4A => X"00000061000000000000007c000000000000006b000000000000008e00000000",
            INIT_4B => X"00000049000000000000004e0000000000000049000000000000004400000000",
            INIT_4C => X"0000001c0000000000000026000000000000002b000000000000003e00000000",
            INIT_4D => X"00000014000000000000000b000000000000000e000000000000001600000000",
            INIT_4E => X"000000140000000000000030000000000000002a000000000000001400000000",
            INIT_4F => X"0000006400000000000000580000000000000038000000000000002500000000",
            INIT_50 => X"000000620000000000000061000000000000005e000000000000005b00000000",
            INIT_51 => X"0000004c000000000000005b000000000000006f000000000000007100000000",
            INIT_52 => X"000000510000000000000050000000000000006e000000000000008400000000",
            INIT_53 => X"000000540000000000000063000000000000005f000000000000004700000000",
            INIT_54 => X"000000330000000000000038000000000000003d000000000000004800000000",
            INIT_55 => X"0000002b0000000000000020000000000000002b000000000000003500000000",
            INIT_56 => X"0000002800000000000000250000000000000028000000000000002e00000000",
            INIT_57 => X"000000420000000000000030000000000000005a000000000000004000000000",
            INIT_58 => X"0000005200000000000000500000000000000060000000000000005700000000",
            INIT_59 => X"000000480000000000000062000000000000006d000000000000007100000000",
            INIT_5A => X"0000004600000000000000450000000000000073000000000000005c00000000",
            INIT_5B => X"000000580000000000000060000000000000005e000000000000004a00000000",
            INIT_5C => X"0000004a000000000000004c0000000000000047000000000000004500000000",
            INIT_5D => X"0000004b000000000000003d000000000000003c000000000000004200000000",
            INIT_5E => X"00000041000000000000003f0000000000000040000000000000004900000000",
            INIT_5F => X"0000003a0000000000000036000000000000005e000000000000004c00000000",
            INIT_60 => X"0000004c00000000000000430000000000000061000000000000006000000000",
            INIT_61 => X"00000050000000000000004e000000000000005a000000000000006900000000",
            INIT_62 => X"00000062000000000000004c0000000000000048000000000000005700000000",
            INIT_63 => X"0000005a000000000000005d000000000000005c000000000000005700000000",
            INIT_64 => X"0000004600000000000000550000000000000054000000000000004f00000000",
            INIT_65 => X"00000057000000000000004d0000000000000048000000000000004200000000",
            INIT_66 => X"0000004f00000000000000500000000000000052000000000000005300000000",
            INIT_67 => X"0000005e00000000000000460000000000000035000000000000004300000000",
            INIT_68 => X"0000006500000000000000510000000000000054000000000000004900000000",
            INIT_69 => X"0000005b0000000000000058000000000000005b000000000000006100000000",
            INIT_6A => X"00000063000000000000005b0000000000000059000000000000006900000000",
            INIT_6B => X"0000005a000000000000005d000000000000005d000000000000005900000000",
            INIT_6C => X"0000003c00000000000000490000000000000055000000000000005800000000",
            INIT_6D => X"0000005b00000000000000540000000000000052000000000000004900000000",
            INIT_6E => X"0000005500000000000000570000000000000056000000000000005d00000000",
            INIT_6F => X"0000006400000000000000570000000000000044000000000000004300000000",
            INIT_70 => X"00000071000000000000006a0000000000000060000000000000005300000000",
            INIT_71 => X"0000005f0000000000000060000000000000005f000000000000006000000000",
            INIT_72 => X"00000068000000000000006d0000000000000069000000000000006600000000",
            INIT_73 => X"0000004a0000000000000052000000000000005a000000000000005b00000000",
            INIT_74 => X"0000004a000000000000004d000000000000004e000000000000005200000000",
            INIT_75 => X"0000005c00000000000000570000000000000055000000000000004d00000000",
            INIT_76 => X"00000054000000000000005a0000000000000059000000000000006400000000",
            INIT_77 => X"0000005a0000000000000057000000000000004d000000000000004e00000000",
            INIT_78 => X"000000680000000000000071000000000000006b000000000000005c00000000",
            INIT_79 => X"0000005c000000000000004d0000000000000042000000000000005200000000",
            INIT_7A => X"0000005a000000000000005b0000000000000051000000000000005f00000000",
            INIT_7B => X"0000003d000000000000004d000000000000005b000000000000005800000000",
            INIT_7C => X"000000520000000000000056000000000000004d000000000000004600000000",
            INIT_7D => X"00000060000000000000005b000000000000005c000000000000005300000000",
            INIT_7E => X"0000005b0000000000000057000000000000005c000000000000006500000000",
            INIT_7F => X"00000057000000000000005b000000000000005a000000000000005c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "sampleifmap_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000024000000000000001a000000000000003d000000000000005300000000",
            INIT_01 => X"00000036000000000000003a0000000000000043000000000000004100000000",
            INIT_02 => X"0000003b00000000000000340000000000000041000000000000003f00000000",
            INIT_03 => X"00000034000000000000002e0000000000000035000000000000003e00000000",
            INIT_04 => X"00000027000000000000002b0000000000000041000000000000004700000000",
            INIT_05 => X"00000026000000000000002d000000000000002f000000000000002f00000000",
            INIT_06 => X"00000032000000000000002a000000000000002d000000000000002f00000000",
            INIT_07 => X"000000290000000000000029000000000000002e000000000000004500000000",
            INIT_08 => X"00000046000000000000003a0000000000000035000000000000006100000000",
            INIT_09 => X"0000004d00000000000000440000000000000043000000000000004600000000",
            INIT_0A => X"0000003900000000000000380000000000000041000000000000004400000000",
            INIT_0B => X"0000002e00000000000000320000000000000039000000000000003400000000",
            INIT_0C => X"00000026000000000000002b0000000000000034000000000000003c00000000",
            INIT_0D => X"00000028000000000000002c000000000000002f000000000000002f00000000",
            INIT_0E => X"00000038000000000000002b000000000000001e000000000000002000000000",
            INIT_0F => X"0000003100000000000000330000000000000035000000000000004300000000",
            INIT_10 => X"00000051000000000000005c0000000000000047000000000000006400000000",
            INIT_11 => X"0000004e00000000000000440000000000000039000000000000004400000000",
            INIT_12 => X"0000003b000000000000003f0000000000000047000000000000004000000000",
            INIT_13 => X"0000003000000000000000310000000000000030000000000000003400000000",
            INIT_14 => X"0000001e00000000000000210000000000000032000000000000003b00000000",
            INIT_15 => X"0000003800000000000000350000000000000030000000000000002b00000000",
            INIT_16 => X"0000003800000000000000390000000000000038000000000000003300000000",
            INIT_17 => X"00000031000000000000002f0000000000000035000000000000003900000000",
            INIT_18 => X"000000590000000000000061000000000000005f000000000000006000000000",
            INIT_19 => X"0000004800000000000000490000000000000037000000000000004900000000",
            INIT_1A => X"000000420000000000000042000000000000004e000000000000004100000000",
            INIT_1B => X"0000003f00000000000000360000000000000037000000000000004300000000",
            INIT_1C => X"00000012000000000000001a000000000000002e000000000000002f00000000",
            INIT_1D => X"00000035000000000000002f0000000000000029000000000000002200000000",
            INIT_1E => X"0000003e00000000000000400000000000000044000000000000003d00000000",
            INIT_1F => X"0000003c000000000000003a000000000000002d000000000000003000000000",
            INIT_20 => X"0000005700000000000000540000000000000061000000000000005c00000000",
            INIT_21 => X"0000004b000000000000004c000000000000003f000000000000004900000000",
            INIT_22 => X"0000004b000000000000004b000000000000004a000000000000004a00000000",
            INIT_23 => X"0000003b0000000000000035000000000000003b000000000000004300000000",
            INIT_24 => X"0000001e00000000000000330000000000000034000000000000003b00000000",
            INIT_25 => X"00000027000000000000002e0000000000000029000000000000001f00000000",
            INIT_26 => X"0000003d000000000000003d000000000000003b000000000000002e00000000",
            INIT_27 => X"0000003c000000000000003a0000000000000030000000000000003400000000",
            INIT_28 => X"0000005900000000000000470000000000000066000000000000006500000000",
            INIT_29 => X"0000004c000000000000004c0000000000000046000000000000005100000000",
            INIT_2A => X"00000047000000000000004e0000000000000051000000000000004c00000000",
            INIT_2B => X"0000003100000000000000350000000000000043000000000000004400000000",
            INIT_2C => X"0000003900000000000000480000000000000041000000000000004300000000",
            INIT_2D => X"000000320000000000000042000000000000003e000000000000002b00000000",
            INIT_2E => X"0000003a00000000000000380000000000000036000000000000003800000000",
            INIT_2F => X"00000041000000000000003c000000000000003d000000000000003c00000000",
            INIT_30 => X"0000006300000000000000490000000000000059000000000000007800000000",
            INIT_31 => X"0000004b00000000000000510000000000000050000000000000005300000000",
            INIT_32 => X"0000004200000000000000550000000000000057000000000000005100000000",
            INIT_33 => X"000000350000000000000043000000000000004f000000000000004c00000000",
            INIT_34 => X"0000004d000000000000004a0000000000000040000000000000003c00000000",
            INIT_35 => X"0000002f00000000000000410000000000000040000000000000004100000000",
            INIT_36 => X"00000030000000000000002d0000000000000036000000000000003500000000",
            INIT_37 => X"00000042000000000000003f000000000000003d000000000000003a00000000",
            INIT_38 => X"0000005b000000000000005b000000000000003b000000000000007500000000",
            INIT_39 => X"00000054000000000000004f0000000000000051000000000000005100000000",
            INIT_3A => X"0000004800000000000000560000000000000056000000000000005700000000",
            INIT_3B => X"0000003f000000000000004a000000000000004c000000000000004d00000000",
            INIT_3C => X"00000049000000000000004c0000000000000049000000000000004200000000",
            INIT_3D => X"0000002f0000000000000038000000000000002f000000000000004700000000",
            INIT_3E => X"0000002a00000000000000230000000000000031000000000000002c00000000",
            INIT_3F => X"00000040000000000000003e0000000000000039000000000000003700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000051000000000000005b0000000000000054000000000000005c00000000",
            INIT_41 => X"000000500000000000000050000000000000004f000000000000005300000000",
            INIT_42 => X"0000004600000000000000490000000000000053000000000000005800000000",
            INIT_43 => X"0000003d00000000000000430000000000000048000000000000005100000000",
            INIT_44 => X"0000004600000000000000460000000000000041000000000000004300000000",
            INIT_45 => X"0000003c000000000000004f0000000000000040000000000000004f00000000",
            INIT_46 => X"0000003b0000000000000034000000000000002d000000000000002c00000000",
            INIT_47 => X"00000040000000000000003d000000000000003d000000000000003a00000000",
            INIT_48 => X"0000005a000000000000004c0000000000000058000000000000006100000000",
            INIT_49 => X"0000004700000000000000530000000000000056000000000000005b00000000",
            INIT_4A => X"0000005300000000000000540000000000000052000000000000004f00000000",
            INIT_4B => X"00000055000000000000004d0000000000000053000000000000005800000000",
            INIT_4C => X"000000460000000000000039000000000000003e000000000000005100000000",
            INIT_4D => X"0000004b00000000000000590000000000000048000000000000005000000000",
            INIT_4E => X"0000003c000000000000003a0000000000000031000000000000002b00000000",
            INIT_4F => X"000000400000000000000039000000000000003f000000000000003a00000000",
            INIT_50 => X"0000006200000000000000560000000000000030000000000000005100000000",
            INIT_51 => X"000000540000000000000052000000000000005b000000000000005900000000",
            INIT_52 => X"0000005000000000000000500000000000000054000000000000005b00000000",
            INIT_53 => X"0000007e00000000000000670000000000000065000000000000005e00000000",
            INIT_54 => X"0000004300000000000000370000000000000049000000000000006b00000000",
            INIT_55 => X"000000440000000000000051000000000000004c000000000000004b00000000",
            INIT_56 => X"0000002d000000000000002f0000000000000031000000000000002000000000",
            INIT_57 => X"00000041000000000000003e000000000000003a000000000000003300000000",
            INIT_58 => X"0000004d0000000000000063000000000000001f000000000000001400000000",
            INIT_59 => X"0000005a000000000000005a0000000000000056000000000000004000000000",
            INIT_5A => X"0000005f00000000000000450000000000000045000000000000005f00000000",
            INIT_5B => X"0000007900000000000000670000000000000088000000000000008f00000000",
            INIT_5C => X"00000050000000000000003f0000000000000052000000000000007600000000",
            INIT_5D => X"000000210000000000000042000000000000004d000000000000005200000000",
            INIT_5E => X"0000002e00000000000000300000000000000030000000000000002100000000",
            INIT_5F => X"0000003f000000000000003b0000000000000036000000000000003000000000",
            INIT_60 => X"0000005c00000000000000700000000000000032000000000000000000000000",
            INIT_61 => X"000000620000000000000069000000000000007a000000000000006e00000000",
            INIT_62 => X"0000007700000000000000540000000000000048000000000000006000000000",
            INIT_63 => X"00000049000000000000005f000000000000007d000000000000009d00000000",
            INIT_64 => X"0000005400000000000000410000000000000047000000000000003400000000",
            INIT_65 => X"0000002a0000000000000041000000000000004f000000000000006000000000",
            INIT_66 => X"0000002900000000000000290000000000000025000000000000002500000000",
            INIT_67 => X"0000003a00000000000000390000000000000038000000000000002d00000000",
            INIT_68 => X"0000005c0000000000000061000000000000003c000000000000001400000000",
            INIT_69 => X"0000006f00000000000000700000000000000078000000000000007d00000000",
            INIT_6A => X"00000080000000000000006e000000000000004c000000000000005900000000",
            INIT_6B => X"0000006c00000000000000620000000000000064000000000000007f00000000",
            INIT_6C => X"0000005b00000000000000620000000000000063000000000000004400000000",
            INIT_6D => X"00000029000000000000003a000000000000004c000000000000006a00000000",
            INIT_6E => X"0000002600000000000000250000000000000023000000000000002100000000",
            INIT_6F => X"0000003500000000000000320000000000000034000000000000002e00000000",
            INIT_70 => X"00000058000000000000003a0000000000000046000000000000003b00000000",
            INIT_71 => X"00000073000000000000006a0000000000000075000000000000007b00000000",
            INIT_72 => X"0000007d00000000000000820000000000000067000000000000006600000000",
            INIT_73 => X"0000008900000000000000660000000000000050000000000000005f00000000",
            INIT_74 => X"00000084000000000000007e000000000000008c000000000000008300000000",
            INIT_75 => X"0000002a0000000000000040000000000000004e000000000000006f00000000",
            INIT_76 => X"00000032000000000000002a0000000000000028000000000000002b00000000",
            INIT_77 => X"00000031000000000000002e0000000000000032000000000000002f00000000",
            INIT_78 => X"0000005e00000000000000320000000000000035000000000000004900000000",
            INIT_79 => X"00000062000000000000006c000000000000007c000000000000007e00000000",
            INIT_7A => X"00000088000000000000008a000000000000007d000000000000007200000000",
            INIT_7B => X"0000008c00000000000000710000000000000062000000000000007b00000000",
            INIT_7C => X"0000008c000000000000008a0000000000000089000000000000008f00000000",
            INIT_7D => X"0000003300000000000000490000000000000069000000000000007500000000",
            INIT_7E => X"0000004d00000000000000320000000000000023000000000000002f00000000",
            INIT_7F => X"00000032000000000000002d000000000000002d000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "sampleifmap_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000056000000000000003a0000000000000041000000000000004800000000",
            INIT_01 => X"0000005300000000000000690000000000000075000000000000007700000000",
            INIT_02 => X"0000008200000000000000930000000000000089000000000000006e00000000",
            INIT_03 => X"00000087000000000000006d000000000000006b000000000000008200000000",
            INIT_04 => X"00000083000000000000007e000000000000007f000000000000008400000000",
            INIT_05 => X"0000002a000000000000003d0000000000000077000000000000008700000000",
            INIT_06 => X"00000055000000000000003c000000000000001b000000000000001a00000000",
            INIT_07 => X"0000003300000000000000240000000000000033000000000000006100000000",
            INIT_08 => X"0000006600000000000000510000000000000048000000000000004700000000",
            INIT_09 => X"00000050000000000000007a000000000000007c000000000000007800000000",
            INIT_0A => X"00000054000000000000006a0000000000000097000000000000006300000000",
            INIT_0B => X"0000005c00000000000000650000000000000079000000000000007c00000000",
            INIT_0C => X"0000006500000000000000680000000000000073000000000000006300000000",
            INIT_0D => X"00000011000000000000001f0000000000000048000000000000005e00000000",
            INIT_0E => X"00000055000000000000003a0000000000000015000000000000000e00000000",
            INIT_0F => X"00000029000000000000001f0000000000000046000000000000006800000000",
            INIT_10 => X"000000640000000000000044000000000000004e000000000000004f00000000",
            INIT_11 => X"0000004b000000000000007d0000000000000088000000000000008600000000",
            INIT_12 => X"00000061000000000000005b0000000000000093000000000000004700000000",
            INIT_13 => X"0000004800000000000000370000000000000071000000000000008e00000000",
            INIT_14 => X"000000320000000000000045000000000000004f000000000000003500000000",
            INIT_15 => X"00000016000000000000000d0000000000000014000000000000002a00000000",
            INIT_16 => X"0000006000000000000000370000000000000023000000000000001400000000",
            INIT_17 => X"00000023000000000000001e000000000000005b000000000000006f00000000",
            INIT_18 => X"0000005800000000000000320000000000000048000000000000005100000000",
            INIT_19 => X"0000005d000000000000008a0000000000000099000000000000008700000000",
            INIT_1A => X"00000071000000000000007f000000000000006f000000000000001f00000000",
            INIT_1B => X"0000008d0000000000000047000000000000005c000000000000007c00000000",
            INIT_1C => X"0000002100000000000000330000000000000041000000000000006700000000",
            INIT_1D => X"0000002c00000000000000240000000000000019000000000000002400000000",
            INIT_1E => X"000000600000000000000036000000000000002b000000000000001a00000000",
            INIT_1F => X"0000001a000000000000001e0000000000000073000000000000008900000000",
            INIT_20 => X"0000005f000000000000004f0000000000000052000000000000005300000000",
            INIT_21 => X"0000006200000000000000860000000000000096000000000000008200000000",
            INIT_22 => X"0000006300000000000000560000000000000017000000000000000a00000000",
            INIT_23 => X"000000740000000000000042000000000000004c000000000000006500000000",
            INIT_24 => X"000000170000000000000027000000000000004e000000000000007a00000000",
            INIT_25 => X"0000002e000000000000002f000000000000002f000000000000002e00000000",
            INIT_26 => X"000000670000000000000034000000000000001b000000000000001400000000",
            INIT_27 => X"00000019000000000000002f0000000000000089000000000000009200000000",
            INIT_28 => X"00000053000000000000004e000000000000005c000000000000005c00000000",
            INIT_29 => X"00000046000000000000006e0000000000000087000000000000007b00000000",
            INIT_2A => X"0000001d00000000000000100000000000000008000000000000000c00000000",
            INIT_2B => X"0000003800000000000000250000000000000034000000000000002f00000000",
            INIT_2C => X"00000012000000000000002b0000000000000039000000000000004600000000",
            INIT_2D => X"0000002c000000000000001d000000000000001c000000000000001900000000",
            INIT_2E => X"0000005e00000000000000310000000000000026000000000000002100000000",
            INIT_2F => X"00000018000000000000003d000000000000008d000000000000008c00000000",
            INIT_30 => X"0000004e0000000000000046000000000000005d000000000000006100000000",
            INIT_31 => X"0000003000000000000000600000000000000076000000000000006b00000000",
            INIT_32 => X"000000130000000000000022000000000000003a000000000000002500000000",
            INIT_33 => X"0000003b0000000000000026000000000000001f000000000000001300000000",
            INIT_34 => X"00000012000000000000001b0000000000000013000000000000002700000000",
            INIT_35 => X"00000018000000000000000a0000000000000011000000000000001100000000",
            INIT_36 => X"000000400000000000000030000000000000002c000000000000002a00000000",
            INIT_37 => X"0000001800000000000000460000000000000080000000000000007800000000",
            INIT_38 => X"000000580000000000000052000000000000004d000000000000005e00000000",
            INIT_39 => X"0000004b000000000000005f000000000000006b000000000000005b00000000",
            INIT_3A => X"0000003900000000000000300000000000000037000000000000004a00000000",
            INIT_3B => X"0000003300000000000000430000000000000035000000000000003a00000000",
            INIT_3C => X"0000000800000000000000030000000000000004000000000000001000000000",
            INIT_3D => X"0000000600000000000000070000000000000013000000000000000e00000000",
            INIT_3E => X"0000002f00000000000000300000000000000017000000000000001100000000",
            INIT_3F => X"0000001b00000000000000570000000000000073000000000000005100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000690000000000000057000000000000003b000000000000004b00000000",
            INIT_41 => X"0000007e00000000000000750000000000000052000000000000005300000000",
            INIT_42 => X"0000003e00000000000000390000000000000022000000000000005500000000",
            INIT_43 => X"0000002e0000000000000039000000000000003d000000000000004200000000",
            INIT_44 => X"0000000d00000000000000120000000000000017000000000000002400000000",
            INIT_45 => X"0000000e000000000000000c000000000000000e000000000000000f00000000",
            INIT_46 => X"0000001e0000000000000036000000000000001c000000000000000700000000",
            INIT_47 => X"0000003e00000000000000680000000000000055000000000000002800000000",
            INIT_48 => X"000000560000000000000051000000000000004d000000000000004d00000000",
            INIT_49 => X"0000007000000000000000570000000000000045000000000000005500000000",
            INIT_4A => X"0000004f0000000000000064000000000000004f000000000000006f00000000",
            INIT_4B => X"0000003a00000000000000450000000000000043000000000000003b00000000",
            INIT_4C => X"0000001500000000000000200000000000000026000000000000003300000000",
            INIT_4D => X"0000000e0000000000000006000000000000000c000000000000001100000000",
            INIT_4E => X"0000000f00000000000000290000000000000022000000000000000f00000000",
            INIT_4F => X"0000005a000000000000004c000000000000002e000000000000001f00000000",
            INIT_50 => X"0000005500000000000000520000000000000051000000000000004f00000000",
            INIT_51 => X"00000039000000000000004a0000000000000060000000000000006500000000",
            INIT_52 => X"0000003e000000000000003a0000000000000057000000000000006d00000000",
            INIT_53 => X"00000044000000000000005a0000000000000058000000000000003d00000000",
            INIT_54 => X"0000002a000000000000002f0000000000000035000000000000003b00000000",
            INIT_55 => X"0000002300000000000000180000000000000023000000000000002c00000000",
            INIT_56 => X"0000001f000000000000001b000000000000001d000000000000002600000000",
            INIT_57 => X"0000003800000000000000270000000000000052000000000000003900000000",
            INIT_58 => X"0000004a000000000000004a0000000000000057000000000000004c00000000",
            INIT_59 => X"000000390000000000000053000000000000005f000000000000006600000000",
            INIT_5A => X"0000003a00000000000000370000000000000063000000000000004d00000000",
            INIT_5B => X"0000004d00000000000000570000000000000054000000000000003f00000000",
            INIT_5C => X"000000440000000000000043000000000000003c000000000000003900000000",
            INIT_5D => X"0000003f00000000000000310000000000000031000000000000003b00000000",
            INIT_5E => X"0000003300000000000000300000000000000031000000000000003c00000000",
            INIT_5F => X"0000002f000000000000002d0000000000000054000000000000003f00000000",
            INIT_60 => X"000000450000000000000040000000000000005a000000000000005500000000",
            INIT_61 => X"000000440000000000000041000000000000004e000000000000005e00000000",
            INIT_62 => X"0000005a0000000000000042000000000000003c000000000000004c00000000",
            INIT_63 => X"000000510000000000000053000000000000004e000000000000004a00000000",
            INIT_64 => X"00000040000000000000004c0000000000000047000000000000004300000000",
            INIT_65 => X"00000048000000000000003e0000000000000039000000000000003b00000000",
            INIT_66 => X"0000003e00000000000000400000000000000042000000000000004400000000",
            INIT_67 => X"00000053000000000000003d0000000000000029000000000000003200000000",
            INIT_68 => X"0000005c0000000000000049000000000000004b000000000000003d00000000",
            INIT_69 => X"00000050000000000000004e0000000000000051000000000000005700000000",
            INIT_6A => X"000000590000000000000050000000000000004c000000000000005d00000000",
            INIT_6B => X"00000050000000000000004e000000000000004c000000000000004a00000000",
            INIT_6C => X"00000035000000000000003e0000000000000045000000000000004a00000000",
            INIT_6D => X"0000004b00000000000000440000000000000042000000000000004000000000",
            INIT_6E => X"0000004400000000000000480000000000000048000000000000004d00000000",
            INIT_6F => X"00000059000000000000004e0000000000000038000000000000003200000000",
            INIT_70 => X"00000064000000000000005a0000000000000051000000000000004600000000",
            INIT_71 => X"0000005500000000000000570000000000000055000000000000005600000000",
            INIT_72 => X"0000005a000000000000005d0000000000000057000000000000005600000000",
            INIT_73 => X"0000003c000000000000003f0000000000000046000000000000004a00000000",
            INIT_74 => X"0000003e000000000000003e000000000000003c000000000000004200000000",
            INIT_75 => X"0000004c00000000000000470000000000000046000000000000004100000000",
            INIT_76 => X"00000047000000000000004e000000000000004d000000000000005500000000",
            INIT_77 => X"0000004f000000000000004d0000000000000041000000000000003e00000000",
            INIT_78 => X"00000059000000000000005f000000000000005d000000000000004f00000000",
            INIT_79 => X"0000005100000000000000460000000000000039000000000000004600000000",
            INIT_7A => X"0000004700000000000000470000000000000040000000000000005300000000",
            INIT_7B => X"0000002f000000000000003d000000000000004c000000000000004a00000000",
            INIT_7C => X"000000460000000000000048000000000000003f000000000000003800000000",
            INIT_7D => X"00000050000000000000004b000000000000004c000000000000004500000000",
            INIT_7E => X"0000004e0000000000000049000000000000004f000000000000005600000000",
            INIT_7F => X"00000049000000000000004f000000000000004c000000000000004f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "sampleifmap_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000d900000000000000d100000000000000b900000000000000a000000000",
            INIT_01 => X"000000f600000000000000f900000000000000f600000000000000e600000000",
            INIT_02 => X"000000dd00000000000000e600000000000000f300000000000000f800000000",
            INIT_03 => X"000000c700000000000000d800000000000000dd00000000000000da00000000",
            INIT_04 => X"000000b400000000000000b800000000000000bb00000000000000bc00000000",
            INIT_05 => X"0000008b0000000000000079000000000000009000000000000000a600000000",
            INIT_06 => X"0000004f00000000000000660000000000000066000000000000006a00000000",
            INIT_07 => X"0000005e000000000000005b0000000000000065000000000000005e00000000",
            INIT_08 => X"000000e600000000000000f200000000000000ef00000000000000e100000000",
            INIT_09 => X"000000eb00000000000000f300000000000000f500000000000000e800000000",
            INIT_0A => X"000000cd00000000000000d800000000000000e600000000000000ed00000000",
            INIT_0B => X"000000ba00000000000000c800000000000000cb00000000000000c900000000",
            INIT_0C => X"0000007f00000000000000a100000000000000ab00000000000000af00000000",
            INIT_0D => X"00000087000000000000007a000000000000008d000000000000008e00000000",
            INIT_0E => X"0000003400000000000000250000000000000052000000000000007600000000",
            INIT_0F => X"000000640000000000000061000000000000006b000000000000005f00000000",
            INIT_10 => X"000000dc00000000000000f100000000000000f900000000000000fc00000000",
            INIT_11 => X"000000d600000000000000df00000000000000e200000000000000d900000000",
            INIT_12 => X"000000b800000000000000c300000000000000cf00000000000000d500000000",
            INIT_13 => X"000000a700000000000000b300000000000000b600000000000000b300000000",
            INIT_14 => X"0000008100000000000000940000000000000098000000000000009f00000000",
            INIT_15 => X"000000720000000000000080000000000000008c000000000000008000000000",
            INIT_16 => X"0000002600000000000000040000000000000028000000000000005700000000",
            INIT_17 => X"0000006900000000000000690000000000000073000000000000006300000000",
            INIT_18 => X"000000d300000000000000de00000000000000e100000000000000e900000000",
            INIT_19 => X"000000c000000000000000c800000000000000cb00000000000000d300000000",
            INIT_1A => X"000000a400000000000000ae00000000000000b700000000000000bb00000000",
            INIT_1B => X"0000009900000000000000a000000000000000a500000000000000a000000000",
            INIT_1C => X"0000008a000000000000008c000000000000008d000000000000009100000000",
            INIT_1D => X"00000069000000000000007f000000000000007d000000000000007d00000000",
            INIT_1E => X"00000037000000000000001a0000000000000025000000000000003b00000000",
            INIT_1F => X"0000006d00000000000000700000000000000078000000000000007000000000",
            INIT_20 => X"000000c900000000000000cf00000000000000c300000000000000cf00000000",
            INIT_21 => X"000000ab00000000000000b300000000000000b400000000000000be00000000",
            INIT_22 => X"000000920000000000000099000000000000009f00000000000000a300000000",
            INIT_23 => X"0000008d00000000000000930000000000000097000000000000009100000000",
            INIT_24 => X"0000008700000000000000830000000000000088000000000000008700000000",
            INIT_25 => X"0000005a0000000000000084000000000000007a000000000000008100000000",
            INIT_26 => X"000000560000000000000030000000000000003d000000000000003a00000000",
            INIT_27 => X"0000006d00000000000000720000000000000078000000000000007500000000",
            INIT_28 => X"000000a200000000000000aa00000000000000ab00000000000000b600000000",
            INIT_29 => X"00000097000000000000009f000000000000009c000000000000009900000000",
            INIT_2A => X"0000008a000000000000008c000000000000008d000000000000009000000000",
            INIT_2B => X"0000008a000000000000008a000000000000008d000000000000008b00000000",
            INIT_2C => X"0000008a0000000000000086000000000000008c000000000000008700000000",
            INIT_2D => X"0000004500000000000000660000000000000089000000000000008c00000000",
            INIT_2E => X"000000740000000000000043000000000000003e000000000000004b00000000",
            INIT_2F => X"0000006e00000000000000700000000000000080000000000000008100000000",
            INIT_30 => X"0000008600000000000000880000000000000088000000000000008d00000000",
            INIT_31 => X"00000085000000000000008c0000000000000086000000000000008800000000",
            INIT_32 => X"0000008d000000000000008b0000000000000089000000000000008700000000",
            INIT_33 => X"00000091000000000000008e0000000000000092000000000000008f00000000",
            INIT_34 => X"0000008f000000000000008a0000000000000091000000000000009100000000",
            INIT_35 => X"00000021000000000000002f000000000000006b000000000000008e00000000",
            INIT_36 => X"0000007f000000000000006c000000000000004b000000000000004800000000",
            INIT_37 => X"00000070000000000000006f0000000000000084000000000000008400000000",
            INIT_38 => X"000000810000000000000080000000000000007d000000000000007600000000",
            INIT_39 => X"00000084000000000000008a0000000000000083000000000000008800000000",
            INIT_3A => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_3B => X"00000099000000000000009a000000000000009e000000000000009600000000",
            INIT_3C => X"0000009400000000000000930000000000000095000000000000009200000000",
            INIT_3D => X"00000011000000000000000d0000000000000042000000000000008000000000",
            INIT_3E => X"0000007a00000000000000800000000000000075000000000000005000000000",
            INIT_3F => X"0000007000000000000000720000000000000080000000000000007b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000850000000000000084000000000000007e000000000000007300000000",
            INIT_41 => X"00000089000000000000008f0000000000000087000000000000008b00000000",
            INIT_42 => X"0000009800000000000000950000000000000091000000000000008b00000000",
            INIT_43 => X"000000aa00000000000000a3000000000000009a000000000000009400000000",
            INIT_44 => X"00000094000000000000009d00000000000000a2000000000000009e00000000",
            INIT_45 => X"0000001e000000000000000e000000000000002c000000000000007300000000",
            INIT_46 => X"0000007e0000000000000088000000000000008b000000000000006900000000",
            INIT_47 => X"0000006f0000000000000074000000000000007a000000000000007700000000",
            INIT_48 => X"0000008800000000000000880000000000000080000000000000007600000000",
            INIT_49 => X"0000008d00000000000000910000000000000088000000000000008d00000000",
            INIT_4A => X"000000a5000000000000009a0000000000000093000000000000008d00000000",
            INIT_4B => X"000000a700000000000000a2000000000000009a000000000000009d00000000",
            INIT_4C => X"0000008a00000000000000910000000000000093000000000000009b00000000",
            INIT_4D => X"00000037000000000000002e0000000000000038000000000000006300000000",
            INIT_4E => X"0000007e000000000000007a000000000000007c000000000000006d00000000",
            INIT_4F => X"0000006e00000000000000750000000000000074000000000000007300000000",
            INIT_50 => X"00000089000000000000008b0000000000000084000000000000007d00000000",
            INIT_51 => X"0000008c00000000000000900000000000000088000000000000008e00000000",
            INIT_52 => X"0000009900000000000000960000000000000090000000000000008b00000000",
            INIT_53 => X"000000980000000000000090000000000000008b000000000000008300000000",
            INIT_54 => X"000000d600000000000000d300000000000000ba00000000000000a600000000",
            INIT_55 => X"0000002a0000000000000045000000000000005c000000000000008000000000",
            INIT_56 => X"000000730000000000000063000000000000005f000000000000005500000000",
            INIT_57 => X"0000006b0000000000000071000000000000006f000000000000007000000000",
            INIT_58 => X"0000008a000000000000008e0000000000000089000000000000008500000000",
            INIT_59 => X"0000008a000000000000008e0000000000000088000000000000008d00000000",
            INIT_5A => X"000000840000000000000088000000000000008f000000000000008900000000",
            INIT_5B => X"000000cb00000000000000c900000000000000b6000000000000008e00000000",
            INIT_5C => X"000000c000000000000000cf00000000000000ce00000000000000d200000000",
            INIT_5D => X"0000002a000000000000009200000000000000bd00000000000000a200000000",
            INIT_5E => X"0000007200000000000000670000000000000028000000000000001b00000000",
            INIT_5F => X"00000068000000000000006c000000000000006a000000000000006d00000000",
            INIT_60 => X"0000008b000000000000008f000000000000008b000000000000008c00000000",
            INIT_61 => X"00000089000000000000008a000000000000008c000000000000008f00000000",
            INIT_62 => X"000000a400000000000000900000000000000085000000000000008700000000",
            INIT_63 => X"00000073000000000000008900000000000000a000000000000000ab00000000",
            INIT_64 => X"0000003b000000000000004b000000000000005d000000000000006a00000000",
            INIT_65 => X"0000005f00000000000000c900000000000000dc000000000000006f00000000",
            INIT_66 => X"00000074000000000000003e0000000000000007000000000000000d00000000",
            INIT_67 => X"0000006400000000000000690000000000000065000000000000006300000000",
            INIT_68 => X"0000008c000000000000008f000000000000008a000000000000009000000000",
            INIT_69 => X"0000008700000000000000820000000000000092000000000000009200000000",
            INIT_6A => X"0000006e000000000000008c0000000000000091000000000000008200000000",
            INIT_6B => X"000000130000000000000031000000000000005c000000000000005e00000000",
            INIT_6C => X"0000001200000000000000190000000000000032000000000000001d00000000",
            INIT_6D => X"0000009d00000000000000d200000000000000d1000000000000007800000000",
            INIT_6E => X"0000004400000000000000130000000000000006000000000000002600000000",
            INIT_6F => X"0000005f00000000000000630000000000000052000000000000004500000000",
            INIT_70 => X"0000008e0000000000000092000000000000008b000000000000009100000000",
            INIT_71 => X"000000800000000000000079000000000000008e000000000000009000000000",
            INIT_72 => X"000000440000000000000054000000000000007f000000000000008500000000",
            INIT_73 => X"00000016000000000000002e0000000000000052000000000000005600000000",
            INIT_74 => X"00000041000000000000001e0000000000000032000000000000001300000000",
            INIT_75 => X"000000cb00000000000000cd00000000000000c900000000000000af00000000",
            INIT_76 => X"0000001600000000000000120000000000000010000000000000006600000000",
            INIT_77 => X"00000058000000000000004f0000000000000038000000000000002300000000",
            INIT_78 => X"000000900000000000000094000000000000008b000000000000008f00000000",
            INIT_79 => X"00000083000000000000008b0000000000000084000000000000008a00000000",
            INIT_7A => X"0000005600000000000000480000000000000042000000000000007500000000",
            INIT_7B => X"000000220000000000000028000000000000004e000000000000006a00000000",
            INIT_7C => X"000000b600000000000000730000000000000046000000000000002400000000",
            INIT_7D => X"000000c300000000000000cd00000000000000c500000000000000cb00000000",
            INIT_7E => X"000000120000000000000025000000000000003d000000000000006c00000000",
            INIT_7F => X"000000530000000000000064000000000000004f000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "sampleifmap_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000900000000000000093000000000000008b000000000000008e00000000",
            INIT_01 => X"0000007900000000000000840000000000000072000000000000008500000000",
            INIT_02 => X"00000045000000000000003c0000000000000059000000000000005100000000",
            INIT_03 => X"0000009b00000000000000530000000000000044000000000000005500000000",
            INIT_04 => X"000000eb00000000000000ed00000000000000db00000000000000c000000000",
            INIT_05 => X"0000007200000000000000d300000000000000d700000000000000d700000000",
            INIT_06 => X"000000140000000000000035000000000000005d000000000000003000000000",
            INIT_07 => X"00000054000000000000008f000000000000008b000000000000004100000000",
            INIT_08 => X"00000089000000000000008e000000000000008d000000000000008f00000000",
            INIT_09 => X"00000043000000000000003a0000000000000045000000000000007400000000",
            INIT_0A => X"0000001c000000000000001d000000000000004b000000000000005100000000",
            INIT_0B => X"000000f2000000000000008c0000000000000019000000000000002400000000",
            INIT_0C => X"000000dc00000000000000e300000000000000eb00000000000000ec00000000",
            INIT_0D => X"0000003a000000000000009500000000000000df00000000000000db00000000",
            INIT_0E => X"0000004e000000000000004e0000000000000054000000000000003900000000",
            INIT_0F => X"0000005b00000000000000a700000000000000a1000000000000008500000000",
            INIT_10 => X"000000860000000000000088000000000000008c000000000000008f00000000",
            INIT_11 => X"00000034000000000000002d0000000000000047000000000000008d00000000",
            INIT_12 => X"0000001600000000000000170000000000000021000000000000004300000000",
            INIT_13 => X"000000d9000000000000009b0000000000000029000000000000002f00000000",
            INIT_14 => X"000000d000000000000000bf00000000000000be00000000000000c700000000",
            INIT_15 => X"0000006700000000000000ad00000000000000df00000000000000dc00000000",
            INIT_16 => X"0000009500000000000000870000000000000073000000000000005d00000000",
            INIT_17 => X"0000005900000000000000a50000000000000094000000000000009800000000",
            INIT_18 => X"000000b5000000000000007e000000000000008c000000000000008f00000000",
            INIT_19 => X"0000002b0000000000000021000000000000004c00000000000000bd00000000",
            INIT_1A => X"0000001700000000000000100000000000000015000000000000003900000000",
            INIT_1B => X"000000c2000000000000009e0000000000000042000000000000003900000000",
            INIT_1C => X"000000c900000000000000c400000000000000b300000000000000b600000000",
            INIT_1D => X"000000b300000000000000de00000000000000ce00000000000000c200000000",
            INIT_1E => X"000000970000000000000095000000000000009c000000000000009700000000",
            INIT_1F => X"0000004200000000000000880000000000000092000000000000009600000000",
            INIT_20 => X"000000ea000000000000009a0000000000000085000000000000008c00000000",
            INIT_21 => X"0000002a0000000000000026000000000000005a00000000000000b500000000",
            INIT_22 => X"0000000b000000000000000b000000000000000b000000000000003400000000",
            INIT_23 => X"000000ba00000000000000a00000000000000031000000000000001400000000",
            INIT_24 => X"0000007300000000000000b900000000000000b900000000000000b000000000",
            INIT_25 => X"000000c400000000000000a1000000000000005a000000000000004500000000",
            INIT_26 => X"0000009900000000000000a000000000000000aa00000000000000b700000000",
            INIT_27 => X"00000026000000000000004d0000000000000088000000000000009300000000",
            INIT_28 => X"000000a300000000000000a30000000000000080000000000000008200000000",
            INIT_29 => X"0000002e000000000000002d000000000000006a000000000000008b00000000",
            INIT_2A => X"0000000f00000000000000090000000000000003000000000000001c00000000",
            INIT_2B => X"000000b400000000000000a20000000000000036000000000000001e00000000",
            INIT_2C => X"00000015000000000000007100000000000000be00000000000000ac00000000",
            INIT_2D => X"0000009500000000000000300000000000000015000000000000001400000000",
            INIT_2E => X"00000085000000000000008e00000000000000ab00000000000000bb00000000",
            INIT_2F => X"0000002700000000000000150000000000000043000000000000008000000000",
            INIT_30 => X"0000001a00000000000000670000000000000084000000000000007c00000000",
            INIT_31 => X"000000300000000000000034000000000000006c000000000000004800000000",
            INIT_32 => X"0000003b000000000000000b0000000000000007000000000000001200000000",
            INIT_33 => X"000000b000000000000000a50000000000000063000000000000005a00000000",
            INIT_34 => X"0000001d000000000000002a00000000000000a900000000000000b100000000",
            INIT_35 => X"00000046000000000000000e0000000000000026000000000000002f00000000",
            INIT_36 => X"0000007500000000000000750000000000000088000000000000009500000000",
            INIT_37 => X"000000300000000000000015000000000000000e000000000000003c00000000",
            INIT_38 => X"0000001e0000000000000049000000000000007c000000000000007900000000",
            INIT_39 => X"0000001f00000000000000440000000000000072000000000000003b00000000",
            INIT_3A => X"000000480000000000000018000000000000000e000000000000000d00000000",
            INIT_3B => X"000000bb00000000000000bb000000000000006c000000000000004f00000000",
            INIT_3C => X"0000002b000000000000001b000000000000008b00000000000000bf00000000",
            INIT_3D => X"0000001b000000000000001c000000000000001b000000000000001e00000000",
            INIT_3E => X"00000059000000000000007b0000000000000084000000000000006c00000000",
            INIT_3F => X"0000003b000000000000002a0000000000000015000000000000001600000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003f00000000000000470000000000000066000000000000006d00000000",
            INIT_41 => X"0000001c000000000000004d0000000000000071000000000000003c00000000",
            INIT_42 => X"000000470000000000000030000000000000001f000000000000001000000000",
            INIT_43 => X"000000b300000000000000bd0000000000000088000000000000004600000000",
            INIT_44 => X"00000036000000000000001f000000000000007400000000000000b400000000",
            INIT_45 => X"0000000e000000000000001b0000000000000029000000000000003500000000",
            INIT_46 => X"0000003c000000000000007c0000000000000085000000000000004800000000",
            INIT_47 => X"0000003b00000000000000320000000000000022000000000000001200000000",
            INIT_48 => X"0000003c000000000000003d0000000000000051000000000000005700000000",
            INIT_49 => X"00000015000000000000004b0000000000000069000000000000003a00000000",
            INIT_4A => X"00000060000000000000004c000000000000002e000000000000001400000000",
            INIT_4B => X"000000a300000000000000a40000000000000091000000000000006100000000",
            INIT_4C => X"000000390000000000000020000000000000007100000000000000aa00000000",
            INIT_4D => X"0000001100000000000000250000000000000031000000000000004700000000",
            INIT_4E => X"000000210000000000000060000000000000006c000000000000002900000000",
            INIT_4F => X"000000320000000000000028000000000000001d000000000000000c00000000",
            INIT_50 => X"0000003c00000000000000400000000000000049000000000000004900000000",
            INIT_51 => X"0000002f0000000000000057000000000000005f000000000000003900000000",
            INIT_52 => X"000000a500000000000000890000000000000062000000000000003d00000000",
            INIT_53 => X"000000b600000000000000b700000000000000b000000000000000a900000000",
            INIT_54 => X"000000360000000000000022000000000000007c00000000000000b600000000",
            INIT_55 => X"0000001b0000000000000033000000000000005c000000000000006000000000",
            INIT_56 => X"0000000c000000000000003b0000000000000046000000000000001100000000",
            INIT_57 => X"00000028000000000000001d0000000000000012000000000000000600000000",
            INIT_58 => X"0000004e00000000000000450000000000000049000000000000004900000000",
            INIT_59 => X"0000002f00000000000000450000000000000059000000000000004100000000",
            INIT_5A => X"00000056000000000000004a000000000000003c000000000000003400000000",
            INIT_5B => X"0000006000000000000000620000000000000060000000000000005b00000000",
            INIT_5C => X"0000003c00000000000000200000000000000053000000000000006200000000",
            INIT_5D => X"00000014000000000000001d000000000000003e000000000000003b00000000",
            INIT_5E => X"00000003000000000000000a0000000000000011000000000000000400000000",
            INIT_5F => X"000000210000000000000011000000000000000a000000000000000700000000",
            INIT_60 => X"0000003600000000000000480000000000000053000000000000004b00000000",
            INIT_61 => X"00000004000000000000000f0000000000000027000000000000002d00000000",
            INIT_62 => X"0000000700000000000000050000000000000002000000000000000300000000",
            INIT_63 => X"0000000b000000000000000a0000000000000008000000000000000700000000",
            INIT_64 => X"000000420000000000000008000000000000000d000000000000000b00000000",
            INIT_65 => X"0000000f0000000000000038000000000000002f000000000000004300000000",
            INIT_66 => X"0000000300000000000000010000000000000002000000000000000200000000",
            INIT_67 => X"00000020000000000000000f000000000000000a000000000000000600000000",
            INIT_68 => X"0000002f00000000000000510000000000000059000000000000005000000000",
            INIT_69 => X"000000190000000000000010000000000000000a000000000000001500000000",
            INIT_6A => X"0000000e000000000000000e000000000000000a000000000000000e00000000",
            INIT_6B => X"0000000c000000000000000e000000000000000e000000000000000e00000000",
            INIT_6C => X"0000001700000000000000060000000000000009000000000000000a00000000",
            INIT_6D => X"00000007000000000000002a0000000000000048000000000000003e00000000",
            INIT_6E => X"0000000500000000000000050000000000000004000000000000000300000000",
            INIT_6F => X"000000210000000000000015000000000000000b000000000000000700000000",
            INIT_70 => X"000000370000000000000049000000000000004f000000000000004900000000",
            INIT_71 => X"0000003a000000000000003b000000000000002f000000000000002e00000000",
            INIT_72 => X"0000001c00000000000000190000000000000011000000000000001a00000000",
            INIT_73 => X"0000001c000000000000001d0000000000000020000000000000001f00000000",
            INIT_74 => X"0000000c00000000000000100000000000000015000000000000001800000000",
            INIT_75 => X"0000000600000000000000080000000000000016000000000000001400000000",
            INIT_76 => X"0000000800000000000000080000000000000007000000000000000800000000",
            INIT_77 => X"0000001f000000000000001b000000000000000f000000000000000b00000000",
            INIT_78 => X"0000004e000000000000004c0000000000000048000000000000004500000000",
            INIT_79 => X"0000003800000000000000480000000000000053000000000000005800000000",
            INIT_7A => X"0000002a000000000000002b0000000000000026000000000000002000000000",
            INIT_7B => X"0000003100000000000000320000000000000033000000000000002f00000000",
            INIT_7C => X"0000001c000000000000001e0000000000000026000000000000002c00000000",
            INIT_7D => X"0000000c00000000000000130000000000000022000000000000002200000000",
            INIT_7E => X"0000000d000000000000000f0000000000000010000000000000000e00000000",
            INIT_7F => X"0000001d000000000000001e000000000000001a000000000000001200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "sampleifmap_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003a00000000000000390000000000000031000000000000002500000000",
            INIT_01 => X"000000510000000000000050000000000000004e000000000000004200000000",
            INIT_02 => X"0000004200000000000000490000000000000052000000000000005600000000",
            INIT_03 => X"0000003800000000000000430000000000000043000000000000004100000000",
            INIT_04 => X"0000007300000000000000400000000000000032000000000000003200000000",
            INIT_05 => X"0000002700000000000000320000000000000038000000000000003400000000",
            INIT_06 => X"00000024000000000000002e0000000000000022000000000000001600000000",
            INIT_07 => X"0000001300000000000000150000000000000012000000000000001d00000000",
            INIT_08 => X"00000044000000000000004d0000000000000048000000000000004300000000",
            INIT_09 => X"000000420000000000000048000000000000004a000000000000004300000000",
            INIT_0A => X"0000003400000000000000390000000000000040000000000000004400000000",
            INIT_0B => X"0000002e00000000000000370000000000000036000000000000003200000000",
            INIT_0C => X"000000290000000000000027000000000000002a000000000000002900000000",
            INIT_0D => X"00000021000000000000001e0000000000000023000000000000002800000000",
            INIT_0E => X"0000001b000000000000001e000000000000002e000000000000002200000000",
            INIT_0F => X"0000001200000000000000160000000000000015000000000000001c00000000",
            INIT_10 => X"0000003e00000000000000480000000000000044000000000000004800000000",
            INIT_11 => X"000000310000000000000038000000000000003d000000000000003a00000000",
            INIT_12 => X"00000028000000000000002b000000000000002d000000000000003000000000",
            INIT_13 => X"00000026000000000000002b000000000000002a000000000000002600000000",
            INIT_14 => X"0000001c000000000000001e0000000000000023000000000000002200000000",
            INIT_15 => X"00000022000000000000001f0000000000000021000000000000002300000000",
            INIT_16 => X"0000000e000000000000000d0000000000000022000000000000003000000000",
            INIT_17 => X"0000001100000000000000130000000000000014000000000000001500000000",
            INIT_18 => X"0000003c000000000000003d0000000000000036000000000000003800000000",
            INIT_19 => X"00000024000000000000002b0000000000000030000000000000003e00000000",
            INIT_1A => X"0000002000000000000000220000000000000023000000000000002300000000",
            INIT_1B => X"0000002000000000000000220000000000000021000000000000001f00000000",
            INIT_1C => X"0000001d000000000000001b000000000000001e000000000000001d00000000",
            INIT_1D => X"00000025000000000000001d000000000000001c000000000000002000000000",
            INIT_1E => X"0000000f000000000000000b0000000000000012000000000000002a00000000",
            INIT_1F => X"0000001100000000000000100000000000000013000000000000001600000000",
            INIT_20 => X"0000003b00000000000000420000000000000039000000000000003900000000",
            INIT_21 => X"0000001b00000000000000200000000000000024000000000000003400000000",
            INIT_22 => X"0000001a000000000000001c000000000000001d000000000000001c00000000",
            INIT_23 => X"0000001e000000000000001c000000000000001a000000000000001a00000000",
            INIT_24 => X"0000001c000000000000001c000000000000001c000000000000001c00000000",
            INIT_25 => X"0000002a00000000000000430000000000000030000000000000001c00000000",
            INIT_26 => X"00000019000000000000000d0000000000000012000000000000001900000000",
            INIT_27 => X"000000110000000000000013000000000000001f000000000000001b00000000",
            INIT_28 => X"00000021000000000000002f000000000000003a000000000000003b00000000",
            INIT_29 => X"000000160000000000000019000000000000001a000000000000001a00000000",
            INIT_2A => X"00000019000000000000001a0000000000000019000000000000001700000000",
            INIT_2B => X"0000001f000000000000001b0000000000000018000000000000001800000000",
            INIT_2C => X"0000001e0000000000000021000000000000001e000000000000001d00000000",
            INIT_2D => X"0000003c000000000000005e000000000000005d000000000000002100000000",
            INIT_2E => X"0000002c000000000000001e000000000000001b000000000000002900000000",
            INIT_2F => X"000000130000000000000018000000000000002d000000000000002b00000000",
            INIT_30 => X"000000140000000000000017000000000000001c000000000000002200000000",
            INIT_31 => X"0000001500000000000000160000000000000017000000000000001600000000",
            INIT_32 => X"0000001a00000000000000190000000000000016000000000000001600000000",
            INIT_33 => X"00000023000000000000001d0000000000000019000000000000001800000000",
            INIT_34 => X"0000001e0000000000000023000000000000001f000000000000002000000000",
            INIT_35 => X"0000002500000000000000370000000000000059000000000000003300000000",
            INIT_36 => X"0000002d000000000000002b0000000000000028000000000000003800000000",
            INIT_37 => X"000000150000000000000017000000000000001e000000000000002400000000",
            INIT_38 => X"0000001200000000000000100000000000000011000000000000001100000000",
            INIT_39 => X"0000001600000000000000160000000000000017000000000000001600000000",
            INIT_3A => X"0000001b000000000000001a0000000000000017000000000000001800000000",
            INIT_3B => X"00000027000000000000001d000000000000001b000000000000001900000000",
            INIT_3C => X"000000300000000000000033000000000000002d000000000000002800000000",
            INIT_3D => X"0000000b00000000000000120000000000000040000000000000004100000000",
            INIT_3E => X"00000020000000000000001f0000000000000025000000000000002200000000",
            INIT_3F => X"0000001500000000000000160000000000000016000000000000001900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000000000120000000000000012000000000000001100000000",
            INIT_41 => X"0000001700000000000000170000000000000016000000000000001500000000",
            INIT_42 => X"0000001e000000000000001c0000000000000018000000000000001900000000",
            INIT_43 => X"0000003b00000000000000330000000000000038000000000000002500000000",
            INIT_44 => X"000000360000000000000037000000000000003a000000000000003b00000000",
            INIT_45 => X"0000001000000000000000110000000000000028000000000000003d00000000",
            INIT_46 => X"0000001b00000000000000180000000000000019000000000000001a00000000",
            INIT_47 => X"0000001400000000000000150000000000000017000000000000001a00000000",
            INIT_48 => X"0000001200000000000000120000000000000012000000000000001300000000",
            INIT_49 => X"0000001800000000000000160000000000000014000000000000001500000000",
            INIT_4A => X"0000003100000000000000200000000000000019000000000000001800000000",
            INIT_4B => X"000000340000000000000039000000000000004c000000000000003e00000000",
            INIT_4C => X"0000003a0000000000000032000000000000002e000000000000003100000000",
            INIT_4D => X"0000002c00000000000000300000000000000031000000000000003800000000",
            INIT_4E => X"0000001900000000000000190000000000000023000000000000002900000000",
            INIT_4F => X"0000001400000000000000140000000000000018000000000000001900000000",
            INIT_50 => X"0000001200000000000000130000000000000012000000000000001400000000",
            INIT_51 => X"0000001700000000000000150000000000000015000000000000001500000000",
            INIT_52 => X"0000003500000000000000240000000000000019000000000000001900000000",
            INIT_53 => X"0000004a000000000000003e0000000000000042000000000000003100000000",
            INIT_54 => X"000000b800000000000000a60000000000000089000000000000006800000000",
            INIT_55 => X"00000021000000000000004b0000000000000068000000000000007c00000000",
            INIT_56 => X"000000190000000000000026000000000000003d000000000000003800000000",
            INIT_57 => X"0000001300000000000000120000000000000019000000000000001800000000",
            INIT_58 => X"0000001300000000000000140000000000000012000000000000001500000000",
            INIT_59 => X"0000001800000000000000160000000000000018000000000000001800000000",
            INIT_5A => X"00000030000000000000001f000000000000001d000000000000001900000000",
            INIT_5B => X"000000be00000000000000b20000000000000097000000000000005500000000",
            INIT_5C => X"000000c500000000000000ca00000000000000cd00000000000000cd00000000",
            INIT_5D => X"00000016000000000000009800000000000000d000000000000000b200000000",
            INIT_5E => X"0000002800000000000000460000000000000025000000000000001800000000",
            INIT_5F => X"0000001100000000000000110000000000000016000000000000001500000000",
            INIT_60 => X"0000001500000000000000160000000000000014000000000000001400000000",
            INIT_61 => X"0000001a00000000000000190000000000000018000000000000001800000000",
            INIT_62 => X"0000007000000000000000420000000000000020000000000000001900000000",
            INIT_63 => X"00000075000000000000008c000000000000009b000000000000009000000000",
            INIT_64 => X"0000003d00000000000000470000000000000058000000000000006400000000",
            INIT_65 => X"0000004e00000000000000d500000000000000e8000000000000007500000000",
            INIT_66 => X"000000460000000000000032000000000000000a000000000000000f00000000",
            INIT_67 => X"0000001000000000000000110000000000000015000000000000001a00000000",
            INIT_68 => X"0000001600000000000000190000000000000016000000000000001400000000",
            INIT_69 => X"0000001a00000000000000190000000000000017000000000000001700000000",
            INIT_6A => X"0000005b00000000000000670000000000000048000000000000001a00000000",
            INIT_6B => X"0000001200000000000000340000000000000056000000000000005000000000",
            INIT_6C => X"00000010000000000000000f0000000000000022000000000000001100000000",
            INIT_6D => X"0000009b00000000000000e000000000000000dd000000000000007c00000000",
            INIT_6E => X"0000003b00000000000000160000000000000007000000000000002400000000",
            INIT_6F => X"0000001000000000000000120000000000000013000000000000002100000000",
            INIT_70 => X"00000016000000000000001b0000000000000017000000000000001800000000",
            INIT_71 => X"0000001500000000000000130000000000000019000000000000001800000000",
            INIT_72 => X"00000029000000000000003a0000000000000055000000000000003700000000",
            INIT_73 => X"000000180000000000000032000000000000004e000000000000003d00000000",
            INIT_74 => X"00000049000000000000001e000000000000002b000000000000000b00000000",
            INIT_75 => X"000000cd00000000000000d100000000000000d800000000000000bf00000000",
            INIT_76 => X"000000170000000000000010000000000000000e000000000000006700000000",
            INIT_77 => X"0000001200000000000000140000000000000016000000000000001b00000000",
            INIT_78 => X"00000017000000000000001a0000000000000016000000000000001a00000000",
            INIT_79 => X"00000034000000000000003c0000000000000025000000000000001900000000",
            INIT_7A => X"0000003b00000000000000380000000000000034000000000000004c00000000",
            INIT_7B => X"00000026000000000000002e000000000000004d000000000000005000000000",
            INIT_7C => X"000000c4000000000000007c0000000000000049000000000000002300000000",
            INIT_7D => X"000000d200000000000000d900000000000000d800000000000000df00000000",
            INIT_7E => X"0000000e00000000000000150000000000000039000000000000007600000000",
            INIT_7F => X"00000011000000000000003e0000000000000047000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "sampleifmap_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001700000000000000190000000000000014000000000000001900000000",
            INIT_01 => X"0000005c00000000000000600000000000000035000000000000002100000000",
            INIT_02 => X"00000042000000000000003e000000000000005d000000000000004900000000",
            INIT_03 => X"000000a2000000000000005a0000000000000047000000000000005100000000",
            INIT_04 => X"000000f500000000000000f500000000000000df00000000000000c400000000",
            INIT_05 => X"0000007900000000000000de00000000000000e400000000000000e300000000",
            INIT_06 => X"000000090000000000000011000000000000003b000000000000002500000000",
            INIT_07 => X"000000130000000000000075000000000000008c000000000000004800000000",
            INIT_08 => X"0000001a00000000000000180000000000000015000000000000001900000000",
            INIT_09 => X"000000450000000000000035000000000000002c000000000000002800000000",
            INIT_0A => X"0000002900000000000000250000000000000052000000000000005800000000",
            INIT_0B => X"000000fb00000000000000940000000000000020000000000000003100000000",
            INIT_0C => X"000000e200000000000000e900000000000000f200000000000000f600000000",
            INIT_0D => X"0000001f000000000000008b00000000000000e200000000000000e100000000",
            INIT_0E => X"0000004300000000000000280000000000000019000000000000000b00000000",
            INIT_0F => X"00000022000000000000009700000000000000a2000000000000008500000000",
            INIT_10 => X"0000002600000000000000160000000000000013000000000000001600000000",
            INIT_11 => X"00000036000000000000002e0000000000000046000000000000005d00000000",
            INIT_12 => X"0000001b00000000000000180000000000000026000000000000004b00000000",
            INIT_13 => X"000000e300000000000000a30000000000000031000000000000003800000000",
            INIT_14 => X"000000da00000000000000cb00000000000000cd00000000000000d600000000",
            INIT_15 => X"0000004a00000000000000a300000000000000e400000000000000e500000000",
            INIT_16 => X"000000950000000000000080000000000000005a000000000000003900000000",
            INIT_17 => X"0000003300000000000000a00000000000000096000000000000009700000000",
            INIT_18 => X"0000007c0000000000000026000000000000000f000000000000001300000000",
            INIT_19 => X"0000002a0000000000000024000000000000005a00000000000000af00000000",
            INIT_1A => X"00000015000000000000000b0000000000000017000000000000003f00000000",
            INIT_1B => X"000000d000000000000000aa000000000000004f000000000000004000000000",
            INIT_1C => X"000000d600000000000000d300000000000000c500000000000000c700000000",
            INIT_1D => X"000000b100000000000000e300000000000000d900000000000000ce00000000",
            INIT_1E => X"000000a200000000000000a700000000000000a8000000000000009800000000",
            INIT_1F => X"0000002a00000000000000880000000000000097000000000000009a00000000",
            INIT_20 => X"000000dc0000000000000065000000000000000a000000000000001200000000",
            INIT_21 => X"0000002e000000000000002f000000000000006f00000000000000be00000000",
            INIT_22 => X"0000000e0000000000000009000000000000000a000000000000003900000000",
            INIT_23 => X"000000cc00000000000000b10000000000000042000000000000001f00000000",
            INIT_24 => X"0000007c00000000000000c600000000000000ca00000000000000c200000000",
            INIT_25 => X"000000d300000000000000ac0000000000000066000000000000004f00000000",
            INIT_26 => X"000000a900000000000000b100000000000000b800000000000000c800000000",
            INIT_27 => X"00000011000000000000004a000000000000008c000000000000009c00000000",
            INIT_28 => X"000000a500000000000000840000000000000014000000000000000e00000000",
            INIT_29 => X"0000003400000000000000370000000000000080000000000000009600000000",
            INIT_2A => X"00000016000000000000000a0000000000000003000000000000001e00000000",
            INIT_2B => X"000000c600000000000000b40000000000000048000000000000002d00000000",
            INIT_2C => X"00000019000000000000007b00000000000000cd00000000000000be00000000",
            INIT_2D => X"000000a30000000000000038000000000000001e000000000000001a00000000",
            INIT_2E => X"00000093000000000000009e00000000000000b800000000000000ca00000000",
            INIT_2F => X"00000011000000000000000d0000000000000044000000000000008800000000",
            INIT_30 => X"0000002100000000000000530000000000000023000000000000000a00000000",
            INIT_31 => X"00000035000000000000003e0000000000000082000000000000005300000000",
            INIT_32 => X"0000004800000000000000100000000000000007000000000000001300000000",
            INIT_33 => X"000000c200000000000000b70000000000000075000000000000006c00000000",
            INIT_34 => X"0000001e000000000000002f00000000000000b700000000000000c300000000",
            INIT_35 => X"0000004f0000000000000014000000000000002b000000000000003100000000",
            INIT_36 => X"000000810000000000000084000000000000009400000000000000a100000000",
            INIT_37 => X"000000180000000000000009000000000000000a000000000000004000000000",
            INIT_38 => X"0000002300000000000000370000000000000021000000000000000a00000000",
            INIT_39 => X"00000024000000000000004e0000000000000088000000000000004600000000",
            INIT_3A => X"0000005800000000000000220000000000000011000000000000000f00000000",
            INIT_3B => X"000000cd00000000000000cd000000000000007e000000000000006100000000",
            INIT_3C => X"0000002b0000000000000020000000000000009800000000000000d000000000",
            INIT_3D => X"0000001f0000000000000020000000000000001f000000000000002000000000",
            INIT_3E => X"00000063000000000000008a0000000000000091000000000000007500000000",
            INIT_3F => X"000000210000000000000019000000000000000c000000000000001700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004100000000000000360000000000000015000000000000000a00000000",
            INIT_41 => X"0000002100000000000000570000000000000088000000000000004700000000",
            INIT_42 => X"00000057000000000000003f0000000000000027000000000000001500000000",
            INIT_43 => X"000000c500000000000000cf000000000000009a000000000000005600000000",
            INIT_44 => X"000000380000000000000025000000000000008100000000000000c600000000",
            INIT_45 => X"0000000f000000000000001c000000000000002c000000000000003700000000",
            INIT_46 => X"00000043000000000000008b0000000000000093000000000000004d00000000",
            INIT_47 => X"0000001f000000000000001c0000000000000014000000000000000e00000000",
            INIT_48 => X"0000003e000000000000002f000000000000000e000000000000000700000000",
            INIT_49 => X"0000001c00000000000000560000000000000080000000000000004500000000",
            INIT_4A => X"0000006f000000000000005e000000000000003c000000000000001e00000000",
            INIT_4B => X"000000b400000000000000b600000000000000a2000000000000006f00000000",
            INIT_4C => X"0000003c0000000000000029000000000000007f00000000000000bc00000000",
            INIT_4D => X"0000000f00000000000000230000000000000035000000000000004b00000000",
            INIT_4E => X"00000026000000000000006f000000000000007a000000000000002c00000000",
            INIT_4F => X"000000160000000000000010000000000000000d000000000000000700000000",
            INIT_50 => X"0000003b00000000000000270000000000000011000000000000000b00000000",
            INIT_51 => X"0000003d00000000000000680000000000000075000000000000004600000000",
            INIT_52 => X"000000b7000000000000009f0000000000000079000000000000005100000000",
            INIT_53 => X"000000c700000000000000c900000000000000c300000000000000b900000000",
            INIT_54 => X"0000003c000000000000002a000000000000008800000000000000c600000000",
            INIT_55 => X"0000001c00000000000000340000000000000062000000000000006600000000",
            INIT_56 => X"000000100000000000000045000000000000004f000000000000001500000000",
            INIT_57 => X"00000016000000000000000c0000000000000007000000000000000300000000",
            INIT_58 => X"00000043000000000000001d0000000000000014000000000000001300000000",
            INIT_59 => X"0000003c00000000000000550000000000000067000000000000004900000000",
            INIT_5A => X"00000064000000000000005b0000000000000050000000000000004500000000",
            INIT_5B => X"0000006d00000000000000710000000000000071000000000000006800000000",
            INIT_5C => X"0000004100000000000000250000000000000059000000000000006d00000000",
            INIT_5D => X"00000017000000000000001f0000000000000042000000000000004000000000",
            INIT_5E => X"00000005000000000000000e0000000000000014000000000000000800000000",
            INIT_5F => X"00000018000000000000000b0000000000000006000000000000000600000000",
            INIT_60 => X"00000025000000000000001d000000000000001c000000000000001700000000",
            INIT_61 => X"000000070000000000000016000000000000002c000000000000002c00000000",
            INIT_62 => X"0000000c000000000000000c000000000000000a000000000000000a00000000",
            INIT_63 => X"0000001000000000000000110000000000000010000000000000000d00000000",
            INIT_64 => X"000000430000000000000009000000000000000f000000000000000f00000000",
            INIT_65 => X"0000001000000000000000380000000000000030000000000000004400000000",
            INIT_66 => X"0000000400000000000000030000000000000003000000000000000400000000",
            INIT_67 => X"00000019000000000000000e0000000000000009000000000000000600000000",
            INIT_68 => X"0000002000000000000000270000000000000025000000000000002100000000",
            INIT_69 => X"0000002000000000000000190000000000000012000000000000001700000000",
            INIT_6A => X"0000001700000000000000170000000000000015000000000000001700000000",
            INIT_6B => X"0000000f00000000000000130000000000000015000000000000001700000000",
            INIT_6C => X"000000180000000000000007000000000000000a000000000000000b00000000",
            INIT_6D => X"0000000800000000000000290000000000000047000000000000003e00000000",
            INIT_6E => X"0000000600000000000000050000000000000005000000000000000400000000",
            INIT_6F => X"0000001d0000000000000018000000000000000e000000000000000900000000",
            INIT_70 => X"0000003200000000000000290000000000000025000000000000002300000000",
            INIT_71 => X"0000004d00000000000000510000000000000043000000000000003c00000000",
            INIT_72 => X"00000030000000000000002d0000000000000024000000000000002c00000000",
            INIT_73 => X"000000230000000000000027000000000000002c000000000000003100000000",
            INIT_74 => X"000000100000000000000015000000000000001b000000000000001d00000000",
            INIT_75 => X"00000009000000000000000a0000000000000019000000000000001700000000",
            INIT_76 => X"0000000b000000000000000a0000000000000009000000000000000b00000000",
            INIT_77 => X"0000001e000000000000001f0000000000000014000000000000000e00000000",
            INIT_78 => X"00000057000000000000003b000000000000002a000000000000002a00000000",
            INIT_79 => X"000000520000000000000066000000000000006f000000000000006d00000000",
            INIT_7A => X"000000470000000000000045000000000000003e000000000000003700000000",
            INIT_7B => X"0000004300000000000000460000000000000048000000000000004a00000000",
            INIT_7C => X"00000029000000000000002b0000000000000033000000000000003b00000000",
            INIT_7D => X"000000120000000000000018000000000000002c000000000000002f00000000",
            INIT_7E => X"0000001300000000000000150000000000000016000000000000001400000000",
            INIT_7F => X"0000001e0000000000000020000000000000001c000000000000001600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "sampleifmap_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000a000000000000000e000000000000000b000000000000000d00000000",
            INIT_01 => X"000000020000000000000005000000000000000a000000000000000900000000",
            INIT_02 => X"0000000200000000000000010000000000000003000000000000000300000000",
            INIT_03 => X"0000000000000000000000050000000000000006000000000000000400000000",
            INIT_04 => X"0000005600000000000000230000000000000000000000000000000100000000",
            INIT_05 => X"00000008000000000000001d0000000000000017000000000000001600000000",
            INIT_06 => X"0000001d0000000000000027000000000000001b000000000000000d00000000",
            INIT_07 => X"0000000500000000000000060000000000000008000000000000001300000000",
            INIT_08 => X"00000004000000000000000a000000000000000c000000000000000d00000000",
            INIT_09 => X"0000000000000000000000030000000000000008000000000000000700000000",
            INIT_0A => X"0000000100000000000000010000000000000002000000000000000400000000",
            INIT_0B => X"0000000100000000000000040000000000000004000000000000000200000000",
            INIT_0C => X"0000001300000000000000100000000000000001000000000000000100000000",
            INIT_0D => X"0000000700000000000000060000000000000006000000000000000700000000",
            INIT_0E => X"000000160000000000000017000000000000002e000000000000002100000000",
            INIT_0F => X"0000000600000000000000040000000000000008000000000000001300000000",
            INIT_10 => X"0000000000000000000000030000000000000004000000000000000700000000",
            INIT_11 => X"0000000000000000000000010000000000000004000000000000000400000000",
            INIT_12 => X"0000000400000000000000040000000000000004000000000000000400000000",
            INIT_13 => X"0000000300000000000000050000000000000006000000000000000400000000",
            INIT_14 => X"00000009000000000000000c0000000000000003000000000000000400000000",
            INIT_15 => X"0000000a00000000000000060000000000000007000000000000000400000000",
            INIT_16 => X"0000000c000000000000000d0000000000000023000000000000002800000000",
            INIT_17 => X"0000000600000000000000030000000000000006000000000000000f00000000",
            INIT_18 => X"0000000b00000000000000080000000000000003000000000000000100000000",
            INIT_19 => X"0000000300000000000000030000000000000004000000000000001200000000",
            INIT_1A => X"0000000700000000000000080000000000000006000000000000000500000000",
            INIT_1B => X"0000000600000000000000060000000000000009000000000000000800000000",
            INIT_1C => X"00000009000000000000000a0000000000000005000000000000000700000000",
            INIT_1D => X"000000170000000000000010000000000000000a000000000000000400000000",
            INIT_1E => X"0000000e00000000000000110000000000000016000000000000001e00000000",
            INIT_1F => X"0000000800000000000000050000000000000006000000000000000f00000000",
            INIT_20 => X"0000001a000000000000001d0000000000000013000000000000000c00000000",
            INIT_21 => X"0000000800000000000000070000000000000006000000000000001700000000",
            INIT_22 => X"0000000800000000000000090000000000000008000000000000000700000000",
            INIT_23 => X"000000080000000000000007000000000000000a000000000000000900000000",
            INIT_24 => X"0000000700000000000000080000000000000007000000000000000900000000",
            INIT_25 => X"0000002700000000000000400000000000000025000000000000000800000000",
            INIT_26 => X"00000015000000000000000e0000000000000010000000000000001000000000",
            INIT_27 => X"00000009000000000000000d000000000000000f000000000000000e00000000",
            INIT_28 => X"0000000c0000000000000016000000000000001e000000000000001800000000",
            INIT_29 => X"0000000800000000000000090000000000000006000000000000000900000000",
            INIT_2A => X"0000000a00000000000000090000000000000005000000000000000500000000",
            INIT_2B => X"000000090000000000000007000000000000000a000000000000000b00000000",
            INIT_2C => X"00000007000000000000000b000000000000000b000000000000000a00000000",
            INIT_2D => X"0000003b000000000000005d0000000000000055000000000000001400000000",
            INIT_2E => X"000000200000000000000013000000000000000e000000000000002200000000",
            INIT_2F => X"000000090000000000000010000000000000001b000000000000001700000000",
            INIT_30 => X"00000007000000000000000a000000000000000b000000000000000c00000000",
            INIT_31 => X"00000007000000000000000a0000000000000008000000000000000800000000",
            INIT_32 => X"0000000e000000000000000a0000000000000005000000000000000600000000",
            INIT_33 => X"0000000c000000000000000a000000000000000c000000000000000d00000000",
            INIT_34 => X"00000007000000000000000e000000000000000e000000000000000900000000",
            INIT_35 => X"00000028000000000000003c0000000000000056000000000000002500000000",
            INIT_36 => X"0000001c000000000000001c000000000000001c000000000000003500000000",
            INIT_37 => X"0000000700000000000000060000000000000010000000000000001400000000",
            INIT_38 => X"0000000700000000000000060000000000000006000000000000000300000000",
            INIT_39 => X"00000009000000000000000c000000000000000a000000000000000b00000000",
            INIT_3A => X"0000000e000000000000000c0000000000000008000000000000000900000000",
            INIT_3B => X"0000001300000000000000100000000000000012000000000000000e00000000",
            INIT_3C => X"00000016000000000000001a0000000000000015000000000000001000000000",
            INIT_3D => X"0000000a0000000000000014000000000000003e000000000000003100000000",
            INIT_3E => X"0000000d0000000000000010000000000000001a000000000000001e00000000",
            INIT_3F => X"0000000700000000000000040000000000000008000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000080000000000000009000000000000000a000000000000000700000000",
            INIT_41 => X"0000000b000000000000000e000000000000000a000000000000000b00000000",
            INIT_42 => X"0000000f000000000000000e000000000000000c000000000000000d00000000",
            INIT_43 => X"0000002800000000000000220000000000000024000000000000001300000000",
            INIT_44 => X"0000002200000000000000220000000000000020000000000000002400000000",
            INIT_45 => X"00000009000000000000000f000000000000002b000000000000003300000000",
            INIT_46 => X"0000000a0000000000000009000000000000000c000000000000001400000000",
            INIT_47 => X"0000000800000000000000080000000000000008000000000000000800000000",
            INIT_48 => X"00000008000000000000000b000000000000000c000000000000000c00000000",
            INIT_49 => X"0000000d000000000000000e000000000000000a000000000000000c00000000",
            INIT_4A => X"000000220000000000000014000000000000000e000000000000000e00000000",
            INIT_4B => X"0000002600000000000000280000000000000031000000000000002700000000",
            INIT_4C => X"000000320000000000000027000000000000001b000000000000002000000000",
            INIT_4D => X"000000260000000000000034000000000000003b000000000000003600000000",
            INIT_4E => X"0000000c000000000000000b0000000000000015000000000000002300000000",
            INIT_4F => X"0000000a000000000000000b0000000000000009000000000000000600000000",
            INIT_50 => X"00000009000000000000000b000000000000000b000000000000000c00000000",
            INIT_51 => X"0000000d000000000000000d000000000000000a000000000000000c00000000",
            INIT_52 => X"00000028000000000000001b0000000000000010000000000000000d00000000",
            INIT_53 => X"0000003f00000000000000320000000000000032000000000000002000000000",
            INIT_54 => X"000000b400000000000000a10000000000000077000000000000005800000000",
            INIT_55 => X"0000002200000000000000540000000000000071000000000000007900000000",
            INIT_56 => X"00000011000000000000001d0000000000000031000000000000003200000000",
            INIT_57 => X"0000000a000000000000000c000000000000000a000000000000000900000000",
            INIT_58 => X"0000000b000000000000000e000000000000000a000000000000000900000000",
            INIT_59 => X"0000000c000000000000000d000000000000000c000000000000000e00000000",
            INIT_5A => X"0000002700000000000000180000000000000012000000000000000c00000000",
            INIT_5B => X"000000ba00000000000000af0000000000000093000000000000004d00000000",
            INIT_5C => X"000000ca00000000000000d200000000000000c800000000000000c800000000",
            INIT_5D => X"0000001c000000000000009e00000000000000d500000000000000b100000000",
            INIT_5E => X"0000002500000000000000460000000000000022000000000000001300000000",
            INIT_5F => X"00000009000000000000000b0000000000000009000000000000000a00000000",
            INIT_60 => X"0000000d000000000000000f000000000000000a000000000000000800000000",
            INIT_61 => X"0000000e000000000000000d000000000000000e000000000000001000000000",
            INIT_62 => X"0000006c000000000000003e0000000000000018000000000000000c00000000",
            INIT_63 => X"0000007d000000000000009300000000000000a2000000000000008e00000000",
            INIT_64 => X"0000004a0000000000000054000000000000005e000000000000006e00000000",
            INIT_65 => X"0000005400000000000000d700000000000000f1000000000000007e00000000",
            INIT_66 => X"0000004900000000000000340000000000000009000000000000000c00000000",
            INIT_67 => X"000000080000000000000009000000000000000d000000000000001900000000",
            INIT_68 => X"0000000e000000000000000f000000000000000b000000000000000b00000000",
            INIT_69 => X"0000000e000000000000000c0000000000000010000000000000001100000000",
            INIT_6A => X"0000005d00000000000000670000000000000044000000000000001400000000",
            INIT_6B => X"00000019000000000000003d000000000000005f000000000000005600000000",
            INIT_6C => X"0000001700000000000000110000000000000023000000000000001600000000",
            INIT_6D => X"000000a700000000000000eb00000000000000eb000000000000008900000000",
            INIT_6E => X"0000004200000000000000170000000000000007000000000000002a00000000",
            INIT_6F => X"0000000700000000000000090000000000000011000000000000002800000000",
            INIT_70 => X"0000000e0000000000000012000000000000000d000000000000000f00000000",
            INIT_71 => X"00000012000000000000000b0000000000000012000000000000001000000000",
            INIT_72 => X"0000002e000000000000003b0000000000000053000000000000003600000000",
            INIT_73 => X"0000001b00000000000000370000000000000053000000000000004400000000",
            INIT_74 => X"0000004c000000000000001c0000000000000027000000000000000c00000000",
            INIT_75 => X"000000e000000000000000e700000000000000e800000000000000c800000000",
            INIT_76 => X"0000001a00000000000000130000000000000016000000000000007300000000",
            INIT_77 => X"00000008000000000000000d0000000000000016000000000000001f00000000",
            INIT_78 => X"0000000e0000000000000013000000000000000d000000000000001000000000",
            INIT_79 => X"000000370000000000000039000000000000001e000000000000000e00000000",
            INIT_7A => X"0000003c00000000000000390000000000000035000000000000004f00000000",
            INIT_7B => X"000000290000000000000032000000000000004e000000000000005200000000",
            INIT_7C => X"000000c8000000000000007c0000000000000047000000000000002300000000",
            INIT_7D => X"000000dd00000000000000ec00000000000000e600000000000000e700000000",
            INIT_7E => X"0000000e000000000000001a0000000000000044000000000000007e00000000",
            INIT_7F => X"00000009000000000000003f0000000000000049000000000000002000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "sampleifmap_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000110000000000000013000000000000000e000000000000001100000000",
            INIT_01 => X"0000005c000000000000005d000000000000002f000000000000001800000000",
            INIT_02 => X"0000003d000000000000003c0000000000000062000000000000004f00000000",
            INIT_03 => X"000000a6000000000000005e0000000000000047000000000000004c00000000",
            INIT_04 => X"000000fc00000000000000fa00000000000000e200000000000000c600000000",
            INIT_05 => X"0000007c00000000000000e700000000000000f000000000000000ed00000000",
            INIT_06 => X"0000000c000000000000001c000000000000004a000000000000002a00000000",
            INIT_07 => X"00000011000000000000007e0000000000000095000000000000004c00000000",
            INIT_08 => X"0000001500000000000000120000000000000010000000000000001200000000",
            INIT_09 => X"000000480000000000000038000000000000002a000000000000002400000000",
            INIT_0A => X"0000002400000000000000240000000000000058000000000000006000000000",
            INIT_0B => X"00000100000000000000009a0000000000000022000000000000002d00000000",
            INIT_0C => X"000000ed00000000000000f400000000000000f900000000000000fa00000000",
            INIT_0D => X"00000027000000000000009600000000000000ee00000000000000ed00000000",
            INIT_0E => X"0000004d000000000000003b000000000000002e000000000000001500000000",
            INIT_0F => X"0000002600000000000000a300000000000000ae000000000000008e00000000",
            INIT_10 => X"0000002200000000000000100000000000000010000000000000001100000000",
            INIT_11 => X"00000042000000000000003c0000000000000049000000000000005c00000000",
            INIT_12 => X"00000021000000000000001c000000000000002c000000000000005400000000",
            INIT_13 => X"000000f000000000000000ae0000000000000037000000000000003e00000000",
            INIT_14 => X"000000e700000000000000d900000000000000d900000000000000e100000000",
            INIT_15 => X"0000005600000000000000b100000000000000ee00000000000000ef00000000",
            INIT_16 => X"000000a40000000000000092000000000000006a000000000000004500000000",
            INIT_17 => X"0000003700000000000000a900000000000000a100000000000000a400000000",
            INIT_18 => X"0000007d0000000000000020000000000000000a000000000000000d00000000",
            INIT_19 => X"000000380000000000000035000000000000006200000000000000b400000000",
            INIT_1A => X"0000001b000000000000000e000000000000001c000000000000004800000000",
            INIT_1B => X"000000e000000000000000b90000000000000059000000000000004900000000",
            INIT_1C => X"000000e300000000000000e400000000000000d500000000000000d500000000",
            INIT_1D => X"000000c000000000000000f200000000000000e100000000000000d700000000",
            INIT_1E => X"000000b000000000000000b500000000000000b400000000000000a500000000",
            INIT_1F => X"0000002a000000000000008d000000000000009f00000000000000a600000000",
            INIT_20 => X"000000e500000000000000650000000000000007000000000000000c00000000",
            INIT_21 => X"00000039000000000000003e000000000000007b00000000000000c900000000",
            INIT_22 => X"0000000f0000000000000009000000000000000f000000000000004100000000",
            INIT_23 => X"000000da00000000000000bf000000000000004f000000000000002600000000",
            INIT_24 => X"0000008a00000000000000d800000000000000db00000000000000d000000000",
            INIT_25 => X"000000e400000000000000b8000000000000006d000000000000005800000000",
            INIT_26 => X"000000b500000000000000bf00000000000000c900000000000000da00000000",
            INIT_27 => X"0000000e000000000000004d000000000000009300000000000000a600000000",
            INIT_28 => X"000000b3000000000000008b0000000000000018000000000000000d00000000",
            INIT_29 => X"0000003d0000000000000045000000000000008d00000000000000a200000000",
            INIT_2A => X"0000001b000000000000000b0000000000000004000000000000002300000000",
            INIT_2B => X"000000d400000000000000c20000000000000056000000000000003600000000",
            INIT_2C => X"00000024000000000000008800000000000000db00000000000000cc00000000",
            INIT_2D => X"000000b100000000000000400000000000000022000000000000002000000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000cc00000000000000dd00000000",
            INIT_2F => X"0000000d000000000000000f0000000000000049000000000000009000000000",
            INIT_30 => X"00000031000000000000005b0000000000000027000000000000000900000000",
            INIT_31 => X"0000003e000000000000004c000000000000008f000000000000006000000000",
            INIT_32 => X"0000005100000000000000150000000000000007000000000000001500000000",
            INIT_33 => X"000000d000000000000000c50000000000000083000000000000007900000000",
            INIT_34 => X"00000026000000000000003800000000000000c100000000000000d100000000",
            INIT_35 => X"000000590000000000000019000000000000002e000000000000003700000000",
            INIT_36 => X"0000008d000000000000009500000000000000a900000000000000b200000000",
            INIT_37 => X"000000140000000000000008000000000000000e000000000000004800000000",
            INIT_38 => X"00000030000000000000003b0000000000000022000000000000000500000000",
            INIT_39 => X"0000002d000000000000005c0000000000000095000000000000005300000000",
            INIT_3A => X"00000064000000000000002a0000000000000013000000000000000f00000000",
            INIT_3B => X"000000db00000000000000db000000000000008c000000000000006f00000000",
            INIT_3C => X"00000033000000000000002600000000000000a000000000000000de00000000",
            INIT_3D => X"0000002700000000000000240000000000000023000000000000002500000000",
            INIT_3E => X"0000006e000000000000009b00000000000000a4000000000000008200000000",
            INIT_3F => X"0000001e0000000000000016000000000000000c000000000000001d00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d000000000000003a0000000000000017000000000000000700000000",
            INIT_41 => X"0000002a00000000000000650000000000000094000000000000005400000000",
            INIT_42 => X"00000065000000000000004a000000000000002b000000000000001600000000",
            INIT_43 => X"000000d300000000000000dd00000000000000a8000000000000006400000000",
            INIT_44 => X"00000040000000000000002b000000000000008900000000000000d400000000",
            INIT_45 => X"0000001500000000000000230000000000000034000000000000003f00000000",
            INIT_46 => X"0000004e000000000000009a00000000000000a2000000000000005600000000",
            INIT_47 => X"0000001c00000000000000180000000000000012000000000000001300000000",
            INIT_48 => X"0000004c00000000000000370000000000000015000000000000000900000000",
            INIT_49 => X"000000250000000000000065000000000000008c000000000000005200000000",
            INIT_4A => X"0000007f000000000000006c0000000000000043000000000000002100000000",
            INIT_4B => X"000000c200000000000000c300000000000000b0000000000000007e00000000",
            INIT_4C => X"000000460000000000000030000000000000008700000000000000c900000000",
            INIT_4D => X"00000015000000000000002e0000000000000041000000000000005600000000",
            INIT_4E => X"00000031000000000000007b0000000000000083000000000000003200000000",
            INIT_4F => X"00000014000000000000000b000000000000000a000000000000000b00000000",
            INIT_50 => X"0000004900000000000000310000000000000017000000000000000b00000000",
            INIT_51 => X"0000004b00000000000000780000000000000084000000000000005700000000",
            INIT_52 => X"000000c800000000000000b10000000000000086000000000000005d00000000",
            INIT_53 => X"000000d500000000000000d400000000000000cf00000000000000c800000000",
            INIT_54 => X"000000480000000000000035000000000000009400000000000000d600000000",
            INIT_55 => X"000000220000000000000040000000000000006e000000000000007100000000",
            INIT_56 => X"00000016000000000000004c0000000000000055000000000000001800000000",
            INIT_57 => X"00000016000000000000000d0000000000000009000000000000000700000000",
            INIT_58 => X"0000004e00000000000000250000000000000016000000000000000f00000000",
            INIT_59 => X"0000004800000000000000600000000000000073000000000000005700000000",
            INIT_5A => X"000000720000000000000069000000000000005d000000000000005200000000",
            INIT_5B => X"0000007b000000000000007e000000000000007d000000000000007700000000",
            INIT_5C => X"0000004c00000000000000300000000000000066000000000000007c00000000",
            INIT_5D => X"0000001b0000000000000029000000000000004e000000000000004b00000000",
            INIT_5E => X"0000000600000000000000100000000000000018000000000000000900000000",
            INIT_5F => X"00000019000000000000000f000000000000000a000000000000000800000000",
            INIT_60 => X"0000002b0000000000000023000000000000001f000000000000001500000000",
            INIT_61 => X"0000000c00000000000000190000000000000030000000000000003200000000",
            INIT_62 => X"000000110000000000000011000000000000000e000000000000000e00000000",
            INIT_63 => X"00000019000000000000001a0000000000000018000000000000001400000000",
            INIT_64 => X"0000004a000000000000000d0000000000000014000000000000001800000000",
            INIT_65 => X"000000120000000000000041000000000000003b000000000000004e00000000",
            INIT_66 => X"0000000300000000000000040000000000000005000000000000000300000000",
            INIT_67 => X"0000001a000000000000000d0000000000000009000000000000000500000000",
            INIT_68 => X"00000025000000000000002c0000000000000028000000000000002100000000",
            INIT_69 => X"00000025000000000000001e0000000000000017000000000000001e00000000",
            INIT_6A => X"0000001c000000000000001c0000000000000019000000000000001c00000000",
            INIT_6B => X"0000001300000000000000170000000000000018000000000000001b00000000",
            INIT_6C => X"0000001c00000000000000060000000000000009000000000000000f00000000",
            INIT_6D => X"00000008000000000000002f0000000000000053000000000000004700000000",
            INIT_6E => X"0000000400000000000000050000000000000005000000000000000200000000",
            INIT_6F => X"0000001c0000000000000015000000000000000b000000000000000600000000",
            INIT_70 => X"0000003b00000000000000300000000000000029000000000000002500000000",
            INIT_71 => X"00000059000000000000005c000000000000004f000000000000004900000000",
            INIT_72 => X"0000003b0000000000000038000000000000002f000000000000003800000000",
            INIT_73 => X"00000028000000000000002b0000000000000030000000000000003900000000",
            INIT_74 => X"000000150000000000000015000000000000001b000000000000002300000000",
            INIT_75 => X"0000000800000000000000100000000000000025000000000000002100000000",
            INIT_76 => X"0000000a000000000000000a0000000000000009000000000000000800000000",
            INIT_77 => X"0000001c000000000000001d0000000000000012000000000000000d00000000",
            INIT_78 => X"0000006500000000000000460000000000000031000000000000002c00000000",
            INIT_79 => X"0000006300000000000000760000000000000080000000000000008000000000",
            INIT_7A => X"000000550000000000000054000000000000004e000000000000004700000000",
            INIT_7B => X"0000004f00000000000000510000000000000053000000000000005700000000",
            INIT_7C => X"000000310000000000000031000000000000003c000000000000004700000000",
            INIT_7D => X"0000001300000000000000200000000000000038000000000000003a00000000",
            INIT_7E => X"0000001500000000000000180000000000000018000000000000001300000000",
            INIT_7F => X"0000001c0000000000000022000000000000001f000000000000001900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "sampleifmap_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004d00000000000000510000000000000052000000000000005300000000",
            INIT_01 => X"0000005c000000000000005b0000000000000055000000000000005100000000",
            INIT_02 => X"0000005c0000000000000065000000000000005f000000000000005c00000000",
            INIT_03 => X"0000004c00000000000000500000000000000052000000000000005700000000",
            INIT_04 => X"0000003e000000000000003f0000000000000041000000000000004400000000",
            INIT_05 => X"0000002f00000000000000340000000000000038000000000000003c00000000",
            INIT_06 => X"0000002200000000000000230000000000000025000000000000002a00000000",
            INIT_07 => X"000000150000000000000019000000000000001d000000000000002400000000",
            INIT_08 => X"0000004d00000000000000530000000000000053000000000000005400000000",
            INIT_09 => X"0000005d000000000000005a0000000000000054000000000000005000000000",
            INIT_0A => X"00000061000000000000005f0000000000000058000000000000005a00000000",
            INIT_0B => X"0000004c000000000000004e0000000000000052000000000000005800000000",
            INIT_0C => X"0000004200000000000000400000000000000044000000000000004700000000",
            INIT_0D => X"0000002e00000000000000340000000000000036000000000000003d00000000",
            INIT_0E => X"0000002300000000000000240000000000000026000000000000002a00000000",
            INIT_0F => X"0000001f000000000000001d000000000000001e000000000000002400000000",
            INIT_10 => X"0000004b00000000000000500000000000000051000000000000005200000000",
            INIT_11 => X"0000004c00000000000000580000000000000054000000000000004b00000000",
            INIT_12 => X"0000006300000000000000570000000000000056000000000000005200000000",
            INIT_13 => X"0000004c000000000000004d0000000000000058000000000000006500000000",
            INIT_14 => X"0000004000000000000000400000000000000044000000000000004900000000",
            INIT_15 => X"0000002d00000000000000340000000000000037000000000000003a00000000",
            INIT_16 => X"0000002c00000000000000290000000000000028000000000000002b00000000",
            INIT_17 => X"0000003500000000000000310000000000000030000000000000003100000000",
            INIT_18 => X"0000004e00000000000000500000000000000051000000000000005300000000",
            INIT_19 => X"0000003200000000000000500000000000000057000000000000004a00000000",
            INIT_1A => X"0000005b00000000000000570000000000000061000000000000005500000000",
            INIT_1B => X"0000005000000000000000580000000000000066000000000000006800000000",
            INIT_1C => X"0000003f000000000000003f0000000000000040000000000000004900000000",
            INIT_1D => X"0000003a00000000000000390000000000000038000000000000003b00000000",
            INIT_1E => X"000000470000000000000044000000000000003f000000000000003d00000000",
            INIT_1F => X"0000004500000000000000450000000000000047000000000000004900000000",
            INIT_20 => X"0000004f000000000000004f000000000000004f000000000000004f00000000",
            INIT_21 => X"00000037000000000000004c0000000000000053000000000000004a00000000",
            INIT_22 => X"0000004b000000000000004b0000000000000054000000000000005300000000",
            INIT_23 => X"00000057000000000000005a0000000000000059000000000000004e00000000",
            INIT_24 => X"0000004600000000000000430000000000000042000000000000005300000000",
            INIT_25 => X"0000005700000000000000540000000000000050000000000000004e00000000",
            INIT_26 => X"0000005900000000000000590000000000000056000000000000005700000000",
            INIT_27 => X"00000049000000000000004f0000000000000054000000000000005800000000",
            INIT_28 => X"0000004d000000000000004b000000000000004a000000000000004c00000000",
            INIT_29 => X"0000004600000000000000460000000000000049000000000000004900000000",
            INIT_2A => X"0000004900000000000000470000000000000045000000000000004600000000",
            INIT_2B => X"00000051000000000000004e000000000000004e000000000000004b00000000",
            INIT_2C => X"0000006200000000000000600000000000000059000000000000005a00000000",
            INIT_2D => X"0000006800000000000000660000000000000068000000000000006400000000",
            INIT_2E => X"0000005e0000000000000061000000000000005f000000000000006300000000",
            INIT_2F => X"0000004200000000000000490000000000000050000000000000005700000000",
            INIT_30 => X"0000004900000000000000470000000000000048000000000000004a00000000",
            INIT_31 => X"00000033000000000000002b000000000000003e000000000000004a00000000",
            INIT_32 => X"0000004700000000000000440000000000000040000000000000004400000000",
            INIT_33 => X"0000005e0000000000000051000000000000004a000000000000004b00000000",
            INIT_34 => X"00000072000000000000006e0000000000000062000000000000006000000000",
            INIT_35 => X"0000006d00000000000000680000000000000064000000000000006600000000",
            INIT_36 => X"000000500000000000000055000000000000005b000000000000006300000000",
            INIT_37 => X"0000004300000000000000460000000000000049000000000000004c00000000",
            INIT_38 => X"0000004800000000000000470000000000000048000000000000004700000000",
            INIT_39 => X"00000029000000000000002a000000000000003a000000000000004700000000",
            INIT_3A => X"0000003f000000000000003a0000000000000036000000000000003900000000",
            INIT_3B => X"0000006000000000000000520000000000000047000000000000004100000000",
            INIT_3C => X"00000067000000000000005d000000000000005e000000000000006900000000",
            INIT_3D => X"00000061000000000000006c000000000000006a000000000000006700000000",
            INIT_3E => X"000000500000000000000054000000000000005b000000000000005d00000000",
            INIT_3F => X"0000004d000000000000004f0000000000000050000000000000005000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000052000000000000004b0000000000000049000000000000004900000000",
            INIT_41 => X"0000002e00000000000000570000000000000067000000000000005800000000",
            INIT_42 => X"0000005200000000000000450000000000000038000000000000003800000000",
            INIT_43 => X"00000057000000000000005a0000000000000057000000000000005100000000",
            INIT_44 => X"0000005b000000000000005e0000000000000063000000000000006200000000",
            INIT_45 => X"00000066000000000000006a0000000000000066000000000000006100000000",
            INIT_46 => X"0000005c00000000000000610000000000000063000000000000005e00000000",
            INIT_47 => X"0000005f000000000000005b0000000000000059000000000000005900000000",
            INIT_48 => X"0000007b000000000000006d000000000000005f000000000000005600000000",
            INIT_49 => X"0000003300000000000000680000000000000099000000000000008800000000",
            INIT_4A => X"000000610000000000000049000000000000003b000000000000003c00000000",
            INIT_4B => X"0000005a0000000000000066000000000000006c000000000000006500000000",
            INIT_4C => X"0000005d00000000000000610000000000000061000000000000005f00000000",
            INIT_4D => X"0000006e00000000000000690000000000000063000000000000005d00000000",
            INIT_4E => X"0000006c000000000000006c0000000000000069000000000000006700000000",
            INIT_4F => X"0000006e000000000000006e000000000000006e000000000000006d00000000",
            INIT_50 => X"0000009d0000000000000096000000000000008b000000000000007f00000000",
            INIT_51 => X"00000032000000000000005700000000000000a200000000000000a000000000",
            INIT_52 => X"0000005800000000000000350000000000000038000000000000004300000000",
            INIT_53 => X"0000005a000000000000006b0000000000000070000000000000006500000000",
            INIT_54 => X"00000060000000000000005e0000000000000060000000000000005e00000000",
            INIT_55 => X"000000650000000000000060000000000000005f000000000000006000000000",
            INIT_56 => X"0000007e000000000000007d0000000000000071000000000000006800000000",
            INIT_57 => X"0000007000000000000000740000000000000077000000000000007b00000000",
            INIT_58 => X"000000a2000000000000009f000000000000009d000000000000009800000000",
            INIT_59 => X"0000002c000000000000005a000000000000009f00000000000000a000000000",
            INIT_5A => X"00000056000000000000003a0000000000000045000000000000004800000000",
            INIT_5B => X"0000005c0000000000000061000000000000005a000000000000006700000000",
            INIT_5C => X"0000005e000000000000005f0000000000000060000000000000005a00000000",
            INIT_5D => X"0000005c00000000000000570000000000000062000000000000006300000000",
            INIT_5E => X"0000008300000000000000830000000000000070000000000000006100000000",
            INIT_5F => X"0000006c00000000000000740000000000000079000000000000007f00000000",
            INIT_60 => X"0000009d00000000000000a0000000000000009e000000000000009b00000000",
            INIT_61 => X"0000003000000000000000720000000000000094000000000000009800000000",
            INIT_62 => X"00000067000000000000005e0000000000000058000000000000004400000000",
            INIT_63 => X"0000005d00000000000000580000000000000060000000000000007300000000",
            INIT_64 => X"0000005e00000000000000620000000000000065000000000000005900000000",
            INIT_65 => X"0000005500000000000000540000000000000065000000000000006300000000",
            INIT_66 => X"00000084000000000000007d000000000000006e000000000000006900000000",
            INIT_67 => X"0000005f000000000000006b0000000000000076000000000000007f00000000",
            INIT_68 => X"0000009200000000000000950000000000000094000000000000009400000000",
            INIT_69 => X"000000500000000000000088000000000000008e000000000000009000000000",
            INIT_6A => X"00000068000000000000005e0000000000000048000000000000002f00000000",
            INIT_6B => X"0000005e000000000000005c0000000000000071000000000000007200000000",
            INIT_6C => X"0000005d00000000000000610000000000000067000000000000005d00000000",
            INIT_6D => X"0000005200000000000000550000000000000061000000000000006000000000",
            INIT_6E => X"00000079000000000000006f000000000000006b000000000000006b00000000",
            INIT_6F => X"0000004d00000000000000570000000000000064000000000000007000000000",
            INIT_70 => X"0000008c000000000000008a0000000000000087000000000000008600000000",
            INIT_71 => X"0000008900000000000000970000000000000093000000000000008e00000000",
            INIT_72 => X"0000003e00000000000000320000000000000049000000000000005d00000000",
            INIT_73 => X"00000062000000000000005a000000000000005e000000000000005900000000",
            INIT_74 => X"0000006100000000000000670000000000000069000000000000006600000000",
            INIT_75 => X"000000530000000000000056000000000000005e000000000000005e00000000",
            INIT_76 => X"00000066000000000000005c0000000000000065000000000000005f00000000",
            INIT_77 => X"0000004b000000000000004a0000000000000052000000000000005f00000000",
            INIT_78 => X"00000090000000000000008b0000000000000086000000000000008300000000",
            INIT_79 => X"00000098000000000000009a000000000000009f000000000000009800000000",
            INIT_7A => X"0000003900000000000000350000000000000076000000000000009e00000000",
            INIT_7B => X"00000066000000000000005f0000000000000064000000000000006700000000",
            INIT_7C => X"0000006a000000000000006f0000000000000074000000000000006e00000000",
            INIT_7D => X"000000550000000000000057000000000000005b000000000000006100000000",
            INIT_7E => X"0000005300000000000000550000000000000062000000000000005400000000",
            INIT_7F => X"0000005f000000000000005a0000000000000055000000000000005300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "sampleifmap_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a000000000000000980000000000000090000000000000008700000000",
            INIT_01 => X"00000073000000000000008900000000000000a100000000000000a400000000",
            INIT_02 => X"0000006e00000000000000800000000000000091000000000000009d00000000",
            INIT_03 => X"000000670000000000000068000000000000007a000000000000007b00000000",
            INIT_04 => X"00000068000000000000006c000000000000006d000000000000006900000000",
            INIT_05 => X"000000570000000000000058000000000000005a000000000000006100000000",
            INIT_06 => X"000000550000000000000057000000000000005c000000000000004f00000000",
            INIT_07 => X"0000005e00000000000000690000000000000069000000000000006500000000",
            INIT_08 => X"000000a4000000000000009f000000000000009a000000000000009400000000",
            INIT_09 => X"0000007f00000000000000b000000000000000b300000000000000aa00000000",
            INIT_0A => X"00000098000000000000009d00000000000000c500000000000000b000000000",
            INIT_0B => X"0000006700000000000000800000000000000091000000000000007100000000",
            INIT_0C => X"0000006600000000000000680000000000000065000000000000006700000000",
            INIT_0D => X"00000059000000000000005b000000000000005f000000000000006100000000",
            INIT_0E => X"0000005b000000000000005b0000000000000056000000000000004f00000000",
            INIT_0F => X"0000004600000000000000560000000000000068000000000000006d00000000",
            INIT_10 => X"000000c500000000000000b200000000000000a4000000000000009b00000000",
            INIT_11 => X"000000c400000000000000f800000000000000ee00000000000000dd00000000",
            INIT_12 => X"000000b800000000000000b000000000000000c8000000000000009c00000000",
            INIT_13 => X"0000006a0000000000000089000000000000008e000000000000006c00000000",
            INIT_14 => X"0000006500000000000000640000000000000063000000000000006400000000",
            INIT_15 => X"00000059000000000000005f0000000000000063000000000000006500000000",
            INIT_16 => X"00000053000000000000005c0000000000000051000000000000005000000000",
            INIT_17 => X"0000004700000000000000490000000000000052000000000000005800000000",
            INIT_18 => X"000000f900000000000000eb00000000000000d600000000000000bf00000000",
            INIT_19 => X"000000f400000000000000fb00000000000000f600000000000000fd00000000",
            INIT_1A => X"000000c300000000000000ac000000000000009e00000000000000a000000000",
            INIT_1B => X"0000006e000000000000008b0000000000000072000000000000007100000000",
            INIT_1C => X"0000006300000000000000610000000000000062000000000000006200000000",
            INIT_1D => X"0000005c00000000000000660000000000000068000000000000006700000000",
            INIT_1E => X"000000490000000000000055000000000000004e000000000000005300000000",
            INIT_1F => X"00000048000000000000004a0000000000000050000000000000004b00000000",
            INIT_20 => X"000000fe00000000000000fd00000000000000fc00000000000000f500000000",
            INIT_21 => X"000000c900000000000000ba00000000000000bb00000000000000f300000000",
            INIT_22 => X"0000009c00000000000000970000000000000080000000000000009100000000",
            INIT_23 => X"000000720000000000000080000000000000006a000000000000007400000000",
            INIT_24 => X"0000006700000000000000650000000000000067000000000000006800000000",
            INIT_25 => X"0000005c0000000000000069000000000000006e000000000000006c00000000",
            INIT_26 => X"000000550000000000000054000000000000004c000000000000005200000000",
            INIT_27 => X"00000049000000000000004d0000000000000053000000000000004e00000000",
            INIT_28 => X"0000010000000000000000fc00000000000000fc00000000000000fb00000000",
            INIT_29 => X"00000072000000000000006b000000000000007e00000000000000e900000000",
            INIT_2A => X"0000006e00000000000000780000000000000073000000000000006900000000",
            INIT_2B => X"0000006700000000000000680000000000000063000000000000006300000000",
            INIT_2C => X"0000006b000000000000006b000000000000006e000000000000006d00000000",
            INIT_2D => X"000000560000000000000060000000000000006e000000000000007000000000",
            INIT_2E => X"00000068000000000000005a000000000000004c000000000000004e00000000",
            INIT_2F => X"0000004f00000000000000520000000000000052000000000000005b00000000",
            INIT_30 => X"000000eb00000000000000f600000000000000f800000000000000f800000000",
            INIT_31 => X"000000760000000000000072000000000000007c00000000000000c800000000",
            INIT_32 => X"0000004f00000000000000530000000000000057000000000000005d00000000",
            INIT_33 => X"00000044000000000000004b0000000000000056000000000000005000000000",
            INIT_34 => X"0000006100000000000000620000000000000064000000000000005f00000000",
            INIT_35 => X"0000006100000000000000610000000000000061000000000000006200000000",
            INIT_36 => X"0000006f000000000000005b0000000000000057000000000000005b00000000",
            INIT_37 => X"0000005200000000000000520000000000000055000000000000006e00000000",
            INIT_38 => X"0000009600000000000000b500000000000000d600000000000000eb00000000",
            INIT_39 => X"0000008400000000000000850000000000000088000000000000008a00000000",
            INIT_3A => X"0000003c0000000000000039000000000000003d000000000000006400000000",
            INIT_3B => X"0000003a00000000000000600000000000000059000000000000004300000000",
            INIT_3C => X"0000005000000000000000470000000000000045000000000000003300000000",
            INIT_3D => X"0000006500000000000000680000000000000065000000000000005e00000000",
            INIT_3E => X"0000006d000000000000005e0000000000000057000000000000005d00000000",
            INIT_3F => X"0000005100000000000000510000000000000062000000000000007700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009900000000",
            INIT_41 => X"00000067000000000000006f000000000000007a000000000000007c00000000",
            INIT_42 => X"000000340000000000000039000000000000005a000000000000006a00000000",
            INIT_43 => X"00000053000000000000006a0000000000000066000000000000004500000000",
            INIT_44 => X"00000055000000000000004d0000000000000047000000000000004000000000",
            INIT_45 => X"0000006d00000000000000660000000000000067000000000000006400000000",
            INIT_46 => X"00000063000000000000005d0000000000000057000000000000006a00000000",
            INIT_47 => X"00000050000000000000005c0000000000000073000000000000007100000000",
            INIT_48 => X"0000006d0000000000000072000000000000006f000000000000006d00000000",
            INIT_49 => X"0000006d00000000000000660000000000000061000000000000006500000000",
            INIT_4A => X"0000005500000000000000670000000000000078000000000000007500000000",
            INIT_4B => X"00000059000000000000005f0000000000000065000000000000005d00000000",
            INIT_4C => X"0000005a0000000000000052000000000000004b000000000000004a00000000",
            INIT_4D => X"0000006600000000000000690000000000000077000000000000007200000000",
            INIT_4E => X"00000062000000000000005e000000000000006b000000000000006f00000000",
            INIT_4F => X"0000004f000000000000006b0000000000000075000000000000006500000000",
            INIT_50 => X"0000005b000000000000005d0000000000000062000000000000006900000000",
            INIT_51 => X"00000071000000000000006f000000000000006a000000000000006300000000",
            INIT_52 => X"0000005f00000000000000610000000000000068000000000000007000000000",
            INIT_53 => X"0000005c0000000000000054000000000000004c000000000000005000000000",
            INIT_54 => X"00000059000000000000004f0000000000000048000000000000005100000000",
            INIT_55 => X"0000005e0000000000000069000000000000007b000000000000007500000000",
            INIT_56 => X"0000006500000000000000670000000000000067000000000000006000000000",
            INIT_57 => X"0000005a000000000000006f0000000000000069000000000000006000000000",
            INIT_58 => X"00000065000000000000005e0000000000000057000000000000005700000000",
            INIT_59 => X"00000064000000000000006b000000000000006e000000000000006c00000000",
            INIT_5A => X"0000006800000000000000560000000000000051000000000000005b00000000",
            INIT_5B => X"0000005c000000000000004c0000000000000049000000000000005d00000000",
            INIT_5C => X"0000004f000000000000004f000000000000004d000000000000005800000000",
            INIT_5D => X"00000056000000000000005d0000000000000064000000000000005b00000000",
            INIT_5E => X"000000600000000000000061000000000000005c000000000000005700000000",
            INIT_5F => X"0000006500000000000000660000000000000060000000000000006000000000",
            INIT_60 => X"0000006900000000000000670000000000000060000000000000005a00000000",
            INIT_61 => X"000000500000000000000056000000000000005f000000000000006500000000",
            INIT_62 => X"0000006a00000000000000600000000000000055000000000000005100000000",
            INIT_63 => X"0000005d00000000000000600000000000000055000000000000006200000000",
            INIT_64 => X"0000004c000000000000004f0000000000000051000000000000005800000000",
            INIT_65 => X"0000005b0000000000000054000000000000004c000000000000004700000000",
            INIT_66 => X"0000005a00000000000000530000000000000056000000000000005c00000000",
            INIT_67 => X"00000060000000000000005b0000000000000060000000000000006200000000",
            INIT_68 => X"00000056000000000000005f0000000000000063000000000000006400000000",
            INIT_69 => X"0000004f000000000000004f000000000000004f000000000000005000000000",
            INIT_6A => X"0000006c00000000000000620000000000000053000000000000005200000000",
            INIT_6B => X"0000005900000000000000610000000000000060000000000000006300000000",
            INIT_6C => X"00000051000000000000004f0000000000000054000000000000005c00000000",
            INIT_6D => X"000000590000000000000052000000000000004a000000000000004c00000000",
            INIT_6E => X"0000005600000000000000520000000000000055000000000000005a00000000",
            INIT_6F => X"000000530000000000000053000000000000005c000000000000005d00000000",
            INIT_70 => X"000000470000000000000049000000000000004e000000000000005700000000",
            INIT_71 => X"0000005300000000000000590000000000000057000000000000004d00000000",
            INIT_72 => X"0000006a0000000000000061000000000000004f000000000000005100000000",
            INIT_73 => X"0000005c00000000000000590000000000000067000000000000006400000000",
            INIT_74 => X"0000005900000000000000580000000000000057000000000000006000000000",
            INIT_75 => X"000000530000000000000054000000000000004f000000000000005200000000",
            INIT_76 => X"000000530000000000000056000000000000005a000000000000005600000000",
            INIT_77 => X"00000049000000000000004f0000000000000056000000000000005600000000",
            INIT_78 => X"000000490000000000000046000000000000003f000000000000003e00000000",
            INIT_79 => X"0000005100000000000000530000000000000056000000000000005400000000",
            INIT_7A => X"0000006b000000000000005e000000000000004a000000000000004e00000000",
            INIT_7B => X"00000058000000000000005b0000000000000068000000000000005f00000000",
            INIT_7C => X"0000005900000000000000580000000000000058000000000000005b00000000",
            INIT_7D => X"0000005300000000000000550000000000000050000000000000005500000000",
            INIT_7E => X"0000005000000000000000560000000000000059000000000000005400000000",
            INIT_7F => X"00000048000000000000004c000000000000004d000000000000004c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "sampleifmap_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000059000000000000005d000000000000005e000000000000005e00000000",
            INIT_01 => X"000000600000000000000060000000000000005a000000000000005a00000000",
            INIT_02 => X"00000065000000000000006e0000000000000066000000000000006100000000",
            INIT_03 => X"0000005200000000000000550000000000000058000000000000005e00000000",
            INIT_04 => X"000000480000000000000049000000000000004b000000000000004e00000000",
            INIT_05 => X"00000038000000000000003d0000000000000041000000000000004500000000",
            INIT_06 => X"000000270000000000000029000000000000002e000000000000003300000000",
            INIT_07 => X"00000019000000000000001d0000000000000022000000000000002800000000",
            INIT_08 => X"00000059000000000000005f000000000000005f000000000000006000000000",
            INIT_09 => X"00000062000000000000005f0000000000000059000000000000005900000000",
            INIT_0A => X"0000006b000000000000006a0000000000000060000000000000006100000000",
            INIT_0B => X"0000005200000000000000550000000000000059000000000000006000000000",
            INIT_0C => X"000000490000000000000047000000000000004b000000000000004f00000000",
            INIT_0D => X"00000035000000000000003b000000000000003d000000000000004400000000",
            INIT_0E => X"000000250000000000000027000000000000002c000000000000003100000000",
            INIT_0F => X"0000001f000000000000001f0000000000000020000000000000002600000000",
            INIT_10 => X"00000057000000000000005c000000000000005c000000000000005e00000000",
            INIT_11 => X"00000051000000000000005d000000000000005a000000000000005400000000",
            INIT_12 => X"0000006e00000000000000630000000000000060000000000000005900000000",
            INIT_13 => X"0000005400000000000000560000000000000062000000000000007000000000",
            INIT_14 => X"0000004600000000000000440000000000000049000000000000004f00000000",
            INIT_15 => X"000000300000000000000036000000000000003a000000000000003f00000000",
            INIT_16 => X"0000002b0000000000000029000000000000002b000000000000002e00000000",
            INIT_17 => X"000000310000000000000030000000000000002e000000000000002f00000000",
            INIT_18 => X"0000005a000000000000005c000000000000005d000000000000005f00000000",
            INIT_19 => X"000000390000000000000056000000000000005d000000000000005300000000",
            INIT_1A => X"000000680000000000000063000000000000006b000000000000005d00000000",
            INIT_1B => X"0000005a00000000000000650000000000000072000000000000007400000000",
            INIT_1C => X"0000004200000000000000420000000000000043000000000000004e00000000",
            INIT_1D => X"0000003900000000000000380000000000000038000000000000003e00000000",
            INIT_1E => X"000000420000000000000041000000000000003e000000000000003c00000000",
            INIT_1F => X"0000003d000000000000003f0000000000000041000000000000004300000000",
            INIT_20 => X"0000005b000000000000005b000000000000005b000000000000005c00000000",
            INIT_21 => X"0000003e00000000000000520000000000000059000000000000005300000000",
            INIT_22 => X"000000580000000000000058000000000000005f000000000000005c00000000",
            INIT_23 => X"0000006400000000000000690000000000000068000000000000005c00000000",
            INIT_24 => X"0000004800000000000000450000000000000046000000000000005b00000000",
            INIT_25 => X"000000530000000000000050000000000000004d000000000000005000000000",
            INIT_26 => X"0000005000000000000000510000000000000051000000000000005300000000",
            INIT_27 => X"0000003f0000000000000046000000000000004b000000000000004f00000000",
            INIT_28 => X"0000005900000000000000570000000000000056000000000000005800000000",
            INIT_29 => X"0000004d000000000000004c000000000000004f000000000000005200000000",
            INIT_2A => X"0000005700000000000000550000000000000052000000000000005000000000",
            INIT_2B => X"0000005f000000000000005e000000000000005e000000000000005a00000000",
            INIT_2C => X"000000630000000000000062000000000000005e000000000000006300000000",
            INIT_2D => X"0000006200000000000000600000000000000064000000000000006400000000",
            INIT_2E => X"0000005300000000000000580000000000000058000000000000005d00000000",
            INIT_2F => X"00000037000000000000003e0000000000000045000000000000004c00000000",
            INIT_30 => X"0000005400000000000000520000000000000054000000000000005500000000",
            INIT_31 => X"00000037000000000000002a000000000000003d000000000000005100000000",
            INIT_32 => X"0000005900000000000000580000000000000057000000000000005300000000",
            INIT_33 => X"00000065000000000000005d0000000000000057000000000000005b00000000",
            INIT_34 => X"0000007300000000000000700000000000000064000000000000006200000000",
            INIT_35 => X"0000006700000000000000670000000000000067000000000000006900000000",
            INIT_36 => X"0000004a000000000000004e0000000000000050000000000000005b00000000",
            INIT_37 => X"000000360000000000000039000000000000003f000000000000004400000000",
            INIT_38 => X"0000005400000000000000520000000000000053000000000000005200000000",
            INIT_39 => X"0000002c00000000000000260000000000000037000000000000004c00000000",
            INIT_3A => X"0000005100000000000000520000000000000055000000000000004c00000000",
            INIT_3B => X"00000063000000000000005b0000000000000053000000000000005000000000",
            INIT_3C => X"0000006c00000000000000610000000000000060000000000000006700000000",
            INIT_3D => X"0000005e00000000000000710000000000000072000000000000006d00000000",
            INIT_3E => X"0000004b000000000000004d000000000000004d000000000000005200000000",
            INIT_3F => X"0000003b00000000000000400000000000000044000000000000004700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005b00000000000000540000000000000052000000000000005100000000",
            INIT_41 => X"0000003100000000000000550000000000000068000000000000005e00000000",
            INIT_42 => X"00000063000000000000005b0000000000000054000000000000004900000000",
            INIT_43 => X"0000005e00000000000000650000000000000064000000000000006100000000",
            INIT_44 => X"0000006200000000000000650000000000000068000000000000006500000000",
            INIT_45 => X"000000670000000000000072000000000000006f000000000000006a00000000",
            INIT_46 => X"0000004e00000000000000520000000000000055000000000000005700000000",
            INIT_47 => X"0000004800000000000000470000000000000046000000000000004a00000000",
            INIT_48 => X"0000008000000000000000730000000000000065000000000000005c00000000",
            INIT_49 => X"000000360000000000000068000000000000009d000000000000008e00000000",
            INIT_4A => X"00000071000000000000005d0000000000000054000000000000004b00000000",
            INIT_4B => X"000000650000000000000075000000000000007c000000000000007500000000",
            INIT_4C => X"00000067000000000000006b000000000000006a000000000000006700000000",
            INIT_4D => X"000000760000000000000074000000000000006e000000000000006800000000",
            INIT_4E => X"000000540000000000000055000000000000005a000000000000006400000000",
            INIT_4F => X"0000005200000000000000550000000000000055000000000000005500000000",
            INIT_50 => X"000000a00000000000000099000000000000008e000000000000008200000000",
            INIT_51 => X"00000035000000000000005900000000000000aa00000000000000a600000000",
            INIT_52 => X"000000680000000000000046000000000000004d000000000000005000000000",
            INIT_53 => X"0000006b000000000000007f0000000000000082000000000000007700000000",
            INIT_54 => X"0000006a0000000000000069000000000000006c000000000000006a00000000",
            INIT_55 => X"00000072000000000000006e0000000000000069000000000000006a00000000",
            INIT_56 => X"0000006000000000000000620000000000000062000000000000006900000000",
            INIT_57 => X"000000550000000000000059000000000000005b000000000000005e00000000",
            INIT_58 => X"000000a400000000000000a2000000000000009f000000000000009a00000000",
            INIT_59 => X"0000002e000000000000005d00000000000000a900000000000000a700000000",
            INIT_5A => X"00000067000000000000004a0000000000000056000000000000005100000000",
            INIT_5B => X"00000072000000000000007a0000000000000070000000000000007b00000000",
            INIT_5C => X"00000067000000000000006a000000000000006d000000000000006a00000000",
            INIT_5D => X"0000006e00000000000000670000000000000069000000000000006b00000000",
            INIT_5E => X"0000006300000000000000650000000000000061000000000000006600000000",
            INIT_5F => X"00000055000000000000005a000000000000005e000000000000006000000000",
            INIT_60 => X"0000009e00000000000000a1000000000000009f000000000000009d00000000",
            INIT_61 => X"000000300000000000000075000000000000009f000000000000009e00000000",
            INIT_62 => X"00000078000000000000006c0000000000000065000000000000004900000000",
            INIT_63 => X"0000007500000000000000740000000000000078000000000000008700000000",
            INIT_64 => X"00000066000000000000006c0000000000000073000000000000006b00000000",
            INIT_65 => X"000000690000000000000064000000000000006a000000000000006900000000",
            INIT_66 => X"0000006500000000000000600000000000000060000000000000007000000000",
            INIT_67 => X"0000004c0000000000000055000000000000005d000000000000006200000000",
            INIT_68 => X"0000009300000000000000970000000000000098000000000000009900000000",
            INIT_69 => X"0000004c00000000000000870000000000000093000000000000009300000000",
            INIT_6A => X"0000007500000000000000670000000000000049000000000000002c00000000",
            INIT_6B => X"0000007100000000000000730000000000000085000000000000008300000000",
            INIT_6C => X"0000006b00000000000000710000000000000077000000000000006c00000000",
            INIT_6D => X"000000640000000000000065000000000000006a000000000000006a00000000",
            INIT_6E => X"00000062000000000000005d0000000000000069000000000000007500000000",
            INIT_6F => X"00000040000000000000004a0000000000000055000000000000005d00000000",
            INIT_70 => X"0000008e000000000000008e000000000000008e000000000000008f00000000",
            INIT_71 => X"0000008300000000000000950000000000000094000000000000008f00000000",
            INIT_72 => X"0000004600000000000000350000000000000041000000000000005400000000",
            INIT_73 => X"0000006d0000000000000068000000000000006b000000000000006300000000",
            INIT_74 => X"00000075000000000000007d000000000000007c000000000000007200000000",
            INIT_75 => X"000000620000000000000065000000000000006c000000000000006e00000000",
            INIT_76 => X"0000005a0000000000000058000000000000006f000000000000006c00000000",
            INIT_77 => X"0000003f00000000000000410000000000000048000000000000005500000000",
            INIT_78 => X"00000091000000000000008e000000000000008d000000000000008c00000000",
            INIT_79 => X"00000093000000000000009900000000000000a0000000000000009900000000",
            INIT_7A => X"0000003a0000000000000034000000000000006f000000000000009700000000",
            INIT_7B => X"0000006e00000000000000650000000000000068000000000000006a00000000",
            INIT_7C => X"0000008000000000000000870000000000000089000000000000007b00000000",
            INIT_7D => X"000000650000000000000068000000000000006c000000000000007300000000",
            INIT_7E => X"0000004e0000000000000059000000000000006f000000000000006300000000",
            INIT_7F => X"0000004d000000000000004a0000000000000048000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "sampleifmap_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000000000009b0000000000000095000000000000008f00000000",
            INIT_01 => X"00000072000000000000008800000000000000a000000000000000a400000000",
            INIT_02 => X"00000068000000000000007a000000000000008f000000000000009b00000000",
            INIT_03 => X"0000006c00000000000000660000000000000077000000000000007600000000",
            INIT_04 => X"0000008000000000000000850000000000000084000000000000007800000000",
            INIT_05 => X"0000006a000000000000006b000000000000006d000000000000007500000000",
            INIT_06 => X"000000560000000000000062000000000000006c000000000000006100000000",
            INIT_07 => X"00000044000000000000004f0000000000000054000000000000005a00000000",
            INIT_08 => X"000000a1000000000000009f000000000000009d000000000000009a00000000",
            INIT_09 => X"0000008100000000000000b000000000000000b100000000000000a700000000",
            INIT_0A => X"0000008e000000000000009700000000000000c700000000000000b300000000",
            INIT_0B => X"0000006c000000000000007b0000000000000089000000000000006800000000",
            INIT_0C => X"000000800000000000000083000000000000007e000000000000007900000000",
            INIT_0D => X"0000006e00000000000000700000000000000073000000000000007700000000",
            INIT_0E => X"0000005e000000000000006a0000000000000069000000000000006300000000",
            INIT_0F => X"000000270000000000000034000000000000004a000000000000005c00000000",
            INIT_10 => X"000000c100000000000000b000000000000000a4000000000000009d00000000",
            INIT_11 => X"000000c700000000000000f700000000000000ec00000000000000da00000000",
            INIT_12 => X"000000b100000000000000ad00000000000000ce00000000000000a300000000",
            INIT_13 => X"0000007100000000000000860000000000000088000000000000006500000000",
            INIT_14 => X"000000810000000000000082000000000000007e000000000000007700000000",
            INIT_15 => X"000000710000000000000076000000000000007a000000000000007d00000000",
            INIT_16 => X"00000050000000000000006a0000000000000067000000000000006800000000",
            INIT_17 => X"000000270000000000000025000000000000002c000000000000003e00000000",
            INIT_18 => X"000000f600000000000000e800000000000000d400000000000000c000000000",
            INIT_19 => X"000000f700000000000000fa00000000000000f200000000000000fa00000000",
            INIT_1A => X"000000c100000000000000ae00000000000000aa00000000000000a900000000",
            INIT_1B => X"00000078000000000000008b0000000000000070000000000000006e00000000",
            INIT_1C => X"000000800000000000000080000000000000007e000000000000007600000000",
            INIT_1D => X"00000074000000000000007e000000000000007f000000000000008000000000",
            INIT_1E => X"0000003e00000000000000600000000000000066000000000000006c00000000",
            INIT_1F => X"0000002b00000000000000270000000000000025000000000000002a00000000",
            INIT_20 => X"000000fb00000000000000fa00000000000000fb00000000000000f500000000",
            INIT_21 => X"000000d200000000000000be00000000000000ba00000000000000f100000000",
            INIT_22 => X"000000a0000000000000009c000000000000009200000000000000a100000000",
            INIT_23 => X"0000007a00000000000000870000000000000073000000000000007d00000000",
            INIT_24 => X"000000800000000000000081000000000000007f000000000000007800000000",
            INIT_25 => X"00000074000000000000007d000000000000007f000000000000007f00000000",
            INIT_26 => X"0000004200000000000000570000000000000062000000000000006a00000000",
            INIT_27 => X"000000290000000000000029000000000000002a000000000000002d00000000",
            INIT_28 => X"000000fe00000000000000fb00000000000000fb00000000000000fb00000000",
            INIT_29 => X"000000820000000000000074000000000000008300000000000000ea00000000",
            INIT_2A => X"0000007c0000000000000082000000000000008a000000000000007f00000000",
            INIT_2B => X"0000006b00000000000000720000000000000077000000000000007a00000000",
            INIT_2C => X"0000007f00000000000000820000000000000080000000000000007600000000",
            INIT_2D => X"0000006c000000000000006f0000000000000077000000000000007d00000000",
            INIT_2E => X"000000500000000000000052000000000000005a000000000000006300000000",
            INIT_2F => X"00000029000000000000002c000000000000002f000000000000003d00000000",
            INIT_30 => X"000000ef00000000000000f900000000000000fc00000000000000fc00000000",
            INIT_31 => X"00000083000000000000007b000000000000008000000000000000cb00000000",
            INIT_32 => X"000000670000000000000066000000000000006c000000000000006f00000000",
            INIT_33 => X"0000004400000000000000510000000000000069000000000000006a00000000",
            INIT_34 => X"0000007400000000000000780000000000000075000000000000006600000000",
            INIT_35 => X"000000730000000000000070000000000000006b000000000000006e00000000",
            INIT_36 => X"00000054000000000000004b0000000000000059000000000000006800000000",
            INIT_37 => X"0000002d000000000000002d0000000000000034000000000000005100000000",
            INIT_38 => X"000000a000000000000000bf00000000000000df00000000000000f500000000",
            INIT_39 => X"0000008a00000000000000890000000000000089000000000000009000000000",
            INIT_3A => X"000000570000000000000051000000000000004b000000000000006d00000000",
            INIT_3B => X"0000003a00000000000000630000000000000066000000000000005a00000000",
            INIT_3C => X"00000065000000000000005f0000000000000056000000000000003a00000000",
            INIT_3D => X"00000074000000000000007a0000000000000074000000000000006d00000000",
            INIT_3E => X"000000500000000000000046000000000000004d000000000000006100000000",
            INIT_3F => X"0000002f000000000000002f0000000000000042000000000000005900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000840000000000000086000000000000008d00000000000000a500000000",
            INIT_41 => X"000000690000000000000070000000000000007b000000000000008200000000",
            INIT_42 => X"00000047000000000000004a000000000000005e000000000000006b00000000",
            INIT_43 => X"00000056000000000000006f000000000000006e000000000000005300000000",
            INIT_44 => X"0000006c0000000000000066000000000000005a000000000000004800000000",
            INIT_45 => X"0000007c000000000000007b000000000000007b000000000000007600000000",
            INIT_46 => X"0000004400000000000000420000000000000049000000000000006c00000000",
            INIT_47 => X"00000030000000000000003d0000000000000054000000000000005200000000",
            INIT_48 => X"00000075000000000000007a0000000000000078000000000000007500000000",
            INIT_49 => X"0000006a00000000000000650000000000000061000000000000006a00000000",
            INIT_4A => X"00000057000000000000006a0000000000000073000000000000007000000000",
            INIT_4B => X"0000006100000000000000680000000000000068000000000000005c00000000",
            INIT_4C => X"00000072000000000000006c000000000000005f000000000000005400000000",
            INIT_4D => X"0000007a0000000000000082000000000000008e000000000000008600000000",
            INIT_4E => X"0000004000000000000000450000000000000064000000000000007700000000",
            INIT_4F => X"00000032000000000000004f0000000000000057000000000000004500000000",
            INIT_50 => X"0000005e00000000000000600000000000000066000000000000006c00000000",
            INIT_51 => X"0000006b000000000000006e000000000000006b000000000000006500000000",
            INIT_52 => X"000000510000000000000056000000000000005d000000000000006700000000",
            INIT_53 => X"00000068000000000000005d0000000000000048000000000000004200000000",
            INIT_54 => X"00000071000000000000006b000000000000005f000000000000005e00000000",
            INIT_55 => X"0000007a00000000000000850000000000000094000000000000008900000000",
            INIT_56 => X"000000420000000000000051000000000000006b000000000000007200000000",
            INIT_57 => X"0000003f0000000000000055000000000000004b000000000000004000000000",
            INIT_58 => X"00000063000000000000005d0000000000000057000000000000005800000000",
            INIT_59 => X"000000570000000000000065000000000000006c000000000000006b00000000",
            INIT_5A => X"000000530000000000000041000000000000003c000000000000004900000000",
            INIT_5B => X"0000005e000000000000004e000000000000003f000000000000004a00000000",
            INIT_5C => X"0000005d000000000000005f0000000000000057000000000000005900000000",
            INIT_5D => X"00000072000000000000007a000000000000007b000000000000006900000000",
            INIT_5E => X"0000003b000000000000004e0000000000000068000000000000006d00000000",
            INIT_5F => X"0000004b000000000000004a000000000000003f000000000000003c00000000",
            INIT_60 => X"0000005f0000000000000061000000000000005f000000000000005d00000000",
            INIT_61 => X"0000003800000000000000450000000000000054000000000000005b00000000",
            INIT_62 => X"0000005500000000000000420000000000000031000000000000003200000000",
            INIT_63 => X"0000004800000000000000550000000000000049000000000000005300000000",
            INIT_64 => X"000000440000000000000043000000000000003e000000000000003e00000000",
            INIT_65 => X"0000006800000000000000640000000000000058000000000000004500000000",
            INIT_66 => X"000000330000000000000040000000000000005a000000000000006500000000",
            INIT_67 => X"00000045000000000000003a0000000000000036000000000000003500000000",
            INIT_68 => X"000000440000000000000051000000000000005b000000000000006000000000",
            INIT_69 => X"0000003000000000000000340000000000000037000000000000003b00000000",
            INIT_6A => X"000000520000000000000040000000000000002e000000000000002f00000000",
            INIT_6B => X"00000039000000000000004d000000000000004f000000000000005200000000",
            INIT_6C => X"0000003a00000000000000340000000000000032000000000000003500000000",
            INIT_6D => X"0000004a0000000000000047000000000000003f000000000000003a00000000",
            INIT_6E => X"0000002e00000000000000340000000000000041000000000000004800000000",
            INIT_6F => X"0000003600000000000000300000000000000031000000000000003000000000",
            INIT_70 => X"0000002b0000000000000031000000000000003c000000000000004900000000",
            INIT_71 => X"0000003000000000000000340000000000000030000000000000002c00000000",
            INIT_72 => X"00000049000000000000003a000000000000002c000000000000003000000000",
            INIT_73 => X"00000035000000000000003e000000000000004f000000000000004b00000000",
            INIT_74 => X"000000390000000000000034000000000000002e000000000000003200000000",
            INIT_75 => X"0000002f0000000000000033000000000000002f000000000000003400000000",
            INIT_76 => X"0000002a000000000000002e0000000000000031000000000000002f00000000",
            INIT_77 => X"0000002a000000000000002b000000000000002d000000000000002b00000000",
            INIT_78 => X"0000002500000000000000270000000000000025000000000000002900000000",
            INIT_79 => X"0000002d00000000000000290000000000000029000000000000002a00000000",
            INIT_7A => X"000000470000000000000036000000000000002b000000000000002f00000000",
            INIT_7B => X"0000002e000000000000003b000000000000004c000000000000004300000000",
            INIT_7C => X"00000030000000000000002d000000000000002a000000000000002b00000000",
            INIT_7D => X"0000002d0000000000000031000000000000002d000000000000002f00000000",
            INIT_7E => X"00000027000000000000002a000000000000002d000000000000002b00000000",
            INIT_7F => X"0000002600000000000000280000000000000028000000000000002500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "sampleifmap_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004f00000000000000530000000000000054000000000000005500000000",
            INIT_01 => X"0000005f000000000000005d0000000000000052000000000000005000000000",
            INIT_02 => X"00000048000000000000004f0000000000000055000000000000005a00000000",
            INIT_03 => X"0000004f0000000000000054000000000000004e000000000000004b00000000",
            INIT_04 => X"0000003d000000000000003c000000000000003e000000000000004400000000",
            INIT_05 => X"000000330000000000000038000000000000003b000000000000003c00000000",
            INIT_06 => X"0000002300000000000000250000000000000029000000000000002e00000000",
            INIT_07 => X"000000150000000000000019000000000000001e000000000000002400000000",
            INIT_08 => X"0000004f00000000000000550000000000000055000000000000005600000000",
            INIT_09 => X"0000005d000000000000005a0000000000000050000000000000004e00000000",
            INIT_0A => X"0000004700000000000000460000000000000049000000000000005400000000",
            INIT_0B => X"0000004800000000000000470000000000000045000000000000004400000000",
            INIT_0C => X"0000003e000000000000003e0000000000000043000000000000004600000000",
            INIT_0D => X"0000002e00000000000000340000000000000035000000000000003800000000",
            INIT_0E => X"0000002000000000000000220000000000000025000000000000002900000000",
            INIT_0F => X"0000001b000000000000001a000000000000001b000000000000002100000000",
            INIT_10 => X"0000004e00000000000000520000000000000053000000000000005400000000",
            INIT_11 => X"0000004800000000000000560000000000000050000000000000004900000000",
            INIT_12 => X"0000004300000000000000380000000000000041000000000000004600000000",
            INIT_13 => X"0000003c0000000000000036000000000000003f000000000000004800000000",
            INIT_14 => X"0000003a000000000000003d0000000000000041000000000000004200000000",
            INIT_15 => X"00000026000000000000002d000000000000002f000000000000003000000000",
            INIT_16 => X"0000002500000000000000220000000000000021000000000000002400000000",
            INIT_17 => X"0000002c000000000000002a0000000000000029000000000000002a00000000",
            INIT_18 => X"0000005000000000000000520000000000000053000000000000005500000000",
            INIT_19 => X"0000002b000000000000004d0000000000000052000000000000004800000000",
            INIT_1A => X"0000003400000000000000320000000000000045000000000000004300000000",
            INIT_1B => X"0000002f0000000000000032000000000000003f000000000000004100000000",
            INIT_1C => X"0000003600000000000000390000000000000034000000000000003200000000",
            INIT_1D => X"0000002c000000000000002b000000000000002b000000000000002d00000000",
            INIT_1E => X"0000003b00000000000000380000000000000032000000000000002f00000000",
            INIT_1F => X"000000370000000000000038000000000000003b000000000000003c00000000",
            INIT_20 => X"0000005100000000000000510000000000000051000000000000005200000000",
            INIT_21 => X"0000002c0000000000000046000000000000004c000000000000004800000000",
            INIT_22 => X"0000001d00000000000000220000000000000033000000000000003d00000000",
            INIT_23 => X"0000002300000000000000260000000000000027000000000000001f00000000",
            INIT_24 => X"0000003b0000000000000039000000000000002b000000000000002900000000",
            INIT_25 => X"000000440000000000000041000000000000003d000000000000003d00000000",
            INIT_26 => X"0000004800000000000000470000000000000042000000000000004400000000",
            INIT_27 => X"00000038000000000000003e0000000000000043000000000000004700000000",
            INIT_28 => X"0000004f000000000000004c000000000000004c000000000000004d00000000",
            INIT_29 => X"00000038000000000000003e0000000000000042000000000000004700000000",
            INIT_2A => X"00000017000000000000001a0000000000000021000000000000002c00000000",
            INIT_2B => X"0000000e000000000000000f0000000000000014000000000000001600000000",
            INIT_2C => X"00000054000000000000004f0000000000000035000000000000001f00000000",
            INIT_2D => X"00000050000000000000004e0000000000000052000000000000005300000000",
            INIT_2E => X"0000004b000000000000004d0000000000000048000000000000004c00000000",
            INIT_2F => X"0000002e0000000000000035000000000000003c000000000000004400000000",
            INIT_30 => X"0000004800000000000000460000000000000047000000000000004900000000",
            INIT_31 => X"0000002000000000000000200000000000000037000000000000004700000000",
            INIT_32 => X"0000001300000000000000140000000000000018000000000000002600000000",
            INIT_33 => X"00000015000000000000000e000000000000000b000000000000001200000000",
            INIT_34 => X"0000005900000000000000460000000000000029000000000000001800000000",
            INIT_35 => X"00000052000000000000004f0000000000000050000000000000005600000000",
            INIT_36 => X"0000004300000000000000480000000000000048000000000000004b00000000",
            INIT_37 => X"0000002a000000000000002d0000000000000034000000000000003b00000000",
            INIT_38 => X"0000004500000000000000440000000000000045000000000000004400000000",
            INIT_39 => X"00000011000000000000001c0000000000000033000000000000004300000000",
            INIT_3A => X"0000000b000000000000000a000000000000000c000000000000001700000000",
            INIT_3B => X"000000180000000000000011000000000000000b000000000000000900000000",
            INIT_3C => X"0000003f00000000000000210000000000000016000000000000001c00000000",
            INIT_3D => X"00000040000000000000004d000000000000004f000000000000004d00000000",
            INIT_3E => X"0000004200000000000000480000000000000049000000000000004100000000",
            INIT_3F => X"0000002b000000000000002f0000000000000036000000000000003c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004e00000000000000470000000000000045000000000000004400000000",
            INIT_41 => X"000000130000000000000046000000000000005d000000000000005200000000",
            INIT_42 => X"000000250000000000000019000000000000000c000000000000001200000000",
            INIT_43 => X"0000001400000000000000210000000000000021000000000000002000000000",
            INIT_44 => X"0000002100000000000000190000000000000018000000000000001600000000",
            INIT_45 => X"0000003b000000000000003c0000000000000038000000000000003100000000",
            INIT_46 => X"0000003f0000000000000049000000000000004b000000000000003b00000000",
            INIT_47 => X"0000003500000000000000340000000000000034000000000000003900000000",
            INIT_48 => X"0000007500000000000000670000000000000059000000000000005000000000",
            INIT_49 => X"000000160000000000000055000000000000008d000000000000008000000000",
            INIT_4A => X"000000380000000000000021000000000000000f000000000000001500000000",
            INIT_4B => X"0000001c0000000000000035000000000000003d000000000000003900000000",
            INIT_4C => X"0000001400000000000000160000000000000016000000000000001500000000",
            INIT_4D => X"0000003a000000000000002d0000000000000023000000000000001800000000",
            INIT_4E => X"0000004100000000000000460000000000000048000000000000003d00000000",
            INIT_4F => X"0000003d000000000000003f0000000000000040000000000000004100000000",
            INIT_50 => X"00000095000000000000008e0000000000000083000000000000007700000000",
            INIT_51 => X"0000001800000000000000470000000000000098000000000000009800000000",
            INIT_52 => X"0000003100000000000000150000000000000011000000000000001e00000000",
            INIT_53 => X"00000021000000000000003f0000000000000044000000000000003c00000000",
            INIT_54 => X"000000110000000000000015000000000000001b000000000000001900000000",
            INIT_55 => X"0000002b000000000000001c0000000000000014000000000000000f00000000",
            INIT_56 => X"0000004a000000000000004d0000000000000046000000000000003700000000",
            INIT_57 => X"0000004100000000000000440000000000000047000000000000004900000000",
            INIT_58 => X"0000009900000000000000960000000000000094000000000000008f00000000",
            INIT_59 => X"00000017000000000000004f0000000000000099000000000000009900000000",
            INIT_5A => X"0000002e00000000000000190000000000000022000000000000002800000000",
            INIT_5B => X"0000002700000000000000370000000000000030000000000000003d00000000",
            INIT_5C => X"00000015000000000000001f0000000000000024000000000000001d00000000",
            INIT_5D => X"0000001f00000000000000120000000000000015000000000000001300000000",
            INIT_5E => X"0000004d000000000000004c000000000000003b000000000000002a00000000",
            INIT_5F => X"00000045000000000000004a000000000000004c000000000000004d00000000",
            INIT_60 => X"0000009400000000000000970000000000000095000000000000009200000000",
            INIT_61 => X"00000020000000000000006b0000000000000092000000000000009200000000",
            INIT_62 => X"0000003b00000000000000340000000000000037000000000000002b00000000",
            INIT_63 => X"00000029000000000000002c0000000000000034000000000000004700000000",
            INIT_64 => X"0000001e000000000000002c0000000000000032000000000000002200000000",
            INIT_65 => X"000000190000000000000012000000000000001c000000000000001a00000000",
            INIT_66 => X"0000005100000000000000450000000000000032000000000000002e00000000",
            INIT_67 => X"000000420000000000000049000000000000004f000000000000005100000000",
            INIT_68 => X"0000008b000000000000008f000000000000008f000000000000009000000000",
            INIT_69 => X"00000040000000000000007e0000000000000089000000000000008a00000000",
            INIT_6A => X"00000041000000000000003d000000000000002e000000000000001a00000000",
            INIT_6B => X"0000002400000000000000280000000000000040000000000000004600000000",
            INIT_6C => X"0000002800000000000000330000000000000036000000000000002400000000",
            INIT_6D => X"000000130000000000000012000000000000001d000000000000002100000000",
            INIT_6E => X"0000004e000000000000003c0000000000000033000000000000002f00000000",
            INIT_6F => X"000000370000000000000040000000000000004a000000000000004f00000000",
            INIT_70 => X"0000008600000000000000860000000000000084000000000000008500000000",
            INIT_71 => X"0000007700000000000000890000000000000088000000000000008600000000",
            INIT_72 => X"00000021000000000000001b0000000000000031000000000000004700000000",
            INIT_73 => X"000000220000000000000020000000000000002a000000000000002e00000000",
            INIT_74 => X"00000032000000000000003d0000000000000039000000000000002800000000",
            INIT_75 => X"000000110000000000000011000000000000001c000000000000002700000000",
            INIT_76 => X"0000004100000000000000300000000000000033000000000000002400000000",
            INIT_77 => X"000000320000000000000036000000000000003e000000000000004600000000",
            INIT_78 => X"000000850000000000000081000000000000007f000000000000007d00000000",
            INIT_79 => X"0000008100000000000000880000000000000091000000000000008c00000000",
            INIT_7A => X"0000001e000000000000001e000000000000005a000000000000008400000000",
            INIT_7B => X"0000002700000000000000270000000000000033000000000000004000000000",
            INIT_7C => X"0000003d00000000000000450000000000000045000000000000003100000000",
            INIT_7D => X"000000130000000000000014000000000000001c000000000000002c00000000",
            INIT_7E => X"0000002d00000000000000290000000000000030000000000000001900000000",
            INIT_7F => X"0000003d000000000000003c0000000000000039000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "sampleifmap_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000091000000000000008b0000000000000084000000000000007d00000000",
            INIT_01 => X"0000005a00000000000000750000000000000091000000000000009500000000",
            INIT_02 => X"0000005000000000000000620000000000000072000000000000008000000000",
            INIT_03 => X"000000280000000000000031000000000000004d000000000000005700000000",
            INIT_04 => X"0000003c0000000000000044000000000000003f000000000000002e00000000",
            INIT_05 => X"000000170000000000000019000000000000001f000000000000002d00000000",
            INIT_06 => X"0000002d000000000000002b000000000000002a000000000000001500000000",
            INIT_07 => X"00000032000000000000003e0000000000000042000000000000004000000000",
            INIT_08 => X"000000930000000000000090000000000000008c000000000000008800000000",
            INIT_09 => X"00000068000000000000009e00000000000000a4000000000000009a00000000",
            INIT_0A => X"00000077000000000000007a00000000000000a6000000000000009500000000",
            INIT_0B => X"00000029000000000000004b0000000000000067000000000000005000000000",
            INIT_0C => X"0000003c00000000000000410000000000000038000000000000002d00000000",
            INIT_0D => X"0000001b000000000000001f0000000000000028000000000000003000000000",
            INIT_0E => X"00000032000000000000002f0000000000000023000000000000001500000000",
            INIT_0F => X"0000001400000000000000230000000000000039000000000000004100000000",
            INIT_10 => X"000000b600000000000000a40000000000000097000000000000009000000000",
            INIT_11 => X"000000b200000000000000eb00000000000000e600000000000000d200000000",
            INIT_12 => X"00000095000000000000008a00000000000000ab000000000000008500000000",
            INIT_13 => X"0000002d00000000000000550000000000000067000000000000004d00000000",
            INIT_14 => X"0000003c000000000000003f0000000000000038000000000000002b00000000",
            INIT_15 => X"0000001d00000000000000270000000000000030000000000000003500000000",
            INIT_16 => X"00000027000000000000002f000000000000001d000000000000001700000000",
            INIT_17 => X"000000150000000000000016000000000000001f000000000000002700000000",
            INIT_18 => X"000000f000000000000000e100000000000000cd00000000000000b700000000",
            INIT_19 => X"000000e600000000000000f200000000000000f200000000000000f800000000",
            INIT_1A => X"0000009f00000000000000840000000000000084000000000000008d00000000",
            INIT_1B => X"000000310000000000000056000000000000004d000000000000005300000000",
            INIT_1C => X"0000003a000000000000003c0000000000000037000000000000002a00000000",
            INIT_1D => X"00000021000000000000002f0000000000000037000000000000003900000000",
            INIT_1E => X"0000001c0000000000000027000000000000001a000000000000001900000000",
            INIT_1F => X"0000001b000000000000001c000000000000001d000000000000001900000000",
            INIT_20 => X"000000f900000000000000f700000000000000f800000000000000f100000000",
            INIT_21 => X"000000b500000000000000ab00000000000000b000000000000000ec00000000",
            INIT_22 => X"0000007600000000000000720000000000000062000000000000007800000000",
            INIT_23 => X"000000340000000000000047000000000000003c000000000000004d00000000",
            INIT_24 => X"0000003a00000000000000390000000000000036000000000000002e00000000",
            INIT_25 => X"0000002000000000000000300000000000000039000000000000003b00000000",
            INIT_26 => X"0000002500000000000000250000000000000017000000000000001800000000",
            INIT_27 => X"0000001a000000000000001f0000000000000020000000000000001c00000000",
            INIT_28 => X"000000fd00000000000000f900000000000000f900000000000000f800000000",
            INIT_29 => X"000000550000000000000053000000000000006a00000000000000e000000000",
            INIT_2A => X"000000410000000000000051000000000000004e000000000000004700000000",
            INIT_2B => X"000000310000000000000034000000000000002e000000000000003000000000",
            INIT_2C => X"0000003900000000000000360000000000000037000000000000003300000000",
            INIT_2D => X"0000001b00000000000000240000000000000033000000000000003d00000000",
            INIT_2E => X"0000003600000000000000270000000000000016000000000000001500000000",
            INIT_2F => X"0000001c000000000000001f000000000000001f000000000000002800000000",
            INIT_30 => X"000000eb00000000000000f500000000000000f800000000000000f700000000",
            INIT_31 => X"0000005e0000000000000060000000000000006d00000000000000c200000000",
            INIT_32 => X"0000001900000000000000230000000000000035000000000000004100000000",
            INIT_33 => X"00000020000000000000002d000000000000002b000000000000001c00000000",
            INIT_34 => X"0000002f000000000000002f0000000000000033000000000000002e00000000",
            INIT_35 => X"00000029000000000000002b000000000000002d000000000000003000000000",
            INIT_36 => X"0000003a0000000000000024000000000000001e000000000000002200000000",
            INIT_37 => X"0000001e000000000000001d0000000000000021000000000000003900000000",
            INIT_38 => X"0000009800000000000000b600000000000000d700000000000000ec00000000",
            INIT_39 => X"00000074000000000000007a0000000000000081000000000000008800000000",
            INIT_3A => X"00000009000000000000000d0000000000000023000000000000005100000000",
            INIT_3B => X"0000002200000000000000490000000000000034000000000000001400000000",
            INIT_3C => X"00000020000000000000001a000000000000001c000000000000001100000000",
            INIT_3D => X"00000031000000000000003b000000000000003b000000000000002f00000000",
            INIT_3E => X"000000340000000000000022000000000000001a000000000000002300000000",
            INIT_3F => X"0000001d000000000000001c000000000000002c000000000000003f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000078000000000000007a0000000000000082000000000000009a00000000",
            INIT_41 => X"0000005c00000000000000680000000000000076000000000000007b00000000",
            INIT_42 => X"00000012000000000000001f0000000000000046000000000000005a00000000",
            INIT_43 => X"000000340000000000000045000000000000003d000000000000001d00000000",
            INIT_44 => X"0000002800000000000000240000000000000024000000000000002200000000",
            INIT_45 => X"0000003d00000000000000410000000000000047000000000000003a00000000",
            INIT_46 => X"00000028000000000000001f0000000000000017000000000000003000000000",
            INIT_47 => X"0000001c0000000000000027000000000000003c000000000000003800000000",
            INIT_48 => X"00000068000000000000006d000000000000006b000000000000006900000000",
            INIT_49 => X"0000005d000000000000005b0000000000000058000000000000005f00000000",
            INIT_4A => X"0000003e00000000000000560000000000000062000000000000006000000000",
            INIT_4B => X"00000031000000000000002f0000000000000038000000000000003800000000",
            INIT_4C => X"00000030000000000000002a0000000000000025000000000000002800000000",
            INIT_4D => X"000000390000000000000048000000000000005b000000000000004c00000000",
            INIT_4E => X"00000023000000000000001d000000000000002c000000000000003600000000",
            INIT_4F => X"0000001d0000000000000037000000000000003d000000000000002a00000000",
            INIT_50 => X"0000005100000000000000530000000000000059000000000000005f00000000",
            INIT_51 => X"00000058000000000000005b0000000000000058000000000000005600000000",
            INIT_52 => X"0000003e00000000000000440000000000000049000000000000005300000000",
            INIT_53 => X"00000034000000000000002c0000000000000023000000000000002800000000",
            INIT_54 => X"000000310000000000000027000000000000001e000000000000002800000000",
            INIT_55 => X"000000320000000000000047000000000000005f000000000000005100000000",
            INIT_56 => X"000000230000000000000025000000000000002a000000000000002900000000",
            INIT_57 => X"00000028000000000000003a0000000000000030000000000000002200000000",
            INIT_58 => X"00000055000000000000004f0000000000000049000000000000004b00000000",
            INIT_59 => X"00000040000000000000004c0000000000000053000000000000005700000000",
            INIT_5A => X"0000003b000000000000002a0000000000000027000000000000003300000000",
            INIT_5B => X"0000003100000000000000290000000000000022000000000000003200000000",
            INIT_5C => X"000000270000000000000024000000000000001e000000000000002600000000",
            INIT_5D => X"0000002d000000000000003c0000000000000045000000000000003700000000",
            INIT_5E => X"0000001d00000000000000220000000000000026000000000000002600000000",
            INIT_5F => X"0000003300000000000000300000000000000024000000000000002000000000",
            INIT_60 => X"0000004d000000000000004f000000000000004e000000000000004c00000000",
            INIT_61 => X"00000021000000000000002c0000000000000039000000000000004400000000",
            INIT_62 => X"0000003d000000000000002e000000000000001e000000000000001d00000000",
            INIT_63 => X"0000002600000000000000320000000000000029000000000000003700000000",
            INIT_64 => X"0000001e000000000000001d000000000000001a000000000000001d00000000",
            INIT_65 => X"00000030000000000000002e0000000000000025000000000000001d00000000",
            INIT_66 => X"0000001800000000000000190000000000000025000000000000002e00000000",
            INIT_67 => X"0000002f00000000000000240000000000000020000000000000001e00000000",
            INIT_68 => X"000000320000000000000040000000000000004a000000000000005000000000",
            INIT_69 => X"0000001b000000000000001e0000000000000020000000000000002600000000",
            INIT_6A => X"0000003c000000000000002d000000000000001b000000000000001b00000000",
            INIT_6B => X"0000001d000000000000002c000000000000002f000000000000003500000000",
            INIT_6C => X"0000001c00000000000000170000000000000017000000000000001c00000000",
            INIT_6D => X"0000002500000000000000200000000000000018000000000000001900000000",
            INIT_6E => X"000000150000000000000015000000000000001d000000000000002300000000",
            INIT_6F => X"00000022000000000000001c000000000000001e000000000000001a00000000",
            INIT_70 => X"0000001a0000000000000021000000000000002d000000000000003a00000000",
            INIT_71 => X"0000001c0000000000000021000000000000001d000000000000001a00000000",
            INIT_72 => X"0000003300000000000000270000000000000018000000000000001b00000000",
            INIT_73 => X"0000001c00000000000000210000000000000032000000000000003100000000",
            INIT_74 => X"0000001d00000000000000190000000000000015000000000000001b00000000",
            INIT_75 => X"0000001700000000000000190000000000000015000000000000001800000000",
            INIT_76 => X"000000120000000000000016000000000000001a000000000000001700000000",
            INIT_77 => X"000000170000000000000019000000000000001a000000000000001500000000",
            INIT_78 => X"0000001500000000000000180000000000000017000000000000001b00000000",
            INIT_79 => X"0000001900000000000000180000000000000019000000000000001a00000000",
            INIT_7A => X"0000003000000000000000210000000000000016000000000000001a00000000",
            INIT_7B => X"0000001800000000000000230000000000000033000000000000002a00000000",
            INIT_7C => X"0000001800000000000000150000000000000014000000000000001500000000",
            INIT_7D => X"00000019000000000000001d0000000000000017000000000000001700000000",
            INIT_7E => X"000000120000000000000016000000000000001b000000000000001800000000",
            INIT_7F => X"0000001600000000000000180000000000000016000000000000001100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "sampleifmap_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004100000000000000150000000000000013000000000000001700000000",
            INIT_01 => X"000000b200000000000000b700000000000000bc00000000000000a400000000",
            INIT_02 => X"000000ba00000000000000ba00000000000000ac00000000000000aa00000000",
            INIT_03 => X"000000b700000000000000b600000000000000b700000000000000b800000000",
            INIT_04 => X"0000005c000000000000007f00000000000000a400000000000000b400000000",
            INIT_05 => X"000000c20000000000000099000000000000006e000000000000006b00000000",
            INIT_06 => X"000000c600000000000000c500000000000000c900000000000000c300000000",
            INIT_07 => X"000000c500000000000000c700000000000000c800000000000000c900000000",
            INIT_08 => X"0000002e00000000000000150000000000000013000000000000001700000000",
            INIT_09 => X"000000b200000000000000bf00000000000000ca000000000000009900000000",
            INIT_0A => X"000000b700000000000000a9000000000000009e00000000000000a400000000",
            INIT_0B => X"000000b200000000000000b400000000000000b800000000000000ba00000000",
            INIT_0C => X"00000056000000000000008a00000000000000ad00000000000000b400000000",
            INIT_0D => X"000000ce00000000000000b4000000000000006a000000000000004a00000000",
            INIT_0E => X"000000ce00000000000000d000000000000000d500000000000000cf00000000",
            INIT_0F => X"000000ca00000000000000cc00000000000000cd00000000000000cf00000000",
            INIT_10 => X"0000001f00000000000000170000000000000014000000000000001700000000",
            INIT_11 => X"000000a800000000000000b900000000000000c8000000000000007f00000000",
            INIT_12 => X"000000a2000000000000009a000000000000009e000000000000009f00000000",
            INIT_13 => X"000000b200000000000000b300000000000000b200000000000000b200000000",
            INIT_14 => X"0000007d00000000000000b600000000000000be00000000000000b500000000",
            INIT_15 => X"000000d100000000000000c50000000000000072000000000000004700000000",
            INIT_16 => X"000000d300000000000000d500000000000000d800000000000000d500000000",
            INIT_17 => X"000000ce00000000000000d000000000000000d300000000000000d400000000",
            INIT_18 => X"0000001700000000000000180000000000000015000000000000001700000000",
            INIT_19 => X"000000a000000000000000af00000000000000bd000000000000006300000000",
            INIT_1A => X"0000009500000000000000a600000000000000a800000000000000a800000000",
            INIT_1B => X"000000c300000000000000bf00000000000000ba00000000000000aa00000000",
            INIT_1C => X"0000008d00000000000000bc00000000000000c800000000000000c300000000",
            INIT_1D => X"000000d600000000000000d20000000000000092000000000000006300000000",
            INIT_1E => X"000000d500000000000000d400000000000000d400000000000000d500000000",
            INIT_1F => X"000000d600000000000000d700000000000000d900000000000000d900000000",
            INIT_20 => X"0000001500000000000000170000000000000017000000000000001900000000",
            INIT_21 => X"0000009700000000000000a500000000000000aa000000000000004800000000",
            INIT_22 => X"0000009b00000000000000b900000000000000b700000000000000af00000000",
            INIT_23 => X"000000bc00000000000000a9000000000000009d000000000000009200000000",
            INIT_24 => X"0000008d00000000000000b200000000000000c400000000000000c500000000",
            INIT_25 => X"000000db00000000000000d300000000000000ac000000000000007900000000",
            INIT_26 => X"000000d900000000000000d900000000000000d900000000000000dd00000000",
            INIT_27 => X"000000ce00000000000000d100000000000000d400000000000000d600000000",
            INIT_28 => X"00000017000000000000001a000000000000001b000000000000001a00000000",
            INIT_29 => X"0000009a00000000000000a4000000000000008f000000000000003100000000",
            INIT_2A => X"000000a600000000000000c800000000000000c200000000000000a900000000",
            INIT_2B => X"000000970000000000000080000000000000007d000000000000008200000000",
            INIT_2C => X"0000008f000000000000009400000000000000a500000000000000a500000000",
            INIT_2D => X"000000c900000000000000bc00000000000000b6000000000000009300000000",
            INIT_2E => X"000000db00000000000000d500000000000000d900000000000000d400000000",
            INIT_2F => X"000000d300000000000000d700000000000000d700000000000000dc00000000",
            INIT_30 => X"00000019000000000000001b000000000000001a000000000000001e00000000",
            INIT_31 => X"000000ab00000000000000b4000000000000007d000000000000002500000000",
            INIT_32 => X"000000b300000000000000ca00000000000000c500000000000000a900000000",
            INIT_33 => X"00000082000000000000007a0000000000000071000000000000008b00000000",
            INIT_34 => X"0000008c000000000000007a0000000000000085000000000000007700000000",
            INIT_35 => X"000000c900000000000000bf00000000000000cb00000000000000b900000000",
            INIT_36 => X"000000db00000000000000d700000000000000da00000000000000d700000000",
            INIT_37 => X"000000e000000000000000dc00000000000000da00000000000000dc00000000",
            INIT_38 => X"00000024000000000000001f0000000000000030000000000000005e00000000",
            INIT_39 => X"000000a800000000000000c100000000000000af000000000000006400000000",
            INIT_3A => X"000000c300000000000000c600000000000000c000000000000000a300000000",
            INIT_3B => X"00000084000000000000008e000000000000009100000000000000ae00000000",
            INIT_3C => X"0000008b000000000000007a0000000000000079000000000000006a00000000",
            INIT_3D => X"000000d500000000000000bd00000000000000d100000000000000c000000000",
            INIT_3E => X"000000e800000000000000ef00000000000000ed00000000000000f200000000",
            INIT_3F => X"000000e500000000000000de00000000000000d500000000000000d000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007a0000000000000072000000000000009e00000000000000b400000000",
            INIT_41 => X"000000a000000000000000be00000000000000be00000000000000b100000000",
            INIT_42 => X"000000c800000000000000c500000000000000ad000000000000008500000000",
            INIT_43 => X"0000009200000000000000a700000000000000b900000000000000c200000000",
            INIT_44 => X"0000008d00000000000000850000000000000081000000000000008100000000",
            INIT_45 => X"000000dc00000000000000bd00000000000000c900000000000000b100000000",
            INIT_46 => X"000000d500000000000000e800000000000000eb00000000000000f100000000",
            INIT_47 => X"000000ea00000000000000e100000000000000c700000000000000bd00000000",
            INIT_48 => X"000000ba00000000000000b200000000000000c000000000000000c500000000",
            INIT_49 => X"0000009d00000000000000c500000000000000c300000000000000c100000000",
            INIT_4A => X"000000bf00000000000000b900000000000000a3000000000000008000000000",
            INIT_4B => X"0000009700000000000000b200000000000000c300000000000000c100000000",
            INIT_4C => X"0000008600000000000000830000000000000081000000000000007200000000",
            INIT_4D => X"000000ea00000000000000d000000000000000c200000000000000aa00000000",
            INIT_4E => X"000000c900000000000000eb00000000000000f000000000000000ec00000000",
            INIT_4F => X"000000eb00000000000000d000000000000000bb00000000000000b900000000",
            INIT_50 => X"000000c000000000000000bb00000000000000c400000000000000ca00000000",
            INIT_51 => X"0000009700000000000000c500000000000000cd00000000000000c800000000",
            INIT_52 => X"000000bd00000000000000b800000000000000af000000000000009500000000",
            INIT_53 => X"0000008800000000000000a800000000000000bb00000000000000c100000000",
            INIT_54 => X"0000008100000000000000800000000000000080000000000000007500000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b500000000000000a700000000",
            INIT_56 => X"000000ce00000000000000ee00000000000000f300000000000000f300000000",
            INIT_57 => X"000000dd00000000000000c100000000000000bb00000000000000ba00000000",
            INIT_58 => X"000000c000000000000000c500000000000000cd00000000000000cd00000000",
            INIT_59 => X"000000a000000000000000c200000000000000d000000000000000cb00000000",
            INIT_5A => X"000000bf00000000000000c100000000000000bf00000000000000a800000000",
            INIT_5B => X"00000077000000000000009200000000000000ac00000000000000c100000000",
            INIT_5C => X"000000870000000000000085000000000000008e000000000000007c00000000",
            INIT_5D => X"000000ea00000000000000bf00000000000000b000000000000000a700000000",
            INIT_5E => X"000000d700000000000000ec00000000000000f100000000000000f300000000",
            INIT_5F => X"000000c400000000000000b900000000000000b800000000000000ba00000000",
            INIT_60 => X"000000c100000000000000c800000000000000cc00000000000000ce00000000",
            INIT_61 => X"000000b400000000000000bf00000000000000c700000000000000c500000000",
            INIT_62 => X"000000ad00000000000000b700000000000000b300000000000000ac00000000",
            INIT_63 => X"00000083000000000000009800000000000000ae00000000000000ae00000000",
            INIT_64 => X"0000009a000000000000008e00000000000000a6000000000000008d00000000",
            INIT_65 => X"000000e600000000000000bf00000000000000ac00000000000000a900000000",
            INIT_66 => X"000000e400000000000000ef00000000000000f100000000000000f000000000",
            INIT_67 => X"000000c000000000000000b800000000000000ba00000000000000c800000000",
            INIT_68 => X"000000bf00000000000000c600000000000000ca00000000000000d200000000",
            INIT_69 => X"000000ca00000000000000b100000000000000b400000000000000c900000000",
            INIT_6A => X"0000008e000000000000008e000000000000009a00000000000000ab00000000",
            INIT_6B => X"0000009c000000000000009300000000000000a800000000000000a800000000",
            INIT_6C => X"000000a4000000000000009600000000000000a900000000000000af00000000",
            INIT_6D => X"000000e600000000000000c500000000000000a0000000000000009e00000000",
            INIT_6E => X"000000f200000000000000f400000000000000f100000000000000f100000000",
            INIT_6F => X"000000d700000000000000c300000000000000bf00000000000000e200000000",
            INIT_70 => X"000000c000000000000000c700000000000000c900000000000000d300000000",
            INIT_71 => X"000000d700000000000000a100000000000000aa00000000000000cf00000000",
            INIT_72 => X"000000ac00000000000000ad00000000000000ba00000000000000bd00000000",
            INIT_73 => X"0000007f000000000000008900000000000000b100000000000000be00000000",
            INIT_74 => X"000000a0000000000000009600000000000000ae00000000000000b400000000",
            INIT_75 => X"000000ec00000000000000c100000000000000b000000000000000af00000000",
            INIT_76 => X"000000fb00000000000000f300000000000000f200000000000000f500000000",
            INIT_77 => X"000000e100000000000000d400000000000000c900000000000000ef00000000",
            INIT_78 => X"000000c100000000000000c500000000000000c400000000000000d300000000",
            INIT_79 => X"000000d9000000000000009a00000000000000b500000000000000d100000000",
            INIT_7A => X"000000b900000000000000c300000000000000c500000000000000ce00000000",
            INIT_7B => X"0000009800000000000000a600000000000000ad00000000000000aa00000000",
            INIT_7C => X"0000009800000000000000a600000000000000b800000000000000a300000000",
            INIT_7D => X"000000cc00000000000000af00000000000000b500000000000000c000000000",
            INIT_7E => X"000000f700000000000000f400000000000000f300000000000000ee00000000",
            INIT_7F => X"000000e200000000000000e200000000000000d500000000000000df00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "sampleifmap_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b500000000000000b400000000000000c200000000000000d600000000",
            INIT_01 => X"000000c6000000000000009b00000000000000c400000000000000c500000000",
            INIT_02 => X"000000b700000000000000ae00000000000000c000000000000000d600000000",
            INIT_03 => X"000000b200000000000000ae00000000000000a100000000000000ad00000000",
            INIT_04 => X"0000009300000000000000bd00000000000000a4000000000000008000000000",
            INIT_05 => X"00000076000000000000009c00000000000000b400000000000000a700000000",
            INIT_06 => X"000000eb00000000000000ef00000000000000d7000000000000009d00000000",
            INIT_07 => X"000000e400000000000000ea00000000000000d600000000000000ce00000000",
            INIT_08 => X"000000a300000000000000a600000000000000c600000000000000d700000000",
            INIT_09 => X"000000b900000000000000be00000000000000ca00000000000000b400000000",
            INIT_0A => X"000000d600000000000000cd00000000000000d200000000000000cf00000000",
            INIT_0B => X"000000ad00000000000000b000000000000000ae00000000000000c100000000",
            INIT_0C => X"0000009900000000000000bf0000000000000089000000000000008100000000",
            INIT_0D => X"0000008700000000000000ab00000000000000c800000000000000a300000000",
            INIT_0E => X"000000c100000000000000b80000000000000090000000000000007400000000",
            INIT_0F => X"000000eb00000000000000ef00000000000000d200000000000000bb00000000",
            INIT_10 => X"000000a400000000000000ae00000000000000cd00000000000000d800000000",
            INIT_11 => X"000000c200000000000000d200000000000000cb00000000000000b900000000",
            INIT_12 => X"000000e200000000000000da00000000000000d300000000000000bf00000000",
            INIT_13 => X"000000b300000000000000be00000000000000cb00000000000000e100000000",
            INIT_14 => X"0000009e00000000000000a80000000000000079000000000000009700000000",
            INIT_15 => X"000000ac00000000000000aa00000000000000c200000000000000a700000000",
            INIT_16 => X"000000a900000000000000990000000000000083000000000000009a00000000",
            INIT_17 => X"000000ec00000000000000de00000000000000b800000000000000a200000000",
            INIT_18 => X"000000b400000000000000c000000000000000d000000000000000d800000000",
            INIT_19 => X"000000d200000000000000d100000000000000ca00000000000000c500000000",
            INIT_1A => X"000000cc00000000000000c500000000000000bd00000000000000ba00000000",
            INIT_1B => X"000000b500000000000000cf00000000000000d500000000000000d100000000",
            INIT_1C => X"000000af0000000000000092000000000000009500000000000000b200000000",
            INIT_1D => X"000000ab000000000000009c00000000000000ae00000000000000b700000000",
            INIT_1E => X"000000b400000000000000a9000000000000009400000000000000a300000000",
            INIT_1F => X"000000cc00000000000000ac00000000000000a000000000000000a600000000",
            INIT_20 => X"000000b600000000000000ca00000000000000d500000000000000da00000000",
            INIT_21 => X"000000ca00000000000000c900000000000000cb00000000000000bf00000000",
            INIT_22 => X"000000c000000000000000c100000000000000c300000000000000ca00000000",
            INIT_23 => X"000000c700000000000000cf00000000000000c600000000000000b200000000",
            INIT_24 => X"000000bb00000000000000a600000000000000cb00000000000000d300000000",
            INIT_25 => X"000000a60000000000000093000000000000009b00000000000000b100000000",
            INIT_26 => X"000000af00000000000000b600000000000000ab00000000000000a700000000",
            INIT_27 => X"000000a7000000000000009f000000000000009c000000000000009c00000000",
            INIT_28 => X"000000ba00000000000000d100000000000000d700000000000000d900000000",
            INIT_29 => X"000000c800000000000000d000000000000000c800000000000000b300000000",
            INIT_2A => X"000000ba00000000000000d200000000000000d700000000000000d100000000",
            INIT_2B => X"000000c200000000000000c400000000000000b600000000000000a100000000",
            INIT_2C => X"000000b900000000000000be00000000000000cf00000000000000cb00000000",
            INIT_2D => X"000000a6000000000000009b000000000000008e000000000000009b00000000",
            INIT_2E => X"0000009f00000000000000ad00000000000000b300000000000000ac00000000",
            INIT_2F => X"0000008f000000000000009e000000000000009e000000000000009600000000",
            INIT_30 => X"000000c000000000000000d600000000000000d500000000000000d600000000",
            INIT_31 => X"000000d900000000000000da00000000000000c500000000000000a900000000",
            INIT_32 => X"000000c300000000000000d400000000000000d900000000000000d700000000",
            INIT_33 => X"000000bf00000000000000c300000000000000b300000000000000aa00000000",
            INIT_34 => X"000000aa00000000000000c000000000000000c000000000000000be00000000",
            INIT_35 => X"000000aa00000000000000a7000000000000008e000000000000008400000000",
            INIT_36 => X"0000009d00000000000000ad00000000000000b300000000000000aa00000000",
            INIT_37 => X"0000007d00000000000000860000000000000093000000000000009d00000000",
            INIT_38 => X"000000ca00000000000000d300000000000000d100000000000000d500000000",
            INIT_39 => X"000000de00000000000000d800000000000000c100000000000000a800000000",
            INIT_3A => X"000000cd00000000000000d300000000000000de00000000000000df00000000",
            INIT_3B => X"000000c600000000000000c900000000000000c200000000000000c200000000",
            INIT_3C => X"0000009900000000000000bc00000000000000c400000000000000c600000000",
            INIT_3D => X"000000a700000000000000ab000000000000009b000000000000008600000000",
            INIT_3E => X"000000a500000000000000b200000000000000bd00000000000000a600000000",
            INIT_3F => X"000000890000000000000085000000000000008e00000000000000a300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000ca00000000000000ce00000000000000ce00000000000000d300000000",
            INIT_41 => X"000000d500000000000000d300000000000000bf00000000000000af00000000",
            INIT_42 => X"000000ab00000000000000c600000000000000d800000000000000d600000000",
            INIT_43 => X"000000c900000000000000c900000000000000ce00000000000000c200000000",
            INIT_44 => X"0000009600000000000000b100000000000000c500000000000000c800000000",
            INIT_45 => X"0000009d00000000000000a7000000000000009e000000000000009000000000",
            INIT_46 => X"000000a800000000000000b000000000000000b5000000000000009f00000000",
            INIT_47 => X"0000009000000000000000950000000000000096000000000000009800000000",
            INIT_48 => X"000000c100000000000000c900000000000000cc00000000000000d200000000",
            INIT_49 => X"000000d200000000000000d000000000000000bc00000000000000b500000000",
            INIT_4A => X"0000007a00000000000000a000000000000000ce00000000000000cd00000000",
            INIT_4B => X"000000c200000000000000c600000000000000d000000000000000b100000000",
            INIT_4C => X"0000009600000000000000a600000000000000b800000000000000c100000000",
            INIT_4D => X"0000009900000000000000a0000000000000009c000000000000008b00000000",
            INIT_4E => X"0000009b000000000000009f00000000000000a0000000000000009b00000000",
            INIT_4F => X"00000083000000000000008c0000000000000098000000000000009800000000",
            INIT_50 => X"000000bb00000000000000c600000000000000ca00000000000000d200000000",
            INIT_51 => X"000000d600000000000000cd00000000000000b200000000000000ae00000000",
            INIT_52 => X"0000008300000000000000a400000000000000cb00000000000000d100000000",
            INIT_53 => X"000000b600000000000000bb00000000000000ca00000000000000b400000000",
            INIT_54 => X"0000008b000000000000009d00000000000000a900000000000000b600000000",
            INIT_55 => X"00000090000000000000009a0000000000000099000000000000008600000000",
            INIT_56 => X"0000008d0000000000000083000000000000008d000000000000009700000000",
            INIT_57 => X"000000930000000000000096000000000000009b000000000000009d00000000",
            INIT_58 => X"000000b500000000000000c200000000000000c800000000000000d200000000",
            INIT_59 => X"000000d700000000000000c400000000000000a800000000000000a800000000",
            INIT_5A => X"000000b800000000000000bd00000000000000c700000000000000d400000000",
            INIT_5B => X"000000ac00000000000000ad00000000000000b900000000000000cb00000000",
            INIT_5C => X"000000760000000000000093000000000000009b00000000000000a300000000",
            INIT_5D => X"0000008d00000000000000910000000000000094000000000000008300000000",
            INIT_5E => X"00000085000000000000007f0000000000000084000000000000009000000000",
            INIT_5F => X"0000009c00000000000000a200000000000000a3000000000000009500000000",
            INIT_60 => X"000000b400000000000000bd00000000000000c200000000000000d000000000",
            INIT_61 => X"000000d300000000000000bd000000000000009e00000000000000a200000000",
            INIT_62 => X"000000c700000000000000c200000000000000c500000000000000d300000000",
            INIT_63 => X"000000a400000000000000a300000000000000ac00000000000000bf00000000",
            INIT_64 => X"0000006d00000000000000820000000000000093000000000000009e00000000",
            INIT_65 => X"0000009100000000000000900000000000000090000000000000008900000000",
            INIT_66 => X"00000086000000000000007c0000000000000084000000000000009000000000",
            INIT_67 => X"00000093000000000000009f00000000000000a2000000000000009700000000",
            INIT_68 => X"000000b500000000000000b000000000000000b100000000000000c200000000",
            INIT_69 => X"000000cd00000000000000b3000000000000008f000000000000009f00000000",
            INIT_6A => X"000000be00000000000000c200000000000000c700000000000000d000000000",
            INIT_6B => X"000000a1000000000000009c00000000000000a500000000000000b500000000",
            INIT_6C => X"0000007200000000000000700000000000000088000000000000009500000000",
            INIT_6D => X"00000092000000000000008a0000000000000085000000000000008900000000",
            INIT_6E => X"0000009000000000000000830000000000000083000000000000009200000000",
            INIT_6F => X"0000008d00000000000000940000000000000095000000000000009600000000",
            INIT_70 => X"000000b200000000000000a5000000000000009d00000000000000ac00000000",
            INIT_71 => X"000000c7000000000000009c000000000000008500000000000000a700000000",
            INIT_72 => X"000000c200000000000000c700000000000000c700000000000000ce00000000",
            INIT_73 => X"0000008b0000000000000084000000000000008500000000000000a000000000",
            INIT_74 => X"0000007e000000000000006b000000000000007e000000000000008c00000000",
            INIT_75 => X"00000095000000000000008a0000000000000081000000000000008200000000",
            INIT_76 => X"0000008e0000000000000091000000000000008c000000000000008d00000000",
            INIT_77 => X"000000980000000000000095000000000000008c000000000000008800000000",
            INIT_78 => X"0000009b00000000000000900000000000000086000000000000009700000000",
            INIT_79 => X"000000b70000000000000082000000000000007d000000000000009e00000000",
            INIT_7A => X"000000a500000000000000b700000000000000bf00000000000000c500000000",
            INIT_7B => X"00000069000000000000005e0000000000000067000000000000008000000000",
            INIT_7C => X"0000007c00000000000000750000000000000070000000000000007700000000",
            INIT_7D => X"0000008f000000000000008b000000000000007d000000000000007900000000",
            INIT_7E => X"0000007d0000000000000081000000000000008c000000000000008b00000000",
            INIT_7F => X"00000096000000000000009b0000000000000095000000000000008400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "sampleifmap_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002f00000000000000100000000000000015000000000000001300000000",
            INIT_01 => X"0000008e00000000000000930000000000000093000000000000008300000000",
            INIT_02 => X"0000008e00000000000000900000000000000089000000000000008700000000",
            INIT_03 => X"0000008f000000000000008c000000000000008c000000000000008d00000000",
            INIT_04 => X"000000490000000000000060000000000000007e000000000000008c00000000",
            INIT_05 => X"000000a40000000000000082000000000000005d000000000000005f00000000",
            INIT_06 => X"0000009d000000000000009b000000000000009c000000000000009b00000000",
            INIT_07 => X"000000970000000000000098000000000000009b000000000000009e00000000",
            INIT_08 => X"0000001f00000000000000110000000000000014000000000000001400000000",
            INIT_09 => X"00000092000000000000009b00000000000000a1000000000000007a00000000",
            INIT_0A => X"00000095000000000000008b0000000000000088000000000000008a00000000",
            INIT_0B => X"0000009700000000000000920000000000000096000000000000009800000000",
            INIT_0C => X"0000004900000000000000750000000000000096000000000000009f00000000",
            INIT_0D => X"000000af000000000000009c0000000000000058000000000000004100000000",
            INIT_0E => X"000000ad00000000000000ab00000000000000a900000000000000a800000000",
            INIT_0F => X"000000a300000000000000a400000000000000a800000000000000ac00000000",
            INIT_10 => X"0000001500000000000000140000000000000014000000000000001400000000",
            INIT_11 => X"0000008c000000000000009700000000000000a2000000000000006600000000",
            INIT_12 => X"0000008b00000000000000880000000000000095000000000000008d00000000",
            INIT_13 => X"0000009f00000000000000980000000000000099000000000000009a00000000",
            INIT_14 => X"0000006d00000000000000a100000000000000ab00000000000000a600000000",
            INIT_15 => X"000000b700000000000000b10000000000000061000000000000003a00000000",
            INIT_16 => X"000000b200000000000000b100000000000000b200000000000000b300000000",
            INIT_17 => X"000000a600000000000000a900000000000000ad00000000000000b100000000",
            INIT_18 => X"0000001100000000000000150000000000000014000000000000001400000000",
            INIT_19 => X"00000082000000000000008c0000000000000099000000000000004f00000000",
            INIT_1A => X"00000087000000000000009d00000000000000a4000000000000009700000000",
            INIT_1B => X"000000b000000000000000a900000000000000a6000000000000009900000000",
            INIT_1C => X"0000007600000000000000a100000000000000af00000000000000b000000000",
            INIT_1D => X"000000c300000000000000c40000000000000085000000000000005200000000",
            INIT_1E => X"000000b300000000000000b400000000000000b700000000000000bd00000000",
            INIT_1F => X"000000ab00000000000000ad00000000000000b100000000000000b300000000",
            INIT_20 => X"0000001300000000000000150000000000000014000000000000001500000000",
            INIT_21 => X"0000007700000000000000820000000000000089000000000000003800000000",
            INIT_22 => X"0000009200000000000000b300000000000000b2000000000000009c00000000",
            INIT_23 => X"000000a70000000000000094000000000000008b000000000000008400000000",
            INIT_24 => X"00000078000000000000009800000000000000a900000000000000af00000000",
            INIT_25 => X"000000d200000000000000ce00000000000000a7000000000000006d00000000",
            INIT_26 => X"000000bf00000000000000c300000000000000c900000000000000d100000000",
            INIT_27 => X"000000ac00000000000000b100000000000000b600000000000000ba00000000",
            INIT_28 => X"0000001600000000000000170000000000000016000000000000001600000000",
            INIT_29 => X"0000007800000000000000820000000000000073000000000000002600000000",
            INIT_2A => X"0000009e00000000000000c300000000000000b9000000000000009200000000",
            INIT_2B => X"00000084000000000000006b000000000000006c000000000000007600000000",
            INIT_2C => X"000000840000000000000081000000000000008f000000000000009200000000",
            INIT_2D => X"000000c700000000000000be00000000000000b7000000000000008f00000000",
            INIT_2E => X"000000d100000000000000cc00000000000000d100000000000000cf00000000",
            INIT_2F => X"000000c200000000000000c700000000000000ca00000000000000d100000000",
            INIT_30 => X"0000001400000000000000150000000000000013000000000000001800000000",
            INIT_31 => X"0000009400000000000000a10000000000000071000000000000001e00000000",
            INIT_32 => X"000000aa00000000000000c200000000000000ba000000000000009700000000",
            INIT_33 => X"0000007100000000000000690000000000000062000000000000008000000000",
            INIT_34 => X"00000080000000000000006b0000000000000074000000000000006800000000",
            INIT_35 => X"000000c500000000000000c000000000000000ca00000000000000b200000000",
            INIT_36 => X"000000d700000000000000d100000000000000cf00000000000000ce00000000",
            INIT_37 => X"000000da00000000000000d700000000000000d600000000000000d800000000",
            INIT_38 => X"0000001d00000000000000180000000000000029000000000000005800000000",
            INIT_39 => X"0000009c00000000000000ba00000000000000ae000000000000006000000000",
            INIT_3A => X"000000ba00000000000000bd00000000000000b5000000000000009500000000",
            INIT_3B => X"000000760000000000000081000000000000008400000000000000a400000000",
            INIT_3C => X"0000007c000000000000006c000000000000006b000000000000005c00000000",
            INIT_3D => X"000000ce00000000000000bb00000000000000cc00000000000000b400000000",
            INIT_3E => X"000000e400000000000000e700000000000000e000000000000000e600000000",
            INIT_3F => X"000000e200000000000000dc00000000000000d300000000000000cd00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000075000000000000006d000000000000009900000000000000b100000000",
            INIT_41 => X"0000009300000000000000b700000000000000bd00000000000000af00000000",
            INIT_42 => X"000000c000000000000000bc00000000000000a1000000000000007800000000",
            INIT_43 => X"00000083000000000000009a00000000000000ad00000000000000b800000000",
            INIT_44 => X"0000007f00000000000000770000000000000073000000000000007300000000",
            INIT_45 => X"000000d800000000000000bc00000000000000c500000000000000a600000000",
            INIT_46 => X"000000d300000000000000e300000000000000e200000000000000e900000000",
            INIT_47 => X"000000e800000000000000e000000000000000c600000000000000bc00000000",
            INIT_48 => X"000000b600000000000000af00000000000000bc00000000000000c200000000",
            INIT_49 => X"0000009000000000000000be00000000000000c200000000000000bf00000000",
            INIT_4A => X"000000b600000000000000b10000000000000098000000000000007300000000",
            INIT_4B => X"0000008a00000000000000a400000000000000b600000000000000b700000000",
            INIT_4C => X"0000007b00000000000000770000000000000076000000000000006600000000",
            INIT_4D => X"000000e900000000000000d000000000000000bd00000000000000a000000000",
            INIT_4E => X"000000cb00000000000000ea00000000000000eb00000000000000e800000000",
            INIT_4F => X"000000eb00000000000000d100000000000000bd00000000000000bb00000000",
            INIT_50 => X"000000bb00000000000000b700000000000000c000000000000000c700000000",
            INIT_51 => X"0000008a00000000000000bf00000000000000cd00000000000000c600000000",
            INIT_52 => X"000000b500000000000000b000000000000000a5000000000000008800000000",
            INIT_53 => X"0000007c000000000000009a00000000000000af00000000000000b800000000",
            INIT_54 => X"0000007800000000000000770000000000000076000000000000006b00000000",
            INIT_55 => X"000000f000000000000000cd00000000000000b0000000000000009e00000000",
            INIT_56 => X"000000d400000000000000f200000000000000f400000000000000f300000000",
            INIT_57 => X"000000e000000000000000c600000000000000c000000000000000c000000000",
            INIT_58 => X"000000bb00000000000000c100000000000000c900000000000000c900000000",
            INIT_59 => X"0000009200000000000000bc00000000000000d100000000000000c900000000",
            INIT_5A => X"000000b700000000000000b900000000000000b6000000000000009b00000000",
            INIT_5B => X"0000006b0000000000000084000000000000009f00000000000000b700000000",
            INIT_5C => X"0000007e000000000000007c0000000000000085000000000000007300000000",
            INIT_5D => X"000000eb00000000000000bd00000000000000aa000000000000009e00000000",
            INIT_5E => X"000000de00000000000000f200000000000000f600000000000000f600000000",
            INIT_5F => X"000000ca00000000000000c000000000000000c000000000000000c200000000",
            INIT_60 => X"000000bd00000000000000c500000000000000c900000000000000cb00000000",
            INIT_61 => X"000000a500000000000000b700000000000000c600000000000000c400000000",
            INIT_62 => X"000000a500000000000000b000000000000000aa000000000000009f00000000",
            INIT_63 => X"00000078000000000000008a00000000000000a200000000000000a400000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008500000000",
            INIT_65 => X"000000e700000000000000bd00000000000000a500000000000000a100000000",
            INIT_66 => X"000000ea00000000000000f700000000000000f800000000000000f400000000",
            INIT_67 => X"000000c700000000000000c100000000000000c300000000000000d000000000",
            INIT_68 => X"000000b900000000000000c400000000000000ca00000000000000d000000000",
            INIT_69 => X"000000b9000000000000009c00000000000000a700000000000000c100000000",
            INIT_6A => X"000000870000000000000087000000000000009100000000000000a100000000",
            INIT_6B => X"0000008f0000000000000089000000000000009e00000000000000a100000000",
            INIT_6C => X"000000a2000000000000009500000000000000a400000000000000a400000000",
            INIT_6D => X"000000e400000000000000c3000000000000009d000000000000009900000000",
            INIT_6E => X"000000f500000000000000f900000000000000f700000000000000f200000000",
            INIT_6F => X"000000de00000000000000cc00000000000000c700000000000000e800000000",
            INIT_70 => X"000000b600000000000000c500000000000000cc00000000000000d200000000",
            INIT_71 => X"000000c1000000000000007d000000000000008e00000000000000bf00000000",
            INIT_72 => X"000000a700000000000000a600000000000000b100000000000000b500000000",
            INIT_73 => X"00000072000000000000008200000000000000aa00000000000000b800000000",
            INIT_74 => X"0000009e000000000000009800000000000000aa00000000000000a500000000",
            INIT_75 => X"000000e700000000000000bd00000000000000ae00000000000000ab00000000",
            INIT_76 => X"000000fb00000000000000f500000000000000f400000000000000f200000000",
            INIT_77 => X"000000e900000000000000dd00000000000000cf00000000000000f200000000",
            INIT_78 => X"000000b900000000000000c500000000000000c800000000000000d400000000",
            INIT_79 => X"000000c00000000000000070000000000000009100000000000000bd00000000",
            INIT_7A => X"000000b400000000000000bd00000000000000be00000000000000c700000000",
            INIT_7B => X"0000008900000000000000a000000000000000a700000000000000a400000000",
            INIT_7C => X"0000009100000000000000a200000000000000b0000000000000009200000000",
            INIT_7D => X"000000c300000000000000a800000000000000b100000000000000b800000000",
            INIT_7E => X"000000f900000000000000f500000000000000f100000000000000e800000000",
            INIT_7F => X"000000eb00000000000000ec00000000000000dd00000000000000e400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "sampleifmap_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ae00000000000000b600000000000000c700000000000000d800000000",
            INIT_01 => X"000000ad000000000000006e000000000000009b00000000000000b000000000",
            INIT_02 => X"000000b200000000000000a800000000000000ba00000000000000d000000000",
            INIT_03 => X"000000a400000000000000a7000000000000009b00000000000000a800000000",
            INIT_04 => X"0000008600000000000000b10000000000000096000000000000006e00000000",
            INIT_05 => X"00000068000000000000009000000000000000ab000000000000009a00000000",
            INIT_06 => X"000000ed00000000000000ee00000000000000d1000000000000009100000000",
            INIT_07 => X"000000ed00000000000000f300000000000000dd00000000000000d200000000",
            INIT_08 => X"0000009e00000000000000a900000000000000ce00000000000000db00000000",
            INIT_09 => X"000000a2000000000000009500000000000000a700000000000000a300000000",
            INIT_0A => X"000000d100000000000000c800000000000000cd00000000000000ca00000000",
            INIT_0B => X"000000a100000000000000aa00000000000000a800000000000000bc00000000",
            INIT_0C => X"0000008700000000000000ad0000000000000078000000000000007000000000",
            INIT_0D => X"00000073000000000000009b00000000000000ba000000000000009300000000",
            INIT_0E => X"000000bc00000000000000b20000000000000084000000000000006200000000",
            INIT_0F => X"000000ef00000000000000f300000000000000d400000000000000b900000000",
            INIT_10 => X"000000a100000000000000b300000000000000d600000000000000dd00000000",
            INIT_11 => X"000000b100000000000000b300000000000000b500000000000000af00000000",
            INIT_12 => X"000000dd00000000000000d400000000000000cf00000000000000bd00000000",
            INIT_13 => X"000000ab00000000000000b800000000000000c500000000000000dc00000000",
            INIT_14 => X"0000008c00000000000000950000000000000067000000000000008b00000000",
            INIT_15 => X"00000093000000000000009400000000000000b1000000000000009700000000",
            INIT_16 => X"0000009c000000000000008a0000000000000070000000000000008300000000",
            INIT_17 => X"000000ea00000000000000d900000000000000b1000000000000009700000000",
            INIT_18 => X"000000b200000000000000c600000000000000da00000000000000df00000000",
            INIT_19 => X"000000c800000000000000be00000000000000c200000000000000c200000000",
            INIT_1A => X"000000c700000000000000bf00000000000000b800000000000000ba00000000",
            INIT_1B => X"000000b100000000000000c800000000000000d000000000000000cb00000000",
            INIT_1C => X"0000009e000000000000007f000000000000008700000000000000ab00000000",
            INIT_1D => X"0000008f0000000000000083000000000000009b00000000000000a800000000",
            INIT_1E => X"0000009f0000000000000094000000000000007e000000000000008900000000",
            INIT_1F => X"000000c5000000000000009e0000000000000090000000000000009300000000",
            INIT_20 => X"000000b700000000000000d000000000000000dd00000000000000e100000000",
            INIT_21 => X"000000c200000000000000be00000000000000c700000000000000bf00000000",
            INIT_22 => X"000000ba00000000000000be00000000000000bc00000000000000c600000000",
            INIT_23 => X"000000bf00000000000000c600000000000000c100000000000000ab00000000",
            INIT_24 => X"000000a9000000000000009400000000000000bf00000000000000cf00000000",
            INIT_25 => X"0000008d000000000000007b000000000000008700000000000000a000000000",
            INIT_26 => X"00000098000000000000009f0000000000000095000000000000008e00000000",
            INIT_27 => X"0000009a000000000000008c0000000000000088000000000000008700000000",
            INIT_28 => X"000000be00000000000000d600000000000000dd00000000000000de00000000",
            INIT_29 => X"000000be00000000000000c800000000000000c300000000000000b300000000",
            INIT_2A => X"000000b200000000000000d100000000000000cd00000000000000c600000000",
            INIT_2B => X"000000b500000000000000b600000000000000b3000000000000009700000000",
            INIT_2C => X"000000a500000000000000ae00000000000000c400000000000000c500000000",
            INIT_2D => X"000000930000000000000089000000000000007c000000000000008600000000",
            INIT_2E => X"0000008b000000000000009900000000000000a1000000000000009900000000",
            INIT_2F => X"0000007d000000000000008b000000000000008b000000000000008300000000",
            INIT_30 => X"000000c600000000000000db00000000000000da00000000000000db00000000",
            INIT_31 => X"000000cf00000000000000d200000000000000bf00000000000000aa00000000",
            INIT_32 => X"000000b400000000000000cf00000000000000ce00000000000000cb00000000",
            INIT_33 => X"000000b000000000000000b400000000000000ae000000000000009c00000000",
            INIT_34 => X"0000009600000000000000b000000000000000b500000000000000b600000000",
            INIT_35 => X"000000980000000000000096000000000000007d000000000000006f00000000",
            INIT_36 => X"0000008a000000000000009a00000000000000a1000000000000009800000000",
            INIT_37 => X"0000006a00000000000000730000000000000080000000000000008a00000000",
            INIT_38 => X"000000cf00000000000000d900000000000000d600000000000000da00000000",
            INIT_39 => X"000000d500000000000000d200000000000000bc00000000000000aa00000000",
            INIT_3A => X"000000b600000000000000c700000000000000d300000000000000d400000000",
            INIT_3B => X"000000b500000000000000ba00000000000000ba00000000000000ae00000000",
            INIT_3C => X"0000008500000000000000ab00000000000000b600000000000000ba00000000",
            INIT_3D => X"00000095000000000000009a0000000000000089000000000000007200000000",
            INIT_3E => X"00000092000000000000009f00000000000000ab000000000000009400000000",
            INIT_3F => X"000000760000000000000073000000000000007b000000000000009000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000d100000000000000d400000000000000d400000000000000d800000000",
            INIT_41 => X"000000cd00000000000000cf00000000000000bd00000000000000b300000000",
            INIT_42 => X"0000008a00000000000000b100000000000000cd00000000000000cd00000000",
            INIT_43 => X"000000b600000000000000bb00000000000000c300000000000000a700000000",
            INIT_44 => X"00000082000000000000009e00000000000000b500000000000000b900000000",
            INIT_45 => X"0000008c0000000000000096000000000000008d000000000000007d00000000",
            INIT_46 => X"00000095000000000000009d00000000000000a3000000000000008d00000000",
            INIT_47 => X"0000007c00000000000000820000000000000083000000000000008500000000",
            INIT_48 => X"000000c800000000000000d000000000000000d200000000000000d700000000",
            INIT_49 => X"000000cc00000000000000ce00000000000000be00000000000000bb00000000",
            INIT_4A => X"00000050000000000000008300000000000000c400000000000000c600000000",
            INIT_4B => X"000000ae00000000000000b800000000000000c2000000000000009100000000",
            INIT_4C => X"00000083000000000000009300000000000000a500000000000000ae00000000",
            INIT_4D => X"00000088000000000000008f000000000000008b000000000000007800000000",
            INIT_4E => X"00000088000000000000008c000000000000008e000000000000008900000000",
            INIT_4F => X"0000007000000000000000790000000000000085000000000000008500000000",
            INIT_50 => X"000000c200000000000000cd00000000000000d000000000000000d700000000",
            INIT_51 => X"000000d100000000000000cd00000000000000b700000000000000b500000000",
            INIT_52 => X"00000051000000000000008100000000000000c200000000000000cc00000000",
            INIT_53 => X"000000a100000000000000ab00000000000000ba000000000000008e00000000",
            INIT_54 => X"000000780000000000000089000000000000009500000000000000a100000000",
            INIT_55 => X"0000007e00000000000000890000000000000087000000000000007300000000",
            INIT_56 => X"0000007a0000000000000070000000000000007b000000000000008500000000",
            INIT_57 => X"0000008000000000000000830000000000000088000000000000008a00000000",
            INIT_58 => X"000000bc00000000000000c800000000000000cd00000000000000d600000000",
            INIT_59 => X"000000d400000000000000c600000000000000af00000000000000b000000000",
            INIT_5A => X"0000008e00000000000000a000000000000000c000000000000000d000000000",
            INIT_5B => X"00000095000000000000009b00000000000000a800000000000000aa00000000",
            INIT_5C => X"00000064000000000000007f0000000000000085000000000000008d00000000",
            INIT_5D => X"0000007b00000000000000800000000000000083000000000000007100000000",
            INIT_5E => X"00000072000000000000006c0000000000000072000000000000007e00000000",
            INIT_5F => X"0000008900000000000000900000000000000090000000000000008200000000",
            INIT_60 => X"000000b700000000000000c000000000000000c400000000000000d200000000",
            INIT_61 => X"000000d200000000000000c000000000000000a600000000000000a900000000",
            INIT_62 => X"000000b400000000000000b600000000000000c000000000000000d100000000",
            INIT_63 => X"0000008c000000000000008d000000000000009900000000000000ab00000000",
            INIT_64 => X"0000005c000000000000006f000000000000007d000000000000008600000000",
            INIT_65 => X"0000007f000000000000007e000000000000007e000000000000007800000000",
            INIT_66 => X"0000007400000000000000690000000000000072000000000000007e00000000",
            INIT_67 => X"00000081000000000000008d0000000000000090000000000000008500000000",
            INIT_68 => X"000000b900000000000000b300000000000000b300000000000000c400000000",
            INIT_69 => X"000000cc00000000000000b5000000000000009700000000000000a600000000",
            INIT_6A => X"000000b300000000000000ba00000000000000c200000000000000cd00000000",
            INIT_6B => X"000000880000000000000085000000000000009200000000000000a600000000",
            INIT_6C => X"00000061000000000000005d0000000000000072000000000000007e00000000",
            INIT_6D => X"0000008000000000000000780000000000000073000000000000007800000000",
            INIT_6E => X"0000007e00000000000000710000000000000071000000000000008000000000",
            INIT_6F => X"0000007b00000000000000820000000000000083000000000000008400000000",
            INIT_70 => X"000000b800000000000000aa00000000000000a100000000000000b100000000",
            INIT_71 => X"000000c3000000000000009c000000000000008c00000000000000ae00000000",
            INIT_72 => X"000000b600000000000000bf00000000000000c100000000000000c900000000",
            INIT_73 => X"00000073000000000000006c0000000000000071000000000000009100000000",
            INIT_74 => X"0000006e0000000000000059000000000000006a000000000000007600000000",
            INIT_75 => X"0000008300000000000000780000000000000070000000000000007200000000",
            INIT_76 => X"0000007c000000000000007f000000000000007a000000000000007b00000000",
            INIT_77 => X"000000860000000000000082000000000000007a000000000000007500000000",
            INIT_78 => X"000000a10000000000000097000000000000008c000000000000009d00000000",
            INIT_79 => X"000000b10000000000000080000000000000008200000000000000a600000000",
            INIT_7A => X"0000009a00000000000000af00000000000000b700000000000000bf00000000",
            INIT_7B => X"0000005300000000000000470000000000000053000000000000007000000000",
            INIT_7C => X"0000006e0000000000000065000000000000005e000000000000006300000000",
            INIT_7D => X"0000007e0000000000000079000000000000006c000000000000006c00000000",
            INIT_7E => X"0000006b000000000000006f000000000000007a000000000000007900000000",
            INIT_7F => X"0000008400000000000000890000000000000084000000000000007300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "sampleifmap_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000280000000000000013000000000000001c000000000000001700000000",
            INIT_01 => X"00000074000000000000006d0000000000000073000000000000007100000000",
            INIT_02 => X"00000069000000000000006a0000000000000067000000000000007100000000",
            INIT_03 => X"0000006b00000000000000690000000000000069000000000000006900000000",
            INIT_04 => X"0000003a000000000000004c0000000000000063000000000000006a00000000",
            INIT_05 => X"0000008900000000000000720000000000000056000000000000005400000000",
            INIT_06 => X"0000007d000000000000007c000000000000007d000000000000007c00000000",
            INIT_07 => X"00000078000000000000007a000000000000007d000000000000007f00000000",
            INIT_08 => X"0000001a0000000000000014000000000000001b000000000000001800000000",
            INIT_09 => X"0000007c00000000000000760000000000000082000000000000006a00000000",
            INIT_0A => X"00000075000000000000006d0000000000000072000000000000007d00000000",
            INIT_0B => X"0000007900000000000000720000000000000076000000000000007800000000",
            INIT_0C => X"00000044000000000000006a0000000000000083000000000000008500000000",
            INIT_0D => X"00000096000000000000008c0000000000000051000000000000003e00000000",
            INIT_0E => X"000000880000000000000089000000000000008c000000000000008a00000000",
            INIT_0F => X"0000008000000000000000810000000000000085000000000000008800000000",
            INIT_10 => X"000000120000000000000017000000000000001a000000000000001800000000",
            INIT_11 => X"0000007b00000000000000740000000000000083000000000000005800000000",
            INIT_12 => X"000000740000000000000074000000000000008d000000000000008b00000000",
            INIT_13 => X"00000084000000000000007d000000000000007f000000000000008100000000",
            INIT_14 => X"000000690000000000000098000000000000009a000000000000008e00000000",
            INIT_15 => X"0000009e000000000000009f0000000000000059000000000000003700000000",
            INIT_16 => X"0000008e00000000000000920000000000000097000000000000009700000000",
            INIT_17 => X"000000840000000000000088000000000000008b000000000000008e00000000",
            INIT_18 => X"0000001200000000000000190000000000000019000000000000001800000000",
            INIT_19 => X"00000073000000000000006a000000000000007c000000000000004500000000",
            INIT_1A => X"00000078000000000000009200000000000000a6000000000000009c00000000",
            INIT_1B => X"0000009700000000000000950000000000000094000000000000008900000000",
            INIT_1C => X"0000006d0000000000000094000000000000009c000000000000009600000000",
            INIT_1D => X"000000a900000000000000b1000000000000007a000000000000004a00000000",
            INIT_1E => X"000000950000000000000098000000000000009d00000000000000a100000000",
            INIT_1F => X"0000008e00000000000000910000000000000094000000000000009600000000",
            INIT_20 => X"0000001700000000000000190000000000000018000000000000001900000000",
            INIT_21 => X"000000680000000000000060000000000000006d000000000000003300000000",
            INIT_22 => X"0000008d00000000000000b200000000000000b800000000000000a100000000",
            INIT_23 => X"0000009300000000000000860000000000000080000000000000007c00000000",
            INIT_24 => X"0000006c00000000000000890000000000000096000000000000009700000000",
            INIT_25 => X"000000b500000000000000b70000000000000098000000000000006000000000",
            INIT_26 => X"000000a400000000000000a800000000000000ae00000000000000b300000000",
            INIT_27 => X"000000930000000000000098000000000000009c00000000000000a000000000",
            INIT_28 => X"0000001c000000000000001b000000000000001a000000000000001a00000000",
            INIT_29 => X"00000066000000000000005f0000000000000059000000000000002300000000",
            INIT_2A => X"0000009f00000000000000c700000000000000c1000000000000009600000000",
            INIT_2B => X"0000007600000000000000620000000000000066000000000000007400000000",
            INIT_2C => X"0000007a00000000000000770000000000000083000000000000008200000000",
            INIT_2D => X"000000aa00000000000000a600000000000000a7000000000000008400000000",
            INIT_2E => X"000000b700000000000000b300000000000000b700000000000000b200000000",
            INIT_2F => X"000000a900000000000000af00000000000000b100000000000000b700000000",
            INIT_30 => X"0000001a00000000000000190000000000000016000000000000001a00000000",
            INIT_31 => X"0000007b0000000000000080000000000000005c000000000000001d00000000",
            INIT_32 => X"000000ab00000000000000c700000000000000c3000000000000009300000000",
            INIT_33 => X"0000006a0000000000000063000000000000005e000000000000007e00000000",
            INIT_34 => X"0000007a0000000000000065000000000000006d000000000000006000000000",
            INIT_35 => X"000000b000000000000000aa00000000000000c000000000000000ac00000000",
            INIT_36 => X"000000ca00000000000000c500000000000000c400000000000000c300000000",
            INIT_37 => X"000000c200000000000000bf00000000000000bf00000000000000c500000000",
            INIT_38 => X"0000001900000000000000110000000000000021000000000000004d00000000",
            INIT_39 => X"0000007e000000000000009b000000000000009a000000000000005800000000",
            INIT_3A => X"000000b900000000000000c100000000000000be000000000000008c00000000",
            INIT_3B => X"00000071000000000000007b000000000000008100000000000000a300000000",
            INIT_3C => X"0000007900000000000000680000000000000067000000000000005800000000",
            INIT_3D => X"000000bd00000000000000a500000000000000c600000000000000b100000000",
            INIT_3E => X"000000da00000000000000e000000000000000db00000000000000e400000000",
            INIT_3F => X"000000cd00000000000000c400000000000000bb00000000000000ba00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006000000000000000560000000000000080000000000000009500000000",
            INIT_41 => X"00000077000000000000009900000000000000a7000000000000009b00000000",
            INIT_42 => X"000000bf00000000000000bf00000000000000a8000000000000006f00000000",
            INIT_43 => X"0000007f000000000000009400000000000000aa00000000000000b700000000",
            INIT_44 => X"0000007c00000000000000740000000000000070000000000000007000000000",
            INIT_45 => X"000000c100000000000000a200000000000000bb00000000000000a300000000",
            INIT_46 => X"000000bb00000000000000cf00000000000000d500000000000000df00000000",
            INIT_47 => X"000000d200000000000000c400000000000000a6000000000000009d00000000",
            INIT_48 => X"0000009b0000000000000092000000000000009e00000000000000a100000000",
            INIT_49 => X"00000075000000000000009f00000000000000a900000000000000a700000000",
            INIT_4A => X"000000b500000000000000b3000000000000009b000000000000006800000000",
            INIT_4B => X"00000087000000000000009f00000000000000b400000000000000b600000000",
            INIT_4C => X"0000007900000000000000750000000000000074000000000000006400000000",
            INIT_4D => X"000000cc00000000000000b200000000000000b2000000000000009e00000000",
            INIT_4E => X"000000a700000000000000cb00000000000000d600000000000000d800000000",
            INIT_4F => X"000000cf00000000000000b00000000000000096000000000000009300000000",
            INIT_50 => X"000000a5000000000000009e00000000000000a500000000000000aa00000000",
            INIT_51 => X"0000007000000000000000a000000000000000b000000000000000af00000000",
            INIT_52 => X"000000b400000000000000b100000000000000a4000000000000007b00000000",
            INIT_53 => X"00000079000000000000009500000000000000ac00000000000000b600000000",
            INIT_54 => X"0000007600000000000000750000000000000074000000000000006a00000000",
            INIT_55 => X"000000d100000000000000af00000000000000a6000000000000009c00000000",
            INIT_56 => X"000000a900000000000000cd00000000000000d800000000000000de00000000",
            INIT_57 => X"000000ba000000000000009f0000000000000093000000000000009100000000",
            INIT_58 => X"000000a600000000000000a900000000000000ae00000000000000ac00000000",
            INIT_59 => X"0000007a000000000000009d00000000000000b000000000000000b000000000",
            INIT_5A => X"000000b600000000000000b900000000000000b1000000000000008d00000000",
            INIT_5B => X"00000068000000000000007f000000000000009d00000000000000b600000000",
            INIT_5C => X"0000007d000000000000007b0000000000000084000000000000007300000000",
            INIT_5D => X"000000ce00000000000000a300000000000000a4000000000000009f00000000",
            INIT_5E => X"000000b500000000000000cd00000000000000d900000000000000e000000000",
            INIT_5F => X"0000009c0000000000000093000000000000008e000000000000009200000000",
            INIT_60 => X"000000a000000000000000a500000000000000a700000000000000a700000000",
            INIT_61 => X"0000008f000000000000009900000000000000a400000000000000a500000000",
            INIT_62 => X"000000a400000000000000ae00000000000000a3000000000000009100000000",
            INIT_63 => X"000000760000000000000085000000000000009f00000000000000a300000000",
            INIT_64 => X"000000920000000000000087000000000000009f000000000000008600000000",
            INIT_65 => X"000000cd00000000000000a800000000000000a300000000000000a300000000",
            INIT_66 => X"000000c700000000000000d600000000000000dc00000000000000df00000000",
            INIT_67 => X"000000980000000000000090000000000000009000000000000000a300000000",
            INIT_68 => X"0000009b00000000000000a000000000000000a200000000000000a900000000",
            INIT_69 => X"000000a40000000000000083000000000000008800000000000000a300000000",
            INIT_6A => X"0000008500000000000000840000000000000088000000000000009200000000",
            INIT_6B => X"000000920000000000000087000000000000009e000000000000009f00000000",
            INIT_6C => X"0000009e000000000000009000000000000000a200000000000000a700000000",
            INIT_6D => X"000000cb00000000000000b00000000000000098000000000000009800000000",
            INIT_6E => X"000000da00000000000000dd00000000000000d800000000000000d700000000",
            INIT_6F => X"000000b600000000000000a2000000000000009f00000000000000c500000000",
            INIT_70 => X"0000009d00000000000000a200000000000000a400000000000000ae00000000",
            INIT_71 => X"000000b2000000000000006d000000000000007800000000000000a800000000",
            INIT_72 => X"000000a300000000000000a100000000000000a700000000000000a600000000",
            INIT_73 => X"00000078000000000000008400000000000000ab00000000000000b600000000",
            INIT_74 => X"00000095000000000000008c00000000000000a300000000000000a900000000",
            INIT_75 => X"000000cc00000000000000aa00000000000000a400000000000000a600000000",
            INIT_76 => X"000000e400000000000000da00000000000000d500000000000000d300000000",
            INIT_77 => X"000000c700000000000000bb00000000000000b000000000000000d600000000",
            INIT_78 => X"0000009f00000000000000a100000000000000a000000000000000af00000000",
            INIT_79 => X"000000b70000000000000068000000000000008400000000000000aa00000000",
            INIT_7A => X"000000b000000000000000b800000000000000b600000000000000bc00000000",
            INIT_7B => X"0000008d00000000000000a300000000000000a800000000000000a200000000",
            INIT_7C => X"00000085000000000000009200000000000000a5000000000000009100000000",
            INIT_7D => X"000000a9000000000000009600000000000000a500000000000000af00000000",
            INIT_7E => X"000000dd00000000000000d900000000000000d400000000000000ca00000000",
            INIT_7F => X"000000c700000000000000c700000000000000ba00000000000000c400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "sampleifmap_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000940000000000000092000000000000009f00000000000000b300000000",
            INIT_01 => X"000000a8000000000000006d000000000000009700000000000000a100000000",
            INIT_02 => X"000000ae00000000000000a400000000000000b500000000000000c700000000",
            INIT_03 => X"000000a600000000000000aa000000000000009c00000000000000a500000000",
            INIT_04 => X"00000077000000000000009f0000000000000088000000000000006900000000",
            INIT_05 => X"00000050000000000000007e000000000000009e000000000000008f00000000",
            INIT_06 => X"000000cd00000000000000d100000000000000b7000000000000007600000000",
            INIT_07 => X"000000c500000000000000c900000000000000b700000000000000af00000000",
            INIT_08 => X"00000083000000000000008500000000000000a400000000000000b500000000",
            INIT_09 => X"0000009f000000000000009700000000000000a5000000000000009500000000",
            INIT_0A => X"000000cd00000000000000c400000000000000c700000000000000c200000000",
            INIT_0B => X"000000a200000000000000ac00000000000000a800000000000000b900000000",
            INIT_0C => X"00000077000000000000009b0000000000000069000000000000006800000000",
            INIT_0D => X"0000005c000000000000008800000000000000ad000000000000008600000000",
            INIT_0E => X"0000009e0000000000000098000000000000006f000000000000004b00000000",
            INIT_0F => X"000000c800000000000000cb00000000000000b0000000000000009800000000",
            INIT_10 => X"00000085000000000000008e00000000000000ac00000000000000b700000000",
            INIT_11 => X"000000aa00000000000000b100000000000000b0000000000000009f00000000",
            INIT_12 => X"000000d900000000000000cf00000000000000c500000000000000b100000000",
            INIT_13 => X"000000aa00000000000000bb00000000000000c600000000000000d900000000",
            INIT_14 => X"0000007e0000000000000085000000000000005a000000000000008300000000",
            INIT_15 => X"0000007e000000000000008200000000000000a2000000000000008b00000000",
            INIT_16 => X"0000008400000000000000760000000000000060000000000000006f00000000",
            INIT_17 => X"000000c700000000000000b80000000000000092000000000000007c00000000",
            INIT_18 => X"0000009500000000000000a100000000000000b000000000000000b900000000",
            INIT_19 => X"000000bc00000000000000b600000000000000b700000000000000af00000000",
            INIT_1A => X"000000c200000000000000b900000000000000aa00000000000000aa00000000",
            INIT_1B => X"000000af00000000000000ca00000000000000d000000000000000c900000000",
            INIT_1C => X"000000910000000000000071000000000000007b00000000000000a400000000",
            INIT_1D => X"0000007b0000000000000071000000000000008c000000000000009d00000000",
            INIT_1E => X"0000008e00000000000000860000000000000070000000000000007700000000",
            INIT_1F => X"000000a600000000000000840000000000000079000000000000007f00000000",
            INIT_20 => X"0000009b00000000000000ad00000000000000b700000000000000bd00000000",
            INIT_21 => X"000000b200000000000000b100000000000000ba00000000000000ab00000000",
            INIT_22 => X"000000b100000000000000b200000000000000ac00000000000000b400000000",
            INIT_23 => X"000000bd00000000000000c300000000000000bc00000000000000a400000000",
            INIT_24 => X"0000009d000000000000008800000000000000b600000000000000c900000000",
            INIT_25 => X"0000007c000000000000006a0000000000000078000000000000009300000000",
            INIT_26 => X"0000008a0000000000000094000000000000008a000000000000008000000000",
            INIT_27 => X"00000082000000000000007a0000000000000077000000000000007800000000",
            INIT_28 => X"000000a100000000000000b700000000000000bc00000000000000bd00000000",
            INIT_29 => X"000000b000000000000000bb00000000000000b7000000000000009e00000000",
            INIT_2A => X"000000a400000000000000c000000000000000bf00000000000000b800000000",
            INIT_2B => X"000000b100000000000000ad00000000000000a6000000000000008b00000000",
            INIT_2C => X"0000009600000000000000a200000000000000bc00000000000000c000000000",
            INIT_2D => X"000000850000000000000079000000000000006b000000000000007600000000",
            INIT_2E => X"0000007d000000000000008d0000000000000096000000000000008e00000000",
            INIT_2F => X"0000006c000000000000007d000000000000007c000000000000007500000000",
            INIT_30 => X"000000a600000000000000bb00000000000000ba00000000000000ba00000000",
            INIT_31 => X"000000c500000000000000c700000000000000b4000000000000009400000000",
            INIT_32 => X"000000a800000000000000c000000000000000c300000000000000c100000000",
            INIT_33 => X"000000aa00000000000000a9000000000000009f000000000000009100000000",
            INIT_34 => X"0000008600000000000000a300000000000000ac00000000000000af00000000",
            INIT_35 => X"0000008b0000000000000086000000000000006c000000000000005d00000000",
            INIT_36 => X"0000007c000000000000008e0000000000000097000000000000008d00000000",
            INIT_37 => X"0000005b00000000000000650000000000000072000000000000007c00000000",
            INIT_38 => X"000000ac00000000000000b700000000000000b500000000000000ba00000000",
            INIT_39 => X"000000cf00000000000000c900000000000000b0000000000000008f00000000",
            INIT_3A => X"000000af00000000000000bd00000000000000cb00000000000000ce00000000",
            INIT_3B => X"000000ac00000000000000ae00000000000000ab00000000000000a500000000",
            INIT_3C => X"00000075000000000000009e00000000000000ab00000000000000b200000000",
            INIT_3D => X"00000088000000000000008a0000000000000078000000000000006100000000",
            INIT_3E => X"00000084000000000000009200000000000000a1000000000000008a00000000",
            INIT_3F => X"000000680000000000000064000000000000006d000000000000008200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000a900000000000000af00000000000000b200000000000000b800000000",
            INIT_41 => X"000000ca00000000000000c600000000000000aa000000000000009200000000",
            INIT_42 => X"0000008800000000000000ab00000000000000c500000000000000c800000000",
            INIT_43 => X"000000aa00000000000000ab00000000000000b400000000000000a100000000",
            INIT_44 => X"00000073000000000000009000000000000000a800000000000000ad00000000",
            INIT_45 => X"0000007e0000000000000086000000000000007c000000000000006c00000000",
            INIT_46 => X"0000008700000000000000910000000000000099000000000000008200000000",
            INIT_47 => X"0000006f00000000000000740000000000000075000000000000007700000000",
            INIT_48 => X"0000009d00000000000000a800000000000000b000000000000000b800000000",
            INIT_49 => X"000000c800000000000000c000000000000000a2000000000000009300000000",
            INIT_4A => X"00000052000000000000008100000000000000b900000000000000bf00000000",
            INIT_4B => X"0000009f00000000000000a600000000000000b3000000000000008d00000000",
            INIT_4C => X"0000007400000000000000840000000000000096000000000000009f00000000",
            INIT_4D => X"0000007a000000000000007f000000000000007a000000000000006900000000",
            INIT_4E => X"0000007a00000000000000800000000000000084000000000000007f00000000",
            INIT_4F => X"00000062000000000000006b0000000000000077000000000000007700000000",
            INIT_50 => X"0000009400000000000000a300000000000000ac00000000000000b800000000",
            INIT_51 => X"000000ca00000000000000ba0000000000000092000000000000008600000000",
            INIT_52 => X"00000058000000000000008200000000000000b200000000000000c000000000",
            INIT_53 => X"00000090000000000000009800000000000000ac000000000000008c00000000",
            INIT_54 => X"00000069000000000000007a0000000000000084000000000000009100000000",
            INIT_55 => X"0000007000000000000000790000000000000077000000000000006400000000",
            INIT_56 => X"0000006c00000000000000640000000000000071000000000000007a00000000",
            INIT_57 => X"000000720000000000000075000000000000007a000000000000007c00000000",
            INIT_58 => X"0000008e000000000000009e00000000000000a900000000000000b700000000",
            INIT_59 => X"000000cc00000000000000b20000000000000084000000000000007e00000000",
            INIT_5A => X"00000090000000000000009d00000000000000af00000000000000c300000000",
            INIT_5B => X"000000830000000000000087000000000000009800000000000000a400000000",
            INIT_5C => X"00000054000000000000006f0000000000000074000000000000007c00000000",
            INIT_5D => X"0000006d00000000000000710000000000000073000000000000006100000000",
            INIT_5E => X"00000064000000000000005f0000000000000066000000000000007200000000",
            INIT_5F => X"0000007b00000000000000820000000000000082000000000000007400000000",
            INIT_60 => X"0000008e000000000000009900000000000000a100000000000000b100000000",
            INIT_61 => X"000000cc00000000000000b2000000000000007a000000000000007700000000",
            INIT_62 => X"000000a800000000000000aa00000000000000b400000000000000c500000000",
            INIT_63 => X"0000007b000000000000007a0000000000000087000000000000009d00000000",
            INIT_64 => X"0000004b000000000000005e000000000000006d000000000000007700000000",
            INIT_65 => X"000000710000000000000070000000000000006f000000000000006800000000",
            INIT_66 => X"00000066000000000000005c0000000000000064000000000000007000000000",
            INIT_67 => X"00000073000000000000007e0000000000000082000000000000007700000000",
            INIT_68 => X"00000091000000000000008d000000000000009000000000000000a300000000",
            INIT_69 => X"000000c800000000000000a9000000000000006b000000000000007400000000",
            INIT_6A => X"000000a300000000000000ac00000000000000b700000000000000c200000000",
            INIT_6B => X"0000007900000000000000730000000000000081000000000000009600000000",
            INIT_6C => X"00000051000000000000004e0000000000000064000000000000007000000000",
            INIT_6D => X"00000072000000000000006a0000000000000065000000000000006800000000",
            INIT_6E => X"0000007000000000000000630000000000000063000000000000007200000000",
            INIT_6F => X"0000006e00000000000000740000000000000075000000000000007600000000",
            INIT_70 => X"0000008f0000000000000083000000000000007e000000000000008e00000000",
            INIT_71 => X"000000c00000000000000091000000000000005f000000000000007c00000000",
            INIT_72 => X"000000a800000000000000b200000000000000b700000000000000be00000000",
            INIT_73 => X"00000065000000000000005c0000000000000062000000000000008200000000",
            INIT_74 => X"0000005f000000000000004b000000000000005c000000000000006800000000",
            INIT_75 => X"00000074000000000000006a0000000000000061000000000000006300000000",
            INIT_76 => X"0000006e0000000000000071000000000000006c000000000000006d00000000",
            INIT_77 => X"000000770000000000000074000000000000006c000000000000006700000000",
            INIT_78 => X"0000007800000000000000700000000000000068000000000000007b00000000",
            INIT_79 => X"000000ae00000000000000760000000000000057000000000000007400000000",
            INIT_7A => X"0000008d00000000000000a400000000000000ae00000000000000b500000000",
            INIT_7B => X"0000004600000000000000390000000000000045000000000000006300000000",
            INIT_7C => X"0000006000000000000000580000000000000051000000000000005700000000",
            INIT_7D => X"00000070000000000000006b000000000000005e000000000000005d00000000",
            INIT_7E => X"0000005d0000000000000061000000000000006c000000000000006b00000000",
            INIT_7F => X"00000076000000000000007b0000000000000076000000000000006500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "sampleifmap_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000c700000000000000cd00000000000000d200000000000000d900000000",
            INIT_01 => X"000000bd00000000000000cf00000000000000d600000000000000da00000000",
            INIT_02 => X"000000a900000000000000a600000000000000ae00000000000000bb00000000",
            INIT_03 => X"0000008f000000000000008c000000000000009a000000000000009600000000",
            INIT_04 => X"000000df00000000000000db00000000000000bf00000000000000a700000000",
            INIT_05 => X"000000e100000000000000e200000000000000d700000000000000db00000000",
            INIT_06 => X"000000bb00000000000000af00000000000000be00000000000000db00000000",
            INIT_07 => X"000000a200000000000000a100000000000000aa00000000000000c800000000",
            INIT_08 => X"000000d700000000000000dc00000000000000dd00000000000000de00000000",
            INIT_09 => X"000000b300000000000000d300000000000000e100000000000000d800000000",
            INIT_0A => X"000000bc00000000000000be00000000000000c000000000000000b400000000",
            INIT_0B => X"000000db00000000000000d100000000000000ce00000000000000c700000000",
            INIT_0C => X"000000ec00000000000000ec00000000000000eb00000000000000e500000000",
            INIT_0D => X"000000e500000000000000e100000000000000e200000000000000e900000000",
            INIT_0E => X"000000cd00000000000000d000000000000000d400000000000000e700000000",
            INIT_0F => X"000000c800000000000000ba00000000000000b700000000000000d800000000",
            INIT_10 => X"000000e800000000000000e700000000000000e900000000000000ea00000000",
            INIT_11 => X"000000ad00000000000000d900000000000000ef00000000000000e900000000",
            INIT_12 => X"000000b700000000000000ad00000000000000b400000000000000a400000000",
            INIT_13 => X"000000e000000000000000d400000000000000bc00000000000000be00000000",
            INIT_14 => X"000000e100000000000000e300000000000000eb00000000000000da00000000",
            INIT_15 => X"000000e100000000000000d600000000000000df00000000000000e500000000",
            INIT_16 => X"000000d800000000000000e600000000000000e800000000000000ea00000000",
            INIT_17 => X"000000d300000000000000d000000000000000ca00000000000000d100000000",
            INIT_18 => X"000000f200000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009e00000000000000e400000000000000f300000000000000f400000000",
            INIT_1A => X"0000009f0000000000000083000000000000009d000000000000009200000000",
            INIT_1B => X"0000009f00000000000000a20000000000000088000000000000009100000000",
            INIT_1C => X"000000d300000000000000c300000000000000cb00000000000000a900000000",
            INIT_1D => X"000000e200000000000000d000000000000000cb00000000000000d100000000",
            INIT_1E => X"000000d500000000000000e400000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e000000000000000db00000000000000c700000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000007500000000000000cf00000000000000f100000000000000f500000000",
            INIT_22 => X"0000006b0000000000000059000000000000006c000000000000006300000000",
            INIT_23 => X"0000005c0000000000000064000000000000005b000000000000006400000000",
            INIT_24 => X"00000095000000000000007c000000000000007c000000000000006600000000",
            INIT_25 => X"000000e900000000000000ca00000000000000b900000000000000b600000000",
            INIT_26 => X"000000cd00000000000000e300000000000000e200000000000000e100000000",
            INIT_27 => X"000000de00000000000000e200000000000000d500000000000000c200000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007e00000000000000d800000000000000ed00000000000000f500000000",
            INIT_2A => X"00000066000000000000005b000000000000005a000000000000004800000000",
            INIT_2B => X"00000063000000000000006b0000000000000067000000000000006500000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005900000000",
            INIT_2D => X"000000eb00000000000000d800000000000000be000000000000007e00000000",
            INIT_2E => X"000000c400000000000000d800000000000000df00000000000000e700000000",
            INIT_2F => X"000000ec00000000000000d900000000000000bd00000000000000ae00000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009e00000000000000d900000000000000db00000000000000f100000000",
            INIT_32 => X"0000009700000000000000840000000000000072000000000000005000000000",
            INIT_33 => X"0000008a000000000000008f0000000000000084000000000000008c00000000",
            INIT_34 => X"000000780000000000000072000000000000007a000000000000008200000000",
            INIT_35 => X"000000e900000000000000dd000000000000009b000000000000006e00000000",
            INIT_36 => X"000000c000000000000000c600000000000000e000000000000000eb00000000",
            INIT_37 => X"000000eb00000000000000cc00000000000000ab00000000000000a700000000",
            INIT_38 => X"000000f600000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009900000000000000d700000000000000c700000000000000e300000000",
            INIT_3A => X"000000ca00000000000000bb0000000000000092000000000000005100000000",
            INIT_3B => X"000000830000000000000083000000000000009e00000000000000cf00000000",
            INIT_3C => X"000000840000000000000083000000000000008d000000000000008100000000",
            INIT_3D => X"000000d7000000000000009f0000000000000084000000000000009f00000000",
            INIT_3E => X"000000d100000000000000d400000000000000d700000000000000e500000000",
            INIT_3F => X"000000dd00000000000000b200000000000000ab00000000000000c500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000008200000000000000da00000000000000ce00000000000000e300000000",
            INIT_42 => X"0000008100000000000000800000000000000082000000000000005100000000",
            INIT_43 => X"0000007d0000000000000074000000000000009100000000000000b800000000",
            INIT_44 => X"0000007d000000000000008e0000000000000089000000000000007c00000000",
            INIT_45 => X"000000c600000000000000900000000000000093000000000000009900000000",
            INIT_46 => X"000000dc00000000000000e900000000000000db00000000000000d600000000",
            INIT_47 => X"000000c900000000000000a900000000000000a400000000000000b800000000",
            INIT_48 => X"000000f200000000000000f400000000000000f300000000000000f300000000",
            INIT_49 => X"0000006e00000000000000a800000000000000be00000000000000e400000000",
            INIT_4A => X"0000006e00000000000000770000000000000086000000000000005300000000",
            INIT_4B => X"0000007800000000000000730000000000000080000000000000008f00000000",
            INIT_4C => X"0000007d00000000000000920000000000000083000000000000007d00000000",
            INIT_4D => X"000000c4000000000000008c000000000000009b000000000000009500000000",
            INIT_4E => X"000000e900000000000000f000000000000000f000000000000000e900000000",
            INIT_4F => X"000000dc00000000000000d700000000000000c800000000000000c800000000",
            INIT_50 => X"000000f500000000000000f400000000000000f100000000000000ef00000000",
            INIT_51 => X"0000005f0000000000000082000000000000008500000000000000dc00000000",
            INIT_52 => X"0000006c00000000000000740000000000000074000000000000004e00000000",
            INIT_53 => X"0000006c000000000000006d000000000000006b000000000000006d00000000",
            INIT_54 => X"0000007300000000000000780000000000000078000000000000007300000000",
            INIT_55 => X"000000a7000000000000008f0000000000000096000000000000008800000000",
            INIT_56 => X"000000f300000000000000f500000000000000e400000000000000d000000000",
            INIT_57 => X"000000f400000000000000f500000000000000f500000000000000f400000000",
            INIT_58 => X"000000f400000000000000f200000000000000e900000000000000de00000000",
            INIT_59 => X"0000005900000000000000a500000000000000a900000000000000d800000000",
            INIT_5A => X"00000064000000000000005b0000000000000043000000000000003d00000000",
            INIT_5B => X"000000600000000000000062000000000000005f000000000000005f00000000",
            INIT_5C => X"00000061000000000000005a000000000000005f000000000000006000000000",
            INIT_5D => X"0000007e00000000000000810000000000000079000000000000006900000000",
            INIT_5E => X"000000f300000000000000f800000000000000d8000000000000009b00000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e300000000000000ec00000000000000df00000000000000d000000000",
            INIT_61 => X"0000006400000000000000b500000000000000b700000000000000bf00000000",
            INIT_62 => X"0000006500000000000000580000000000000038000000000000003700000000",
            INIT_63 => X"0000005400000000000000560000000000000063000000000000006f00000000",
            INIT_64 => X"00000071000000000000005d0000000000000054000000000000005200000000",
            INIT_65 => X"0000008100000000000000700000000000000062000000000000006d00000000",
            INIT_66 => X"000000f400000000000000f500000000000000e200000000000000ae00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c300000000000000db00000000000000cc00000000000000c800000000",
            INIT_69 => X"00000066000000000000009c000000000000009a00000000000000aa00000000",
            INIT_6A => X"00000066000000000000006c0000000000000063000000000000006800000000",
            INIT_6B => X"00000055000000000000005e0000000000000075000000000000007300000000",
            INIT_6C => X"0000008c000000000000007a000000000000006a000000000000005a00000000",
            INIT_6D => X"0000007c000000000000006c0000000000000068000000000000008000000000",
            INIT_6E => X"000000d400000000000000c300000000000000b3000000000000009600000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a900000000000000cf00000000000000d200000000000000c800000000",
            INIT_71 => X"0000008a0000000000000093000000000000009400000000000000a400000000",
            INIT_72 => X"0000005d000000000000006a000000000000005c000000000000008100000000",
            INIT_73 => X"0000004d0000000000000054000000000000005d000000000000005900000000",
            INIT_74 => X"0000005100000000000000510000000000000051000000000000004c00000000",
            INIT_75 => X"00000052000000000000004b000000000000004a000000000000004f00000000",
            INIT_76 => X"0000008f000000000000008c000000000000007b000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bf00000000",
            INIT_78 => X"0000007700000000000000c400000000000000e200000000000000d200000000",
            INIT_79 => X"000000c000000000000000ba0000000000000096000000000000007000000000",
            INIT_7A => X"00000037000000000000004d000000000000004d000000000000006c00000000",
            INIT_7B => X"0000003f000000000000003c000000000000002f000000000000002d00000000",
            INIT_7C => X"00000036000000000000003b000000000000003f000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000032000000000000003100000000",
            INIT_7E => X"00000067000000000000005b000000000000004b000000000000004700000000",
            INIT_7F => X"000000f400000000000000f600000000000000e1000000000000008700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "sampleifmap_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006000000000000000b400000000000000c100000000000000c700000000",
            INIT_01 => X"000000a100000000000000c00000000000000091000000000000005d00000000",
            INIT_02 => X"00000062000000000000005c0000000000000049000000000000005600000000",
            INIT_03 => X"00000047000000000000004f000000000000004f000000000000006800000000",
            INIT_04 => X"0000001b000000000000001e000000000000001c000000000000002500000000",
            INIT_05 => X"0000001c00000000000000160000000000000032000000000000003400000000",
            INIT_06 => X"00000068000000000000005b0000000000000035000000000000001800000000",
            INIT_07 => X"000000f300000000000000f700000000000000ce000000000000008000000000",
            INIT_08 => X"0000007100000000000000c200000000000000c700000000000000d300000000",
            INIT_09 => X"00000047000000000000009f000000000000009d000000000000007800000000",
            INIT_0A => X"0000007c0000000000000074000000000000005a000000000000004400000000",
            INIT_0B => X"0000006600000000000000800000000000000079000000000000009500000000",
            INIT_0C => X"0000006400000000000000700000000000000062000000000000004e00000000",
            INIT_0D => X"00000063000000000000005c0000000000000093000000000000009400000000",
            INIT_0E => X"0000008e0000000000000087000000000000006c000000000000005e00000000",
            INIT_0F => X"000000f500000000000000f200000000000000b7000000000000009c00000000",
            INIT_10 => X"0000006600000000000000b700000000000000ca00000000000000dc00000000",
            INIT_11 => X"0000001e000000000000008400000000000000a5000000000000006e00000000",
            INIT_12 => X"00000053000000000000006b0000000000000062000000000000003900000000",
            INIT_13 => X"0000006400000000000000810000000000000065000000000000005200000000",
            INIT_14 => X"0000009f000000000000009e00000000000000ae000000000000009900000000",
            INIT_15 => X"000000a300000000000000a200000000000000a800000000000000ac00000000",
            INIT_16 => X"00000077000000000000009c00000000000000af00000000000000a000000000",
            INIT_17 => X"000000f700000000000000e40000000000000087000000000000007200000000",
            INIT_18 => X"0000006200000000000000bc00000000000000cf00000000000000db00000000",
            INIT_19 => X"0000002a000000000000006f000000000000008d000000000000005300000000",
            INIT_1A => X"0000003e000000000000004c0000000000000048000000000000003a00000000",
            INIT_1B => X"0000005d00000000000000400000000000000038000000000000003500000000",
            INIT_1C => X"00000065000000000000005b000000000000007c00000000000000a000000000",
            INIT_1D => X"000000670000000000000067000000000000006b000000000000007400000000",
            INIT_1E => X"00000043000000000000007e000000000000009b000000000000006300000000",
            INIT_1F => X"000000f800000000000000d90000000000000076000000000000005100000000",
            INIT_20 => X"0000006500000000000000c700000000000000d200000000000000d900000000",
            INIT_21 => X"0000003c000000000000005d0000000000000058000000000000003800000000",
            INIT_22 => X"00000046000000000000003f000000000000002e000000000000003800000000",
            INIT_23 => X"0000004100000000000000400000000000000036000000000000003c00000000",
            INIT_24 => X"0000006700000000000000690000000000000072000000000000006300000000",
            INIT_25 => X"00000061000000000000005d0000000000000060000000000000006400000000",
            INIT_26 => X"000000490000000000000064000000000000006f000000000000006600000000",
            INIT_27 => X"000000f900000000000000d40000000000000072000000000000005200000000",
            INIT_28 => X"0000007500000000000000ca00000000000000cd00000000000000d100000000",
            INIT_29 => X"0000004400000000000000510000000000000046000000000000005300000000",
            INIT_2A => X"00000033000000000000002b0000000000000023000000000000003200000000",
            INIT_2B => X"0000003f0000000000000057000000000000004d000000000000004400000000",
            INIT_2C => X"0000004800000000000000520000000000000047000000000000003400000000",
            INIT_2D => X"0000005d000000000000003e0000000000000043000000000000004000000000",
            INIT_2E => X"0000006c0000000000000053000000000000003c000000000000005800000000",
            INIT_2F => X"000000fa00000000000000cc000000000000006c000000000000007000000000",
            INIT_30 => X"0000006800000000000000c500000000000000ca00000000000000cd00000000",
            INIT_31 => X"000000490000000000000047000000000000006f000000000000005d00000000",
            INIT_32 => X"0000002200000000000000260000000000000029000000000000003f00000000",
            INIT_33 => X"0000004f000000000000008e0000000000000063000000000000004b00000000",
            INIT_34 => X"0000007600000000000000930000000000000056000000000000001e00000000",
            INIT_35 => X"0000009900000000000000660000000000000072000000000000006300000000",
            INIT_36 => X"0000008d000000000000004a000000000000003f00000000000000b200000000",
            INIT_37 => X"000000f600000000000000c3000000000000005a000000000000007700000000",
            INIT_38 => X"0000005700000000000000b900000000000000c200000000000000c600000000",
            INIT_39 => X"000000630000000000000061000000000000006c000000000000003100000000",
            INIT_3A => X"0000002400000000000000270000000000000033000000000000005f00000000",
            INIT_3B => X"0000003700000000000000570000000000000032000000000000002800000000",
            INIT_3C => X"0000007f0000000000000097000000000000004f000000000000002000000000",
            INIT_3D => X"0000009c00000000000000740000000000000088000000000000007a00000000",
            INIT_3E => X"0000004a00000000000000350000000000000037000000000000009f00000000",
            INIT_3F => X"000000f000000000000000c2000000000000004e000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004d00000000000000a900000000000000b400000000000000b600000000",
            INIT_41 => X"00000090000000000000006c000000000000003b000000000000002500000000",
            INIT_42 => X"00000020000000000000002b000000000000003c000000000000006a00000000",
            INIT_43 => X"00000021000000000000001e000000000000001c000000000000001d00000000",
            INIT_44 => X"00000058000000000000003a000000000000002a000000000000002700000000",
            INIT_45 => X"00000075000000000000007a0000000000000079000000000000006a00000000",
            INIT_46 => X"000000320000000000000033000000000000002f000000000000004300000000",
            INIT_47 => X"000000e100000000000000ba0000000000000050000000000000003300000000",
            INIT_48 => X"0000007d00000000000000a400000000000000a500000000000000a800000000",
            INIT_49 => X"0000008d000000000000006f0000000000000060000000000000005b00000000",
            INIT_4A => X"000000240000000000000037000000000000004a000000000000006000000000",
            INIT_4B => X"0000001f000000000000001d000000000000001e000000000000001e00000000",
            INIT_4C => X"000000ae00000000000000400000000000000018000000000000002300000000",
            INIT_4D => X"000000b500000000000000b300000000000000cb00000000000000cd00000000",
            INIT_4E => X"00000030000000000000002b0000000000000026000000000000005700000000",
            INIT_4F => X"000000d300000000000000ae000000000000005b000000000000004200000000",
            INIT_50 => X"000000b400000000000000af00000000000000a300000000000000a200000000",
            INIT_51 => X"0000008d000000000000006c0000000000000076000000000000009800000000",
            INIT_52 => X"00000030000000000000004e0000000000000053000000000000005b00000000",
            INIT_53 => X"0000001d00000000000000190000000000000018000000000000001900000000",
            INIT_54 => X"000000a400000000000000470000000000000026000000000000002700000000",
            INIT_55 => X"000000a600000000000000a900000000000000b100000000000000b800000000",
            INIT_56 => X"00000031000000000000001e000000000000001e000000000000005100000000",
            INIT_57 => X"000000ce00000000000000a9000000000000005f000000000000004e00000000",
            INIT_58 => X"000000a600000000000000b300000000000000ac000000000000009a00000000",
            INIT_59 => X"0000009200000000000000670000000000000075000000000000009200000000",
            INIT_5A => X"0000003600000000000000520000000000000055000000000000005700000000",
            INIT_5B => X"000000250000000000000021000000000000001e000000000000002000000000",
            INIT_5C => X"000000650000000000000056000000000000004d000000000000003600000000",
            INIT_5D => X"00000089000000000000008e0000000000000079000000000000006b00000000",
            INIT_5E => X"000000360000000000000021000000000000001e000000000000003c00000000",
            INIT_5F => X"000000c700000000000000a5000000000000005b000000000000004e00000000",
            INIT_60 => X"00000094000000000000009e00000000000000a900000000000000a600000000",
            INIT_61 => X"0000007100000000000000670000000000000085000000000000008f00000000",
            INIT_62 => X"0000003c000000000000004b0000000000000051000000000000004f00000000",
            INIT_63 => X"0000002c000000000000002a0000000000000027000000000000002a00000000",
            INIT_64 => X"0000004d00000000000000410000000000000036000000000000003000000000",
            INIT_65 => X"0000008b0000000000000083000000000000006e000000000000005a00000000",
            INIT_66 => X"000000360000000000000026000000000000001d000000000000003500000000",
            INIT_67 => X"000000c400000000000000a9000000000000005b000000000000004600000000",
            INIT_68 => X"0000008d0000000000000093000000000000009700000000000000a200000000",
            INIT_69 => X"0000004e000000000000006b0000000000000085000000000000008900000000",
            INIT_6A => X"0000003c0000000000000046000000000000004e000000000000004800000000",
            INIT_6B => X"00000030000000000000002e000000000000002a000000000000003200000000",
            INIT_6C => X"00000042000000000000003b0000000000000033000000000000003100000000",
            INIT_6D => X"0000007100000000000000650000000000000059000000000000004c00000000",
            INIT_6E => X"000000340000000000000023000000000000001d000000000000004500000000",
            INIT_6F => X"000000ba00000000000000ae0000000000000062000000000000003f00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009400000000",
            INIT_71 => X"0000003c000000000000006a000000000000008c000000000000008f00000000",
            INIT_72 => X"000000370000000000000042000000000000004a000000000000004200000000",
            INIT_73 => X"0000003a00000000000000360000000000000034000000000000003900000000",
            INIT_74 => X"000000460000000000000041000000000000003a000000000000003a00000000",
            INIT_75 => X"0000005d00000000000000570000000000000050000000000000004900000000",
            INIT_76 => X"0000003700000000000000260000000000000025000000000000004d00000000",
            INIT_77 => X"000000b400000000000000b30000000000000083000000000000004a00000000",
            INIT_78 => X"000000a200000000000000a00000000000000095000000000000009000000000",
            INIT_79 => X"0000003d000000000000007e0000000000000092000000000000009e00000000",
            INIT_7A => X"00000043000000000000003a0000000000000039000000000000003900000000",
            INIT_7B => X"0000004800000000000000490000000000000045000000000000004600000000",
            INIT_7C => X"0000006200000000000000590000000000000049000000000000004400000000",
            INIT_7D => X"0000006100000000000000630000000000000061000000000000005e00000000",
            INIT_7E => X"0000004700000000000000400000000000000045000000000000005200000000",
            INIT_7F => X"000000ba00000000000000b600000000000000a4000000000000007700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "sampleifmap_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000ca00000000000000d000000000000000d000000000000000d700000000",
            INIT_01 => X"000000b900000000000000ca00000000000000d100000000000000d700000000",
            INIT_02 => X"000000a0000000000000009800000000000000a800000000000000b800000000",
            INIT_03 => X"0000009d000000000000009a00000000000000a7000000000000009d00000000",
            INIT_04 => X"000000e100000000000000e100000000000000cb00000000000000b500000000",
            INIT_05 => X"000000e400000000000000e500000000000000db00000000000000de00000000",
            INIT_06 => X"000000c400000000000000b800000000000000c500000000000000dd00000000",
            INIT_07 => X"000000a500000000000000b000000000000000b800000000000000d000000000",
            INIT_08 => X"000000d900000000000000e100000000000000e000000000000000e200000000",
            INIT_09 => X"000000ab00000000000000cc00000000000000dd00000000000000d500000000",
            INIT_0A => X"000000b100000000000000b200000000000000bd00000000000000b400000000",
            INIT_0B => X"000000e000000000000000d000000000000000cd00000000000000c400000000",
            INIT_0C => X"000000f300000000000000f200000000000000f000000000000000ec00000000",
            INIT_0D => X"000000e700000000000000e400000000000000e500000000000000ee00000000",
            INIT_0E => X"000000d200000000000000d400000000000000d600000000000000e700000000",
            INIT_0F => X"000000c500000000000000bf00000000000000be00000000000000de00000000",
            INIT_10 => X"000000eb00000000000000ea00000000000000ea00000000000000eb00000000",
            INIT_11 => X"000000a600000000000000d600000000000000ef00000000000000ea00000000",
            INIT_12 => X"000000b100000000000000a800000000000000b100000000000000a600000000",
            INIT_13 => X"000000df00000000000000ce00000000000000b700000000000000b800000000",
            INIT_14 => X"000000e800000000000000e300000000000000ec00000000000000dc00000000",
            INIT_15 => X"000000e000000000000000d900000000000000e400000000000000eb00000000",
            INIT_16 => X"000000dd00000000000000e600000000000000e900000000000000e900000000",
            INIT_17 => X"000000d200000000000000d100000000000000ce00000000000000d900000000",
            INIT_18 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"0000009900000000000000e300000000000000f400000000000000f400000000",
            INIT_1A => X"0000009f0000000000000082000000000000009b000000000000009200000000",
            INIT_1B => X"000000a000000000000000a2000000000000008a000000000000009000000000",
            INIT_1C => X"000000dc00000000000000c200000000000000cd00000000000000ac00000000",
            INIT_1D => X"000000e000000000000000d300000000000000d300000000000000de00000000",
            INIT_1E => X"000000db00000000000000e500000000000000e900000000000000e600000000",
            INIT_1F => X"000000d400000000000000e200000000000000df00000000000000cf00000000",
            INIT_20 => X"000000f400000000000000f400000000000000f400000000000000f500000000",
            INIT_21 => X"0000007000000000000000cd00000000000000f000000000000000f500000000",
            INIT_22 => X"0000006d000000000000005b000000000000006d000000000000006200000000",
            INIT_23 => X"0000005c0000000000000064000000000000005c000000000000006500000000",
            INIT_24 => X"0000009a000000000000007c000000000000007d000000000000006800000000",
            INIT_25 => X"000000e300000000000000c900000000000000c200000000000000c200000000",
            INIT_26 => X"000000d300000000000000e300000000000000de00000000000000dc00000000",
            INIT_27 => X"000000e100000000000000e800000000000000dc00000000000000cb00000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000007b00000000000000d400000000000000eb00000000000000f600000000",
            INIT_2A => X"00000069000000000000005f000000000000005d000000000000004700000000",
            INIT_2B => X"00000066000000000000006e000000000000006a000000000000006700000000",
            INIT_2C => X"0000005d000000000000005b0000000000000059000000000000005b00000000",
            INIT_2D => X"000000e600000000000000d900000000000000c5000000000000008100000000",
            INIT_2E => X"000000c600000000000000d600000000000000da00000000000000dd00000000",
            INIT_2F => X"000000ed00000000000000e200000000000000c500000000000000b400000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"0000009c00000000000000d500000000000000d600000000000000f000000000",
            INIT_32 => X"0000009a00000000000000890000000000000077000000000000004f00000000",
            INIT_33 => X"00000096000000000000009b000000000000008b000000000000009000000000",
            INIT_34 => X"0000007e00000000000000790000000000000080000000000000008e00000000",
            INIT_35 => X"000000e900000000000000e100000000000000a0000000000000007200000000",
            INIT_36 => X"000000ba00000000000000c000000000000000da00000000000000e900000000",
            INIT_37 => X"000000ec00000000000000d400000000000000b000000000000000a500000000",
            INIT_38 => X"000000f700000000000000f300000000000000f300000000000000f400000000",
            INIT_39 => X"0000009600000000000000d300000000000000c100000000000000e200000000",
            INIT_3A => X"000000c800000000000000bc0000000000000098000000000000005100000000",
            INIT_3B => X"00000090000000000000008d00000000000000a500000000000000cd00000000",
            INIT_3C => X"0000008f000000000000008d0000000000000096000000000000008e00000000",
            INIT_3D => X"000000d600000000000000a3000000000000008c00000000000000a700000000",
            INIT_3E => X"000000d200000000000000d300000000000000d100000000000000e000000000",
            INIT_3F => X"000000dc00000000000000af00000000000000ae00000000000000c700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f400000000000000f300000000000000f400000000",
            INIT_41 => X"0000007f00000000000000d800000000000000ca00000000000000e100000000",
            INIT_42 => X"0000008700000000000000840000000000000086000000000000005100000000",
            INIT_43 => X"00000087000000000000007c000000000000009700000000000000b900000000",
            INIT_44 => X"0000008800000000000000960000000000000091000000000000008600000000",
            INIT_45 => X"000000c0000000000000008e000000000000009e00000000000000a400000000",
            INIT_46 => X"000000d700000000000000e700000000000000d800000000000000cf00000000",
            INIT_47 => X"000000c4000000000000009c000000000000009e00000000000000b100000000",
            INIT_48 => X"000000f200000000000000f400000000000000f200000000000000f200000000",
            INIT_49 => X"0000006e00000000000000a800000000000000bd00000000000000e300000000",
            INIT_4A => X"000000760000000000000080000000000000008c000000000000005300000000",
            INIT_4B => X"00000081000000000000007c0000000000000087000000000000009300000000",
            INIT_4C => X"000000860000000000000097000000000000008b000000000000008500000000",
            INIT_4D => X"000000c1000000000000009100000000000000a4000000000000009e00000000",
            INIT_4E => X"000000e600000000000000ef00000000000000ef00000000000000e500000000",
            INIT_4F => X"000000d700000000000000cc00000000000000be00000000000000c100000000",
            INIT_50 => X"000000f400000000000000f300000000000000ef00000000000000e800000000",
            INIT_51 => X"0000005e0000000000000080000000000000008100000000000000da00000000",
            INIT_52 => X"00000070000000000000007a000000000000007a000000000000004f00000000",
            INIT_53 => X"0000007300000000000000730000000000000070000000000000007100000000",
            INIT_54 => X"0000007e000000000000007f0000000000000080000000000000007c00000000",
            INIT_55 => X"000000aa0000000000000099000000000000009e000000000000009000000000",
            INIT_56 => X"000000f400000000000000f600000000000000e300000000000000ce00000000",
            INIT_57 => X"000000f400000000000000f500000000000000f300000000000000f300000000",
            INIT_58 => X"000000f200000000000000f200000000000000e300000000000000cd00000000",
            INIT_59 => X"00000058000000000000009f00000000000000a100000000000000d300000000",
            INIT_5A => X"00000066000000000000005e0000000000000045000000000000003c00000000",
            INIT_5B => X"0000006600000000000000670000000000000061000000000000006200000000",
            INIT_5C => X"00000067000000000000005f0000000000000064000000000000006800000000",
            INIT_5D => X"000000800000000000000089000000000000007f000000000000007100000000",
            INIT_5E => X"000000f300000000000000f800000000000000d7000000000000009900000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000dc00000000000000e400000000000000d500000000000000bc00000000",
            INIT_61 => X"0000006300000000000000ad00000000000000aa00000000000000b400000000",
            INIT_62 => X"00000066000000000000005a0000000000000039000000000000003700000000",
            INIT_63 => X"0000005500000000000000580000000000000067000000000000007200000000",
            INIT_64 => X"00000073000000000000005d0000000000000055000000000000005500000000",
            INIT_65 => X"0000008600000000000000760000000000000065000000000000007000000000",
            INIT_66 => X"000000f400000000000000f500000000000000e100000000000000b000000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000b500000000000000ca00000000000000bc00000000000000b800000000",
            INIT_69 => X"00000063000000000000008d0000000000000086000000000000009800000000",
            INIT_6A => X"00000067000000000000006f0000000000000066000000000000006700000000",
            INIT_6B => X"0000005600000000000000600000000000000078000000000000007600000000",
            INIT_6C => X"00000092000000000000007d000000000000006b000000000000005c00000000",
            INIT_6D => X"0000007f000000000000006e000000000000006a000000000000008400000000",
            INIT_6E => X"000000d200000000000000c300000000000000b3000000000000009800000000",
            INIT_6F => X"000000f400000000000000f400000000000000f500000000000000ee00000000",
            INIT_70 => X"0000009800000000000000bd00000000000000c200000000000000b600000000",
            INIT_71 => X"0000007e000000000000007f000000000000007b000000000000009200000000",
            INIT_72 => X"0000005e0000000000000069000000000000005d000000000000007c00000000",
            INIT_73 => X"0000004f0000000000000055000000000000005d000000000000005a00000000",
            INIT_74 => X"0000005500000000000000540000000000000053000000000000004e00000000",
            INIT_75 => X"00000053000000000000004c000000000000004b000000000000005100000000",
            INIT_76 => X"0000008a000000000000008a000000000000007a000000000000006500000000",
            INIT_77 => X"000000f400000000000000f400000000000000f400000000000000bc00000000",
            INIT_78 => X"0000006500000000000000a700000000000000cc00000000000000bd00000000",
            INIT_79 => X"000000ae00000000000000a9000000000000007d000000000000006500000000",
            INIT_7A => X"00000036000000000000004f000000000000004d000000000000006700000000",
            INIT_7B => X"0000003e000000000000003b000000000000002f000000000000002b00000000",
            INIT_7C => X"000000340000000000000039000000000000003e000000000000003b00000000",
            INIT_7D => X"00000040000000000000003d0000000000000030000000000000002f00000000",
            INIT_7E => X"00000061000000000000005a000000000000004a000000000000004600000000",
            INIT_7F => X"000000f400000000000000f600000000000000df000000000000008000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "sampleifmap_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000054000000000000009700000000000000a400000000000000ae00000000",
            INIT_01 => X"0000009200000000000000ac000000000000007c000000000000005200000000",
            INIT_02 => X"0000005a00000000000000570000000000000049000000000000005300000000",
            INIT_03 => X"00000044000000000000004c000000000000004b000000000000006400000000",
            INIT_04 => X"00000017000000000000001a0000000000000017000000000000002100000000",
            INIT_05 => X"000000190000000000000014000000000000002f000000000000003000000000",
            INIT_06 => X"0000006400000000000000560000000000000032000000000000001500000000",
            INIT_07 => X"000000f300000000000000f700000000000000ca000000000000007800000000",
            INIT_08 => X"0000006800000000000000b300000000000000b400000000000000c000000000",
            INIT_09 => X"00000040000000000000008e0000000000000087000000000000006800000000",
            INIT_0A => X"00000078000000000000006c0000000000000057000000000000004100000000",
            INIT_0B => X"00000062000000000000007d0000000000000076000000000000009500000000",
            INIT_0C => X"00000060000000000000006a0000000000000059000000000000004600000000",
            INIT_0D => X"0000006000000000000000590000000000000090000000000000009000000000",
            INIT_0E => X"0000008b00000000000000820000000000000067000000000000005a00000000",
            INIT_0F => X"000000f400000000000000f100000000000000b2000000000000009700000000",
            INIT_10 => X"0000005e00000000000000ab00000000000000bd00000000000000d100000000",
            INIT_11 => X"0000001c00000000000000760000000000000092000000000000006200000000",
            INIT_12 => X"0000004f0000000000000067000000000000005f000000000000003600000000",
            INIT_13 => X"0000005f00000000000000800000000000000064000000000000005300000000",
            INIT_14 => X"0000009e000000000000009b00000000000000aa000000000000009200000000",
            INIT_15 => X"000000a100000000000000a000000000000000a800000000000000ab00000000",
            INIT_16 => X"00000077000000000000009b00000000000000ac000000000000009e00000000",
            INIT_17 => X"000000f700000000000000e20000000000000080000000000000006f00000000",
            INIT_18 => X"0000005b00000000000000b000000000000000c100000000000000d000000000",
            INIT_19 => X"000000280000000000000064000000000000007f000000000000004c00000000",
            INIT_1A => X"0000003900000000000000490000000000000044000000000000003500000000",
            INIT_1B => X"00000059000000000000003d0000000000000035000000000000003200000000",
            INIT_1C => X"0000006200000000000000570000000000000077000000000000009c00000000",
            INIT_1D => X"0000006400000000000000630000000000000068000000000000007100000000",
            INIT_1E => X"0000003f000000000000007a0000000000000098000000000000006000000000",
            INIT_1F => X"000000f800000000000000d60000000000000070000000000000004d00000000",
            INIT_20 => X"0000005f00000000000000be00000000000000c300000000000000ca00000000",
            INIT_21 => X"000000380000000000000053000000000000004e000000000000003300000000",
            INIT_22 => X"00000044000000000000003c0000000000000027000000000000003300000000",
            INIT_23 => X"0000003d000000000000003b0000000000000033000000000000003900000000",
            INIT_24 => X"000000650000000000000066000000000000006e000000000000005f00000000",
            INIT_25 => X"00000060000000000000005c000000000000005f000000000000006300000000",
            INIT_26 => X"000000460000000000000060000000000000006c000000000000006400000000",
            INIT_27 => X"000000f900000000000000d0000000000000006c000000000000004f00000000",
            INIT_28 => X"0000006e00000000000000c000000000000000c000000000000000c200000000",
            INIT_29 => X"0000003f0000000000000049000000000000003e000000000000004c00000000",
            INIT_2A => X"000000300000000000000028000000000000001d000000000000002e00000000",
            INIT_2B => X"0000003b00000000000000530000000000000048000000000000004100000000",
            INIT_2C => X"00000043000000000000004d0000000000000043000000000000003000000000",
            INIT_2D => X"00000058000000000000003b0000000000000040000000000000003c00000000",
            INIT_2E => X"00000069000000000000004e0000000000000036000000000000005200000000",
            INIT_2F => X"000000f900000000000000c90000000000000065000000000000006b00000000",
            INIT_30 => X"0000006100000000000000bb00000000000000be00000000000000c300000000",
            INIT_31 => X"0000004300000000000000410000000000000063000000000000005500000000",
            INIT_32 => X"0000002000000000000000230000000000000026000000000000003a00000000",
            INIT_33 => X"0000004c000000000000008d0000000000000060000000000000004800000000",
            INIT_34 => X"00000071000000000000008c000000000000004f000000000000001900000000",
            INIT_35 => X"000000920000000000000061000000000000006d000000000000005e00000000",
            INIT_36 => X"0000008a0000000000000045000000000000003a00000000000000ab00000000",
            INIT_37 => X"000000f400000000000000c00000000000000053000000000000007400000000",
            INIT_38 => X"0000005200000000000000b000000000000000b700000000000000bd00000000",
            INIT_39 => X"0000005e00000000000000590000000000000063000000000000002c00000000",
            INIT_3A => X"0000002100000000000000240000000000000030000000000000005a00000000",
            INIT_3B => X"000000340000000000000055000000000000002f000000000000002600000000",
            INIT_3C => X"0000007b0000000000000091000000000000004a000000000000001c00000000",
            INIT_3D => X"0000009700000000000000710000000000000086000000000000007700000000",
            INIT_3E => X"0000004700000000000000320000000000000033000000000000009c00000000",
            INIT_3F => X"000000ee00000000000000c00000000000000047000000000000003b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004800000000000000a300000000000000ad00000000000000ae00000000",
            INIT_41 => X"0000008b00000000000000650000000000000036000000000000002200000000",
            INIT_42 => X"0000001e0000000000000028000000000000003a000000000000006600000000",
            INIT_43 => X"0000001e000000000000001a0000000000000019000000000000001a00000000",
            INIT_44 => X"0000005600000000000000350000000000000026000000000000002500000000",
            INIT_45 => X"0000007200000000000000760000000000000075000000000000006800000000",
            INIT_46 => X"0000002e0000000000000030000000000000002b000000000000003e00000000",
            INIT_47 => X"000000df00000000000000b8000000000000004b000000000000002f00000000",
            INIT_48 => X"00000078000000000000009e00000000000000a000000000000000a200000000",
            INIT_49 => X"0000008800000000000000670000000000000059000000000000005700000000",
            INIT_4A => X"0000002200000000000000340000000000000048000000000000005c00000000",
            INIT_4B => X"0000001d000000000000001b000000000000001b000000000000001c00000000",
            INIT_4C => X"000000af000000000000003d0000000000000015000000000000002000000000",
            INIT_4D => X"000000b400000000000000b100000000000000ca00000000000000cf00000000",
            INIT_4E => X"0000002c00000000000000280000000000000022000000000000005400000000",
            INIT_4F => X"000000d100000000000000ab0000000000000057000000000000003e00000000",
            INIT_50 => X"000000b000000000000000a8000000000000009c000000000000009c00000000",
            INIT_51 => X"0000008800000000000000660000000000000070000000000000009300000000",
            INIT_52 => X"0000002d000000000000004b0000000000000051000000000000005600000000",
            INIT_53 => X"0000001a00000000000000170000000000000016000000000000001600000000",
            INIT_54 => X"000000a400000000000000450000000000000022000000000000002300000000",
            INIT_55 => X"000000a500000000000000a900000000000000b100000000000000b900000000",
            INIT_56 => X"0000002d000000000000001a0000000000000019000000000000004e00000000",
            INIT_57 => X"000000cc00000000000000a7000000000000005c000000000000004b00000000",
            INIT_58 => X"000000a100000000000000ad00000000000000a7000000000000009500000000",
            INIT_59 => X"0000008e00000000000000630000000000000071000000000000008d00000000",
            INIT_5A => X"00000033000000000000004f0000000000000053000000000000005300000000",
            INIT_5B => X"00000022000000000000001f000000000000001c000000000000001d00000000",
            INIT_5C => X"0000006100000000000000510000000000000048000000000000003200000000",
            INIT_5D => X"00000085000000000000008a0000000000000074000000000000006600000000",
            INIT_5E => X"00000032000000000000001d000000000000001b000000000000003700000000",
            INIT_5F => X"000000c600000000000000a40000000000000059000000000000004c00000000",
            INIT_60 => X"00000090000000000000009b00000000000000a600000000000000a400000000",
            INIT_61 => X"0000006c00000000000000630000000000000082000000000000008b00000000",
            INIT_62 => X"0000003800000000000000480000000000000050000000000000004c00000000",
            INIT_63 => X"0000002900000000000000270000000000000024000000000000002600000000",
            INIT_64 => X"00000048000000000000003d0000000000000033000000000000002d00000000",
            INIT_65 => X"00000083000000000000007c0000000000000067000000000000005400000000",
            INIT_66 => X"000000320000000000000021000000000000001a000000000000003100000000",
            INIT_67 => X"000000c300000000000000a90000000000000059000000000000004500000000",
            INIT_68 => X"0000008d0000000000000092000000000000009400000000000000a000000000",
            INIT_69 => X"0000004900000000000000660000000000000082000000000000008700000000",
            INIT_6A => X"000000380000000000000042000000000000004d000000000000004500000000",
            INIT_6B => X"0000002d000000000000002b0000000000000028000000000000002f00000000",
            INIT_6C => X"0000003d00000000000000360000000000000030000000000000002e00000000",
            INIT_6D => X"0000006a000000000000005e0000000000000054000000000000004600000000",
            INIT_6E => X"00000030000000000000001f000000000000001a000000000000004000000000",
            INIT_6F => X"000000ba00000000000000af0000000000000062000000000000003d00000000",
            INIT_70 => X"0000008c000000000000008e000000000000008d000000000000009300000000",
            INIT_71 => X"000000390000000000000068000000000000008b000000000000008f00000000",
            INIT_72 => X"00000034000000000000003f000000000000004a000000000000004000000000",
            INIT_73 => X"0000003600000000000000330000000000000031000000000000003700000000",
            INIT_74 => X"00000042000000000000003d0000000000000036000000000000003600000000",
            INIT_75 => X"000000570000000000000051000000000000004a000000000000004400000000",
            INIT_76 => X"0000003400000000000000230000000000000021000000000000004800000000",
            INIT_77 => X"000000b500000000000000b60000000000000084000000000000004800000000",
            INIT_78 => X"000000a300000000000000a10000000000000096000000000000009200000000",
            INIT_79 => X"0000003a000000000000007c0000000000000091000000000000009d00000000",
            INIT_7A => X"0000004100000000000000390000000000000038000000000000003700000000",
            INIT_7B => X"0000004500000000000000460000000000000042000000000000004300000000",
            INIT_7C => X"0000005f00000000000000570000000000000048000000000000004300000000",
            INIT_7D => X"0000005e0000000000000060000000000000005f000000000000005c00000000",
            INIT_7E => X"00000046000000000000003e0000000000000044000000000000005100000000",
            INIT_7F => X"000000b900000000000000b600000000000000a3000000000000007600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "sampleifmap_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000b600000000000000bf00000000000000ca00000000000000d100000000",
            INIT_01 => X"000000af00000000000000c600000000000000d100000000000000d100000000",
            INIT_02 => X"000000a0000000000000009d00000000000000a500000000000000ab00000000",
            INIT_03 => X"0000008f000000000000008d000000000000009a000000000000009500000000",
            INIT_04 => X"000000db00000000000000d600000000000000bc00000000000000a400000000",
            INIT_05 => X"000000d600000000000000d900000000000000ca00000000000000d100000000",
            INIT_06 => X"000000ad00000000000000a100000000000000b100000000000000d000000000",
            INIT_07 => X"000000950000000000000095000000000000009d00000000000000b700000000",
            INIT_08 => X"000000cd00000000000000d200000000000000d400000000000000d400000000",
            INIT_09 => X"000000a300000000000000c800000000000000db00000000000000cf00000000",
            INIT_0A => X"000000b600000000000000b800000000000000b600000000000000a500000000",
            INIT_0B => X"000000d700000000000000cd00000000000000c900000000000000c200000000",
            INIT_0C => X"000000e400000000000000e300000000000000e300000000000000df00000000",
            INIT_0D => X"000000d700000000000000d300000000000000d400000000000000dd00000000",
            INIT_0E => X"000000bb00000000000000c300000000000000cd00000000000000df00000000",
            INIT_0F => X"000000ba00000000000000ad00000000000000aa00000000000000c600000000",
            INIT_10 => X"000000e200000000000000e300000000000000e500000000000000e600000000",
            INIT_11 => X"000000a400000000000000d300000000000000ec00000000000000e300000000",
            INIT_12 => X"000000b800000000000000b700000000000000ad000000000000009f00000000",
            INIT_13 => X"000000e000000000000000cf00000000000000bf00000000000000bc00000000",
            INIT_14 => X"000000d600000000000000e000000000000000e500000000000000db00000000",
            INIT_15 => X"000000d300000000000000c800000000000000d000000000000000d600000000",
            INIT_16 => X"000000c500000000000000db00000000000000e000000000000000de00000000",
            INIT_17 => X"000000c600000000000000c500000000000000bc00000000000000b900000000",
            INIT_18 => X"000000f100000000000000f400000000000000f400000000000000f500000000",
            INIT_19 => X"000000af00000000000000e300000000000000f100000000000000f200000000",
            INIT_1A => X"000000bb00000000000000a100000000000000b000000000000000a800000000",
            INIT_1B => X"000000b600000000000000b800000000000000a000000000000000ae00000000",
            INIT_1C => X"000000ca00000000000000d000000000000000d500000000000000b900000000",
            INIT_1D => X"000000d400000000000000c400000000000000ba00000000000000b900000000",
            INIT_1E => X"000000bb00000000000000d500000000000000dc00000000000000d700000000",
            INIT_1F => X"000000c800000000000000d400000000000000c500000000000000a900000000",
            INIT_20 => X"000000f400000000000000f400000000000000f300000000000000f500000000",
            INIT_21 => X"0000008400000000000000cd00000000000000f100000000000000f500000000",
            INIT_22 => X"000000a7000000000000008a00000000000000a1000000000000008b00000000",
            INIT_23 => X"0000008d000000000000009b000000000000008b000000000000009f00000000",
            INIT_24 => X"000000a4000000000000009900000000000000a6000000000000008e00000000",
            INIT_25 => X"000000e000000000000000c400000000000000a900000000000000a900000000",
            INIT_26 => X"000000b100000000000000d400000000000000d100000000000000d100000000",
            INIT_27 => X"000000d200000000000000cc00000000000000b800000000000000a000000000",
            INIT_28 => X"000000f300000000000000f400000000000000f400000000000000f500000000",
            INIT_29 => X"0000008100000000000000d700000000000000ee00000000000000f600000000",
            INIT_2A => X"000000aa00000000000000a0000000000000009c000000000000007100000000",
            INIT_2B => X"000000a700000000000000b100000000000000aa00000000000000aa00000000",
            INIT_2C => X"0000008f0000000000000098000000000000009d000000000000009d00000000",
            INIT_2D => X"000000e400000000000000cd00000000000000b3000000000000009400000000",
            INIT_2E => X"000000aa00000000000000c100000000000000ce00000000000000da00000000",
            INIT_2F => X"000000df00000000000000c000000000000000a0000000000000009300000000",
            INIT_30 => X"000000f400000000000000f300000000000000f300000000000000f500000000",
            INIT_31 => X"000000b400000000000000dd00000000000000dd00000000000000f100000000",
            INIT_32 => X"000000cf00000000000000c400000000000000b4000000000000008300000000",
            INIT_33 => X"000000d300000000000000d900000000000000cb00000000000000c800000000",
            INIT_34 => X"000000bf00000000000000c000000000000000c300000000000000cc00000000",
            INIT_35 => X"000000e100000000000000cd00000000000000a600000000000000a300000000",
            INIT_36 => X"000000a900000000000000b100000000000000d500000000000000e300000000",
            INIT_37 => X"000000da00000000000000b20000000000000092000000000000009100000000",
            INIT_38 => X"000000f700000000000000f200000000000000f200000000000000f400000000",
            INIT_39 => X"000000c000000000000000d900000000000000ca00000000000000e600000000",
            INIT_3A => X"000000e800000000000000e000000000000000c2000000000000008600000000",
            INIT_3B => X"000000d100000000000000ce00000000000000d700000000000000ea00000000",
            INIT_3C => X"000000cf00000000000000ca00000000000000d000000000000000cf00000000",
            INIT_3D => X"000000cc000000000000009a00000000000000b400000000000000e000000000",
            INIT_3E => X"000000bc00000000000000c400000000000000c900000000000000dc00000000",
            INIT_3F => X"000000c7000000000000009a000000000000009200000000000000ab00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000f500000000000000f300000000000000f300000000000000f500000000",
            INIT_41 => X"000000ae00000000000000df00000000000000d100000000000000e300000000",
            INIT_42 => X"000000c100000000000000c100000000000000ba000000000000008700000000",
            INIT_43 => X"000000c900000000000000c100000000000000cc00000000000000dd00000000",
            INIT_44 => X"000000c600000000000000cd00000000000000cd00000000000000ca00000000",
            INIT_45 => X"000000bc00000000000000a300000000000000d000000000000000dc00000000",
            INIT_46 => X"000000cb00000000000000df00000000000000d100000000000000cb00000000",
            INIT_47 => X"000000b20000000000000094000000000000008b00000000000000a100000000",
            INIT_48 => X"000000f200000000000000f300000000000000f100000000000000f200000000",
            INIT_49 => X"000000a400000000000000c200000000000000cd00000000000000e500000000",
            INIT_4A => X"000000b800000000000000bd00000000000000c1000000000000008c00000000",
            INIT_4B => X"000000c400000000000000c000000000000000c400000000000000ca00000000",
            INIT_4C => X"000000c600000000000000d000000000000000ca00000000000000c700000000",
            INIT_4D => X"000000c800000000000000bc00000000000000e000000000000000d700000000",
            INIT_4E => X"000000e300000000000000ed00000000000000ee00000000000000e600000000",
            INIT_4F => X"000000d300000000000000ca00000000000000ba00000000000000bc00000000",
            INIT_50 => X"000000f400000000000000f300000000000000ee00000000000000ea00000000",
            INIT_51 => X"0000009c00000000000000a900000000000000a000000000000000df00000000",
            INIT_52 => X"000000ac00000000000000b300000000000000b1000000000000008600000000",
            INIT_53 => X"000000b700000000000000b400000000000000ae00000000000000ae00000000",
            INIT_54 => X"000000be00000000000000bc00000000000000be00000000000000bb00000000",
            INIT_55 => X"000000c400000000000000d000000000000000dc00000000000000cd00000000",
            INIT_56 => X"000000f400000000000000f600000000000000e600000000000000d900000000",
            INIT_57 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_58 => X"000000f200000000000000f200000000000000e600000000000000d300000000",
            INIT_59 => X"0000009700000000000000be00000000000000b600000000000000d800000000",
            INIT_5A => X"000000a00000000000000093000000000000006e000000000000006a00000000",
            INIT_5B => X"000000aa00000000000000a6000000000000009f000000000000009e00000000",
            INIT_5C => X"000000a6000000000000009e00000000000000a300000000000000a900000000",
            INIT_5D => X"000000af00000000000000c600000000000000bd00000000000000ad00000000",
            INIT_5E => X"000000f300000000000000f800000000000000e000000000000000b700000000",
            INIT_5F => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_60 => X"000000e100000000000000e900000000000000da00000000000000c400000000",
            INIT_61 => X"0000009f00000000000000c300000000000000b400000000000000bd00000000",
            INIT_62 => X"000000a0000000000000008d000000000000005c000000000000005d00000000",
            INIT_63 => X"0000008c000000000000008f00000000000000a800000000000000ba00000000",
            INIT_64 => X"000000a700000000000000920000000000000089000000000000008b00000000",
            INIT_65 => X"00000096000000000000008f0000000000000083000000000000009800000000",
            INIT_66 => X"000000f400000000000000f300000000000000e300000000000000bc00000000",
            INIT_67 => X"000000f400000000000000f400000000000000f400000000000000f400000000",
            INIT_68 => X"000000c100000000000000d300000000000000c700000000000000c300000000",
            INIT_69 => X"0000008900000000000000a2000000000000009500000000000000a400000000",
            INIT_6A => X"000000a600000000000000b200000000000000aa000000000000009600000000",
            INIT_6B => X"0000009200000000000000a600000000000000cd00000000000000bd00000000",
            INIT_6C => X"000000d300000000000000c000000000000000ac000000000000009900000000",
            INIT_6D => X"0000008a0000000000000080000000000000008000000000000000af00000000",
            INIT_6E => X"000000d300000000000000bf00000000000000b100000000000000a000000000",
            INIT_6F => X"000000f300000000000000f300000000000000f500000000000000ef00000000",
            INIT_70 => X"000000a200000000000000c800000000000000cf00000000000000c200000000",
            INIT_71 => X"00000089000000000000008e0000000000000088000000000000009c00000000",
            INIT_72 => X"0000009f00000000000000b100000000000000b200000000000000a200000000",
            INIT_73 => X"0000008b000000000000009500000000000000a3000000000000009600000000",
            INIT_74 => X"0000009300000000000000920000000000000092000000000000008d00000000",
            INIT_75 => X"00000085000000000000007f000000000000007c000000000000008600000000",
            INIT_76 => X"000000a600000000000000ad00000000000000a3000000000000009500000000",
            INIT_77 => X"000000f400000000000000f300000000000000f500000000000000cc00000000",
            INIT_78 => X"0000006e00000000000000ad00000000000000d000000000000000c300000000",
            INIT_79 => X"000000b900000000000000b4000000000000008b000000000000007100000000",
            INIT_7A => X"00000057000000000000007f000000000000009a000000000000008500000000",
            INIT_7B => X"0000005f0000000000000059000000000000004c000000000000004900000000",
            INIT_7C => X"00000058000000000000005e0000000000000060000000000000005c00000000",
            INIT_7D => X"0000006700000000000000630000000000000056000000000000005600000000",
            INIT_7E => X"0000009b000000000000008f0000000000000074000000000000006d00000000",
            INIT_7F => X"000000f500000000000000f500000000000000e800000000000000af00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "sampleifmap_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000006500000000000000a100000000000000aa00000000000000b700000000",
            INIT_01 => X"000000a100000000000000b50000000000000088000000000000006000000000",
            INIT_02 => X"0000008700000000000000810000000000000084000000000000008000000000",
            INIT_03 => X"0000006a000000000000007d000000000000007d000000000000008c00000000",
            INIT_04 => X"00000027000000000000002c000000000000002b000000000000003500000000",
            INIT_05 => X"0000002800000000000000230000000000000047000000000000004d00000000",
            INIT_06 => X"0000009700000000000000910000000000000050000000000000002000000000",
            INIT_07 => X"000000f300000000000000f600000000000000db00000000000000a700000000",
            INIT_08 => X"0000007c00000000000000c200000000000000c100000000000000ca00000000",
            INIT_09 => X"0000004900000000000000990000000000000092000000000000007800000000",
            INIT_0A => X"0000009400000000000000830000000000000087000000000000006900000000",
            INIT_0B => X"0000008300000000000000a9000000000000009f00000000000000b800000000",
            INIT_0C => X"0000007a00000000000000840000000000000076000000000000006600000000",
            INIT_0D => X"00000073000000000000006f00000000000000aa00000000000000af00000000",
            INIT_0E => X"000000b500000000000000b20000000000000091000000000000006f00000000",
            INIT_0F => X"000000f400000000000000f200000000000000c500000000000000bb00000000",
            INIT_10 => X"0000007200000000000000b800000000000000c800000000000000d800000000",
            INIT_11 => X"000000240000000000000082000000000000009d000000000000007300000000",
            INIT_12 => X"0000006300000000000000810000000000000095000000000000004f00000000",
            INIT_13 => X"00000084000000000000009d0000000000000081000000000000006f00000000",
            INIT_14 => X"000000b900000000000000b700000000000000c100000000000000b100000000",
            INIT_15 => X"000000bd00000000000000ba00000000000000c100000000000000c800000000",
            INIT_16 => X"0000009700000000000000b600000000000000c700000000000000b500000000",
            INIT_17 => X"000000f600000000000000e800000000000000a2000000000000009400000000",
            INIT_18 => X"0000007100000000000000bb00000000000000cc00000000000000d900000000",
            INIT_19 => X"0000003d0000000000000071000000000000008b000000000000006000000000",
            INIT_1A => X"0000005d00000000000000730000000000000070000000000000004e00000000",
            INIT_1B => X"0000007d000000000000005e0000000000000053000000000000005500000000",
            INIT_1C => X"0000008a000000000000007f000000000000009f00000000000000bf00000000",
            INIT_1D => X"0000008f000000000000008c000000000000009500000000000000a000000000",
            INIT_1E => X"00000063000000000000009f00000000000000bd000000000000008a00000000",
            INIT_1F => X"000000f700000000000000e2000000000000009a000000000000007300000000",
            INIT_20 => X"0000007500000000000000c700000000000000d000000000000000d500000000",
            INIT_21 => X"000000540000000000000063000000000000005c000000000000004900000000",
            INIT_22 => X"0000006900000000000000610000000000000041000000000000004b00000000",
            INIT_23 => X"0000005f00000000000000670000000000000057000000000000005f00000000",
            INIT_24 => X"00000097000000000000009900000000000000a2000000000000008600000000",
            INIT_25 => X"0000008f00000000000000890000000000000090000000000000009600000000",
            INIT_26 => X"0000006f000000000000008f0000000000000099000000000000009300000000",
            INIT_27 => X"000000f700000000000000de0000000000000092000000000000007300000000",
            INIT_28 => X"0000008300000000000000cc00000000000000ce00000000000000cc00000000",
            INIT_29 => X"0000005a000000000000005c0000000000000051000000000000006500000000",
            INIT_2A => X"000000450000000000000039000000000000002d000000000000004600000000",
            INIT_2B => X"00000057000000000000007d000000000000006f000000000000006200000000",
            INIT_2C => X"0000006700000000000000700000000000000066000000000000004a00000000",
            INIT_2D => X"0000007d000000000000005e0000000000000065000000000000006200000000",
            INIT_2E => X"0000009500000000000000710000000000000052000000000000007300000000",
            INIT_2F => X"000000f800000000000000d40000000000000089000000000000009a00000000",
            INIT_30 => X"0000007500000000000000ce00000000000000d000000000000000d100000000",
            INIT_31 => X"0000005e0000000000000056000000000000007a000000000000006900000000",
            INIT_32 => X"0000002f00000000000000330000000000000036000000000000005600000000",
            INIT_33 => X"0000006300000000000000ad0000000000000083000000000000006600000000",
            INIT_34 => X"00000082000000000000009e0000000000000064000000000000002d00000000",
            INIT_35 => X"000000ab000000000000007c000000000000008a000000000000007900000000",
            INIT_36 => X"000000ab000000000000005f000000000000004b00000000000000bb00000000",
            INIT_37 => X"000000fa00000000000000cf0000000000000075000000000000009800000000",
            INIT_38 => X"0000006800000000000000cc00000000000000d600000000000000dd00000000",
            INIT_39 => X"0000008000000000000000720000000000000074000000000000003b00000000",
            INIT_3A => X"0000003000000000000000340000000000000041000000000000007c00000000",
            INIT_3B => X"0000004b000000000000006c0000000000000046000000000000003800000000",
            INIT_3C => X"0000008f00000000000000a6000000000000005f000000000000003000000000",
            INIT_3D => X"000000af000000000000008f00000000000000a7000000000000009100000000",
            INIT_3E => X"000000620000000000000048000000000000004a00000000000000af00000000",
            INIT_3F => X"000000fb00000000000000d60000000000000068000000000000005400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006300000000000000c900000000000000d400000000000000d700000000",
            INIT_41 => X"000000b000000000000000800000000000000044000000000000002f00000000",
            INIT_42 => X"0000002d00000000000000380000000000000050000000000000008700000000",
            INIT_43 => X"0000002f000000000000002b0000000000000027000000000000002800000000",
            INIT_44 => X"0000006e0000000000000050000000000000003c000000000000003700000000",
            INIT_45 => X"0000008b00000000000000900000000000000093000000000000007d00000000",
            INIT_46 => X"0000004300000000000000460000000000000043000000000000005c00000000",
            INIT_47 => X"000000fb00000000000000d9000000000000006d000000000000004500000000",
            INIT_48 => X"0000009d00000000000000cb00000000000000cf00000000000000cf00000000",
            INIT_49 => X"000000aa00000000000000850000000000000075000000000000007300000000",
            INIT_4A => X"0000003000000000000000480000000000000065000000000000007e00000000",
            INIT_4B => X"0000002d00000000000000290000000000000029000000000000002800000000",
            INIT_4C => X"000000c000000000000000530000000000000027000000000000003200000000",
            INIT_4D => X"000000c900000000000000c700000000000000dc00000000000000da00000000",
            INIT_4E => X"0000003f00000000000000380000000000000034000000000000006b00000000",
            INIT_4F => X"000000f700000000000000d2000000000000007e000000000000005a00000000",
            INIT_50 => X"000000d800000000000000ce00000000000000c000000000000000bc00000000",
            INIT_51 => X"000000a10000000000000086000000000000009a00000000000000bf00000000",
            INIT_52 => X"0000003e00000000000000680000000000000073000000000000007900000000",
            INIT_53 => X"0000002900000000000000230000000000000022000000000000002100000000",
            INIT_54 => X"000000b300000000000000550000000000000031000000000000003300000000",
            INIT_55 => X"000000bb00000000000000be00000000000000c000000000000000c700000000",
            INIT_56 => X"0000004200000000000000260000000000000027000000000000006000000000",
            INIT_57 => X"000000f500000000000000d10000000000000085000000000000006f00000000",
            INIT_58 => X"000000c600000000000000cd00000000000000c600000000000000bf00000000",
            INIT_59 => X"000000a00000000000000084000000000000009e00000000000000b500000000",
            INIT_5A => X"00000046000000000000006f0000000000000076000000000000007200000000",
            INIT_5B => X"00000031000000000000002c0000000000000026000000000000002700000000",
            INIT_5C => X"0000007e0000000000000069000000000000005d000000000000004400000000",
            INIT_5D => X"000000a600000000000000ad0000000000000096000000000000008700000000",
            INIT_5E => X"00000047000000000000002a0000000000000028000000000000004800000000",
            INIT_5F => X"000000f200000000000000cf0000000000000082000000000000007100000000",
            INIT_60 => X"000000b800000000000000c600000000000000d100000000000000ce00000000",
            INIT_61 => X"00000085000000000000008200000000000000a300000000000000ab00000000",
            INIT_62 => X"0000004d0000000000000068000000000000006f000000000000006b00000000",
            INIT_63 => X"000000390000000000000035000000000000002f000000000000003200000000",
            INIT_64 => X"0000006800000000000000570000000000000048000000000000003f00000000",
            INIT_65 => X"000000b000000000000000a80000000000000091000000000000007800000000",
            INIT_66 => X"0000004700000000000000300000000000000028000000000000004500000000",
            INIT_67 => X"000000ee00000000000000d4000000000000007e000000000000006600000000",
            INIT_68 => X"000000bd00000000000000c200000000000000c200000000000000c700000000",
            INIT_69 => X"00000065000000000000008600000000000000a600000000000000b200000000",
            INIT_6A => X"0000004f00000000000000600000000000000069000000000000006300000000",
            INIT_6B => X"0000003e000000000000003b0000000000000036000000000000003e00000000",
            INIT_6C => X"00000057000000000000004e0000000000000045000000000000004100000000",
            INIT_6D => X"0000008f00000000000000810000000000000074000000000000006400000000",
            INIT_6E => X"00000047000000000000002c0000000000000027000000000000005700000000",
            INIT_6F => X"000000e800000000000000df0000000000000085000000000000005900000000",
            INIT_70 => X"000000bc00000000000000be00000000000000bc00000000000000c100000000",
            INIT_71 => X"00000050000000000000009000000000000000bc00000000000000bd00000000",
            INIT_72 => X"0000004600000000000000580000000000000063000000000000005a00000000",
            INIT_73 => X"0000004e000000000000004a0000000000000045000000000000004900000000",
            INIT_74 => X"0000005d0000000000000056000000000000004e000000000000004e00000000",
            INIT_75 => X"00000072000000000000006d0000000000000066000000000000006100000000",
            INIT_76 => X"0000004a00000000000000300000000000000030000000000000005e00000000",
            INIT_77 => X"000000e700000000000000e800000000000000ad000000000000006400000000",
            INIT_78 => X"000000cd00000000000000d000000000000000c700000000000000c400000000",
            INIT_79 => X"0000005500000000000000a500000000000000bb00000000000000c800000000",
            INIT_7A => X"00000054000000000000004e000000000000004c000000000000004c00000000",
            INIT_7B => X"0000006300000000000000620000000000000059000000000000005400000000",
            INIT_7C => X"0000007c00000000000000720000000000000063000000000000005e00000000",
            INIT_7D => X"0000007f00000000000000800000000000000081000000000000007d00000000",
            INIT_7E => X"000000600000000000000054000000000000005b000000000000007000000000",
            INIT_7F => X"000000df00000000000000e100000000000000cc000000000000009400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEIFMAP_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0 : if BRAM_NAME = "samplegold_layersamples_instance0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000014000000000000000f0000000000000012000000000000001200000000",
            INIT_01 => X"0000001d000000000000000f000000000000000d000000000000001700000000",
            INIT_02 => X"000000010000000000000000000000000000000a000000000000001d00000000",
            INIT_03 => X"000000160000000000000015000000000000000c000000000000000600000000",
            INIT_04 => X"000000130000000000000013000000000000000f000000000000001200000000",
            INIT_05 => X"0000000000000000000000030000000000000008000000000000000400000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_07 => X"0000000b0000000000000000000000000000000b000000000000000500000000",
            INIT_08 => X"0000001b0000000000000012000000000000001b000000000000001300000000",
            INIT_09 => X"000000000000000000000000000000000000001e000000000000002000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000c00000000000000000000000000000001000000000000000100000000",
            INIT_0C => X"000000000000000000000011000000000000000b000000000000001900000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000300000000000000030000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"000000000000000000000000000000000000001c000000000000000400000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_20 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000007000000000000000400000000",
            INIT_5A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000a000000000000003f000000000000000f000000000000001a00000000",
            INIT_62 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000002000000000000000250000000000000038000000000000003a00000000",
            INIT_64 => X"0000002700000000000000250000000000000029000000000000002200000000",
            INIT_65 => X"00000000000000000000003a000000000000002c000000000000002000000000",
            INIT_66 => X"0000001d000000000000001d000000000000001e000000000000000000000000",
            INIT_67 => X"00000024000000000000001f0000000000000020000000000000002000000000",
            INIT_68 => X"0000002100000000000000280000000000000022000000000000001e00000000",
            INIT_69 => X"0000000e000000000000002f000000000000002f000000000000003000000000",
            INIT_6A => X"0000001d00000000000000190000000000000021000000000000000f00000000",
            INIT_6B => X"00000033000000000000002f0000000000000023000000000000002200000000",
            INIT_6C => X"00000029000000000000003a0000000000000028000000000000003400000000",
            INIT_6D => X"0000002a00000000000000410000000000000031000000000000003300000000",
            INIT_6E => X"00000017000000000000001f000000000000002a000000000000003000000000",
            INIT_6F => X"0000001a000000000000002d0000000000000021000000000000001c00000000",
            INIT_70 => X"0000000000000000000000000000000000000029000000000000001c00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000006000000000000000e0000000000000018000000000000000300000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_7D => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_7E => X"0000000000000000000000060000000000000000000000000000001b00000000",
            INIT_7F => X"0000001e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE0;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1 : if BRAM_NAME = "samplegold_layersamples_instance1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001400000000000000110000000000000000000000000000000000000000",
            INIT_01 => X"0000001d00000000000000000000000000000003000000000000000500000000",
            INIT_02 => X"0000000000000000000000080000000000000000000000000000001000000000",
            INIT_03 => X"000000000000000000000017000000000000000f000000000000000300000000",
            INIT_04 => X"00000006000000000000000a000000000000001a000000000000000000000000",
            INIT_05 => X"0000000300000000000000440000000000000000000000000000000400000000",
            INIT_06 => X"000000020000000000000000000000000000000b000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000000b000000000000001700000000",
            INIT_08 => X"00000000000000000000000b000000000000001e000000000000000c00000000",
            INIT_09 => X"0000000400000000000000000000000000000037000000000000000000000000",
            INIT_0A => X"0000002000000000000000020000000000000011000000000000000a00000000",
            INIT_0B => X"0000000600000000000000000000000000000006000000000000001400000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_0D => X"0000001100000000000000000000000000000000000000000000002000000000",
            INIT_0E => X"00000028000000000000001d0000000000000000000000000000000800000000",
            INIT_0F => X"0000000000000000000000080000000000000011000000000000000400000000",
            INIT_10 => X"00000000000000000000000b000000000000000b000000000000000000000000",
            INIT_11 => X"0000000000000000000000060000000000000000000000000000001000000000",
            INIT_12 => X"0000000000000000000000240000000000000018000000000000000000000000",
            INIT_13 => X"000000120000000000000009000000000000000e000000000000002700000000",
            INIT_14 => X"0000000000000000000000000000000000000015000000000000001200000000",
            INIT_15 => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_16 => X"0000005800000000000000000000000000000023000000000000002b00000000",
            INIT_17 => X"00000011000000000000002d0000000000000028000000000000000d00000000",
            INIT_18 => X"00000022000000000000001b0000000000000000000000000000000000000000",
            INIT_19 => X"000000360000000000000000000000000000000b000000000000001f00000000",
            INIT_1A => X"0000000000000000000000450000000000000012000000000000002300000000",
            INIT_1B => X"0000001a0000000000000021000000000000001f000000000000000700000000",
            INIT_1C => X"0000002e00000000000000280000000000000022000000000000001e00000000",
            INIT_1D => X"00000038000000000000002a000000000000002f000000000000002f00000000",
            INIT_1E => X"0000002700000000000000000000000000000025000000000000003300000000",
            INIT_1F => X"0000002a00000000000000240000000000000024000000000000002500000000",
            INIT_20 => X"0000002e000000000000002f0000000000000036000000000000002f00000000",
            INIT_21 => X"00000052000000000000002e000000000000002c000000000000003a00000000",
            INIT_22 => X"00000026000000000000002b0000000000000013000000000000000000000000",
            INIT_23 => X"0000002e000000000000002f000000000000002a000000000000002a00000000",
            INIT_24 => X"000000280000000000000045000000000000002a000000000000002f00000000",
            INIT_25 => X"00000019000000000000002c0000000000000033000000000000002b00000000",
            INIT_26 => X"0000002400000000000000230000000000000028000000000000001900000000",
            INIT_27 => X"0000002e000000000000002d0000000000000031000000000000002e00000000",
            INIT_28 => X"00000000000000000000001f000000000000003a000000000000004300000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000000000000000000000a000000000000000200000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000170000000000000008000000000000001000000000",
            INIT_2F => X"000000000000000000000003000000000000001c000000000000001f00000000",
            INIT_30 => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_31 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000004200000000000000000000000000000000000000000000001100000000",
            INIT_33 => X"000000000000000000000000000000000000003f000000000000002d00000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000007100000000",
            INIT_35 => X"0000002c00000000000000280000000000000000000000000000000e00000000",
            INIT_36 => X"00000026000000000000005a0000000000000000000000000000002500000000",
            INIT_37 => X"0000006c0000000000000000000000000000002a000000000000003b00000000",
            INIT_38 => X"0000003400000000000000000000000000000023000000000000000500000000",
            INIT_39 => X"0000003c0000000000000048000000000000005d000000000000002400000000",
            INIT_3A => X"0000001e0000000000000052000000000000002f000000000000000000000000",
            INIT_3B => X"0000003100000000000000590000000000000000000000000000003e00000000",
            INIT_3C => X"0000002c00000000000000000000000000000000000000000000003700000000",
            INIT_3D => X"000000000000000000000060000000000000003e000000000000006100000000",
            INIT_3E => X"000000310000000000000012000000000000005c000000000000007300000000",
            INIT_3F => X"0000001500000000000000730000000000000048000000000000002500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005a00000000000000000000000000000000000000000000003800000000",
            INIT_41 => X"000000750000000000000000000000000000006a000000000000004a00000000",
            INIT_42 => X"00000037000000000000000c0000000000000012000000000000004700000000",
            INIT_43 => X"0000003100000000000000280000000000000065000000000000004d00000000",
            INIT_44 => X"00000038000000000000008b0000000000000006000000000000000000000000",
            INIT_45 => X"00000050000000000000004f0000000000000000000000000000004600000000",
            INIT_46 => X"0000006800000000000000130000000000000025000000000000000600000000",
            INIT_47 => X"0000002a000000000000000b0000000000000084000000000000004200000000",
            INIT_48 => X"00000000000000000000002c000000000000002e000000000000001300000000",
            INIT_49 => X"00000004000000000000005b0000000000000016000000000000002900000000",
            INIT_4A => X"0000003a000000000000004a0000000000000000000000000000000000000000",
            INIT_4B => X"0000001800000000000000640000000000000000000000000000009f00000000",
            INIT_4C => X"0000003b0000000000000030000000000000004d000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000017000000000000005a00000000",
            INIT_4E => X"00000094000000000000003c000000000000000f000000000000000c00000000",
            INIT_4F => X"00000020000000000000004c0000000000000093000000000000000000000000",
            INIT_50 => X"0000001a00000000000000410000000000000083000000000000007100000000",
            INIT_51 => X"0000003100000000000000200000000000000023000000000000001d00000000",
            INIT_52 => X"00000000000000000000004e000000000000002b000000000000001d00000000",
            INIT_53 => X"0000003c000000000000003a000000000000007300000000000000d800000000",
            INIT_54 => X"0000003c000000000000003d0000000000000038000000000000004700000000",
            INIT_55 => X"0000005f000000000000004f0000000000000040000000000000003e00000000",
            INIT_56 => X"000000af00000000000000820000000000000000000000000000001200000000",
            INIT_57 => X"0000003e000000000000003f0000000000000049000000000000004200000000",
            INIT_58 => X"0000005000000000000000400000000000000038000000000000003900000000",
            INIT_59 => X"00000045000000000000006a000000000000003d000000000000004800000000",
            INIT_5A => X"00000039000000000000005a00000000000000cb000000000000000000000000",
            INIT_5B => X"00000041000000000000003c0000000000000042000000000000004d00000000",
            INIT_5C => X"00000038000000000000004e000000000000004d000000000000004800000000",
            INIT_5D => X"0000003e000000000000004b0000000000000076000000000000007b00000000",
            INIT_5E => X"0000004300000000000000350000000000000048000000000000005400000000",
            INIT_5F => X"0000005500000000000000440000000000000038000000000000004400000000",
            INIT_60 => X"00000080000000000000006f000000000000001a000000000000003a00000000",
            INIT_61 => X"0000000800000000000000080000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000050000000000000003000000000000000600000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_64 => X"0000000700000000000000050000000000000006000000000000000000000000",
            INIT_65 => X"0000000a0000000000000007000000000000000c000000000000000a00000000",
            INIT_66 => X"000000000000000000000000000000000000001a000000000000004900000000",
            INIT_67 => X"0000000000000000000000060000000000000024000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_69 => X"0000000000000000000000070000000000000004000000000000000400000000",
            INIT_6A => X"0000001a000000000000000d0000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000170000000000000007000000000000001500000000",
            INIT_6C => X"0000000900000000000000250000000000000028000000000000000000000000",
            INIT_6D => X"000000370000000000000000000000000000000d000000000000000500000000",
            INIT_6E => X"0000000000000000000000000000000000000005000000000000001b00000000",
            INIT_6F => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_70 => X"0000000b0000000000000013000000000000005a000000000000002600000000",
            INIT_71 => X"0000000e00000000000000060000000000000056000000000000008000000000",
            INIT_72 => X"0000002500000000000000250000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000018000000000000000f00000000",
            INIT_74 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_75 => X"0000001f000000000000001a000000000000002a000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_77 => X"0000000700000000000000060000000000000027000000000000000900000000",
            INIT_78 => X"0000002100000000000000000000000000000004000000000000000000000000",
            INIT_79 => X"000000110000000000000009000000000000000a000000000000000000000000",
            INIT_7A => X"000000170000000000000000000000000000000b000000000000000000000000",
            INIT_7B => X"0000001c00000000000000070000000000000015000000000000001d00000000",
            INIT_7C => X"0000000000000000000000160000000000000019000000000000001000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000004000000000000000b0000000000000004000000000000001000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE1;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2 : if BRAM_NAME = "samplegold_layersamples_instance2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001a00000000000000000000000000000000000000000000001c00000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_02 => X"00000000000000000000002f0000000000000003000000000000000000000000",
            INIT_03 => X"0000001100000000000000040000000000000009000000000000000000000000",
            INIT_04 => X"0000000c000000000000004a0000000000000000000000000000000000000000",
            INIT_05 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_07 => X"00000085000000000000009c0000000000000046000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_09 => X"00000000000000000000001b0000000000000041000000000000002000000000",
            INIT_0A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000004600000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000001200000000000000070000000000000004000000000000000000000000",
            INIT_11 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000001300000000000000140000000000000000000000000000000000000000",
            INIT_18 => X"0000002200000000000000280000000000000000000000000000000400000000",
            INIT_19 => X"000000a200000000000000a3000000000000009d000000000000000000000000",
            INIT_1A => X"000000ac000000000000009d00000000000000a400000000000000a500000000",
            INIT_1B => X"0000007c000000000000009400000000000000ad00000000000000b700000000",
            INIT_1C => X"0000009200000000000000920000000000000084000000000000007c00000000",
            INIT_1D => X"000000ac00000000000000a800000000000000ad00000000000000a200000000",
            INIT_1E => X"000000a000000000000000a9000000000000008c00000000000000a000000000",
            INIT_1F => X"0000003e000000000000002e000000000000003a000000000000007a00000000",
            INIT_20 => X"00000089000000000000008b000000000000006e000000000000004e00000000",
            INIT_21 => X"000000af00000000000000b000000000000000ac000000000000006a00000000",
            INIT_22 => X"0000002d00000000000000480000000000000073000000000000008e00000000",
            INIT_23 => X"00000027000000000000000a000000000000001e000000000000000700000000",
            INIT_24 => X"0000002b000000000000004d0000000000000067000000000000003a00000000",
            INIT_25 => X"0000005900000000000000a200000000000000aa00000000000000a400000000",
            INIT_26 => X"0000000c00000000000000150000000000000027000000000000004d00000000",
            INIT_27 => X"00000025000000000000001b000000000000002d000000000000003300000000",
            INIT_28 => X"00000094000000000000001f0000000000000017000000000000003a00000000",
            INIT_29 => X"000000430000000000000047000000000000004e000000000000006000000000",
            INIT_2A => X"000000310000000000000000000000000000001f000000000000002f00000000",
            INIT_2B => X"0000002f000000000000001c0000000000000017000000000000003900000000",
            INIT_2C => X"00000099000000000000008e0000000000000012000000000000001600000000",
            INIT_2D => X"000000310000000000000045000000000000003b000000000000002500000000",
            INIT_2E => X"0000002a000000000000003e0000000000000000000000000000002d00000000",
            INIT_2F => X"0000000e00000000000000170000000000000012000000000000001000000000",
            INIT_30 => X"0000002f000000000000009f0000000000000062000000000000002a00000000",
            INIT_31 => X"0000002f000000000000002d000000000000003e000000000000003200000000",
            INIT_32 => X"0000001000000000000000280000000000000032000000000000000000000000",
            INIT_33 => X"0000000a000000000000001c0000000000000026000000000000000e00000000",
            INIT_34 => X"0000002600000000000000370000000000000062000000000000002c00000000",
            INIT_35 => X"0000001e00000000000000290000000000000027000000000000002e00000000",
            INIT_36 => X"000000220000000000000009000000000000002d000000000000002f00000000",
            INIT_37 => X"0000002b00000000000000000000000000000014000000000000004100000000",
            INIT_38 => X"0000003600000000000000220000000000000055000000000000000e00000000",
            INIT_39 => X"000000420000000000000054000000000000000d000000000000003000000000",
            INIT_3A => X"00000079000000000000002d000000000000000f000000000000002600000000",
            INIT_3B => X"0000000000000000000000240000000000000005000000000000001000000000",
            INIT_3C => X"0000002800000000000000080000000000000020000000000000003500000000",
            INIT_3D => X"00000006000000000000001d0000000000000034000000000000002d00000000",
            INIT_3E => X"00000000000000000000008a0000000000000062000000000000000900000000",
            INIT_3F => X"0000001700000000000000000000000000000023000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000600000000000000000000000000000000000000000000001a00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"00000000000000000000003a0000000000000006000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000002300000000000000220000000000000000000000000000000000000000",
            INIT_52 => X"00000027000000000000001e0000000000000020000000000000002500000000",
            INIT_53 => X"00000017000000000000001d0000000000000024000000000000002600000000",
            INIT_54 => X"0000001e00000000000000240000000000000026000000000000001a00000000",
            INIT_55 => X"0000002a000000000000002c0000000000000023000000000000001800000000",
            INIT_56 => X"0000000f00000000000000200000000000000028000000000000001f00000000",
            INIT_57 => X"00000000000000000000001d000000000000000e000000000000001d00000000",
            INIT_58 => X"0000001c000000000000002b0000000000000020000000000000000900000000",
            INIT_59 => X"0000002100000000000000280000000000000039000000000000000600000000",
            INIT_5A => X"000000060000000000000000000000000000001a000000000000002700000000",
            INIT_5B => X"000000000000000000000000000000000000002e000000000000002100000000",
            INIT_5C => X"00000000000000000000002c0000000000000025000000000000000000000000",
            INIT_5D => X"0000000f00000000000000290000000000000021000000000000004c00000000",
            INIT_5E => X"0000000000000000000000000000000000000004000000000000002400000000",
            INIT_5F => X"0000000000000000000000090000000000000000000000000000004800000000",
            INIT_60 => X"000000260000000000000000000000000000004a000000000000000000000000",
            INIT_61 => X"0000000b00000000000000090000000000000056000000000000000200000000",
            INIT_62 => X"0000005900000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_64 => X"00000000000000000000000a0000000000000000000000000000002b00000000",
            INIT_65 => X"000000000000000000000013000000000000003e000000000000001a00000000",
            INIT_66 => X"00000000000000000000008e0000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_68 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000036000000000000003f00000000",
            INIT_6A => X"0000000000000000000000000000000000000066000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000015000000000000000a00000000",
            INIT_6C => X"0000003800000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000004200000000",
            INIT_6E => X"0000001d00000000000000000000000000000000000000000000004200000000",
            INIT_6F => X"0000000200000000000000000000000000000008000000000000000f00000000",
            INIT_70 => X"0000001100000000000000040000000000000021000000000000000000000000",
            INIT_71 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_72 => X"00000021000000000000001e0000000000000000000000000000002500000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_74 => X"00000027000000000000000f0000000000000000000000000000002c00000000",
            INIT_75 => X"0000000000000000000000050000000000000002000000000000000000000000",
            INIT_76 => X"0000001400000000000000340000000000000030000000000000000c00000000",
            INIT_77 => X"0000007800000000000000000000000000000004000000000000002a00000000",
            INIT_78 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_79 => X"0000000900000000000000080000000000000000000000000000000000000000",
            INIT_7A => X"0000002000000000000000000000000000000000000000000000000100000000",
            INIT_7B => X"0000000000000000000000400000000000000000000000000000001400000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE2;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3 : if BRAM_NAME = "samplegold_layersamples_instance3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000005d00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000002b00000000000000000000000000000000000000000000000400000000",
            INIT_0A => X"0000002f000000000000002c000000000000002d000000000000003000000000",
            INIT_0B => X"00000037000000000000003a0000000000000030000000000000002900000000",
            INIT_0C => X"0000002700000000000000260000000000000025000000000000002a00000000",
            INIT_0D => X"00000035000000000000002c0000000000000031000000000000002a00000000",
            INIT_0E => X"00000000000000000000002d000000000000002e000000000000003000000000",
            INIT_0F => X"0000000c000000000000003b0000000000000029000000000000001f00000000",
            INIT_10 => X"0000001f000000000000000e0000000000000000000000000000000000000000",
            INIT_11 => X"0000002e0000000000000029000000000000001c000000000000002500000000",
            INIT_12 => X"0000002d000000000000003b0000000000000032000000000000003500000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_14 => X"0000001a00000000000000040000000000000000000000000000000000000000",
            INIT_15 => X"0000003200000000000000230000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000019000000000000002500000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000110000000000000000000000000000000600000000",
            INIT_19 => X"0000000000000000000000180000000000000012000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_1D => X"0000000300000000000000030000000000000038000000000000000b00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000007000000000000003a00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000005000000000000001a00000000",
            INIT_2A => X"0000000400000000000000180000000000000003000000000000000f00000000",
            INIT_2B => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000000000a000000000000001100000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000800000000000000080000000000000011000000000000000a00000000",
            INIT_43 => X"0000000b000000000000000c000000000000000c000000000000000400000000",
            INIT_44 => X"00000023000000000000002d0000000000000021000000000000000b00000000",
            INIT_45 => X"0000000000000000000000060000000000000008000000000000001100000000",
            INIT_46 => X"00000008000000000000000c000000000000000a000000000000000a00000000",
            INIT_47 => X"0000004200000000000000230000000000000005000000000000000000000000",
            INIT_48 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"000000330000000000000035000000000000000a000000000000001700000000",
            INIT_4A => X"0000003700000000000000050000000000000008000000000000000500000000",
            INIT_4B => X"0000000000000000000000000000000000000009000000000000001600000000",
            INIT_4C => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000500000000000000000000000000000000000000000000000c00000000",
            INIT_4E => X"0000000000000000000000000000000000000008000000000000000800000000",
            INIT_4F => X"00000004000000000000001a0000000000000000000000000000000200000000",
            INIT_50 => X"0000000e00000000000000000000000000000006000000000000001000000000",
            INIT_51 => X"0000000e00000000000000020000000000000000000000000000000100000000",
            INIT_52 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_54 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000003e00000000000000030000000000000006000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_57 => X"0000000700000000000000150000000000000014000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000120000000000000018000000000000001c00000000",
            INIT_5A => X"0000000000000000000000110000000000000000000000000000003100000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000003500000000000000350000000000000002000000000000000000000000",
            INIT_5E => X"000000090000000000000000000000000000000e000000000000002100000000",
            INIT_5F => X"00000000000000000000000e0000000000000005000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000026000000000000000000000000",
            INIT_62 => X"0000003000000000000000260000000000000000000000000000000000000000",
            INIT_63 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000002300000000000000000000000000000004000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_66 => X"0000000000000000000000110000000000000036000000000000004e00000000",
            INIT_67 => X"0000000000000000000000030000000000000018000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_69 => X"0000000000000000000000370000000000000051000000000000001e00000000",
            INIT_6A => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000c00000000000000210000000000000035000000000000000a00000000",
            INIT_6C => X"0000000400000000000000280000000000000056000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000003000000000000000500000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000001800000000000000000000000000000016000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000b000000000000004f0000000000000018000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_77 => X"0000000300000000000000000000000000000022000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000a0000000000000013000000000000000d000000000000000000000000",
            INIT_7B => X"0000000800000000000000150000000000000009000000000000000e00000000",
            INIT_7C => X"00000022000000000000001c000000000000000c000000000000000600000000",
            INIT_7D => X"0000000200000000000000060000000000000013000000000000001b00000000",
            INIT_7E => X"0000000d0000000000000009000000000000000b000000000000000800000000",
            INIT_7F => X"0000001a000000000000000f0000000000000036000000000000000f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE3;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4 : if BRAM_NAME = "samplegold_layersamples_instance4" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002400000000000000350000000000000034000000000000001f00000000",
            INIT_01 => X"00000026000000000000000a000000000000001a000000000000002100000000",
            INIT_02 => X"00000008000000000000000a000000000000000b000000000000002400000000",
            INIT_03 => X"0000002000000000000000280000000000000033000000000000005100000000",
            INIT_04 => X"0000002b000000000000004b000000000000005e000000000000005300000000",
            INIT_05 => X"000000140000000000000033000000000000001a000000000000001900000000",
            INIT_06 => X"0000002e00000000000000190000000000000012000000000000000e00000000",
            INIT_07 => X"0000005b0000000000000036000000000000002f000000000000004500000000",
            INIT_08 => X"00000015000000000000003b0000000000000042000000000000005d00000000",
            INIT_09 => X"00000015000000000000005e0000000000000071000000000000001b00000000",
            INIT_0A => X"000000640000000000000044000000000000007e000000000000003500000000",
            INIT_0B => X"00000067000000000000003b0000000000000033000000000000003b00000000",
            INIT_0C => X"0000000100000000000000250000000000000039000000000000003800000000",
            INIT_0D => X"000000130000000000000028000000000000009e000000000000007f00000000",
            INIT_0E => X"0000004b000000000000007d000000000000007e00000000000000bd00000000",
            INIT_0F => X"00000050000000000000007f000000000000005b000000000000002e00000000",
            INIT_10 => X"0000007a0000000000000015000000000000003c000000000000004700000000",
            INIT_11 => X"0000005a00000000000000170000000000000043000000000000009400000000",
            INIT_12 => X"0000004e000000000000006500000000000000a8000000000000007500000000",
            INIT_13 => X"0000003b00000000000000460000000000000081000000000000007800000000",
            INIT_14 => X"000000a5000000000000008e0000000000000033000000000000004c00000000",
            INIT_15 => X"000000a500000000000000390000000000000039000000000000004000000000",
            INIT_16 => X"0000005f0000000000000050000000000000006a000000000000008500000000",
            INIT_17 => X"0000004b0000000000000048000000000000004c000000000000007800000000",
            INIT_18 => X"0000006600000000000000b800000000000000b0000000000000002600000000",
            INIT_19 => X"0000005900000000000000660000000000000038000000000000007300000000",
            INIT_1A => X"0000006500000000000000330000000000000051000000000000004e00000000",
            INIT_1B => X"0000000e000000000000002b000000000000002c000000000000004100000000",
            INIT_1C => X"00000075000000000000008600000000000000b300000000000000c000000000",
            INIT_1D => X"00000079000000000000005f0000000000000033000000000000006f00000000",
            INIT_1E => X"000000250000000000000040000000000000005a000000000000004200000000",
            INIT_1F => X"000000c700000000000000270000000000000027000000000000002f00000000",
            INIT_20 => X"0000009e00000000000000a2000000000000008b00000000000000ab00000000",
            INIT_21 => X"0000007900000000000000b90000000000000091000000000000006500000000",
            INIT_22 => X"0000005a00000000000000470000000000000040000000000000003c00000000",
            INIT_23 => X"000000cb00000000000000c10000000000000068000000000000007100000000",
            INIT_24 => X"000000a500000000000000e700000000000000c9000000000000009d00000000",
            INIT_25 => X"0000006f000000000000007c0000000000000085000000000000008a00000000",
            INIT_26 => X"0000008a00000000000000880000000000000080000000000000007800000000",
            INIT_27 => X"000000b100000000000000a1000000000000008c000000000000008e00000000",
            INIT_28 => X"00000075000000000000007a00000000000000af00000000000000e500000000",
            INIT_29 => X"0000008400000000000000760000000000000071000000000000007000000000",
            INIT_2A => X"000000a3000000000000009a0000000000000095000000000000008c00000000",
            INIT_2B => X"000000ef00000000000000a60000000000000085000000000000009d00000000",
            INIT_2C => X"0000007300000000000000790000000000000080000000000000008800000000",
            INIT_2D => X"0000009b000000000000008c0000000000000082000000000000007700000000",
            INIT_2E => X"0000009700000000000000ab00000000000000a3000000000000009300000000",
            INIT_2F => X"0000007400000000000000a7000000000000007f000000000000008f00000000",
            INIT_30 => X"0000007c000000000000007e0000000000000089000000000000007f00000000",
            INIT_31 => X"0000009a00000000000000850000000000000086000000000000008800000000",
            INIT_32 => X"000000000000000000000000000000000000008d00000000000000af00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000000b000000000000001c00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000033000000000000001400000000",
            INIT_39 => X"000000000000000000000000000000000000001e000000000000001400000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_3B => X"00000028000000000000001c000000000000003e000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"000000190000000000000000000000000000001e000000000000000700000000",
            INIT_3E => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000006000000000000001a0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_43 => X"00000000000000000000001d0000000000000004000000000000000f00000000",
            INIT_44 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_45 => X"000000020000000000000000000000000000002f000000000000002500000000",
            INIT_46 => X"0000000000000000000000000000000000000003000000000000004f00000000",
            INIT_47 => X"0000002600000000000000000000000000000006000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_49 => X"0000000d000000000000000d0000000000000018000000000000000000000000",
            INIT_4A => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_4B => X"0000000800000000000000180000000000000000000000000000000900000000",
            INIT_4C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_4E => X"00000000000000000000001e000000000000003d000000000000000000000000",
            INIT_4F => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_51 => X"0000003200000000000000220000000000000000000000000000002e00000000",
            INIT_52 => X"0000003600000000000000000000000000000000000000000000000300000000",
            INIT_53 => X"00000000000000000000000d000000000000003a000000000000002600000000",
            INIT_54 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000150000000000000012000000000000000000000000",
            INIT_56 => X"00000031000000000000001f000000000000002e000000000000000000000000",
            INIT_57 => X"0000000800000000000000000000000000000000000000000000000100000000",
            INIT_58 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_59 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"000000000000000000000000000000000000000d000000000000000f00000000",
            INIT_5B => X"0000004100000000000000210000000000000016000000000000000000000000",
            INIT_5C => X"000000a200000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000c0000000000000037000000000000003f000000000000005200000000",
            INIT_5E => X"0000000000000000000000020000000000000000000000000000000600000000",
            INIT_5F => X"00000036000000000000000d0000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000560000000000000041000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_62 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_63 => X"0000002500000000000000000000000000000002000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000006000000000000003e00000000",
            INIT_65 => X"0000000700000000000000000000000000000000000000000000000100000000",
            INIT_66 => X"0000004200000000000000000000000000000000000000000000000a00000000",
            INIT_67 => X"0000003600000000000000180000000000000000000000000000000c00000000",
            INIT_68 => X"0000000000000000000000090000000000000013000000000000002400000000",
            INIT_69 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000000000000000000001f0000000000000004000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"000000070000000000000000000000000000002d000000000000000500000000",
            INIT_79 => X"0000000000000000000000010000000000000002000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_7B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000300000000000000000000000000000000000000000000003b00000000",
            INIT_7D => X"0000000600000000000000010000000000000010000000000000000000000000",
            INIT_7E => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_7F => X"0000005d00000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE4;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5 : if BRAM_NAME = "samplegold_layersamples_instance5" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000000000000000000000f000000000000001c000000000000000000000000",
            INIT_03 => X"0000000000000000000000520000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000130000000000000012000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_06 => X"0000000500000000000000000000000000000017000000000000000c00000000",
            INIT_07 => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000003000000000000001d00000000",
            INIT_09 => X"0000000000000000000000110000000000000000000000000000001600000000",
            INIT_0A => X"0000000800000000000000000000000000000000000000000000001200000000",
            INIT_0B => X"0000001b00000000000000000000000000000011000000000000000000000000",
            INIT_0C => X"0000001900000000000000090000000000000000000000000000000000000000",
            INIT_0D => X"000000030000000000000000000000000000003b000000000000000000000000",
            INIT_0E => X"0000000000000000000000050000000000000000000000000000001000000000",
            INIT_0F => X"0000000000000000000000120000000000000012000000000000000000000000",
            INIT_10 => X"00000000000000000000000d0000000000000033000000000000000000000000",
            INIT_11 => X"0000002d00000000000000000000000000000000000000000000005800000000",
            INIT_12 => X"0000002800000000000000020000000000000000000000000000000400000000",
            INIT_13 => X"0000001d000000000000002c000000000000003e000000000000003300000000",
            INIT_14 => X"0000003b00000000000000000000000000000036000000000000007000000000",
            INIT_15 => X"0000004e000000000000004e000000000000002e000000000000000000000000",
            INIT_16 => X"00000056000000000000004f0000000000000049000000000000004400000000",
            INIT_17 => X"0000005a0000000000000053000000000000005a000000000000005800000000",
            INIT_18 => X"0000000000000000000000080000000000000048000000000000006f00000000",
            INIT_19 => X"0000004c000000000000004a0000000000000048000000000000004900000000",
            INIT_1A => X"00000057000000000000005b000000000000005b000000000000005400000000",
            INIT_1B => X"00000060000000000000005a000000000000005e000000000000005d00000000",
            INIT_1C => X"0000005000000000000000310000000000000000000000000000008a00000000",
            INIT_1D => X"000000570000000000000053000000000000004d000000000000004500000000",
            INIT_1E => X"0000007400000000000000610000000000000064000000000000006100000000",
            INIT_1F => X"0000006700000000000000670000000000000050000000000000005e00000000",
            INIT_20 => X"00000055000000000000005f0000000000000049000000000000004100000000",
            INIT_21 => X"0000005200000000000000520000000000000052000000000000004900000000",
            INIT_22 => X"000000450000000000000053000000000000006b000000000000005e00000000",
            INIT_23 => X"0000002e0000000000000033000000000000002e000000000000002f00000000",
            INIT_24 => X"0000002f0000000000000031000000000000002f000000000000002f00000000",
            INIT_25 => X"00000027000000000000001c0000000000000023000000000000002b00000000",
            INIT_26 => X"0000003200000000000000240000000000000027000000000000002600000000",
            INIT_27 => X"00000034000000000000002d0000000000000035000000000000003200000000",
            INIT_28 => X"0000000400000000000000250000000000000013000000000000005500000000",
            INIT_29 => X"0000002400000000000000150000000000000013000000000000002100000000",
            INIT_2A => X"0000003b000000000000001a0000000000000028000000000000002d00000000",
            INIT_2B => X"0000002c0000000000000038000000000000002e000000000000003400000000",
            INIT_2C => X"0000004f000000000000001a0000000000000000000000000000000000000000",
            INIT_2D => X"000000270000000000000004000000000000000b000000000000000a00000000",
            INIT_2E => X"0000002c00000000000000790000000000000000000000000000003900000000",
            INIT_2F => X"0000001a00000000000000230000000000000025000000000000003600000000",
            INIT_30 => X"0000000000000000000000530000000000000018000000000000000800000000",
            INIT_31 => X"00000053000000000000000e0000000000000000000000000000001200000000",
            INIT_32 => X"00000049000000000000000a0000000000000063000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000001a000000000000002c00000000",
            INIT_34 => X"00000000000000000000000b000000000000005f000000000000000800000000",
            INIT_35 => X"0000000000000000000000390000000000000000000000000000001e00000000",
            INIT_36 => X"00000049000000000000002e0000000000000000000000000000003800000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000230000000000000000000000000000000000000000000000bf00000000",
            INIT_39 => X"000000150000000000000000000000000000000d000000000000000400000000",
            INIT_3A => X"0000005000000000000000610000000000000000000000000000000c00000000",
            INIT_3B => X"000000a400000000000000000000000000000000000000000000000a00000000",
            INIT_3C => X"00000027000000000000001e0000000000000000000000000000000000000000",
            INIT_3D => X"0000000100000000000000000000000000000000000000000000000d00000000",
            INIT_3E => X"0000000000000000000000680000000000000045000000000000000000000000",
            INIT_3F => X"00000000000000000000007c0000000000000000000000000000000800000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000120000000000000022000000000000002a000000000000000000000000",
            INIT_41 => X"0000003c00000000000000000000000000000017000000000000000000000000",
            INIT_42 => X"0000001c00000000000000000000000000000003000000000000001100000000",
            INIT_43 => X"0000000000000000000000220000000000000006000000000000003100000000",
            INIT_44 => X"0000000a0000000000000044000000000000003a000000000000002600000000",
            INIT_45 => X"00000000000000000000004a0000000000000000000000000000001800000000",
            INIT_46 => X"00000017000000000000000e000000000000002a000000000000001900000000",
            INIT_47 => X"0000004800000000000000050000000000000000000000000000000a00000000",
            INIT_48 => X"000000110000000000000051000000000000001c000000000000005600000000",
            INIT_49 => X"0000000b000000000000000000000000000000a3000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000005600000000",
            INIT_4B => X"0000001e000000000000002d0000000000000028000000000000001400000000",
            INIT_4C => X"0000000000000000000000280000000000000040000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000009800000000",
            INIT_4E => X"0000001000000000000000090000000000000000000000000000000000000000",
            INIT_4F => X"000000000000000000000011000000000000000e000000000000001000000000",
            INIT_50 => X"0000001f00000000000000480000000000000041000000000000000300000000",
            INIT_51 => X"0000000a00000000000000050000000000000009000000000000000000000000",
            INIT_52 => X"0000001700000000000000140000000000000010000000000000000800000000",
            INIT_53 => X"0000000000000000000000170000000000000008000000000000001000000000",
            INIT_54 => X"0000000000000000000000000000000000000074000000000000001000000000",
            INIT_55 => X"0000000d00000000000000090000000000000000000000000000001100000000",
            INIT_56 => X"000000000000000000000009000000000000000d000000000000001000000000",
            INIT_57 => X"0000000d00000000000000000000000000000000000000000000002600000000",
            INIT_58 => X"0000001600000000000000000000000000000000000000000000001900000000",
            INIT_59 => X"0000001000000000000000180000000000000009000000000000000c00000000",
            INIT_5A => X"000000030000000000000031000000000000000b000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_61 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000001200000000000000040000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000270000000000000001000000000000000000000000",
            INIT_6B => X"0000000000000000000000080000000000000038000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000014000000000000000000000000",
            INIT_71 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE5;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6 : if BRAM_NAME = "samplegold_layersamples_instance6" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_01 => X"00000030000000000000001e0000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_03 => X"000000010000000000000024000000000000001c000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000036000000000000002f0000000000000000000000000000000000000000",
            INIT_14 => X"0000003000000000000000350000000000000035000000000000003300000000",
            INIT_15 => X"0000002b0000000000000036000000000000003b000000000000003900000000",
            INIT_16 => X"0000002800000000000000250000000000000020000000000000002000000000",
            INIT_17 => X"0000003600000000000000380000000000000030000000000000002700000000",
            INIT_18 => X"0000003b00000000000000420000000000000033000000000000003900000000",
            INIT_19 => X"0000000200000000000000020000000000000023000000000000003900000000",
            INIT_1A => X"0000002700000000000000110000000000000006000000000000000600000000",
            INIT_1B => X"0000003900000000000000360000000000000013000000000000003000000000",
            INIT_1C => X"00000000000000000000001e000000000000003d000000000000003700000000",
            INIT_1D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_1E => X"0000001500000000000000170000000000000000000000000000000100000000",
            INIT_1F => X"0000004000000000000000370000000000000032000000000000000000000000",
            INIT_20 => X"000000000000000000000000000000000000001e000000000000001200000000",
            INIT_21 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_22 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000003300000000000000440000000000000010000000000000003400000000",
            INIT_24 => X"0000000000000000000000000000000000000006000000000000002500000000",
            INIT_25 => X"0000000000000000000000000000000000000009000000000000001000000000",
            INIT_26 => X"00000031000000000000000f0000000000000000000000000000000000000000",
            INIT_27 => X"0000002b000000000000000d000000000000000b000000000000003800000000",
            INIT_28 => X"0000002a0000000000000000000000000000000b000000000000000800000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000003d0000000000000007000000000000002c000000000000000000000000",
            INIT_2B => X"00000017000000000000002e0000000000000011000000000000000e00000000",
            INIT_2C => X"0000000000000000000000130000000000000003000000000000000800000000",
            INIT_2D => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000250000000000000000000000000000001900000000",
            INIT_2F => X"00000000000000000000000a000000000000002e000000000000002200000000",
            INIT_30 => X"000000000000000000000000000000000000000f000000000000001300000000",
            INIT_31 => X"0000001100000000000000150000000000000000000000000000000200000000",
            INIT_32 => X"00000000000000000000001c0000000000000000000000000000000900000000",
            INIT_33 => X"0000002c0000000000000000000000000000000c000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"00000014000000000000000e0000000000000016000000000000002100000000",
            INIT_36 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_37 => X"0000000000000000000000050000000000000006000000000000001f00000000",
            INIT_38 => X"00000028000000000000001e0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000150000000000000014000000000000000500000000",
            INIT_3A => X"0000001700000000000000110000000000000006000000000000002c00000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000003c00000000000000320000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000002800000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000002c00000000000000290000000000000023000000000000002200000000",
            INIT_4D => X"0000002f000000000000002b0000000000000028000000000000002000000000",
            INIT_4E => X"0000001e000000000000001d0000000000000029000000000000003200000000",
            INIT_4F => X"000000240000000000000028000000000000002e000000000000002900000000",
            INIT_50 => X"0000000e0000000000000021000000000000002c000000000000002400000000",
            INIT_51 => X"00000005000000000000002e0000000000000030000000000000004300000000",
            INIT_52 => X"0000001500000000000000190000000000000029000000000000002100000000",
            INIT_53 => X"000000280000000000000002000000000000003f000000000000002c00000000",
            INIT_54 => X"000000280000000000000020000000000000002a000000000000002900000000",
            INIT_55 => X"0000001c00000000000000000000000000000010000000000000002400000000",
            INIT_56 => X"0000000b000000000000001a0000000000000032000000000000000c00000000",
            INIT_57 => X"00000024000000000000002e0000000000000000000000000000005c00000000",
            INIT_58 => X"000000250000000000000027000000000000000c000000000000003800000000",
            INIT_59 => X"0000001800000000000000230000000000000000000000000000001900000000",
            INIT_5A => X"0000002c00000000000000000000000000000026000000000000001a00000000",
            INIT_5B => X"0000001300000000000000000000000000000041000000000000000500000000",
            INIT_5C => X"000000250000000000000024000000000000002a000000000000002700000000",
            INIT_5D => X"0000001200000000000000380000000000000014000000000000000000000000",
            INIT_5E => X"000000000000000000000024000000000000001a000000000000002b00000000",
            INIT_5F => X"000000000000000000000000000000000000002f000000000000003700000000",
            INIT_60 => X"0000000000000000000000430000000000000025000000000000001600000000",
            INIT_61 => X"0000001d0000000000000007000000000000002a000000000000003400000000",
            INIT_62 => X"0000000e00000000000000240000000000000011000000000000002000000000",
            INIT_63 => X"0000001500000000000000000000000000000000000000000000004600000000",
            INIT_64 => X"0000002b00000000000000000000000000000039000000000000001c00000000",
            INIT_65 => X"000000250000000000000000000000000000000d000000000000002800000000",
            INIT_66 => X"0000003400000000000000290000000000000006000000000000000b00000000",
            INIT_67 => X"0000000b00000000000000350000000000000000000000000000000200000000",
            INIT_68 => X"0000002c00000000000000110000000000000000000000000000001800000000",
            INIT_69 => X"0000000d000000000000000d0000000000000011000000000000000000000000",
            INIT_6A => X"000000340000000000000000000000000000003f000000000000000000000000",
            INIT_6B => X"00000000000000000000001b000000000000000e000000000000000000000000",
            INIT_6C => X"00000000000000000000002b0000000000000005000000000000003f00000000",
            INIT_6D => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_6E => X"00000014000000000000002a0000000000000000000000000000003900000000",
            INIT_6F => X"0000000f000000000000002c000000000000001d000000000000000000000000",
            INIT_70 => X"000000100000000000000000000000000000000f000000000000002f00000000",
            INIT_71 => X"0000003800000000000000000000000000000000000000000000002f00000000",
            INIT_72 => X"0000000000000000000000320000000000000029000000000000000000000000",
            INIT_73 => X"0000000f000000000000002b0000000000000027000000000000000500000000",
            INIT_74 => X"0000002100000000000000110000000000000008000000000000000800000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000005000000000000005200000000",
            INIT_77 => X"0000000000000000000000030000000000000007000000000000000000000000",
            INIT_78 => X"0000001400000000000000030000000000000000000000000000000000000000",
            INIT_79 => X"0000002e00000000000000220000000000000000000000000000000000000000",
            INIT_7A => X"0000000500000000000000020000000000000006000000000000000000000000",
            INIT_7B => X"0000000200000000000000000000000000000000000000000000000100000000",
            INIT_7C => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000000d0000000000000022000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000006000000000000000900000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE6;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7 : if BRAM_NAME = "samplegold_layersamples_instance7" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000013000000000000001500000000",
            INIT_01 => X"0000000000000000000000000000000000000014000000000000000400000000",
            INIT_02 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000001a00000000000000120000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_38 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000000000000000000002f000000000000003d000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000012000000000000001f000000000000001300000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000900000000000000130000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000004200000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"000000000000000000000000000000000000000d000000000000004500000000",
            INIT_54 => X"00000000000000000000000a000000000000001f000000000000000400000000",
            INIT_55 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000250000000000000010000000000000000e00000000",
            INIT_57 => X"0000000000000000000000000000000000000009000000000000000900000000",
            INIT_58 => X"0000001700000000000000190000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"000000200000000000000027000000000000000e000000000000000000000000",
            INIT_5E => X"0000003e00000000000000400000000000000037000000000000001b00000000",
            INIT_5F => X"00000021000000000000002a0000000000000031000000000000003a00000000",
            INIT_60 => X"0000002100000000000000260000000000000014000000000000001c00000000",
            INIT_61 => X"00000037000000000000000b000000000000000a000000000000001200000000",
            INIT_62 => X"00000050000000000000004b000000000000003f000000000000004100000000",
            INIT_63 => X"00000042000000000000004c0000000000000056000000000000005500000000",
            INIT_64 => X"0000001e00000000000000290000000000000032000000000000003e00000000",
            INIT_65 => X"0000000a00000000000000020000000000000000000000000000000000000000",
            INIT_66 => X"0000000b00000000000000030000000000000000000000000000000000000000",
            INIT_67 => X"0000000200000000000000080000000000000000000000000000000100000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000001800000000000000100000000000000000000000000000000000000000",
            INIT_6A => X"0000002200000000000000060000000000000006000000000000000a00000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_6D => X"0000000400000000000000060000000000000003000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000004000000000000000400000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000002b000000000000002b0000000000000000000000000000000000000000",
            INIT_75 => X"0000002b000000000000002c000000000000002b000000000000002b00000000",
            INIT_76 => X"0000002c000000000000002b000000000000002b000000000000002b00000000",
            INIT_77 => X"0000002b000000000000002b000000000000002a000000000000002d00000000",
            INIT_78 => X"0000002b000000000000002b000000000000002b000000000000002c00000000",
            INIT_79 => X"0000002c000000000000002b000000000000002b000000000000002b00000000",
            INIT_7A => X"00000028000000000000001c000000000000002b000000000000002900000000",
            INIT_7B => X"0000002c000000000000002b000000000000002c000000000000003100000000",
            INIT_7C => X"0000002b000000000000002b000000000000002b000000000000002900000000",
            INIT_7D => X"00000023000000000000002b000000000000002c000000000000002d00000000",
            INIT_7E => X"0000002b000000000000002c000000000000001a000000000000001c00000000",
            INIT_7F => X"00000032000000000000002c000000000000002b000000000000002b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE7;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8 : if BRAM_NAME = "samplegold_layersamples_instance8" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002c000000000000002b000000000000002c000000000000002d00000000",
            INIT_01 => X"0000002c0000000000000020000000000000002f000000000000001f00000000",
            INIT_02 => X"0000002b00000000000000460000000000000033000000000000002d00000000",
            INIT_03 => X"000000220000000000000019000000000000002b000000000000002b00000000",
            INIT_04 => X"00000020000000000000002c0000000000000029000000000000002e00000000",
            INIT_05 => X"0000003100000000000000330000000000000029000000000000003200000000",
            INIT_06 => X"0000002900000000000000170000000000000014000000000000002000000000",
            INIT_07 => X"0000002f00000000000000380000000000000032000000000000002b00000000",
            INIT_08 => X"0000001300000000000000120000000000000025000000000000002100000000",
            INIT_09 => X"0000002b000000000000001e000000000000001d000000000000001700000000",
            INIT_0A => X"0000002e000000000000004b0000000000000026000000000000003200000000",
            INIT_0B => X"000000270000000000000029000000000000001f000000000000001600000000",
            INIT_0C => X"0000003b00000000000000210000000000000005000000000000001b00000000",
            INIT_0D => X"000000150000000000000020000000000000002d000000000000005500000000",
            INIT_0E => X"0000001e00000000000000260000000000000014000000000000001900000000",
            INIT_0F => X"0000002700000000000000340000000000000015000000000000003b00000000",
            INIT_10 => X"0000001900000000000000210000000000000043000000000000002e00000000",
            INIT_11 => X"0000002f000000000000002a0000000000000020000000000000001c00000000",
            INIT_12 => X"0000002a000000000000006b000000000000003b000000000000003500000000",
            INIT_13 => X"0000002300000000000000320000000000000037000000000000003000000000",
            INIT_14 => X"0000002300000000000000270000000000000017000000000000002800000000",
            INIT_15 => X"000000140000000000000018000000000000001e000000000000002500000000",
            INIT_16 => X"00000025000000000000001d000000000000002e000000000000001900000000",
            INIT_17 => X"00000027000000000000002b0000000000000029000000000000002700000000",
            INIT_18 => X"0000002800000000000000280000000000000030000000000000002c00000000",
            INIT_19 => X"0000002400000000000000240000000000000029000000000000001f00000000",
            INIT_1A => X"00000017000000000000001a0000000000000017000000000000000c00000000",
            INIT_1B => X"0000002200000000000000210000000000000019000000000000001400000000",
            INIT_1C => X"00000023000000000000001f000000000000001c000000000000001d00000000",
            INIT_1D => X"000000000000000000000025000000000000002c000000000000002900000000",
            INIT_1E => X"0000000000000000000000000000000000000001000000000000001200000000",
            INIT_1F => X"0000002d000000000000002f000000000000002b000000000000000d00000000",
            INIT_20 => X"00000021000000000000003c0000000000000036000000000000003100000000",
            INIT_21 => X"0000000000000000000000000000000000000024000000000000001800000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_23 => X"0000002000000000000000260000000000000021000000000000003f00000000",
            INIT_24 => X"00000019000000000000001f000000000000000e000000000000000e00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_26 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000001500000000000000070000000000000012000000000000002700000000",
            INIT_28 => X"00000023000000000000001a000000000000000d000000000000001700000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000600000000000000030000000000000000000000000000000000000000",
            INIT_2B => X"00000008000000000000000d0000000000000015000000000000000a00000000",
            INIT_2C => X"000000520000000000000024000000000000001a000000000000001100000000",
            INIT_2D => X"0000004e000000000000004f000000000000004f000000000000004f00000000",
            INIT_2E => X"0000004d0000000000000051000000000000004f000000000000004f00000000",
            INIT_2F => X"0000004f000000000000004f0000000000000051000000000000005200000000",
            INIT_30 => X"0000004f0000000000000052000000000000004e000000000000004f00000000",
            INIT_31 => X"0000004f000000000000004e0000000000000050000000000000004f00000000",
            INIT_32 => X"000000800000000000000054000000000000004f000000000000004d00000000",
            INIT_33 => X"0000004e0000000000000050000000000000003a000000000000003100000000",
            INIT_34 => X"0000004e000000000000004e0000000000000051000000000000004e00000000",
            INIT_35 => X"0000004a0000000000000056000000000000004c000000000000004f00000000",
            INIT_36 => X"0000003100000000000000710000000000000064000000000000006f00000000",
            INIT_37 => X"0000004f000000000000004e0000000000000051000000000000002700000000",
            INIT_38 => X"0000004e000000000000004c0000000000000051000000000000004500000000",
            INIT_39 => X"0000006f000000000000002a0000000000000079000000000000005000000000",
            INIT_3A => X"0000001100000000000000370000000000000050000000000000004300000000",
            INIT_3B => X"0000003f000000000000004e000000000000004f000000000000005200000000",
            INIT_3C => X"0000004f000000000000004b0000000000000021000000000000002200000000",
            INIT_3D => X"0000004800000000000000570000000000000035000000000000006400000000",
            INIT_3E => X"0000005b0000000000000068000000000000007a000000000000006a00000000",
            INIT_3F => X"0000003400000000000000490000000000000048000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007f00000000000000540000000000000054000000000000004b00000000",
            INIT_41 => X"00000064000000000000003e0000000000000058000000000000005e00000000",
            INIT_42 => X"0000000000000000000000600000000000000043000000000000004b00000000",
            INIT_43 => X"0000003a000000000000001c0000000000000051000000000000004400000000",
            INIT_44 => X"000000030000000000000080000000000000007c000000000000002900000000",
            INIT_45 => X"0000007400000000000000620000000000000000000000000000000000000000",
            INIT_46 => X"000000250000000000000066000000000000005f000000000000007400000000",
            INIT_47 => X"0000000000000000000000370000000000000014000000000000000000000000",
            INIT_48 => X"000000760000000000000028000000000000004c000000000000003900000000",
            INIT_49 => X"0000002700000000000000400000000000000048000000000000005000000000",
            INIT_4A => X"00000000000000000000002a0000000000000023000000000000001600000000",
            INIT_4B => X"0000004d00000000000000400000000000000045000000000000005d00000000",
            INIT_4C => X"0000005900000000000000850000000000000061000000000000006d00000000",
            INIT_4D => X"00000062000000000000007c0000000000000064000000000000006900000000",
            INIT_4E => X"0000005e00000000000000200000000000000049000000000000005500000000",
            INIT_4F => X"000000540000000000000055000000000000005a000000000000005500000000",
            INIT_50 => X"0000005b000000000000004c000000000000004d000000000000006100000000",
            INIT_51 => X"00000037000000000000003c0000000000000053000000000000004d00000000",
            INIT_52 => X"00000038000000000000000f000000000000002b000000000000002800000000",
            INIT_53 => X"0000004a000000000000002e0000000000000030000000000000003400000000",
            INIT_54 => X"0000004500000000000000540000000000000054000000000000004e00000000",
            INIT_55 => X"0000001c000000000000002b0000000000000018000000000000003300000000",
            INIT_56 => X"00000037000000000000003a0000000000000000000000000000002e00000000",
            INIT_57 => X"0000002c00000000000000000000000000000002000000000000001d00000000",
            INIT_58 => X"0000001d0000000000000000000000000000000f000000000000001700000000",
            INIT_59 => X"000000370000000000000006000000000000002c000000000000003a00000000",
            INIT_5A => X"000000120000000000000023000000000000000a000000000000000000000000",
            INIT_5B => X"0000004400000000000000460000000000000000000000000000000800000000",
            INIT_5C => X"0000000d000000000000001b0000000000000049000000000000005200000000",
            INIT_5D => X"0000000900000000000000750000000000000006000000000000000c00000000",
            INIT_5E => X"000000070000000000000009000000000000000f000000000000000600000000",
            INIT_5F => X"00000006000000000000003d0000000000000022000000000000000000000000",
            INIT_60 => X"0000000b000000000000001c0000000000000001000000000000000000000000",
            INIT_61 => X"00000004000000000000000a0000000000000062000000000000001000000000",
            INIT_62 => X"0000000000000000000000000000000000000002000000000000000500000000",
            INIT_63 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000001500000000000000130000000000000013000000000000001d00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000004a000000000000003a0000000000000028000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000500000000000000190000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000008000000000000001700000000",
            INIT_77 => X"0000007600000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000017000000000000007c00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000062000000000000005f0000000000000032000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000005600000000",
            INIT_7C => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_7D => X"00000000000000000000004e0000000000000023000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000720000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE8;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9 : if BRAM_NAME = "samplegold_layersamples_instance9" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000a300000000000000790000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_02 => X"0000003d00000000000000440000000000000028000000000000001300000000",
            INIT_03 => X"0000004e00000000000000660000000000000024000000000000006f00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000001900000000000000000000000000000000000000000000000900000000",
            INIT_0F => X"0000004d00000000000000000000000000000004000000000000002000000000",
            INIT_10 => X"0000006300000000000000550000000000000053000000000000008e00000000",
            INIT_11 => X"0000001c0000000000000000000000000000001d000000000000007000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000019000000000000001e000000000000001c000000000000001900000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000500000000000000440000000000000042000000000000000000000000",
            INIT_19 => X"0000002200000000000000000000000000000003000000000000000a00000000",
            INIT_1A => X"0000001900000000000000160000000000000014000000000000001d00000000",
            INIT_1B => X"0000005000000000000000490000000000000000000000000000000c00000000",
            INIT_1C => X"00000010000000000000000b0000000000000000000000000000001d00000000",
            INIT_1D => X"0000001500000000000000150000000000000017000000000000000e00000000",
            INIT_1E => X"0000001500000000000000150000000000000015000000000000001500000000",
            INIT_1F => X"0000001000000000000000160000000000000017000000000000001800000000",
            INIT_20 => X"0000001500000000000000150000000000000016000000000000001500000000",
            INIT_21 => X"0000001600000000000000160000000000000016000000000000001700000000",
            INIT_22 => X"0000001700000000000000150000000000000016000000000000001500000000",
            INIT_23 => X"0000000e00000000000000000000000000000021000000000000001a00000000",
            INIT_24 => X"0000001500000000000000160000000000000016000000000000001600000000",
            INIT_25 => X"0000001600000000000000170000000000000015000000000000001600000000",
            INIT_26 => X"00000007000000000000001f000000000000000f000000000000001900000000",
            INIT_27 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000c00000000000000070000000000000015000000000000001600000000",
            INIT_29 => X"0000002700000000000000180000000000000018000000000000001200000000",
            INIT_2A => X"0000000000000000000000000000000000000013000000000000000700000000",
            INIT_2B => X"0000000f000000000000000c0000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_2D => X"0000001100000000000000120000000000000016000000000000001700000000",
            INIT_2E => X"00000001000000000000000a0000000000000008000000000000001100000000",
            INIT_2F => X"0000000900000000000000000000000000000002000000000000000000000000",
            INIT_30 => X"0000001f000000000000000b0000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000019000000000000001100000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_34 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_36 => X"000000000000000000000008000000000000000c000000000000001000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000002000000000000000100000000",
            INIT_39 => X"0000000000000000000000020000000000000014000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000100000000000000050000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000040000000000000007000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_4A => X"00000015000000000000000a0000000000000022000000000000000000000000",
            INIT_4B => X"000000000000000000000009000000000000000a000000000000001600000000",
            INIT_4C => X"0000004400000000000000570000000000000059000000000000005200000000",
            INIT_4D => X"000000000000000000000008000000000000001d000000000000002000000000",
            INIT_4E => X"0000000c000000000000000d000000000000000b000000000000003000000000",
            INIT_4F => X"000000bc00000000000000320000000000000009000000000000000a00000000",
            INIT_50 => X"00000022000000000000002d000000000000004c00000000000000a700000000",
            INIT_51 => X"0000002100000000000000000000000000000007000000000000001300000000",
            INIT_52 => X"0000000b000000000000000a000000000000000d000000000000001400000000",
            INIT_53 => X"000000320000000000000041000000000000001b000000000000000700000000",
            INIT_54 => X"0000000c00000000000000140000000000000027000000000000002800000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000001400000000000000110000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_63 => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_64 => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_67 => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_6B => X"0000000000000000000000310000000000000000000000000000000000000000",
            INIT_6C => X"000000090000000000000012000000000000001b000000000000000000000000",
            INIT_6D => X"0000002000000000000000080000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000003e00000000",
            INIT_6F => X"0000003600000000000000160000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000340000000000000000000000000000001500000000",
            INIT_71 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_72 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000a2000000000000000d000000000000000600000000",
            INIT_74 => X"000000000000000000000001000000000000000c000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000021000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000a00000000000000030000000000000000000000000000000000000000",
            INIT_7B => X"0000000b00000000000000050000000000000013000000000000000000000000",
            INIT_7C => X"0000000700000000000000060000000000000012000000000000001000000000",
            INIT_7D => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"000000000000000000000012000000000000000a000000000000001300000000",
            INIT_7F => X"0000000600000000000000000000000000000000000000000000003500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE9;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10 : if BRAM_NAME = "samplegold_layersamples_instance10" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000038000000000000001f00000000",
            INIT_01 => X"0000000d000000000000001c000000000000001d000000000000000d00000000",
            INIT_02 => X"0000001b0000000000000000000000000000001e000000000000000500000000",
            INIT_03 => X"00000013000000000000000c0000000000000009000000000000002000000000",
            INIT_04 => X"0000002100000000000000320000000000000039000000000000009d00000000",
            INIT_05 => X"000000160000000000000023000000000000001b000000000000001300000000",
            INIT_06 => X"0000001600000000000000100000000000000000000000000000001a00000000",
            INIT_07 => X"0000006c00000000000000120000000000000012000000000000001100000000",
            INIT_08 => X"0000003700000000000000430000000000000057000000000000008100000000",
            INIT_09 => X"0000001100000000000000140000000000000005000000000000002600000000",
            INIT_0A => X"0000000900000000000000090000000000000003000000000000000000000000",
            INIT_0B => X"0000003f0000000000000028000000000000000f000000000000000f00000000",
            INIT_0C => X"00000000000000000000000c0000000000000035000000000000003b00000000",
            INIT_0D => X"00000000000000000000000c000000000000000b000000000000000c00000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000001b000000000000001a000000000000001e000000000000000000000000",
            INIT_34 => X"0000000f00000000000000250000000000000026000000000000002300000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000100000000000000000000000000000000000000000000001300000000",
            INIT_38 => X"0000000000000000000000000000000000000014000000000000001200000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000001d000000000000002e0000000000000030000000000000001700000000",
            INIT_3C => X"000000390000000000000043000000000000000e000000000000001a00000000",
            INIT_3D => X"0000000000000000000000320000000000000040000000000000003800000000",
            INIT_3E => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000019000000000000001a000000000000001e000000000000001c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000005900000000000000a50000000000000099000000000000001f00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000900000000000000070000000000000001000000000000000000000000",
            INIT_43 => X"0000000b000000000000000c000000000000000e000000000000000a00000000",
            INIT_44 => X"000000000000000000000000000000000000000a000000000000004500000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000100000000000000010000000000000001000000000000000200000000",
            INIT_47 => X"0000000200000000000000020000000000000003000000000000000200000000",
            INIT_48 => X"0000000200000000000000040000000000000003000000000000000100000000",
            INIT_49 => X"0000000200000000000000010000000000000001000000000000000200000000",
            INIT_4A => X"0000000100000000000000010000000000000001000000000000000100000000",
            INIT_4B => X"0000000200000000000000000000000000000001000000000000000000000000",
            INIT_4C => X"000000000000000000000000000000000000000e000000000000001c00000000",
            INIT_4D => X"00000007000000000000000a0000000000000000000000000000000000000000",
            INIT_4E => X"0000000400000000000000000000000000000000000000000000000100000000",
            INIT_4F => X"00000024000000000000002a0000000000000011000000000000000600000000",
            INIT_50 => X"0000000100000000000000010000000000000016000000000000002500000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_52 => X"0000000200000000000000080000000000000002000000000000000200000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000009000000000000000c0000000000000031000000000000002a00000000",
            INIT_56 => X"0000000200000000000000000000000000000001000000000000000400000000",
            INIT_57 => X"000000400000000000000039000000000000000c000000000000000000000000",
            INIT_58 => X"000000000000000000000000000000000000002a000000000000004300000000",
            INIT_59 => X"00000028000000000000002d0000000000000000000000000000000000000000",
            INIT_5A => X"0000004700000000000000780000000000000089000000000000008200000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000044000000000000004d0000000000000001000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000002000000000000003400000000",
            INIT_5E => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000005200000000000000690000000000000066000000000000005500000000",
            INIT_60 => X"0000000000000000000000000000000000000008000000000000003900000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"000000000000000000000000000000000000001c000000000000000400000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_65 => X"0000004b00000000000000380000000000000024000000000000001a00000000",
            INIT_66 => X"0000004f00000000000000410000000000000047000000000000002000000000",
            INIT_67 => X"0000003c000000000000001c000000000000003f000000000000005600000000",
            INIT_68 => X"000000350000000000000048000000000000004a000000000000005b00000000",
            INIT_69 => X"0000000800000000000000000000000000000012000000000000002700000000",
            INIT_6A => X"0000000500000000000000120000000000000011000000000000000500000000",
            INIT_6B => X"00000000000000000000000a0000000000000000000000000000000d00000000",
            INIT_6C => X"0000005600000000000000470000000000000032000000000000001800000000",
            INIT_6D => X"00000040000000000000004c000000000000005e000000000000005f00000000",
            INIT_6E => X"0000000000000000000000000000000000000011000000000000002b00000000",
            INIT_6F => X"0000000800000000000000130000000000000012000000000000000000000000",
            INIT_70 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000010000000000000017000000000000000000000000",
            INIT_73 => X"00000017000000000000001c0000000000000000000000000000000000000000",
            INIT_74 => X"0000005d00000000000000240000000000000000000000000000000300000000",
            INIT_75 => X"0000001a00000000000000570000000000000059000000000000004d00000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_78 => X"0000007800000000000000600000000000000005000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_7A => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"000000ef00000000000000ef00000000000000ef000000000000000000000000",
            INIT_7F => X"000000f000000000000000f000000000000000ef00000000000000ef00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE10;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11 : if BRAM_NAME = "samplegold_layersamples_instance11" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000f300000000000000f100000000000000ed00000000000000ef00000000",
            INIT_01 => X"000000f000000000000000ef00000000000000f000000000000000ef00000000",
            INIT_02 => X"000000f000000000000000f000000000000000f000000000000000f100000000",
            INIT_03 => X"000000ef00000000000000f000000000000000f000000000000000f000000000",
            INIT_04 => X"000000f100000000000000ee00000000000000e900000000000000ef00000000",
            INIT_05 => X"000000f100000000000000f100000000000000f000000000000000ef00000000",
            INIT_06 => X"000000f000000000000000f100000000000000f000000000000000f000000000",
            INIT_07 => X"000000ec00000000000000ed00000000000000f200000000000000f000000000",
            INIT_08 => X"000000f200000000000000f300000000000000cf00000000000000de00000000",
            INIT_09 => X"000000f500000000000000f700000000000000f300000000000000f200000000",
            INIT_0A => X"000000eb00000000000000f200000000000000f200000000000000f600000000",
            INIT_0B => X"000000c400000000000000cd00000000000000e500000000000000eb00000000",
            INIT_0C => X"000000f800000000000000fa00000000000000d700000000000000b500000000",
            INIT_0D => X"000000fd00000000000000de00000000000000d200000000000000f800000000",
            INIT_0E => X"000000e000000000000000f200000000000000f100000000000000f000000000",
            INIT_0F => X"000000f000000000000000f300000000000000ea00000000000000f100000000",
            INIT_10 => X"000000fc00000000000000f300000000000000e000000000000000e900000000",
            INIT_11 => X"000000dc00000000000000d300000000000000ac00000000000000aa00000000",
            INIT_12 => X"000000f700000000000000f300000000000000e600000000000000ee00000000",
            INIT_13 => X"000000b900000000000000d200000000000000f500000000000000fc00000000",
            INIT_14 => X"000000bd00000000000000f700000000000000b700000000000000a200000000",
            INIT_15 => X"000000d300000000000000d000000000000000df00000000000000c900000000",
            INIT_16 => X"000000b60000000000000083000000000000006b000000000000007500000000",
            INIT_17 => X"000000e700000000000000e400000000000000ee00000000000000ec00000000",
            INIT_18 => X"00000075000000000000005600000000000000e900000000000000db00000000",
            INIT_19 => X"000000b100000000000000de00000000000000ad000000000000008200000000",
            INIT_1A => X"000000c200000000000000cf00000000000000be00000000000000a900000000",
            INIT_1B => X"000000a3000000000000008e000000000000008f00000000000000a000000000",
            INIT_1C => X"000000b100000000000000d1000000000000005000000000000000ae00000000",
            INIT_1D => X"000000ff00000000000000f400000000000000e400000000000000c000000000",
            INIT_1E => X"000000d400000000000000c600000000000000c100000000000000e900000000",
            INIT_1F => X"000000c200000000000000c700000000000000c600000000000000c900000000",
            INIT_20 => X"000000d500000000000000d100000000000000cb000000000000009200000000",
            INIT_21 => X"000000ae00000000000000c900000000000000d400000000000000d400000000",
            INIT_22 => X"0000008f000000000000009a000000000000009b00000000000000b400000000",
            INIT_23 => X"00000031000000000000008a000000000000007f000000000000008000000000",
            INIT_24 => X"0000005c0000000000000051000000000000004c000000000000004800000000",
            INIT_25 => X"0000008a000000000000008b000000000000008b000000000000007000000000",
            INIT_26 => X"0000006b0000000000000068000000000000006f000000000000007a00000000",
            INIT_27 => X"0000001700000000000000000000000000000075000000000000006800000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_29 => X"000000290000000000000027000000000000001a000000000000003000000000",
            INIT_2A => X"0000006b00000000000000560000000000000042000000000000002e00000000",
            INIT_2B => X"0000000500000000000000000000000000000000000000000000007900000000",
            INIT_2C => X"0000003a00000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000003b00000000000000290000000000000025000000000000004500000000",
            INIT_2E => X"00000097000000000000006a0000000000000053000000000000005100000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000003f000000000000001f000000000000000e000000000000000000000000",
            INIT_32 => X"0000001e00000000000000ad000000000000007f000000000000006700000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_35 => X"00000076000000000000006a000000000000004f000000000000002100000000",
            INIT_36 => X"00000000000000000000000000000000000000b3000000000000008c00000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000350000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000001e00000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000160000000000000017000000000000003500000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000004900000000000000730000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"000000000000000000000061000000000000004f000000000000003200000000",
            INIT_49 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000005400000000000000750000000000000017000000000000002f00000000",
            INIT_4B => X"0000000000000000000000000000000000000009000000000000003b00000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"00000000000000000000001f0000000000000057000000000000007b00000000",
            INIT_4E => X"0000000000000000000000000000000000000034000000000000000300000000",
            INIT_4F => X"00000051000000000000003a0000000000000012000000000000000000000000",
            INIT_50 => X"000000000000000000000018000000000000004c000000000000002700000000",
            INIT_51 => X"000000000000000000000007000000000000001f000000000000000000000000",
            INIT_52 => X"00000046000000000000002b0000000000000000000000000000000000000000",
            INIT_53 => X"000000000000000000000000000000000000000f000000000000002900000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000c00000000000000000000000000000000000000000000002500000000",
            INIT_57 => X"0000004c00000000000000330000000000000024000000000000000000000000",
            INIT_58 => X"000000590000000000000054000000000000002f000000000000002a00000000",
            INIT_59 => X"0000002f00000000000000310000000000000047000000000000005300000000",
            INIT_5A => X"0000002e00000000000000190000000000000020000000000000001e00000000",
            INIT_5B => X"0000000000000000000000020000000000000001000000000000001700000000",
            INIT_5C => X"00000066000000000000005f0000000000000030000000000000005e00000000",
            INIT_5D => X"0000005d0000000000000064000000000000006b000000000000006e00000000",
            INIT_5E => X"00000016000000000000002f0000000000000049000000000000005000000000",
            INIT_5F => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000001800000000000000170000000000000000000000000000000000000000",
            INIT_64 => X"000000030000000000000003000000000000001a000000000000002500000000",
            INIT_65 => X"0000000700000000000000000000000000000000000000000000001400000000",
            INIT_66 => X"0000000000000000000000000000000000000011000000000000003e00000000",
            INIT_67 => X"0000000300000000000000000000000000000018000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_69 => X"0000000000000000000000020000000000000046000000000000001500000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000b000000000000000a000000000000000a000000000000000a00000000",
            INIT_70 => X"0000000a0000000000000008000000000000000a000000000000000a00000000",
            INIT_71 => X"0000000a0000000000000009000000000000000d000000000000000b00000000",
            INIT_72 => X"0000000b0000000000000009000000000000000b000000000000000a00000000",
            INIT_73 => X"0000000b000000000000000b000000000000000a000000000000000b00000000",
            INIT_74 => X"00000006000000000000000b000000000000000a000000000000000c00000000",
            INIT_75 => X"0000000b000000000000000a000000000000001a000000000000002b00000000",
            INIT_76 => X"0000000b000000000000000b000000000000000a000000000000000c00000000",
            INIT_77 => X"000000100000000000000009000000000000000b000000000000000a00000000",
            INIT_78 => X"000000320000000000000010000000000000001a000000000000000900000000",
            INIT_79 => X"0000000c000000000000000c000000000000000a000000000000002a00000000",
            INIT_7A => X"0000000a000000000000000e0000000000000010000000000000001a00000000",
            INIT_7B => X"0000000000000000000000220000000000000000000000000000000a00000000",
            INIT_7C => X"00000036000000000000001b0000000000000010000000000000001500000000",
            INIT_7D => X"00000049000000000000000e000000000000000f000000000000001000000000",
            INIT_7E => X"0000000c000000000000000c0000000000000031000000000000004b00000000",
            INIT_7F => X"0000001400000000000000040000000000000016000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE11;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12 : if BRAM_NAME = "samplegold_layersamples_instance12" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d0000000000000027000000000000001a000000000000000f00000000",
            INIT_01 => X"0000001000000000000000040000000000000015000000000000004300000000",
            INIT_02 => X"0000001500000000000000180000000000000012000000000000001200000000",
            INIT_03 => X"0000000c000000000000002a0000000000000028000000000000002c00000000",
            INIT_04 => X"0000004000000000000000000000000000000009000000000000000c00000000",
            INIT_05 => X"00000036000000000000005c0000000000000049000000000000001800000000",
            INIT_06 => X"0000004500000000000000000000000000000000000000000000001d00000000",
            INIT_07 => X"0000001300000000000000100000000000000044000000000000004600000000",
            INIT_08 => X"0000003e0000000000000020000000000000001d000000000000001800000000",
            INIT_09 => X"00000047000000000000001a0000000000000032000000000000005100000000",
            INIT_0A => X"0000000d00000000000000150000000000000000000000000000001900000000",
            INIT_0B => X"0000002700000000000000240000000000000029000000000000002b00000000",
            INIT_0C => X"0000007f000000000000002d0000000000000021000000000000002b00000000",
            INIT_0D => X"00000019000000000000000c0000000000000002000000000000000200000000",
            INIT_0E => X"0000001300000000000000000000000000000020000000000000001100000000",
            INIT_0F => X"00000030000000000000001d0000000000000023000000000000001e00000000",
            INIT_10 => X"0000004300000000000000590000000000000032000000000000003700000000",
            INIT_11 => X"00000047000000000000004e000000000000004e000000000000005000000000",
            INIT_12 => X"000000330000000000000042000000000000003d000000000000003900000000",
            INIT_13 => X"00000035000000000000003a0000000000000034000000000000004100000000",
            INIT_14 => X"0000004b0000000000000054000000000000003c000000000000003400000000",
            INIT_15 => X"0000006200000000000000610000000000000057000000000000005400000000",
            INIT_16 => X"000000490000000000000048000000000000004e000000000000005b00000000",
            INIT_17 => X"0000002b000000000000002b0000000000000045000000000000004700000000",
            INIT_18 => X"0000000300000000000000000000000000000034000000000000000b00000000",
            INIT_19 => X"0000001f000000000000004a000000000000002a000000000000001300000000",
            INIT_1A => X"0000001e000000000000002e0000000000000034000000000000003400000000",
            INIT_1B => X"0000000000000000000000230000000000000016000000000000001a00000000",
            INIT_1C => X"00000011000000000000000b000000000000001e000000000000002700000000",
            INIT_1D => X"000000000000000000000000000000000000005f000000000000001800000000",
            INIT_1E => X"0000001300000000000000120000000000000000000000000000000000000000",
            INIT_1F => X"0000001200000000000000000000000000000027000000000000001a00000000",
            INIT_20 => X"0000001300000000000000120000000000000011000000000000001600000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_22 => X"00000020000000000000000c000000000000000f000000000000000300000000",
            INIT_23 => X"0000000f00000000000000050000000000000000000000000000002900000000",
            INIT_24 => X"0000002200000000000000140000000000000010000000000000001000000000",
            INIT_25 => X"0000000400000000000000090000000000000000000000000000000300000000",
            INIT_26 => X"00000025000000000000001b0000000000000014000000000000000a00000000",
            INIT_27 => X"0000001300000000000000130000000000000013000000000000001000000000",
            INIT_28 => X"0000001200000000000000130000000000000013000000000000001400000000",
            INIT_29 => X"0000001400000000000000140000000000000013000000000000001400000000",
            INIT_2A => X"0000000f00000000000000150000000000000013000000000000001400000000",
            INIT_2B => X"0000001300000000000000120000000000000013000000000000001300000000",
            INIT_2C => X"0000001000000000000000120000000000000013000000000000001200000000",
            INIT_2D => X"00000012000000000000001f0000000000000021000000000000000000000000",
            INIT_2E => X"0000001200000000000000100000000000000014000000000000001300000000",
            INIT_2F => X"0000001100000000000000140000000000000012000000000000001400000000",
            INIT_30 => X"0000000000000000000000000000000000000001000000000000001400000000",
            INIT_31 => X"0000001300000000000000120000000000000033000000000000003100000000",
            INIT_32 => X"000000170000000000000013000000000000001a000000000000001400000000",
            INIT_33 => X"0000002b00000000000000000000000000000013000000000000001400000000",
            INIT_34 => X"0000001c00000000000000090000000000000011000000000000000000000000",
            INIT_35 => X"0000001600000000000000150000000000000013000000000000004c00000000",
            INIT_36 => X"00000012000000000000003f000000000000000d000000000000000000000000",
            INIT_37 => X"0000000a000000000000002f0000000000000000000000000000001300000000",
            INIT_38 => X"000000000000000000000002000000000000000c000000000000001f00000000",
            INIT_39 => X"00000028000000000000001d000000000000002c000000000000000000000000",
            INIT_3A => X"0000001900000000000000030000000000000031000000000000003f00000000",
            INIT_3B => X"0000001a0000000000000012000000000000000e000000000000000000000000",
            INIT_3C => X"0000000300000000000000190000000000000007000000000000000000000000",
            INIT_3D => X"0000000a0000000000000000000000000000001f000000000000006b00000000",
            INIT_3E => X"0000000000000000000000010000000000000026000000000000001100000000",
            INIT_3F => X"00000014000000000000005c0000000000000035000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000500000000000000070000000000000000000000000000000200000000",
            INIT_41 => X"000000010000000000000062000000000000002c000000000000002100000000",
            INIT_42 => X"00000050000000000000000e000000000000000a000000000000004900000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_44 => X"0000003b0000000000000024000000000000001e000000000000000800000000",
            INIT_45 => X"00000039000000000000002b000000000000001b00000000000000c500000000",
            INIT_46 => X"0000000000000000000000150000000000000008000000000000002a00000000",
            INIT_47 => X"00000008000000000000001c0000000000000012000000000000001e00000000",
            INIT_48 => X"0000006000000000000000000000000000000002000000000000000e00000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000e00000000000000000000000000000021000000000000001500000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000001c00000000000000170000000000000004000000000000000000000000",
            INIT_50 => X"0000000b00000000000000410000000000000000000000000000002d00000000",
            INIT_51 => X"00000058000000000000001d000000000000000b000000000000000400000000",
            INIT_52 => X"000000280000000000000016000000000000000f000000000000000500000000",
            INIT_53 => X"0000003700000000000000110000000000000025000000000000003500000000",
            INIT_54 => X"0000000000000000000000100000000000000027000000000000000000000000",
            INIT_55 => X"0000000000000000000000880000000000000019000000000000000c00000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000470000000000000035000000000000002100000000",
            INIT_58 => X"00000017000000000000000f000000000000001c000000000000001800000000",
            INIT_59 => X"0000000000000000000000070000000000000055000000000000001900000000",
            INIT_5A => X"000000240000000000000044000000000000002c000000000000000000000000",
            INIT_5B => X"0000001a0000000000000000000000000000003e000000000000003500000000",
            INIT_5C => X"0000001e000000000000001d000000000000001c000000000000001f00000000",
            INIT_5D => X"0000005300000000000000260000000000000018000000000000003e00000000",
            INIT_5E => X"00000035000000000000002e000000000000001f000000000000002e00000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000003d00000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000022000000000000002a00000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000200000000000000080000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000003f00000000",
            INIT_7C => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000001a0000000000000000000000000000004d000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE12;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13 : if BRAM_NAME = "samplegold_layersamples_instance13" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000070000000000000012000000000000000b00000000",
            INIT_0A => X"0000003e000000000000003f0000000000000062000000000000004500000000",
            INIT_0B => X"000000000000000000000000000000000000003d000000000000004a00000000",
            INIT_0C => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_0D => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000010000000000000003000000000000000b000000000000000200000000",
            INIT_11 => X"0000000000000000000000000000000000000009000000000000000900000000",
            INIT_12 => X"0000000c00000000000000200000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000001b0000000000000019000000000000001c000000000000002000000000",
            INIT_15 => X"0000002c0000000000000000000000000000000c000000000000001c00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_17 => X"0000002c000000000000002c0000000000000000000000000000000000000000",
            INIT_18 => X"0000002c000000000000002c000000000000002c000000000000002c00000000",
            INIT_19 => X"0000002d000000000000002c000000000000002d000000000000002c00000000",
            INIT_1A => X"0000002c000000000000002c000000000000002c000000000000002a00000000",
            INIT_1B => X"0000002c000000000000002c000000000000002c000000000000002c00000000",
            INIT_1C => X"0000002b000000000000002c000000000000002b000000000000002c00000000",
            INIT_1D => X"000000110000000000000030000000000000002e000000000000002b00000000",
            INIT_1E => X"0000002c000000000000002b000000000000002c000000000000002000000000",
            INIT_1F => X"0000002c000000000000002c000000000000002c000000000000002b00000000",
            INIT_20 => X"000000310000000000000027000000000000002f000000000000002c00000000",
            INIT_21 => X"00000017000000000000000d0000000000000009000000000000001700000000",
            INIT_22 => X"0000001f000000000000002c000000000000002c000000000000002b00000000",
            INIT_23 => X"0000002e000000000000002d0000000000000029000000000000002600000000",
            INIT_24 => X"0000000e00000000000000290000000000000019000000000000003900000000",
            INIT_25 => X"000000270000000000000015000000000000000a000000000000000f00000000",
            INIT_26 => X"000000000000000000000000000000000000002a000000000000002800000000",
            INIT_27 => X"0000002a000000000000002b000000000000002b000000000000001000000000",
            INIT_28 => X"0000002700000000000000260000000000000028000000000000002a00000000",
            INIT_29 => X"0000000000000000000000090000000000000011000000000000001f00000000",
            INIT_2A => X"00000036000000000000001b0000000000000011000000000000002600000000",
            INIT_2B => X"0000000e00000000000000190000000000000024000000000000002000000000",
            INIT_2C => X"0000000b000000000000001f000000000000000f000000000000001000000000",
            INIT_2D => X"000000240000000000000011000000000000001a000000000000001200000000",
            INIT_2E => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000003100000000",
            INIT_30 => X"000000190000000000000022000000000000002b000000000000000000000000",
            INIT_31 => X"000000000000000000000000000000000000001e000000000000000c00000000",
            INIT_32 => X"0000000600000000000000040000000000000000000000000000000300000000",
            INIT_33 => X"0000000c00000000000000310000000000000017000000000000000500000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000260000000000000000000000000000000c000000000000000000000000",
            INIT_36 => X"0000002800000000000000290000000000000029000000000000001400000000",
            INIT_37 => X"0000000c0000000000000011000000000000000c000000000000001d00000000",
            INIT_38 => X"000000000000000000000001000000000000000e000000000000000700000000",
            INIT_39 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000300000000000000038000000000000002c000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000010000000000000034000000000000004a00000000",
            INIT_4B => X"0000000500000000000000000000000000000004000000000000000600000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"00000000000000000000000d0000000000000004000000000000000000000000",
            INIT_4F => X"0000000000000000000000090000000000000003000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000500000000000000000000000000000009000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000001000000000000000000000000000000000000000000000000500000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000039000000000000001e000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_6B => X"0000002a00000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000090000000000000000000000000000000400000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000002b00000000000000130000000000000000000000000000001e00000000",
            INIT_7A => X"000000240000000000000000000000000000000c000000000000002200000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_7C => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000001a00000000000000160000000000000005000000000000001600000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE13;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14 : if BRAM_NAME = "samplegold_layersamples_instance14" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e000000000000005d0000000000000000000000000000000000000000",
            INIT_01 => X"0000001c000000000000001d000000000000001c000000000000001900000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"00000000000000000000000b000000000000000b000000000000000000000000",
            INIT_04 => X"00000027000000000000002c000000000000004b000000000000000000000000",
            INIT_05 => X"0000000b000000000000001f000000000000001f000000000000002400000000",
            INIT_06 => X"0000001200000000000000020000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000003000000000000000d00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000220000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000002e00000000000000180000000000000000000000000000000000000000",
            INIT_4E => X"000000000000000000000016000000000000003d000000000000002e00000000",
            INIT_4F => X"0000001e00000000000000170000000000000020000000000000000000000000",
            INIT_50 => X"00000010000000000000000f0000000000000014000000000000001a00000000",
            INIT_51 => X"0000000f00000000000000040000000000000005000000000000000b00000000",
            INIT_52 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000800000000000000000000000000000000000000000000000a00000000",
            INIT_54 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_56 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000f00000000000000120000000000000013000000000000000700000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000200000000000000020000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_5E => X"000000210000000000000025000000000000000d000000000000000000000000",
            INIT_5F => X"0000001900000000000000150000000000000008000000000000000a00000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000001300000000000000000000000000000000000000000000001200000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_65 => X"0000001b00000000000000160000000000000011000000000000000200000000",
            INIT_66 => X"0000001b000000000000000b0000000000000008000000000000000d00000000",
            INIT_67 => X"00000011000000000000001e0000000000000009000000000000001c00000000",
            INIT_68 => X"0000000900000000000000180000000000000012000000000000000400000000",
            INIT_69 => X"00000015000000000000001e0000000000000007000000000000000d00000000",
            INIT_6A => X"00000007000000000000000f000000000000001e000000000000001500000000",
            INIT_6B => X"0000000f000000000000000f0000000000000003000000000000000700000000",
            INIT_6C => X"0000000f000000000000000a000000000000001b000000000000000a00000000",
            INIT_6D => X"0000001f000000000000001b000000000000001a000000000000000d00000000",
            INIT_6E => X"0000001000000000000000280000000000000024000000000000001900000000",
            INIT_6F => X"00000009000000000000001d0000000000000013000000000000000500000000",
            INIT_70 => X"0000000a000000000000000e000000000000000e000000000000000e00000000",
            INIT_71 => X"0000001200000000000000190000000000000025000000000000002600000000",
            INIT_72 => X"00000014000000000000001b0000000000000015000000000000000f00000000",
            INIT_73 => X"0000000b00000000000000120000000000000000000000000000000500000000",
            INIT_74 => X"000000080000000000000005000000000000000a000000000000000d00000000",
            INIT_75 => X"00000007000000000000000b000000000000000b000000000000000900000000",
            INIT_76 => X"00000014000000000000000c000000000000000a000000000000000300000000",
            INIT_77 => X"0000000b000000000000000b000000000000000b000000000000000a00000000",
            INIT_78 => X"0000003c000000000000002f0000000000000008000000000000000b00000000",
            INIT_79 => X"00000035000000000000003a000000000000003a000000000000003f00000000",
            INIT_7A => X"000000330000000000000033000000000000002a000000000000003200000000",
            INIT_7B => X"0000002f000000000000002d000000000000002f000000000000002800000000",
            INIT_7C => X"0000003800000000000000340000000000000029000000000000003300000000",
            INIT_7D => X"0000002d000000000000002b000000000000002f000000000000002f00000000",
            INIT_7E => X"0000002f0000000000000019000000000000002f000000000000002900000000",
            INIT_7F => X"00000032000000000000002c000000000000002b000000000000003200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE14;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15 : if BRAM_NAME = "samplegold_layersamples_instance15" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000024000000000000002e000000000000002b000000000000002100000000",
            INIT_01 => X"0000002200000000000000200000000000000023000000000000002500000000",
            INIT_02 => X"00000027000000000000003c0000000000000000000000000000002a00000000",
            INIT_03 => X"00000017000000000000002d0000000000000023000000000000001f00000000",
            INIT_04 => X"0000001a00000000000000210000000000000027000000000000002a00000000",
            INIT_05 => X"0000000700000000000000190000000000000017000000000000002100000000",
            INIT_06 => X"00000025000000000000001c000000000000001a000000000000000b00000000",
            INIT_07 => X"0000000f000000000000000f0000000000000019000000000000001500000000",
            INIT_08 => X"00000012000000000000000e0000000000000015000000000000001000000000",
            INIT_09 => X"000000190000000000000016000000000000000e000000000000001500000000",
            INIT_0A => X"0000000d000000000000001e0000000000000027000000000000001900000000",
            INIT_0B => X"0000001100000000000000230000000000000020000000000000001500000000",
            INIT_0C => X"0000002700000000000000260000000000000024000000000000001d00000000",
            INIT_0D => X"00000030000000000000001b000000000000001b000000000000001c00000000",
            INIT_0E => X"000000050000000000000016000000000000000d000000000000002d00000000",
            INIT_0F => X"0000002a0000000000000018000000000000001b000000000000002400000000",
            INIT_10 => X"0000002f0000000000000034000000000000002a000000000000003200000000",
            INIT_11 => X"000000220000000000000036000000000000002d000000000000003100000000",
            INIT_12 => X"0000002e00000000000000000000000000000019000000000000000b00000000",
            INIT_13 => X"0000003b000000000000003f0000000000000038000000000000002e00000000",
            INIT_14 => X"00000029000000000000002e0000000000000035000000000000003700000000",
            INIT_15 => X"0000001b00000000000000200000000000000019000000000000001100000000",
            INIT_16 => X"0000001c00000000000000310000000000000023000000000000000000000000",
            INIT_17 => X"000000280000000000000035000000000000003a000000000000003900000000",
            INIT_18 => X"00000019000000000000002e0000000000000021000000000000002100000000",
            INIT_19 => X"0000001b000000000000001c0000000000000021000000000000002b00000000",
            INIT_1A => X"000000310000000000000042000000000000002d000000000000001200000000",
            INIT_1B => X"0000002d0000000000000032000000000000002e000000000000002c00000000",
            INIT_1C => X"0000002600000000000000210000000000000016000000000000001f00000000",
            INIT_1D => X"000000090000000000000004000000000000000c000000000000001c00000000",
            INIT_1E => X"0000002100000000000000310000000000000031000000000000002e00000000",
            INIT_1F => X"0000000f00000000000000150000000000000023000000000000002400000000",
            INIT_20 => X"00000008000000000000000d000000000000001e000000000000002d00000000",
            INIT_21 => X"0000003500000000000000030000000000000003000000000000000500000000",
            INIT_22 => X"00000026000000000000001e000000000000001a000000000000002a00000000",
            INIT_23 => X"00000014000000000000000d0000000000000011000000000000003700000000",
            INIT_24 => X"0000000c00000000000000010000000000000009000000000000001300000000",
            INIT_25 => X"0000001800000000000000270000000000000002000000000000000500000000",
            INIT_26 => X"00000011000000000000000d0000000000000012000000000000001000000000",
            INIT_27 => X"00000006000000000000000a0000000000000013000000000000001500000000",
            INIT_28 => X"000000080000000000000001000000000000000d000000000000000a00000000",
            INIT_29 => X"0000000a000000000000000c000000000000000d000000000000000700000000",
            INIT_2A => X"000000090000000000000005000000000000000b000000000000000f00000000",
            INIT_2B => X"0000000700000000000000080000000000000015000000000000000900000000",
            INIT_2C => X"00000009000000000000000a0000000000000006000000000000000900000000",
            INIT_2D => X"0000000a00000000000000080000000000000008000000000000000400000000",
            INIT_2E => X"00000003000000000000000a000000000000000c000000000000000c00000000",
            INIT_2F => X"00000009000000000000000a0000000000000000000000000000001500000000",
            INIT_30 => X"000000780000000000000000000000000000000a000000000000000900000000",
            INIT_31 => X"0000005700000000000000550000000000000044000000000000002b00000000",
            INIT_32 => X"0000004200000000000000670000000000000051000000000000005100000000",
            INIT_33 => X"0000005600000000000000480000000000000056000000000000005500000000",
            INIT_34 => X"0000002700000000000000720000000000000043000000000000005700000000",
            INIT_35 => X"0000005100000000000000500000000000000057000000000000003800000000",
            INIT_36 => X"0000008f00000000000000430000000000000053000000000000005400000000",
            INIT_37 => X"0000005a000000000000005a000000000000003c000000000000001100000000",
            INIT_38 => X"0000002c0000000000000022000000000000006f000000000000003e00000000",
            INIT_39 => X"00000067000000000000004b000000000000004a000000000000004e00000000",
            INIT_3A => X"0000000000000000000000ba0000000000000033000000000000004100000000",
            INIT_3B => X"00000037000000000000004e0000000000000061000000000000003400000000",
            INIT_3C => X"0000003c00000000000000440000000000000023000000000000006c00000000",
            INIT_3D => X"00000064000000000000005c000000000000003d000000000000005000000000",
            INIT_3E => X"0000001a0000000000000019000000000000005a000000000000006600000000",
            INIT_3F => X"00000042000000000000002b000000000000004e000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003a00000000000000250000000000000039000000000000002e00000000",
            INIT_41 => X"00000050000000000000006b0000000000000039000000000000003500000000",
            INIT_42 => X"0000000e000000000000001a0000000000000030000000000000004e00000000",
            INIT_43 => X"0000001800000000000000120000000000000020000000000000005600000000",
            INIT_44 => X"0000002f0000000000000027000000000000000e000000000000005000000000",
            INIT_45 => X"0000003d000000000000003e000000000000005c000000000000003e00000000",
            INIT_46 => X"0000001b0000000000000073000000000000001d000000000000000000000000",
            INIT_47 => X"000000400000000000000038000000000000002e000000000000005b00000000",
            INIT_48 => X"0000004100000000000000430000000000000026000000000000000900000000",
            INIT_49 => X"0000000a00000000000000340000000000000033000000000000003e00000000",
            INIT_4A => X"000000710000000000000044000000000000006b000000000000003300000000",
            INIT_4B => X"000000380000000000000031000000000000003b000000000000003a00000000",
            INIT_4C => X"000000630000000000000058000000000000004f000000000000004700000000",
            INIT_4D => X"000000210000000000000018000000000000007c000000000000005300000000",
            INIT_4E => X"0000005600000000000000150000000000000068000000000000004000000000",
            INIT_4F => X"0000006400000000000000420000000000000020000000000000005000000000",
            INIT_50 => X"0000003100000000000000460000000000000051000000000000006000000000",
            INIT_51 => X"000000400000000000000038000000000000001a000000000000005d00000000",
            INIT_52 => X"0000002600000000000000490000000000000044000000000000004c00000000",
            INIT_53 => X"00000042000000000000003f0000000000000054000000000000004500000000",
            INIT_54 => X"0000003e00000000000000380000000000000061000000000000004f00000000",
            INIT_55 => X"00000059000000000000005b000000000000005f000000000000003f00000000",
            INIT_56 => X"00000054000000000000004c0000000000000033000000000000002b00000000",
            INIT_57 => X"000000730000000000000031000000000000004a000000000000006500000000",
            INIT_58 => X"00000056000000000000003f0000000000000000000000000000004d00000000",
            INIT_59 => X"0000003b00000000000000360000000000000047000000000000005600000000",
            INIT_5A => X"00000039000000000000006f0000000000000043000000000000000e00000000",
            INIT_5B => X"0000004c0000000000000073000000000000001c000000000000002700000000",
            INIT_5C => X"0000003300000000000000440000000000000038000000000000002900000000",
            INIT_5D => X"00000022000000000000002d000000000000002a000000000000003400000000",
            INIT_5E => X"0000003800000000000000440000000000000060000000000000005100000000",
            INIT_5F => X"0000003800000000000000330000000000000031000000000000002f00000000",
            INIT_60 => X"0000003e000000000000001f0000000000000030000000000000003100000000",
            INIT_61 => X"000000220000000000000025000000000000001f000000000000002000000000",
            INIT_62 => X"000000260000000000000029000000000000001d000000000000002400000000",
            INIT_63 => X"000000470000000000000004000000000000002a000000000000002100000000",
            INIT_64 => X"0000001a00000000000000230000000000000025000000000000002500000000",
            INIT_65 => X"000000140000000000000011000000000000001e000000000000002100000000",
            INIT_66 => X"00000023000000000000001d0000000000000017000000000000001200000000",
            INIT_67 => X"0000001e00000000000000510000000000000000000000000000003000000000",
            INIT_68 => X"0000003e0000000000000016000000000000001c000000000000002100000000",
            INIT_69 => X"0000000000000000000000080000000000000005000000000000000800000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000a00000000000000000000000000000000000000000000000d00000000",
            INIT_7C => X"000000320000000000000000000000000000000c000000000000001d00000000",
            INIT_7D => X"000000000000000000000000000000000000000f000000000000002100000000",
            INIT_7E => X"000000450000000000000069000000000000002d000000000000000800000000",
            INIT_7F => X"0000000000000000000000030000000000000006000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE15;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16 : if BRAM_NAME = "samplegold_layersamples_instance16" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000040000000000000004f0000000000000032000000000000002000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000003400000000",
            INIT_03 => X"0000005e000000000000003a0000000000000023000000000000000000000000",
            INIT_04 => X"00000016000000000000001f000000000000002f000000000000005900000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_06 => X"0000007200000000000000100000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000c00000000000000400000000000000020000000000000000b00000000",
            INIT_0A => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000017000000000000004300000000",
            INIT_0C => X"0000000000000000000000000000000000000011000000000000001900000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000020000000000000003000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_1D => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_1E => X"0000000b00000000000000050000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000d000000000000000b0000000000000002000000000000000a00000000",
            INIT_24 => X"0000000b000000000000000e000000000000000f000000000000000d00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000090000000000000012000000000000000d000000000000000100000000",
            INIT_27 => X"0000000f00000000000000000000000000000025000000000000000a00000000",
            INIT_28 => X"0000000000000000000000110000000000000016000000000000001900000000",
            INIT_29 => X"0000001a00000000000000130000000000000000000000000000000000000000",
            INIT_2A => X"0000000900000000000000110000000000000021000000000000001700000000",
            INIT_2B => X"0000001d00000000000000000000000000000000000000000000002400000000",
            INIT_2C => X"0000000700000000000000100000000000000016000000000000001e00000000",
            INIT_2D => X"000000240000000000000031000000000000001f000000000000002100000000",
            INIT_2E => X"0000000000000000000000130000000000000024000000000000002300000000",
            INIT_2F => X"0000002300000000000000000000000000000010000000000000000000000000",
            INIT_30 => X"0000000d00000000000000040000000000000001000000000000002400000000",
            INIT_31 => X"00000009000000000000001c000000000000001f000000000000001400000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_33 => X"00000029000000000000002e0000000000000002000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000000000000000000001d0000000000000014000000000000003a00000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000002300000000000000190000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000019000000000000003400000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"00000018000000000000001a0000000000000018000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000001200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000001400000000000000140000000000000008000000000000000d00000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000000000000000000003000000000000000c000000000000000900000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"000000080000000000000000000000000000000a000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"00000004000000000000000c0000000000000000000000000000000100000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000500000000000000000000000000000000000000000000000900000000",
            INIT_61 => X"00000000000000000000000b000000000000000f000000000000000000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000e00000000000000460000000000000000000000000000000d00000000",
            INIT_64 => X"0000000000000000000000090000000000000000000000000000000000000000",
            INIT_65 => X"00000000000000000000000f000000000000000e000000000000001900000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_67 => X"0000004100000000000000150000000000000005000000000000000000000000",
            INIT_68 => X"0000000900000000000000010000000000000017000000000000000000000000",
            INIT_69 => X"00000010000000000000000d0000000000000019000000000000000300000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_6B => X"0000000000000000000000190000000000000015000000000000000000000000",
            INIT_6C => X"000000000000000000000011000000000000000e000000000000001200000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_6E => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000180000000000000000000000000000001200000000",
            INIT_70 => X"0000001700000000000000000000000000000000000000000000000100000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_72 => X"0000000700000000000000210000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_74 => X"0000000000000000000000030000000000000008000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000170000000000000014000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_79 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_7B => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE16;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17 : if BRAM_NAME = "samplegold_layersamples_instance17" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_02 => X"0000001900000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000200000000000000000000000000000002000000000000000000000000",
            INIT_0A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_0C => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_0D => X"0000000300000000000000050000000000000000000000000000000100000000",
            INIT_0E => X"0000000400000000000000030000000000000008000000000000000200000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_10 => X"0000000400000000000000060000000000000000000000000000002200000000",
            INIT_11 => X"0000000000000000000000000000000000000008000000000000000400000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000300000000000000020000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000110000000000000005000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"00000001000000000000000a0000000000000009000000000000000200000000",
            INIT_50 => X"000000050000000000000003000000000000000e000000000000001500000000",
            INIT_51 => X"0000000000000000000000040000000000000000000000000000000800000000",
            INIT_52 => X"0000000400000000000000010000000000000000000000000000000000000000",
            INIT_53 => X"0000001e000000000000001e0000000000000023000000000000000a00000000",
            INIT_54 => X"0000000f0000000000000011000000000000002d000000000000001200000000",
            INIT_55 => X"0000002d000000000000000f0000000000000026000000000000000900000000",
            INIT_56 => X"0000001d00000000000000150000000000000025000000000000002c00000000",
            INIT_57 => X"00000000000000000000001a0000000000000024000000000000000f00000000",
            INIT_58 => X"0000003b000000000000003f000000000000004e000000000000001200000000",
            INIT_59 => X"0000003500000000000000260000000000000027000000000000003f00000000",
            INIT_5A => X"00000039000000000000003a0000000000000047000000000000004200000000",
            INIT_5B => X"0000000000000000000000030000000000000009000000000000001600000000",
            INIT_5C => X"0000000000000000000000170000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"00000001000000000000000d0000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"000000000000000000000000000000000000000c000000000000000d00000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000002f000000000000001b0000000000000005000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000010000000000000001c0000000000000016000000000000000000000000",
            INIT_67 => X"000000000000000000000000000000000000000a000000000000000c00000000",
            INIT_68 => X"0000000100000000000000000000000000000023000000000000001600000000",
            INIT_69 => X"000000000000000000000001000000000000001a000000000000001300000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"00000000000000000000002f000000000000000e000000000000000100000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000002b00000000000000280000000000000000000000000000000000000000",
            INIT_6E => X"00000033000000000000001c0000000000000000000000000000000400000000",
            INIT_6F => X"0000000000000000000000000000000000000018000000000000002e00000000",
            INIT_70 => X"0000001300000000000000300000000000000023000000000000000000000000",
            INIT_71 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000012000000000000001c0000000000000022000000000000003200000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_74 => X"0000004200000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000001c00000000000000040000000000000000000000000000001e00000000",
            INIT_76 => X"0000000400000000000000030000000000000000000000000000000500000000",
            INIT_77 => X"0000002800000000000000430000000000000037000000000000001b00000000",
            INIT_78 => X"0000000700000000000000040000000000000006000000000000001200000000",
            INIT_79 => X"0000000500000000000000020000000000000009000000000000001b00000000",
            INIT_7A => X"0000000400000000000000000000000000000000000000000000000e00000000",
            INIT_7B => X"0000000f00000000000000050000000000000004000000000000000a00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_7D => X"0000000000000000000000010000000000000003000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE17;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18 : if BRAM_NAME = "samplegold_layersamples_instance18" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000700000000000000020000000000000009000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000f300000000000000c300000000000000df000000000000000d00000000",
            INIT_03 => X"000000f800000000000000f100000000000000fb00000000000000f500000000",
            INIT_04 => X"000000f6000000000000010000000000000000f400000000000000f900000000",
            INIT_05 => X"000000f400000000000000fd00000000000000f500000000000000fb00000000",
            INIT_06 => X"000000e900000000000000ec00000000000000bf00000000000000dd00000000",
            INIT_07 => X"000000f900000000000000ef00000000000000e500000000000000f400000000",
            INIT_08 => X"000000f800000000000000de00000000000000ee00000000000000f000000000",
            INIT_09 => X"000000d400000000000000f100000000000000fe00000000000000f300000000",
            INIT_0A => X"000000e400000000000000da00000000000000da00000000000000b000000000",
            INIT_0B => X"000000e600000000000000da00000000000000e000000000000000db00000000",
            INIT_0C => X"000000ed00000000000000f300000000000000bd00000000000000d000000000",
            INIT_0D => X"0000009c00000000000000c300000000000000ec00000000000000ee00000000",
            INIT_0E => X"000000cb00000000000000cc00000000000000cb00000000000000c100000000",
            INIT_0F => X"000000a500000000000000a800000000000000b900000000000000ce00000000",
            INIT_10 => X"000000d200000000000000d3000000000000008c000000000000007a00000000",
            INIT_11 => X"00000093000000000000007e000000000000009700000000000000c800000000",
            INIT_12 => X"000000b200000000000000a900000000000000a4000000000000009700000000",
            INIT_13 => X"000000740000000000000079000000000000008d00000000000000b800000000",
            INIT_14 => X"0000007d000000000000008d0000000000000068000000000000006400000000",
            INIT_15 => X"00000063000000000000006c000000000000005e000000000000006000000000",
            INIT_16 => X"0000009000000000000000910000000000000079000000000000007900000000",
            INIT_17 => X"0000008e0000000000000073000000000000007c000000000000007d00000000",
            INIT_18 => X"000000740000000000000058000000000000009d000000000000006b00000000",
            INIT_19 => X"000000a00000000000000074000000000000006f000000000000006900000000",
            INIT_1A => X"00000086000000000000009200000000000000a200000000000000a000000000",
            INIT_1B => X"000000ad00000000000000b0000000000000008f000000000000008b00000000",
            INIT_1C => X"0000008000000000000000860000000000000053000000000000007300000000",
            INIT_1D => X"000000c600000000000000b80000000000000099000000000000008a00000000",
            INIT_1E => X"000000a500000000000000c400000000000000c200000000000000cf00000000",
            INIT_1F => X"0000006500000000000000a200000000000000a2000000000000009800000000",
            INIT_20 => X"000000b0000000000000009f00000000000000a0000000000000004700000000",
            INIT_21 => X"000000c800000000000000d000000000000000d200000000000000cf00000000",
            INIT_22 => X"00000081000000000000009c00000000000000a800000000000000ba00000000",
            INIT_23 => X"00000096000000000000009100000000000000a1000000000000009600000000",
            INIT_24 => X"000000b500000000000000a90000000000000090000000000000008b00000000",
            INIT_25 => X"000000af00000000000000b500000000000000b500000000000000bb00000000",
            INIT_26 => X"000000a700000000000000aa00000000000000b400000000000000aa00000000",
            INIT_27 => X"000000af0000000000000064000000000000007f000000000000009600000000",
            INIT_28 => X"000000a900000000000000a900000000000000b000000000000000b000000000",
            INIT_29 => X"0000006f000000000000007900000000000000ab00000000000000bb00000000",
            INIT_2A => X"00000068000000000000008b000000000000009e00000000000000a400000000",
            INIT_2B => X"000000a90000000000000094000000000000003d000000000000005000000000",
            INIT_2C => X"0000009000000000000000750000000000000079000000000000009e00000000",
            INIT_2D => X"000000730000000000000066000000000000006e000000000000009d00000000",
            INIT_2E => X"0000003000000000000000410000000000000059000000000000006600000000",
            INIT_2F => X"0000008d000000000000008e000000000000007c000000000000002200000000",
            INIT_30 => X"00000064000000000000006f000000000000006a000000000000006d00000000",
            INIT_31 => X"0000004400000000000000550000000000000058000000000000005700000000",
            INIT_32 => X"0000001b00000000000000220000000000000035000000000000003800000000",
            INIT_33 => X"0000003c000000000000003c000000000000003d000000000000003900000000",
            INIT_34 => X"0000004000000000000000450000000000000041000000000000003f00000000",
            INIT_35 => X"0000002400000000000000310000000000000037000000000000004000000000",
            INIT_36 => X"00000018000000000000001b000000000000001c000000000000002100000000",
            INIT_37 => X"0000002b0000000000000023000000000000001f000000000000001600000000",
            INIT_38 => X"00000037000000000000002c0000000000000032000000000000002c00000000",
            INIT_39 => X"0000001b000000000000001a000000000000001f000000000000003900000000",
            INIT_3A => X"000000000000000000000000000000000000000c000000000000001e00000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000003b0000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000001f00000000000000080000000000000000000000000000000000000000",
            INIT_44 => X"0000000300000000000000000000000000000045000000000000000700000000",
            INIT_45 => X"0000001200000000000000000000000000000000000000000000000b00000000",
            INIT_46 => X"0000000a00000000000000000000000000000012000000000000000100000000",
            INIT_47 => X"0000006e000000000000000b0000000000000001000000000000000000000000",
            INIT_48 => X"00000010000000000000008b0000000000000046000000000000004600000000",
            INIT_49 => X"000000400000000000000046000000000000001f000000000000001d00000000",
            INIT_4A => X"0000004f00000000000000500000000000000051000000000000004a00000000",
            INIT_4B => X"000000030000000000000004000000000000003d000000000000003d00000000",
            INIT_4C => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000004700000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_50 => X"000000270000000000000000000000000000000b000000000000000000000000",
            INIT_51 => X"000000000000000000000011000000000000000a000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000380000000000000050000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000011000000000000003600000000",
            INIT_58 => X"0000002700000000000000140000000000000000000000000000000000000000",
            INIT_59 => X"0000001c00000000000000110000000000000000000000000000000500000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_5B => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_5E => X"000000000000000000000000000000000000000f000000000000002200000000",
            INIT_5F => X"0000002c00000000000000420000000000000036000000000000001700000000",
            INIT_60 => X"0000001700000000000000050000000000000000000000000000000000000000",
            INIT_61 => X"0000002c00000000000000250000000000000000000000000000002e00000000",
            INIT_62 => X"00000036000000000000003a000000000000001c000000000000000200000000",
            INIT_63 => X"0000000000000000000000230000000000000013000000000000002300000000",
            INIT_64 => X"00000000000000000000000e000000000000001c000000000000000200000000",
            INIT_65 => X"0000000f00000000000000050000000000000020000000000000000300000000",
            INIT_66 => X"0000001000000000000000160000000000000024000000000000001600000000",
            INIT_67 => X"0000002d000000000000000e000000000000000b000000000000001300000000",
            INIT_68 => X"00000029000000000000002c000000000000001b000000000000002800000000",
            INIT_69 => X"0000001a00000000000000230000000000000007000000000000000600000000",
            INIT_6A => X"000000030000000000000014000000000000000b000000000000000700000000",
            INIT_6B => X"00000010000000000000001f000000000000002c000000000000000000000000",
            INIT_6C => X"000000150000000000000015000000000000000c000000000000000500000000",
            INIT_6D => X"0000000700000000000000160000000000000000000000000000001000000000",
            INIT_6E => X"0000000000000000000000000000000000000002000000000000000b00000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001200000000000000050000000000000000000000000000000000000000",
            INIT_71 => X"0000000200000000000000050000000000000018000000000000000000000000",
            INIT_72 => X"0000002400000000000000230000000000000000000000000000000000000000",
            INIT_73 => X"00000027000000000000002e000000000000003b000000000000004500000000",
            INIT_74 => X"0000001d00000000000000090000000000000019000000000000002000000000",
            INIT_75 => X"0000000c0000000000000013000000000000000e000000000000001400000000",
            INIT_76 => X"00000039000000000000001a0000000000000014000000000000000e00000000",
            INIT_77 => X"000000140000000000000019000000000000001a000000000000003000000000",
            INIT_78 => X"0000000200000000000000170000000000000011000000000000001400000000",
            INIT_79 => X"0000000a00000000000000070000000000000016000000000000003200000000",
            INIT_7A => X"00000024000000000000002d000000000000000d000000000000001500000000",
            INIT_7B => X"00000003000000000000000a000000000000000b000000000000000900000000",
            INIT_7C => X"0000005300000000000000000000000000000021000000000000001b00000000",
            INIT_7D => X"0000001700000000000000080000000000000002000000000000002500000000",
            INIT_7E => X"0000000900000000000000110000000000000021000000000000000300000000",
            INIT_7F => X"0000000400000000000000000000000000000006000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE18;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19 : if BRAM_NAME = "samplegold_layersamples_instance19" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004b0000000000000049000000000000001e000000000000001f00000000",
            INIT_01 => X"0000002a00000000000000100000000000000007000000000000004700000000",
            INIT_02 => X"0000001f00000000000000320000000000000028000000000000003300000000",
            INIT_03 => X"0000002000000000000000120000000000000026000000000000002400000000",
            INIT_04 => X"00000020000000000000001c0000000000000035000000000000002800000000",
            INIT_05 => X"0000002c00000000000000360000000000000028000000000000000000000000",
            INIT_06 => X"000000260000000000000025000000000000002d000000000000001400000000",
            INIT_07 => X"00000024000000000000002c0000000000000025000000000000003400000000",
            INIT_08 => X"0000000b00000000000000000000000000000011000000000000003300000000",
            INIT_09 => X"00000026000000000000002e000000000000003b000000000000000000000000",
            INIT_0A => X"0000003600000000000000310000000000000041000000000000004d00000000",
            INIT_0B => X"000000330000000000000026000000000000002b000000000000002d00000000",
            INIT_0C => X"0000000000000000000000020000000000000000000000000000001400000000",
            INIT_0D => X"00000035000000000000002b0000000000000026000000000000003200000000",
            INIT_0E => X"0000002e00000000000000310000000000000033000000000000003400000000",
            INIT_0F => X"0000001a00000000000000300000000000000011000000000000003000000000",
            INIT_10 => X"0000004000000000000000040000000000000000000000000000000700000000",
            INIT_11 => X"0000003e00000000000000490000000000000055000000000000003e00000000",
            INIT_12 => X"0000002c000000000000002d000000000000003b000000000000003e00000000",
            INIT_13 => X"000000130000000000000012000000000000001c000000000000000000000000",
            INIT_14 => X"0000004700000000000000350000000000000008000000000000000900000000",
            INIT_15 => X"00000035000000000000003e000000000000003c000000000000003d00000000",
            INIT_16 => X"00000023000000000000002f0000000000000022000000000000002a00000000",
            INIT_17 => X"0000001300000000000000170000000000000010000000000000001f00000000",
            INIT_18 => X"0000003d00000000000000410000000000000050000000000000002300000000",
            INIT_19 => X"0000001f00000000000000440000000000000042000000000000003000000000",
            INIT_1A => X"00000024000000000000002f000000000000004b000000000000002500000000",
            INIT_1B => X"0000001b000000000000001a000000000000001c000000000000001c00000000",
            INIT_1C => X"0000003a000000000000002c0000000000000042000000000000005f00000000",
            INIT_1D => X"000000200000000000000016000000000000004b000000000000003d00000000",
            INIT_1E => X"0000002500000000000000230000000000000028000000000000003100000000",
            INIT_1F => X"0000004b00000000000000170000000000000023000000000000002000000000",
            INIT_20 => X"0000003a0000000000000035000000000000002b000000000000003800000000",
            INIT_21 => X"0000002c000000000000002a000000000000002e000000000000003900000000",
            INIT_22 => X"00000019000000000000002a0000000000000021000000000000002a00000000",
            INIT_23 => X"0000003700000000000000380000000000000020000000000000002400000000",
            INIT_24 => X"0000002c000000000000002c0000000000000033000000000000003100000000",
            INIT_25 => X"0000001600000000000000300000000000000028000000000000003000000000",
            INIT_26 => X"0000002400000000000000210000000000000024000000000000002300000000",
            INIT_27 => X"000000260000000000000025000000000000001d000000000000001f00000000",
            INIT_28 => X"0000002700000000000000250000000000000026000000000000002800000000",
            INIT_29 => X"00000025000000000000000d0000000000000041000000000000001c00000000",
            INIT_2A => X"0000000d00000000000000250000000000000025000000000000002100000000",
            INIT_2B => X"000000120000000000000028000000000000001f000000000000000000000000",
            INIT_2C => X"0000000900000000000000190000000000000011000000000000001900000000",
            INIT_2D => X"0000001a00000000000000070000000000000019000000000000002300000000",
            INIT_2E => X"0000000000000000000000160000000000000016000000000000000900000000",
            INIT_2F => X"0000001e000000000000000c000000000000002a000000000000001e00000000",
            INIT_30 => X"0000001b00000000000000170000000000000017000000000000000e00000000",
            INIT_31 => X"000000050000000000000023000000000000001f000000000000000000000000",
            INIT_32 => X"000000160000000000000000000000000000001b000000000000001400000000",
            INIT_33 => X"0000000e0000000000000021000000000000000c000000000000002d00000000",
            INIT_34 => X"00000000000000000000001e0000000000000013000000000000000c00000000",
            INIT_35 => X"0000001700000000000000030000000000000028000000000000005900000000",
            INIT_36 => X"0000002200000000000000180000000000000000000000000000002200000000",
            INIT_37 => X"000000000000000000000017000000000000000d000000000000001800000000",
            INIT_38 => X"0000001200000000000000000000000000000000000000000000000e00000000",
            INIT_39 => X"00000019000000000000001a0000000000000037000000000000000200000000",
            INIT_3A => X"0000001800000000000000000000000000000007000000000000000000000000",
            INIT_3B => X"000000000000000000000000000000000000000a000000000000000300000000",
            INIT_3C => X"0000002200000000000000120000000000000008000000000000000000000000",
            INIT_3D => X"0000002a0000000000000013000000000000000e000000000000003b00000000",
            INIT_3E => X"00000023000000000000001c000000000000000a000000000000002100000000",
            INIT_3F => X"000000100000000000000000000000000000001c000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000000000000000000046000000000000003e000000000000000f00000000",
            INIT_41 => X"0000000900000000000000230000000000000000000000000000003100000000",
            INIT_42 => X"00000003000000000000001b0000000000000031000000000000000000000000",
            INIT_43 => X"0000001f000000000000001b0000000000000006000000000000000d00000000",
            INIT_44 => X"0000000c00000000000000000000000000000021000000000000004c00000000",
            INIT_45 => X"0000002700000000000000180000000000000014000000000000000000000000",
            INIT_46 => X"0000001300000000000000190000000000000022000000000000003200000000",
            INIT_47 => X"000000220000000000000000000000000000000f000000000000000c00000000",
            INIT_48 => X"0000002500000000000000000000000000000009000000000000002000000000",
            INIT_49 => X"0000001a00000000000000210000000000000000000000000000000b00000000",
            INIT_4A => X"0000000300000000000000040000000000000002000000000000000700000000",
            INIT_4B => X"0000001b000000000000003d0000000000000000000000000000001c00000000",
            INIT_4C => X"00000000000000000000000c0000000000000007000000000000000b00000000",
            INIT_4D => X"0000000a00000000000000070000000000000025000000000000003300000000",
            INIT_4E => X"0000000d000000000000000c000000000000001b000000000000001a00000000",
            INIT_4F => X"0000000000000000000000030000000000000016000000000000001700000000",
            INIT_50 => X"0000000f00000000000000230000000000000004000000000000000000000000",
            INIT_51 => X"0000001c00000000000000150000000000000000000000000000000f00000000",
            INIT_52 => X"0000001f000000000000002f0000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"00000000000000000000000c0000000000000041000000000000000b00000000",
            INIT_55 => X"00000000000000000000003e0000000000000011000000000000000000000000",
            INIT_56 => X"0000000300000000000000080000000000000018000000000000000400000000",
            INIT_57 => X"00000000000000000000000b0000000000000003000000000000000000000000",
            INIT_58 => X"0000000b00000000000000000000000000000008000000000000002f00000000",
            INIT_59 => X"0000001700000000000000040000000000000004000000000000000a00000000",
            INIT_5A => X"0000001b00000000000000050000000000000007000000000000000d00000000",
            INIT_5B => X"0000000a000000000000000f000000000000000f000000000000000000000000",
            INIT_5C => X"00000019000000000000001a000000000000000d000000000000000800000000",
            INIT_5D => X"00000025000000000000000a0000000000000010000000000000001400000000",
            INIT_5E => X"0000000b000000000000000e000000000000000c000000000000000500000000",
            INIT_5F => X"0000001a00000000000000120000000000000017000000000000001700000000",
            INIT_60 => X"0000001d000000000000001a000000000000001a000000000000001a00000000",
            INIT_61 => X"000000000000000000000039000000000000000b000000000000001a00000000",
            INIT_62 => X"0000001a0000000000000015000000000000000d000000000000001400000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_76 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_78 => X"0000002200000000000000180000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000001e000000000000000b0000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_7D => X"0000001200000000000000030000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000016000000000000002c00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE19;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20 : if BRAM_NAME = "samplegold_layersamples_instance20" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000004500000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_1C => X"000000190000000000000019000000000000000f000000000000000800000000",
            INIT_1D => X"0000002a0000000000000024000000000000002c000000000000002400000000",
            INIT_1E => X"0000002f00000000000000280000000000000029000000000000002600000000",
            INIT_1F => X"000000100000000000000000000000000000000d000000000000002400000000",
            INIT_20 => X"0000002a00000000000000210000000000000024000000000000001900000000",
            INIT_21 => X"0000000000000000000000370000000000000024000000000000002900000000",
            INIT_22 => X"000000270000000000000032000000000000002b000000000000002a00000000",
            INIT_23 => X"0000002100000000000000160000000000000000000000000000001600000000",
            INIT_24 => X"0000001c00000000000000310000000000000023000000000000002e00000000",
            INIT_25 => X"0000001b00000000000000000000000000000030000000000000001500000000",
            INIT_26 => X"0000001c0000000000000027000000000000002e000000000000002d00000000",
            INIT_27 => X"0000003300000000000000240000000000000026000000000000000000000000",
            INIT_28 => X"0000001000000000000000270000000000000029000000000000002600000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"000000000000000000000000000000000000001c000000000000002a00000000",
            INIT_2B => X"0000000700000000000000060000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_2D => X"0000002700000000000000080000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000000000000d000000000000002c000000000000000d00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"000000000000000000000000000000000000001d000000000000001700000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000001300000000000000090000000000000000000000000000000b00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000006000000000000000a0000000000000014000000000000000800000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000800000000000000010000000000000000000000000000000400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000003000000000000000d00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_5C => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000380000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_60 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000001000000000000001d00000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_65 => X"0000000100000000000000000000000000000000000000000000000c00000000",
            INIT_66 => X"0000000100000000000000000000000000000000000000000000001300000000",
            INIT_67 => X"0000000b00000000000000000000000000000000000000000000001900000000",
            INIT_68 => X"000000080000000000000004000000000000000a000000000000000000000000",
            INIT_69 => X"0000000000000000000000400000000000000000000000000000000000000000",
            INIT_6A => X"0000000700000000000000070000000000000000000000000000003800000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000060000000000000006000000000000000000000000",
            INIT_6D => X"0000002600000000000000260000000000000007000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_71 => X"0000000000000000000000060000000000000026000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000040000000000000000000000000000000a00000000",
            INIT_75 => X"0000000000000000000000000000000000000007000000000000000500000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_78 => X"00000013000000000000000e0000000000000008000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_7A => X"0000001900000000000000000000000000000000000000000000000100000000",
            INIT_7B => X"0000000700000000000000000000000000000000000000000000000f00000000",
            INIT_7C => X"0000001c00000000000000120000000000000013000000000000000c00000000",
            INIT_7D => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_7E => X"00000008000000000000000c0000000000000000000000000000000000000000",
            INIT_7F => X"0000001100000000000000180000000000000009000000000000000500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE20;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21 : if BRAM_NAME = "samplegold_layersamples_instance21" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000170000000000000016000000000000001600000000",
            INIT_01 => X"0000000500000000000000020000000000000002000000000000000000000000",
            INIT_02 => X"00000014000000000000000e0000000000000000000000000000000000000000",
            INIT_03 => X"0000001b000000000000000f0000000000000012000000000000000b00000000",
            INIT_04 => X"00000002000000000000000a0000000000000015000000000000001100000000",
            INIT_05 => X"0000001000000000000000100000000000000007000000000000000a00000000",
            INIT_06 => X"0000003000000000000000000000000000000012000000000000000d00000000",
            INIT_07 => X"0000001200000000000000130000000000000014000000000000000f00000000",
            INIT_08 => X"0000001400000000000000120000000000000015000000000000001600000000",
            INIT_09 => X"0000001800000000000000150000000000000012000000000000001200000000",
            INIT_0A => X"0000001200000000000000290000000000000000000000000000001b00000000",
            INIT_0B => X"0000002d000000000000000e0000000000000014000000000000001000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000001c000000000000001d0000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000020000000000000014000000000000002900000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_68 => X"000000260000000000000042000000000000002d000000000000000500000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"00000011000000000000000f0000000000000000000000000000000000000000",
            INIT_6E => X"0000000d0000000000000020000000000000001b000000000000001600000000",
            INIT_6F => X"00000004000000000000001f0000000000000013000000000000000100000000",
            INIT_70 => X"0000001f00000000000000140000000000000001000000000000001100000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"00000014000000000000000f0000000000000009000000000000000600000000",
            INIT_74 => X"00000021000000000000001a000000000000001b000000000000001800000000",
            INIT_75 => X"0000000b000000000000000f0000000000000011000000000000000a00000000",
            INIT_76 => X"0000000000000000000000010000000000000006000000000000000400000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"000000350000000000000032000000000000000d000000000000000000000000",
            INIT_7D => X"0000002e0000000000000030000000000000002a000000000000002900000000",
            INIT_7E => X"0000002e000000000000002d000000000000002e000000000000002b00000000",
            INIT_7F => X"000000320000000000000033000000000000002c000000000000002e00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE21;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22 : if BRAM_NAME = "samplegold_layersamples_instance22" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003100000000000000390000000000000034000000000000002e00000000",
            INIT_01 => X"0000002800000000000000320000000000000042000000000000002300000000",
            INIT_02 => X"00000027000000000000002d000000000000002a000000000000003000000000",
            INIT_03 => X"0000003400000000000000340000000000000039000000000000002e00000000",
            INIT_04 => X"0000002600000000000000360000000000000036000000000000003400000000",
            INIT_05 => X"0000002b000000000000001b000000000000002a000000000000001d00000000",
            INIT_06 => X"0000002c00000000000000280000000000000021000000000000002000000000",
            INIT_07 => X"0000003500000000000000360000000000000033000000000000002800000000",
            INIT_08 => X"0000003d00000000000000450000000000000027000000000000003800000000",
            INIT_09 => X"00000043000000000000003c0000000000000034000000000000003b00000000",
            INIT_0A => X"0000004c0000000000000038000000000000003d000000000000003a00000000",
            INIT_0B => X"0000003800000000000000320000000000000037000000000000003700000000",
            INIT_0C => X"0000002800000000000000280000000000000026000000000000003500000000",
            INIT_0D => X"00000026000000000000002b0000000000000030000000000000002a00000000",
            INIT_0E => X"0000003300000000000000340000000000000036000000000000002900000000",
            INIT_0F => X"000000260000000000000031000000000000002e000000000000003500000000",
            INIT_10 => X"0000003900000000000000350000000000000034000000000000002e00000000",
            INIT_11 => X"0000003400000000000000330000000000000035000000000000003800000000",
            INIT_12 => X"0000003700000000000000330000000000000033000000000000003700000000",
            INIT_13 => X"0000002d000000000000001f0000000000000023000000000000002f00000000",
            INIT_14 => X"0000003a000000000000003a000000000000002f000000000000002a00000000",
            INIT_15 => X"0000003400000000000000360000000000000035000000000000003800000000",
            INIT_16 => X"0000003300000000000000350000000000000033000000000000003300000000",
            INIT_17 => X"0000001e000000000000000d000000000000002a000000000000003400000000",
            INIT_18 => X"0000003500000000000000300000000000000029000000000000003000000000",
            INIT_19 => X"0000003500000000000000340000000000000034000000000000003200000000",
            INIT_1A => X"0000003200000000000000320000000000000038000000000000003400000000",
            INIT_1B => X"0000001000000000000000000000000000000029000000000000003000000000",
            INIT_1C => X"00000023000000000000001e0000000000000022000000000000001800000000",
            INIT_1D => X"0000003300000000000000350000000000000037000000000000003200000000",
            INIT_1E => X"0000003200000000000000310000000000000030000000000000003700000000",
            INIT_1F => X"0000000c00000000000000080000000000000000000000000000002b00000000",
            INIT_20 => X"00000020000000000000000c000000000000000b000000000000000c00000000",
            INIT_21 => X"000000340000000000000024000000000000001a000000000000001900000000",
            INIT_22 => X"0000001900000000000000320000000000000033000000000000003300000000",
            INIT_23 => X"0000004500000000000000260000000000000014000000000000002d00000000",
            INIT_24 => X"0000002300000000000000260000000000000021000000000000002500000000",
            INIT_25 => X"0000001b000000000000003b0000000000000039000000000000004700000000",
            INIT_26 => X"0000001100000000000000120000000000000013000000000000001a00000000",
            INIT_27 => X"0000002200000000000000200000000000000014000000000000000a00000000",
            INIT_28 => X"0000002a00000000000000270000000000000026000000000000002300000000",
            INIT_29 => X"000000200000000000000017000000000000002e000000000000003000000000",
            INIT_2A => X"0000001100000000000000130000000000000015000000000000001d00000000",
            INIT_2B => X"000000160000000000000015000000000000001d000000000000001700000000",
            INIT_2C => X"0000001300000000000000170000000000000016000000000000001300000000",
            INIT_2D => X"00000009000000000000000b0000000000000003000000000000001300000000",
            INIT_2E => X"0000000700000000000000040000000000000000000000000000000600000000",
            INIT_2F => X"0000000200000000000000000000000000000003000000000000000600000000",
            INIT_30 => X"0000001500000000000000000000000000000000000000000000000100000000",
            INIT_31 => X"0000000300000000000000030000000000000004000000000000000000000000",
            INIT_32 => X"0000000600000000000000070000000000000009000000000000000000000000",
            INIT_33 => X"0000000000000000000000020000000000000005000000000000000300000000",
            INIT_34 => X"0000001d00000000000000000000000000000018000000000000000400000000",
            INIT_35 => X"0000003200000000000000410000000000000064000000000000004a00000000",
            INIT_36 => X"0000003f00000000000000390000000000000047000000000000004400000000",
            INIT_37 => X"0000003100000000000000400000000000000041000000000000003c00000000",
            INIT_38 => X"0000004500000000000000260000000000000048000000000000004200000000",
            INIT_39 => X"0000004100000000000000390000000000000070000000000000006200000000",
            INIT_3A => X"00000049000000000000004b0000000000000038000000000000004f00000000",
            INIT_3B => X"000000500000000000000044000000000000002d000000000000004800000000",
            INIT_3C => X"0000006700000000000000470000000000000027000000000000004b00000000",
            INIT_3D => X"0000004300000000000000370000000000000054000000000000005400000000",
            INIT_3E => X"00000042000000000000004b0000000000000040000000000000002a00000000",
            INIT_3F => X"0000004c00000000000000540000000000000035000000000000003b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000004200000000000000760000000000000044000000000000003100000000",
            INIT_41 => X"000000380000000000000049000000000000003c000000000000003b00000000",
            INIT_42 => X"0000004200000000000000370000000000000055000000000000003e00000000",
            INIT_43 => X"00000046000000000000004c000000000000004e000000000000001500000000",
            INIT_44 => X"0000004700000000000000700000000000000055000000000000004500000000",
            INIT_45 => X"0000004e00000000000000430000000000000040000000000000004500000000",
            INIT_46 => X"000000510000000000000029000000000000003f000000000000005200000000",
            INIT_47 => X"0000006000000000000000440000000000000050000000000000005000000000",
            INIT_48 => X"0000004e00000000000000530000000000000047000000000000005c00000000",
            INIT_49 => X"0000005200000000000000590000000000000054000000000000004b00000000",
            INIT_4A => X"0000005000000000000000520000000000000049000000000000004c00000000",
            INIT_4B => X"000000630000000000000065000000000000003a000000000000004a00000000",
            INIT_4C => X"0000004e00000000000000430000000000000023000000000000002f00000000",
            INIT_4D => X"00000053000000000000005d0000000000000057000000000000005600000000",
            INIT_4E => X"0000005000000000000000550000000000000055000000000000005900000000",
            INIT_4F => X"0000008400000000000000640000000000000053000000000000003300000000",
            INIT_50 => X"0000004d00000000000000230000000000000007000000000000004400000000",
            INIT_51 => X"000000540000000000000051000000000000005a000000000000005900000000",
            INIT_52 => X"00000033000000000000004f0000000000000055000000000000005300000000",
            INIT_53 => X"000000cd00000000000000620000000000000056000000000000004d00000000",
            INIT_54 => X"00000039000000000000001b0000000000000004000000000000001500000000",
            INIT_55 => X"000000560000000000000055000000000000003e000000000000004e00000000",
            INIT_56 => X"0000004d00000000000000310000000000000050000000000000005400000000",
            INIT_57 => X"0000001600000000000000d2000000000000007e000000000000005300000000",
            INIT_58 => X"0000002800000000000000160000000000000018000000000000000f00000000",
            INIT_59 => X"00000041000000000000003a0000000000000038000000000000000800000000",
            INIT_5A => X"000000500000000000000051000000000000002b000000000000004c00000000",
            INIT_5B => X"0000000000000000000000640000000000000043000000000000007800000000",
            INIT_5C => X"0000001300000000000000340000000000000039000000000000000000000000",
            INIT_5D => X"0000003d00000000000000280000000000000000000000000000001800000000",
            INIT_5E => X"0000006500000000000000680000000000000069000000000000003e00000000",
            INIT_5F => X"0000003c0000000000000059000000000000007a000000000000005e00000000",
            INIT_60 => X"0000005c00000000000000560000000000000060000000000000006100000000",
            INIT_61 => X"0000002900000000000000560000000000000058000000000000005500000000",
            INIT_62 => X"00000039000000000000003e0000000000000042000000000000003b00000000",
            INIT_63 => X"0000004e00000000000000340000000000000038000000000000003a00000000",
            INIT_64 => X"0000004400000000000000400000000000000046000000000000004300000000",
            INIT_65 => X"000000220000000000000025000000000000003f000000000000004e00000000",
            INIT_66 => X"0000001a00000000000000200000000000000019000000000000002800000000",
            INIT_67 => X"0000001c000000000000001f0000000000000018000000000000001a00000000",
            INIT_68 => X"0000000a00000000000000140000000000000017000000000000001400000000",
            INIT_69 => X"0000001800000000000000190000000000000022000000000000000000000000",
            INIT_6A => X"0000001600000000000000080000000000000016000000000000001300000000",
            INIT_6B => X"0000001700000000000000110000000000000013000000000000000800000000",
            INIT_6C => X"0000003b00000000000000050000000000000000000000000000001600000000",
            INIT_6D => X"0000000100000000000000090000000000000007000000000000000100000000",
            INIT_6E => X"0000000500000000000000060000000000000004000000000000000000000000",
            INIT_6F => X"0000000200000000000000080000000000000006000000000000000c00000000",
            INIT_70 => X"00000000000000000000000d0000000000000018000000000000000d00000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000031000000000000000d0000000000000000000000000000000000000000",
            INIT_76 => X"00000034000000000000002e0000000000000024000000000000001200000000",
            INIT_77 => X"0000000000000000000000000000000000000028000000000000002f00000000",
            INIT_78 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_79 => X"0000001200000000000000050000000000000006000000000000002000000000",
            INIT_7A => X"0000000000000000000000000000000000000001000000000000000900000000",
            INIT_7B => X"000000000000000000000000000000000000000f000000000000000600000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000800000000000000000000000000000000000000000000001400000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE22;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23 : if BRAM_NAME = "samplegold_layersamples_instance23" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000002b0000000000000027000000000000002c000000000000002e00000000",
            INIT_02 => X"0000000000000000000000180000000000000022000000000000002700000000",
            INIT_03 => X"0000000800000000000000020000000000000003000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_05 => X"0000000500000000000000050000000000000002000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000002100000000000000030000000000000001000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000014000000000000007e00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_0D => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"000000b7000000000000007e0000000000000000000000000000000000000000",
            INIT_14 => X"0000007400000000000000a3000000000000007d000000000000006700000000",
            INIT_15 => X"0000002f000000000000006d000000000000007500000000000000a300000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000700000000000000090000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000001000000000000000b00000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000000000000000000003b000000000000000000000000",
            INIT_22 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000001800000000000000130000000000000014000000000000001800000000",
            INIT_24 => X"0000004e00000000000000130000000000000004000000000000001000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000700000000000000000000000000000000000000000000000700000000",
            INIT_27 => X"0000000700000000000000050000000000000005000000000000000200000000",
            INIT_28 => X"0000000000000000000000050000000000000000000000000000000500000000",
            INIT_29 => X"0000004800000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"00000037000000000000003b0000000000000033000000000000004600000000",
            INIT_2B => X"0000002000000000000000300000000000000036000000000000003c00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000003900000000000000390000000000000000000000000000000000000000",
            INIT_2E => X"00000032000000000000003d000000000000004a000000000000003c00000000",
            INIT_2F => X"0000000000000000000000310000000000000031000000000000003900000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000002d0000000000000037000000000000005a000000000000000d00000000",
            INIT_32 => X"00000049000000000000003a000000000000003f000000000000003d00000000",
            INIT_33 => X"0000000000000000000000220000000000000037000000000000004100000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000000000000000000001a000000000000001d000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000002b000000000000001a000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"000000150000000000000012000000000000003f000000000000000200000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000001b00000000000000020000000000000006000000000000000000000000",
            INIT_48 => X"00000015000000000000000f0000000000000013000000000000002f00000000",
            INIT_49 => X"000000040000000000000006000000000000001e000000000000001a00000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000c00000000000000070000000000000000000000000000000100000000",
            INIT_4C => X"0000000f0000000000000000000000000000000c000000000000002300000000",
            INIT_4D => X"0000000000000000000000120000000000000006000000000000000f00000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_4F => X"0000000000000000000000000000000000000002000000000000000100000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000001200000000000000120000000000000015000000000000001f00000000",
            INIT_57 => X"0000001300000000000000130000000000000016000000000000001b00000000",
            INIT_58 => X"0000001200000000000000130000000000000015000000000000001500000000",
            INIT_59 => X"0000002000000000000000000000000000000008000000000000001100000000",
            INIT_5A => X"0000001500000000000000140000000000000011000000000000001100000000",
            INIT_5B => X"0000001600000000000000130000000000000015000000000000000d00000000",
            INIT_5C => X"0000000000000000000000180000000000000018000000000000001600000000",
            INIT_5D => X"0000000000000000000000110000000000000002000000000000000000000000",
            INIT_5E => X"0000000000000000000000060000000000000002000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_60 => X"00000005000000000000000b0000000000000000000000000000000000000000",
            INIT_61 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_62 => X"000000150000000000000026000000000000003f000000000000000000000000",
            INIT_63 => X"0000001b000000000000001b000000000000001e000000000000002e00000000",
            INIT_64 => X"0000000000000000000000000000000000000006000000000000002500000000",
            INIT_65 => X"0000001400000000000000000000000000000000000000000000000f00000000",
            INIT_66 => X"000000330000000000000026000000000000002d000000000000000c00000000",
            INIT_67 => X"00000022000000000000001c000000000000001c000000000000001d00000000",
            INIT_68 => X"0000000800000000000000000000000000000000000000000000001000000000",
            INIT_69 => X"0000002b00000000000000390000000000000000000000000000000000000000",
            INIT_6A => X"0000002b00000000000000330000000000000018000000000000002900000000",
            INIT_6B => X"0000004000000000000000210000000000000031000000000000001e00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_6F => X"0000000000000000000000020000000000000015000000000000000300000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000002000000000000002900000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000022000000000000003d00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_7C => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"00000002000000000000001c000000000000002e000000000000002300000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_7F => X"0000000000000000000000000000000000000009000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE23;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24 : if BRAM_NAME = "samplegold_layersamples_instance24" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d00000000000000140000000000000000000000000000000000000000",
            INIT_01 => X"000000340000000000000005000000000000000b000000000000001500000000",
            INIT_02 => X"0000000000000000000000050000000000000016000000000000002100000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_04 => X"0000004f000000000000000f0000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_06 => X"0000000f000000000000000c000000000000000e000000000000004800000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_0A => X"0000000700000000000000060000000000000007000000000000000300000000",
            INIT_0B => X"0000000000000000000000020000000000000001000000000000000200000000",
            INIT_0C => X"000000040000000000000000000000000000000e000000000000000700000000",
            INIT_0D => X"0000000000000000000000050000000000000007000000000000000100000000",
            INIT_0E => X"00000008000000000000000c0000000000000000000000000000000400000000",
            INIT_0F => X"0000000d00000000000000080000000000000003000000000000000b00000000",
            INIT_10 => X"0000000a00000000000000030000000000000005000000000000000c00000000",
            INIT_11 => X"0000001700000000000000080000000000000008000000000000000900000000",
            INIT_12 => X"0000000d000000000000000a0000000000000008000000000000000000000000",
            INIT_13 => X"0000000f00000000000000080000000000000010000000000000000700000000",
            INIT_14 => X"0000000300000000000000060000000000000007000000000000000400000000",
            INIT_15 => X"000000000000000000000000000000000000000e000000000000000f00000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000012000000000000000b0000000000000004000000000000000000000000",
            INIT_1B => X"0000000a000000000000000f0000000000000010000000000000001200000000",
            INIT_1C => X"0000000000000000000000000000000000000007000000000000000a00000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"00000000000000000000000b000000000000000a000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000f00000000000000060000000000000000000000000000000000000000",
            INIT_39 => X"0000001d00000000000000030000000000000000000000000000000300000000",
            INIT_3A => X"000000000000000000000000000000000000000b000000000000001f00000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"000000180000000000000014000000000000000f000000000000000200000000",
            INIT_47 => X"00000010000000000000000f000000000000000f000000000000001400000000",
            INIT_48 => X"000000050000000000000005000000000000000b000000000000000c00000000",
            INIT_49 => X"0000000000000000000000010000000000000000000000000000000400000000",
            INIT_4A => X"0000000000000000000000010000000000000006000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"00000024000000000000000d0000000000000000000000000000000000000000",
            INIT_53 => X"0000003f0000000000000038000000000000003d000000000000004200000000",
            INIT_54 => X"0000000a0000000000000033000000000000003f000000000000004000000000",
            INIT_55 => X"0000000000000000000000000000000000000003000000000000000600000000",
            INIT_56 => X"00000012000000000000001a000000000000003a000000000000000500000000",
            INIT_57 => X"000000100000000000000013000000000000001d000000000000001a00000000",
            INIT_58 => X"00000004000000000000001a0000000000000013000000000000001100000000",
            INIT_59 => X"0000000100000000000000000000000000000000000000000000000400000000",
            INIT_5A => X"0000000100000000000000010000000000000006000000000000000000000000",
            INIT_5B => X"0000000100000000000000040000000000000000000000000000000000000000",
            INIT_5C => X"0000000500000000000000040000000000000000000000000000000000000000",
            INIT_5D => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_5F => X"0000000100000000000000000000000000000006000000000000000b00000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000010000000000000030000000000000001300000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"000000170000000000000061000000000000002a000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000800000000000000070000000000000008000000000000000400000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_69 => X"0000004900000000000000450000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000060000000000000002000000000000000a00000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_6C => X"0000000400000000000000000000000000000001000000000000000000000000",
            INIT_6D => X"0000005a00000000000000090000000000000000000000000000000300000000",
            INIT_6E => X"0000000000000000000000130000000000000045000000000000007500000000",
            INIT_6F => X"0000000000000000000000010000000000000001000000000000000000000000",
            INIT_70 => X"00000034000000000000001a0000000000000003000000000000000500000000",
            INIT_71 => X"000000000000000000000005000000000000000e000000000000001300000000",
            INIT_72 => X"0000007400000000000000820000000000000047000000000000000c00000000",
            INIT_73 => X"0000000100000000000000010000000000000009000000000000003700000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"00000080000000000000007a000000000000006e000000000000000000000000",
            INIT_78 => X"00000070000000000000008b0000000000000084000000000000008300000000",
            INIT_79 => X"0000004800000000000000510000000000000057000000000000005200000000",
            INIT_7A => X"00000040000000000000003a0000000000000034000000000000004a00000000",
            INIT_7B => X"000000180000000000000010000000000000000c000000000000000c00000000",
            INIT_7C => X"000000270000000000000022000000000000001f000000000000001900000000",
            INIT_7D => X"0000003e000000000000003c000000000000003a000000000000003400000000",
            INIT_7E => X"0000000a000000000000003f0000000000000043000000000000004300000000",
            INIT_7F => X"000000040000000000000004000000000000000c000000000000000b00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE24;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25 : if BRAM_NAME = "samplegold_layersamples_instance25" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000200000000000000000000000000000002000000000000000300000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"000000bc00000000000000d500000000000000c0000000000000000d00000000",
            INIT_07 => X"000000bb00000000000000c000000000000000b300000000000000a700000000",
            INIT_08 => X"000000bc00000000000000b900000000000000b500000000000000b800000000",
            INIT_09 => X"000000d400000000000000cb00000000000000bf00000000000000ba00000000",
            INIT_0A => X"0000008500000000000000e000000000000000e100000000000000c500000000",
            INIT_0B => X"0000008d000000000000008e0000000000000092000000000000008a00000000",
            INIT_0C => X"0000009e00000000000000960000000000000098000000000000009100000000",
            INIT_0D => X"000000c300000000000000db00000000000000df00000000000000d200000000",
            INIT_0E => X"00000081000000000000007400000000000000e000000000000000de00000000",
            INIT_0F => X"0000007e000000000000006c0000000000000065000000000000007300000000",
            INIT_10 => X"000000c000000000000000840000000000000081000000000000008300000000",
            INIT_11 => X"000000db00000000000000be00000000000000e400000000000000e200000000",
            INIT_12 => X"000000940000000000000090000000000000007200000000000000cd00000000",
            INIT_13 => X"000000990000000000000097000000000000008d000000000000008e00000000",
            INIT_14 => X"000000e2000000000000009e00000000000000a2000000000000009500000000",
            INIT_15 => X"000000d800000000000000d800000000000000c700000000000000e300000000",
            INIT_16 => X"000000b400000000000000b200000000000000b100000000000000c000000000",
            INIT_17 => X"000000b000000000000000b800000000000000ba00000000000000b500000000",
            INIT_18 => X"000000df00000000000000dc00000000000000cb00000000000000cc00000000",
            INIT_19 => X"000000d600000000000000cf00000000000000d600000000000000d600000000",
            INIT_1A => X"000000ca00000000000000c500000000000000c300000000000000c300000000",
            INIT_1B => X"000000cc00000000000000c600000000000000c500000000000000c600000000",
            INIT_1C => X"000000db00000000000000de00000000000000dd00000000000000df00000000",
            INIT_1D => X"000000d20000000000000098000000000000008b00000000000000c500000000",
            INIT_1E => X"000000de00000000000000e100000000000000dd00000000000000dd00000000",
            INIT_1F => X"000000de00000000000000dd00000000000000da00000000000000da00000000",
            INIT_20 => X"000000e700000000000000e100000000000000e300000000000000e000000000",
            INIT_21 => X"0000009f0000000000000049000000000000007d00000000000000d700000000",
            INIT_22 => X"000000dc00000000000000df00000000000000e200000000000000da00000000",
            INIT_23 => X"000000db00000000000000db00000000000000da00000000000000d900000000",
            INIT_24 => X"000000e600000000000000e900000000000000e100000000000000de00000000",
            INIT_25 => X"0000005d000000000000003c000000000000006400000000000000de00000000",
            INIT_26 => X"000000d800000000000000d400000000000000ce00000000000000a900000000",
            INIT_27 => X"000000df00000000000000dc00000000000000da00000000000000d800000000",
            INIT_28 => X"000000dd00000000000000e700000000000000e300000000000000e100000000",
            INIT_29 => X"0000003700000000000000350000000000000029000000000000007500000000",
            INIT_2A => X"000000bf000000000000008b000000000000005f000000000000003e00000000",
            INIT_2B => X"000000e100000000000000da00000000000000d800000000000000d300000000",
            INIT_2C => X"0000007f00000000000000d100000000000000e400000000000000de00000000",
            INIT_2D => X"000000650000000000000053000000000000002a000000000000002c00000000",
            INIT_2E => X"0000007300000000000000350000000000000040000000000000004300000000",
            INIT_2F => X"000000d000000000000000ce00000000000000ca00000000000000a300000000",
            INIT_30 => X"000000c600000000000000cc00000000000000cd00000000000000cf00000000",
            INIT_31 => X"000000ba00000000000000cb00000000000000ae00000000000000a300000000",
            INIT_32 => X"000000c900000000000000b800000000000000bc00000000000000b900000000",
            INIT_33 => X"00000064000000000000006b000000000000006b00000000000000c800000000",
            INIT_34 => X"0000005800000000000000580000000000000057000000000000005d00000000",
            INIT_35 => X"0000007000000000000000700000000000000071000000000000006500000000",
            INIT_36 => X"00000070000000000000007b000000000000007b000000000000007400000000",
            INIT_37 => X"0000003d00000000000000480000000000000049000000000000004600000000",
            INIT_38 => X"0000003300000000000000330000000000000035000000000000003700000000",
            INIT_39 => X"0000002500000000000000270000000000000028000000000000003300000000",
            INIT_3A => X"0000002400000000000000400000000000000026000000000000002200000000",
            INIT_3B => X"0000002100000000000000210000000000000024000000000000002300000000",
            INIT_3C => X"000000220000000000000020000000000000001e000000000000002300000000",
            INIT_3D => X"0000002d000000000000001d000000000000001c000000000000001e00000000",
            INIT_3E => X"0000000000000000000000000000000000000053000000000000005000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000002000000000000000180000000000000017000000000000002900000000",
            INIT_44 => X"000000160000000000000014000000000000001a000000000000001300000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_46 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000600000000000000000000000000000007000000000000000000000000",
            INIT_4F => X"0000000100000000000000030000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000001c000000000000000b0000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000007400000000000000150000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000004c00000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000003800000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"00000007000000000000002d0000000000000000000000000000000000000000",
            INIT_5E => X"00000008000000000000002a0000000000000061000000000000004d00000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"00000000000000000000001e000000000000004f000000000000002000000000",
            INIT_62 => X"0000007c00000000000000700000000000000024000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000021000000000000005f00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000003f00000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"00000063000000000000005f000000000000005c000000000000005200000000",
            INIT_69 => X"00000048000000000000002b000000000000001f000000000000003c00000000",
            INIT_6A => X"00000030000000000000000d000000000000002a000000000000001a00000000",
            INIT_6B => X"0000000000000000000000000000000000000031000000000000003b00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"00000020000000000000001e0000000000000010000000000000000000000000",
            INIT_6E => X"00000034000000000000002f000000000000002d000000000000002800000000",
            INIT_6F => X"000000290000000000000032000000000000003a000000000000003900000000",
            INIT_70 => X"00000017000000000000001e0000000000000020000000000000001c00000000",
            INIT_71 => X"00000005000000000000000c000000000000000a000000000000001200000000",
            INIT_72 => X"0000000000000000000000000000000000000003000000000000000300000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000036000000000000003e0000000000000000000000000000000000000000",
            INIT_77 => X"0000002700000000000000170000000000000013000000000000002b00000000",
            INIT_78 => X"00000019000000000000001c0000000000000018000000000000001d00000000",
            INIT_79 => X"0000001d0000000000000019000000000000001b000000000000001c00000000",
            INIT_7A => X"0000003b000000000000003b0000000000000017000000000000001600000000",
            INIT_7B => X"0000000500000000000000070000000000000000000000000000001a00000000",
            INIT_7C => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_7D => X"0000001c000000000000001f0000000000000013000000000000000200000000",
            INIT_7E => X"0000001b0000000000000039000000000000003c000000000000001d00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE25;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26 : if BRAM_NAME = "samplegold_layersamples_instance26" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000020000000000000001e0000000000000022000000000000000000000000",
            INIT_02 => X"00000000000000000000000b0000000000000037000000000000003600000000",
            INIT_03 => X"0000000800000000000000000000000000000009000000000000000600000000",
            INIT_04 => X"0000000600000000000000090000000000000000000000000000000d00000000",
            INIT_05 => X"0000002a00000000000000260000000000000024000000000000002600000000",
            INIT_06 => X"0000002500000000000000120000000000000027000000000000003700000000",
            INIT_07 => X"0000002300000000000000230000000000000026000000000000002700000000",
            INIT_08 => X"0000001c000000000000002c0000000000000022000000000000001a00000000",
            INIT_09 => X"0000002400000000000000240000000000000027000000000000002200000000",
            INIT_0A => X"0000001b00000000000000190000000000000024000000000000002a00000000",
            INIT_0B => X"0000001700000000000000160000000000000017000000000000001c00000000",
            INIT_0C => X"0000002100000000000000240000000000000026000000000000001800000000",
            INIT_0D => X"0000000b00000000000000100000000000000025000000000000002600000000",
            INIT_0E => X"00000026000000000000002e000000000000004a000000000000003e00000000",
            INIT_0F => X"00000021000000000000001b000000000000001e000000000000002200000000",
            INIT_10 => X"0000002700000000000000230000000000000022000000000000001f00000000",
            INIT_11 => X"0000000000000000000000000000000000000022000000000000002b00000000",
            INIT_12 => X"00000022000000000000003f0000000000000052000000000000001200000000",
            INIT_13 => X"0000001f000000000000001e000000000000001a000000000000001c00000000",
            INIT_14 => X"0000002700000000000000290000000000000020000000000000002100000000",
            INIT_15 => X"0000000000000000000000020000000000000017000000000000001d00000000",
            INIT_16 => X"000000350000000000000046000000000000003d000000000000001d00000000",
            INIT_17 => X"00000020000000000000001e000000000000002a000000000000002600000000",
            INIT_18 => X"0000001800000000000000230000000000000028000000000000002200000000",
            INIT_19 => X"0000001b00000000000000000000000000000007000000000000001800000000",
            INIT_1A => X"00000032000000000000001e000000000000000f000000000000001700000000",
            INIT_1B => X"0000002900000000000000350000000000000041000000000000005b00000000",
            INIT_1C => X"0000001b0000000000000019000000000000002b000000000000002500000000",
            INIT_1D => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000300000000000000000000000000000000000000000000002600000000",
            INIT_1F => X"0000002800000000000000200000000000000036000000000000000300000000",
            INIT_20 => X"0000002800000000000000250000000000000025000000000000003200000000",
            INIT_21 => X"00000039000000000000001d0000000000000011000000000000002e00000000",
            INIT_22 => X"00000024000000000000002c0000000000000027000000000000002d00000000",
            INIT_23 => X"0000001a00000000000000350000000000000038000000000000003100000000",
            INIT_24 => X"0000001400000000000000120000000000000014000000000000001a00000000",
            INIT_25 => X"00000023000000000000002a000000000000001a000000000000001200000000",
            INIT_26 => X"000000340000000000000033000000000000002c000000000000002b00000000",
            INIT_27 => X"0000002200000000000000160000000000000039000000000000002f00000000",
            INIT_28 => X"000000170000000000000011000000000000001c000000000000001e00000000",
            INIT_29 => X"0000000e00000000000000110000000000000018000000000000001800000000",
            INIT_2A => X"0000001600000000000000110000000000000011000000000000001200000000",
            INIT_2B => X"0000000f00000000000000110000000000000003000000000000002500000000",
            INIT_2C => X"000000090000000000000010000000000000000b000000000000000f00000000",
            INIT_2D => X"0000000600000000000000070000000000000006000000000000000c00000000",
            INIT_2E => X"000000100000000000000020000000000000001e000000000000000700000000",
            INIT_2F => X"0000000b00000000000000000000000000000015000000000000003400000000",
            INIT_30 => X"0000000d0000000000000008000000000000000d000000000000001800000000",
            INIT_31 => X"00000009000000000000000d000000000000000d000000000000000c00000000",
            INIT_32 => X"000000310000000000000015000000000000001b000000000000001700000000",
            INIT_33 => X"0000000e00000000000000000000000000000001000000000000001c00000000",
            INIT_34 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_35 => X"0000001d00000000000000040000000000000000000000000000000000000000",
            INIT_36 => X"0000001a000000000000002f000000000000000e000000000000000c00000000",
            INIT_37 => X"0000001b00000000000000000000000000000000000000000000000500000000",
            INIT_38 => X"00000010000000000000000f0000000000000019000000000000000000000000",
            INIT_39 => X"000000120000000000000021000000000000001c000000000000001700000000",
            INIT_3A => X"0000000000000000000000180000000000000029000000000000001100000000",
            INIT_3B => X"0000000000000000000000020000000000000003000000000000000000000000",
            INIT_3C => X"0000000500000000000000000000000000000000000000000000000600000000",
            INIT_3D => X"0000000f000000000000000f000000000000001f000000000000000500000000",
            INIT_3E => X"00000000000000000000000b000000000000001a000000000000001e00000000",
            INIT_3F => X"0000000e00000000000000080000000000000008000000000000000b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002300000000000000100000000000000001000000000000000700000000",
            INIT_41 => X"0000001f000000000000000d0000000000000010000000000000000e00000000",
            INIT_42 => X"0000001300000000000000150000000000000001000000000000000e00000000",
            INIT_43 => X"0000000d00000000000000110000000000000019000000000000001500000000",
            INIT_44 => X"0000000d000000000000001d0000000000000017000000000000001300000000",
            INIT_45 => X"0000000000000000000000250000000000000011000000000000000d00000000",
            INIT_46 => X"0000001a000000000000001f000000000000000d000000000000000000000000",
            INIT_47 => X"00000008000000000000000a000000000000000b000000000000000f00000000",
            INIT_48 => X"0000000c000000000000000d000000000000000b000000000000000f00000000",
            INIT_49 => X"000000000000000000000010000000000000002f000000000000000c00000000",
            INIT_4A => X"0000002d000000000000003c0000000000000000000000000000000000000000",
            INIT_4B => X"0000000d00000000000000030000000000000005000000000000001200000000",
            INIT_4C => X"0000000e000000000000000a000000000000000e000000000000000b00000000",
            INIT_4D => X"00000000000000000000000d0000000000000016000000000000003400000000",
            INIT_4E => X"0000001f000000000000002e0000000000000026000000000000000000000000",
            INIT_4F => X"0000000900000000000000140000000000000012000000000000001900000000",
            INIT_50 => X"00000032000000000000000c000000000000000b000000000000000900000000",
            INIT_51 => X"000000000000000000000002000000000000000d000000000000001300000000",
            INIT_52 => X"0000001b000000000000001c000000000000001f000000000000000c00000000",
            INIT_53 => X"0000001d0000000000000015000000000000001b000000000000000100000000",
            INIT_54 => X"0000000d00000000000000310000000000000010000000000000001900000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_56 => X"0000000000000000000000210000000000000053000000000000001e00000000",
            INIT_57 => X"0000002b00000000000000620000000000000011000000000000002d00000000",
            INIT_58 => X"0000000000000000000000000000000000000020000000000000001800000000",
            INIT_59 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000800000000000000000000000000000000000000000000002600000000",
            INIT_5B => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_5C => X"00000010000000000000000b000000000000000b000000000000001400000000",
            INIT_5D => X"0000001d00000000000000170000000000000012000000000000001800000000",
            INIT_5E => X"0000000d0000000000000008000000000000000c000000000000000500000000",
            INIT_5F => X"0000000000000000000000040000000000000001000000000000000a00000000",
            INIT_60 => X"00000008000000000000000c0000000000000004000000000000000600000000",
            INIT_61 => X"0000001200000000000000140000000000000010000000000000000b00000000",
            INIT_62 => X"0000001800000000000000180000000000000018000000000000001100000000",
            INIT_63 => X"0000001400000000000000020000000000000045000000000000001c00000000",
            INIT_64 => X"000000200000000000000014000000000000001b000000000000001500000000",
            INIT_65 => X"0000001a00000000000000160000000000000021000000000000001800000000",
            INIT_66 => X"0000004d000000000000002d000000000000001d000000000000001800000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE26;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27 : if BRAM_NAME = "samplegold_layersamples_instance27" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000005100000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000005400000000000000640000000000000048000000000000005e00000000",
            INIT_0F => X"0000003b00000000000000490000000000000065000000000000005100000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000200000000000000030000000000000003000000000000000000000000",
            INIT_1E => X"0000000500000000000000000000000000000000000000000000000700000000",
            INIT_1F => X"0000000e00000000000000070000000000000000000000000000002400000000",
            INIT_20 => X"00000011000000000000000e0000000000000011000000000000001000000000",
            INIT_21 => X"000000120000000000000013000000000000000d000000000000001400000000",
            INIT_22 => X"0000001e00000000000000110000000000000013000000000000001400000000",
            INIT_23 => X"0000000c00000000000000050000000000000001000000000000001c00000000",
            INIT_24 => X"0000002a00000000000000280000000000000027000000000000003000000000",
            INIT_25 => X"00000027000000000000002d000000000000002f000000000000002600000000",
            INIT_26 => X"0000001b000000000000001a000000000000001e000000000000001a00000000",
            INIT_27 => X"0000002500000000000000160000000000000003000000000000000000000000",
            INIT_28 => X"0000003400000000000000380000000000000030000000000000003500000000",
            INIT_29 => X"000000380000000000000037000000000000003a000000000000003300000000",
            INIT_2A => X"0000000100000000000000190000000000000019000000000000001f00000000",
            INIT_2B => X"0000001e000000000000002a0000000000000018000000000000000200000000",
            INIT_2C => X"0000001e00000000000000260000000000000021000000000000001900000000",
            INIT_2D => X"0000001600000000000000220000000000000020000000000000002400000000",
            INIT_2E => X"00000004000000000000000a0000000000000014000000000000001200000000",
            INIT_2F => X"00000007000000000000000a000000000000001c000000000000000700000000",
            INIT_30 => X"0000000d000000000000000d000000000000000e000000000000000400000000",
            INIT_31 => X"00000015000000000000001d0000000000000007000000000000000f00000000",
            INIT_32 => X"000000060000000000000010000000000000000f000000000000001200000000",
            INIT_33 => X"0000001400000000000000100000000000000013000000000000000700000000",
            INIT_34 => X"0000001500000000000000130000000000000015000000000000001800000000",
            INIT_35 => X"0000001200000000000000140000000000000012000000000000001600000000",
            INIT_36 => X"00000000000000000000000d000000000000000d000000000000001400000000",
            INIT_37 => X"000000160000000000000013000000000000000c000000000000000000000000",
            INIT_38 => X"0000001500000000000000150000000000000018000000000000001600000000",
            INIT_39 => X"0000001500000000000000140000000000000015000000000000001500000000",
            INIT_3A => X"0000000b00000000000000250000000000000013000000000000001400000000",
            INIT_3B => X"0000001b00000000000000190000000000000000000000000000000000000000",
            INIT_3C => X"0000001400000000000000150000000000000016000000000000001600000000",
            INIT_3D => X"0000001b00000000000000180000000000000010000000000000001300000000",
            INIT_3E => X"00000000000000000000001d000000000000001d000000000000001e00000000",
            INIT_3F => X"0000001200000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001200000000000000160000000000000018000000000000000f00000000",
            INIT_41 => X"0000001f000000000000001f000000000000001b000000000000001100000000",
            INIT_42 => X"0000000000000000000000000000000000000010000000000000002e00000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"00000016000000000000000d0000000000000000000000000000000000000000",
            INIT_45 => X"0000001f000000000000001c000000000000001d000000000000001a00000000",
            INIT_46 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_48 => X"0000000c0000000000000010000000000000001a000000000000000000000000",
            INIT_49 => X"00000008000000000000000b000000000000000e000000000000001000000000",
            INIT_4A => X"00000007000000000000000c0000000000000005000000000000000000000000",
            INIT_4B => X"0000000f00000000000000010000000000000008000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000002400000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000003900000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000006300000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000c000000000000004f0000000000000007000000000000000000000000",
            INIT_7B => X"0000000d000000000000000e0000000000000001000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"00000010000000000000004c0000000000000000000000000000000200000000",
            INIT_7F => X"0000000f000000000000002a0000000000000017000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE27;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28 : if BRAM_NAME = "samplegold_layersamples_instance28" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000500000000000000030000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000300000000000000140000000000000000000000000000000000000000",
            INIT_09 => X"0000000f00000000000000130000000000000005000000000000000500000000",
            INIT_0A => X"0000001a0000000000000013000000000000000c000000000000000c00000000",
            INIT_0B => X"0000000f00000000000000140000000000000016000000000000001400000000",
            INIT_0C => X"000000120000000000000014000000000000001d000000000000000600000000",
            INIT_0D => X"00000017000000000000000b0000000000000016000000000000001400000000",
            INIT_0E => X"0000001e0000000000000019000000000000001b000000000000001100000000",
            INIT_0F => X"0000003e000000000000001c0000000000000009000000000000001d00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_12 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_14 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_16 => X"0000002c0000000000000000000000000000000e000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_1B => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_1D => X"0000000000000000000000150000000000000000000000000000003200000000",
            INIT_1E => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_1F => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_21 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000001f0000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000400000000000000000000000000000008000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000003000000000000002300000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000700000000000000000000000000000006000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000030000000000000002000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000070000000000000007000000000000000a000000000000000000000000",
            INIT_42 => X"0000000000000000000000210000000000000011000000000000000800000000",
            INIT_43 => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"000000090000000000000009000000000000002b000000000000000000000000",
            INIT_45 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000010000000000000000400000000",
            INIT_47 => X"0000000d000000000000000d0000000000000017000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000090000000000000005000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000020000000000000004000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000000d000000000000001b000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_7D => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE28;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29 : if BRAM_NAME = "samplegold_layersamples_instance29" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_07 => X"00000000000000000000000c0000000000000000000000000000001100000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_0D => X"0000001200000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_0F => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_11 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_14 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_17 => X"0000000000000000000000020000000000000008000000000000000000000000",
            INIT_18 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000a00000000000000060000000000000006000000000000000500000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000007000000000000000200000000",
            INIT_1C => X"00000000000000000000000d0000000000000005000000000000000200000000",
            INIT_1D => X"00000002000000000000000f0000000000000013000000000000000b00000000",
            INIT_1E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_20 => X"0000000b000000000000000b0000000000000008000000000000001400000000",
            INIT_21 => X"000000000000000000000005000000000000000d000000000000000500000000",
            INIT_22 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_23 => X"0000000a00000000000000150000000000000000000000000000000000000000",
            INIT_24 => X"0000000900000000000000080000000000000014000000000000001400000000",
            INIT_25 => X"0000000500000000000000000000000000000000000000000000000400000000",
            INIT_26 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_27 => X"0000000f00000000000000220000000000000000000000000000000700000000",
            INIT_28 => X"000000040000000000000008000000000000000c000000000000000c00000000",
            INIT_29 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_2B => X"00000010000000000000000e000000000000000d000000000000000b00000000",
            INIT_2C => X"000000000000000000000007000000000000000f000000000000000700000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000c00000000000000060000000000000000000000000000000100000000",
            INIT_30 => X"0000000000000000000000000000000000000001000000000000000f00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"00000009000000000000000c0000000000000014000000000000000000000000",
            INIT_34 => X"0000000000000000000000030000000000000000000000000000000100000000",
            INIT_35 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_38 => X"0000001b00000000000000140000000000000000000000000000000000000000",
            INIT_39 => X"0000005200000000000000080000000000000000000000000000001500000000",
            INIT_3A => X"0000000f00000000000000000000000000000018000000000000000000000000",
            INIT_3B => X"000000910000000000000000000000000000003e000000000000000000000000",
            INIT_3C => X"0000001000000000000000100000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000004e000000000000000d000000000000001b00000000",
            INIT_3E => X"00000000000000000000001d0000000000000000000000000000000800000000",
            INIT_3F => X"00000000000000000000007c0000000000000000000000000000003f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000e000000000000000c0000000000000033000000000000002b00000000",
            INIT_41 => X"0000000000000000000000000000000000000039000000000000001e00000000",
            INIT_42 => X"00000000000000000000003d0000000000000000000000000000002200000000",
            INIT_43 => X"00000031000000000000000c0000000000000060000000000000000000000000",
            INIT_44 => X"00000029000000000000002f0000000000000000000000000000003300000000",
            INIT_45 => X"00000025000000000000002c0000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000025000000000000000000000000",
            INIT_47 => X"000000300000000000000084000000000000001b000000000000004600000000",
            INIT_48 => X"00000000000000000000002d000000000000005d000000000000000000000000",
            INIT_49 => X"0000000800000000000000000000000000000056000000000000000600000000",
            INIT_4A => X"000000290000000000000000000000000000001d000000000000000000000000",
            INIT_4B => X"00000000000000000000004700000000000000ab000000000000002500000000",
            INIT_4C => X"000000030000000000000000000000000000004c000000000000002000000000",
            INIT_4D => X"00000009000000000000001a0000000000000000000000000000002b00000000",
            INIT_4E => X"0000001500000000000000410000000000000000000000000000001f00000000",
            INIT_4F => X"000000000000000000000000000000000000003800000000000000a900000000",
            INIT_50 => X"0000001100000000000000100000000000000030000000000000003300000000",
            INIT_51 => X"0000001000000000000000140000000000000019000000000000000e00000000",
            INIT_52 => X"000000840000000000000006000000000000002a000000000000000400000000",
            INIT_53 => X"0000002a00000000000000000000000000000000000000000000002b00000000",
            INIT_54 => X"0000001a00000000000000000000000000000022000000000000002000000000",
            INIT_55 => X"000000030000000000000018000000000000000e000000000000001f00000000",
            INIT_56 => X"0000000100000000000000730000000000000016000000000000005000000000",
            INIT_57 => X"000000060000000000000017000000000000001d000000000000000400000000",
            INIT_58 => X"0000001d00000000000000200000000000000008000000000000004800000000",
            INIT_59 => X"0000005200000000000000170000000000000027000000000000001700000000",
            INIT_5A => X"000000270000000000000021000000000000004a000000000000003200000000",
            INIT_5B => X"0000000000000000000000160000000000000004000000000000002d00000000",
            INIT_5C => X"0000003b0000000000000025000000000000001c000000000000002200000000",
            INIT_5D => X"0000001900000000000000520000000000000032000000000000001f00000000",
            INIT_5E => X"000000320000000000000000000000000000005c000000000000000000000000",
            INIT_5F => X"00000000000000000000001e0000000000000007000000000000000000000000",
            INIT_60 => X"0000002400000000000000400000000000000038000000000000003400000000",
            INIT_61 => X"0000001800000000000000030000000000000036000000000000002900000000",
            INIT_62 => X"0000000000000000000000410000000000000005000000000000000000000000",
            INIT_63 => X"0000002700000000000000070000000000000000000000000000002f00000000",
            INIT_64 => X"00000031000000000000001c0000000000000046000000000000002c00000000",
            INIT_65 => X"0000001700000000000000170000000000000000000000000000003700000000",
            INIT_66 => X"000000260000000000000028000000000000002e000000000000000000000000",
            INIT_67 => X"0000000000000000000000590000000000000022000000000000000000000000",
            INIT_68 => X"00000049000000000000003c0000000000000029000000000000002a00000000",
            INIT_69 => X"000000000000000000000045000000000000001e000000000000000000000000",
            INIT_6A => X"0000001000000000000000350000000000000008000000000000000000000000",
            INIT_6B => X"0000001f00000000000000000000000000000020000000000000000b00000000",
            INIT_6C => X"0000000000000000000000670000000000000049000000000000002100000000",
            INIT_6D => X"000000000000000000000019000000000000005a000000000000000000000000",
            INIT_6E => X"0000001e00000000000000230000000000000015000000000000000000000000",
            INIT_6F => X"0000003200000000000000220000000000000025000000000000000800000000",
            INIT_70 => X"0000000000000000000000000000000000000025000000000000002500000000",
            INIT_71 => X"0000000a00000000000000390000000000000018000000000000001c00000000",
            INIT_72 => X"00000000000000000000000d000000000000001b000000000000000000000000",
            INIT_73 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000a00000000000000120000000000000000000000000000000500000000",
            INIT_75 => X"00000000000000000000000a0000000000000003000000000000003100000000",
            INIT_76 => X"0000000c00000000000000140000000000000000000000000000000000000000",
            INIT_77 => X"0000001900000000000000110000000000000000000000000000001500000000",
            INIT_78 => X"0000000000000000000000000000000000000021000000000000005800000000",
            INIT_79 => X"0000003400000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000013000000000000005200000000",
            INIT_7B => X"00000017000000000000001f0000000000000017000000000000000000000000",
            INIT_7C => X"0000001e00000000000000390000000000000000000000000000001500000000",
            INIT_7D => X"00000000000000000000004c0000000000000017000000000000000100000000",
            INIT_7E => X"000000460000000000000007000000000000001e000000000000000000000000",
            INIT_7F => X"00000000000000000000000e0000000000000000000000000000002800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE29;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30 : if BRAM_NAME = "samplegold_layersamples_instance30" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000250000000000000012000000000000000700000000",
            INIT_01 => X"0000004e0000000000000000000000000000000d000000000000002b00000000",
            INIT_02 => X"0000000000000000000000110000000000000040000000000000002a00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000004800000000000000420000000000000000000000000000000000000000",
            INIT_05 => X"0000001e000000000000003b0000000000000019000000000000000000000000",
            INIT_06 => X"0000000000000000000000370000000000000000000000000000000000000000",
            INIT_07 => X"0000001400000000000000250000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_09 => X"000000000000000000000000000000000000000c000000000000002300000000",
            INIT_0A => X"000000100000000000000000000000000000001b000000000000001000000000",
            INIT_0B => X"0000001300000000000000020000000000000000000000000000000000000000",
            INIT_0C => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_0D => X"0000001f000000000000003a0000000000000019000000000000001000000000",
            INIT_0E => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000023000000000000001d00000000",
            INIT_10 => X"0000000000000000000000110000000000000032000000000000000000000000",
            INIT_11 => X"0000000900000000000000000000000000000000000000000000001700000000",
            INIT_12 => X"00000012000000000000000a0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000100000000000000250000000000000005000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000001000000000000000a00000000",
            INIT_16 => X"000000130000000000000000000000000000000a000000000000001600000000",
            INIT_17 => X"0000000b00000000000000150000000000000005000000000000000d00000000",
            INIT_18 => X"00000000000000000000000e0000000000000003000000000000000200000000",
            INIT_19 => X"0000000b00000000000000110000000000000000000000000000000000000000",
            INIT_1A => X"0000005700000000000000950000000000000037000000000000003d00000000",
            INIT_1B => X"0000000100000000000000000000000000000000000000000000002600000000",
            INIT_1C => X"0000001400000000000000010000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000110000000000000000000000000000000600000000",
            INIT_1E => X"0000003b00000000000000130000000000000000000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000d000000000000001400000000",
            INIT_20 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_22 => X"0000003600000000000000010000000000000000000000000000000000000000",
            INIT_23 => X"0000002d00000000000000190000000000000000000000000000002100000000",
            INIT_24 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_25 => X"0000001900000000000000000000000000000000000000000000001800000000",
            INIT_26 => X"0000003b00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000004000000000000003300000000",
            INIT_28 => X"0000002e000000000000003e0000000000000000000000000000000000000000",
            INIT_29 => X"00000007000000000000000c000000000000000f000000000000004f00000000",
            INIT_2A => X"0000001000000000000000000000000000000011000000000000000000000000",
            INIT_2B => X"0000001e00000000000000080000000000000018000000000000000000000000",
            INIT_2C => X"0000000d0000000000000002000000000000004c000000000000000000000000",
            INIT_2D => X"0000000000000000000000070000000000000014000000000000000200000000",
            INIT_2E => X"0000000300000000000000030000000000000002000000000000001500000000",
            INIT_2F => X"0000000000000000000000190000000000000009000000000000000d00000000",
            INIT_30 => X"0000001f00000000000000110000000000000005000000000000003800000000",
            INIT_31 => X"0000001000000000000000030000000000000003000000000000000700000000",
            INIT_32 => X"0000000000000000000000190000000000000006000000000000000000000000",
            INIT_33 => X"0000003200000000000000000000000000000000000000000000002500000000",
            INIT_34 => X"00000000000000000000000b0000000000000016000000000000000a00000000",
            INIT_35 => X"000000090000000000000001000000000000000f000000000000002200000000",
            INIT_36 => X"00000006000000000000000a000000000000000c000000000000002700000000",
            INIT_37 => X"0000000d000000000000001f0000000000000015000000000000000c00000000",
            INIT_38 => X"000000170000000000000000000000000000000e000000000000003000000000",
            INIT_39 => X"0000002e00000000000000110000000000000000000000000000002600000000",
            INIT_3A => X"000000240000000000000015000000000000000b000000000000000200000000",
            INIT_3B => X"00000031000000000000000a0000000000000025000000000000000700000000",
            INIT_3C => X"0000001100000000000000000000000000000000000000000000001b00000000",
            INIT_3D => X"000000090000000000000033000000000000002e000000000000001800000000",
            INIT_3E => X"00000015000000000000002b0000000000000027000000000000002300000000",
            INIT_3F => X"00000018000000000000003c0000000000000000000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000003e00000000000000150000000000000000000000000000000000000000",
            INIT_41 => X"0000004400000000000000460000000000000046000000000000004600000000",
            INIT_42 => X"0000002d000000000000003c0000000000000035000000000000003f00000000",
            INIT_43 => X"0000000000000000000000110000000000000026000000000000000600000000",
            INIT_44 => X"0000005300000000000000310000000000000015000000000000000900000000",
            INIT_45 => X"0000004c00000000000000430000000000000052000000000000003e00000000",
            INIT_46 => X"00000014000000000000004c000000000000002d000000000000005300000000",
            INIT_47 => X"00000009000000000000000b0000000000000001000000000000002a00000000",
            INIT_48 => X"0000004100000000000000380000000000000028000000000000000200000000",
            INIT_49 => X"0000005000000000000000510000000000000052000000000000004000000000",
            INIT_4A => X"00000014000000000000001b0000000000000044000000000000004700000000",
            INIT_4B => X"0000000b000000000000001b000000000000000a000000000000001200000000",
            INIT_4C => X"0000003f00000000000000320000000000000025000000000000000f00000000",
            INIT_4D => X"0000004f0000000000000045000000000000004c000000000000004700000000",
            INIT_4E => X"0000001e0000000000000000000000000000001d000000000000004300000000",
            INIT_4F => X"0000001300000000000000000000000000000019000000000000000900000000",
            INIT_50 => X"0000004500000000000000400000000000000022000000000000001700000000",
            INIT_51 => X"00000042000000000000004c0000000000000043000000000000004e00000000",
            INIT_52 => X"0000002500000000000000000000000000000006000000000000000500000000",
            INIT_53 => X"0000000c000000000000000c000000000000000e000000000000003a00000000",
            INIT_54 => X"00000045000000000000003d000000000000004e000000000000003000000000",
            INIT_55 => X"0000001900000000000000510000000000000057000000000000004300000000",
            INIT_56 => X"0000002d00000000000000090000000000000020000000000000000000000000",
            INIT_57 => X"0000002c000000000000000b0000000000000025000000000000003c00000000",
            INIT_58 => X"00000047000000000000003b0000000000000020000000000000005c00000000",
            INIT_59 => X"0000000c00000000000000090000000000000059000000000000005000000000",
            INIT_5A => X"0000002400000000000000050000000000000024000000000000002600000000",
            INIT_5B => X"0000001e000000000000002c000000000000002a000000000000003d00000000",
            INIT_5C => X"0000005b00000000000000420000000000000044000000000000002600000000",
            INIT_5D => X"000000270000000000000000000000000000000d000000000000004600000000",
            INIT_5E => X"00000022000000000000000f0000000000000015000000000000001500000000",
            INIT_5F => X"00000045000000000000002c0000000000000030000000000000002f00000000",
            INIT_60 => X"000000280000000000000026000000000000003d000000000000003700000000",
            INIT_61 => X"000000000000000000000000000000000000001e000000000000000200000000",
            INIT_62 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_64 => X"0000001900000000000000000000000000000038000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"00000000000000000000001c0000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_68 => X"00000000000000000000001d0000000000000000000000000000004800000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000000000000000000000000000000000001d000000000000000000000000",
            INIT_6B => X"0000003e00000000000000040000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000800000000000000000000000000000000000000000000002000000000",
            INIT_6E => X"0000002b00000000000000000000000000000000000000000000000800000000",
            INIT_6F => X"000000000000000000000015000000000000000f000000000000000000000000",
            INIT_70 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000250000000000000000000000000000000000000000",
            INIT_72 => X"000000000000000000000000000000000000002a000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_74 => X"0000000000000000000000320000000000000000000000000000000000000000",
            INIT_75 => X"0000000100000000000000020000000000000009000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_78 => X"00000000000000000000000b0000000000000018000000000000000000000000",
            INIT_79 => X"0000000d000000000000000f000000000000000e000000000000000000000000",
            INIT_7A => X"0000001500000000000000160000000000000016000000000000000e00000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000500000000000000000000000000000000000000000000000c00000000",
            INIT_7D => X"00000009000000000000001b0000000000000027000000000000000300000000",
            INIT_7E => X"0000000000000000000000270000000000000012000000000000001200000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE30;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31 : if BRAM_NAME = "samplegold_layersamples_instance31" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_01 => X"00000016000000000000000f0000000000000014000000000000002600000000",
            INIT_02 => X"0000000000000000000000000000000000000015000000000000000e00000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000d00000000000000370000000000000000000000000000000500000000",
            INIT_05 => X"0000001400000000000000000000000000000017000000000000001700000000",
            INIT_06 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000100000000000000000000000000000017000000000000000000000000",
            INIT_08 => X"0000000200000000000000470000000000000000000000000000000000000000",
            INIT_09 => X"0000000a000000000000000e0000000000000005000000000000000300000000",
            INIT_0A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000090000000000000013000000000000001c000000000000000a00000000",
            INIT_0D => X"00000000000000000000000d0000000000000014000000000000000000000000",
            INIT_0E => X"0000001c00000000000000000000000000000000000000000000000900000000",
            INIT_0F => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000c00000000000000340000000000000000000000000000000100000000",
            INIT_11 => X"0000000f00000000000000000000000000000000000000000000001400000000",
            INIT_12 => X"00000024000000000000001d0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000013000000000000001a0000000000000025000000000000000000000000",
            INIT_15 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_16 => X"0000001c000000000000003f0000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"00000000000000000000000e0000000000000013000000000000000000000000",
            INIT_19 => X"0000000000000000000000360000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000009000000000000000f0000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000230000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_56 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000d00000000000000150000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_60 => X"000000100000000000000000000000000000000a000000000000000000000000",
            INIT_61 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000c00000000000000140000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_69 => X"0000000b00000000000000100000000000000000000000000000000000000000",
            INIT_6A => X"0000001500000000000000010000000000000000000000000000000000000000",
            INIT_6B => X"00000000000000000000000a0000000000000000000000000000000100000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_6F => X"0000000f00000000000000000000000000000000000000000000001600000000",
            INIT_70 => X"00000004000000000000000b0000000000000000000000000000000000000000",
            INIT_71 => X"0000000e00000000000000060000000000000000000000000000001800000000",
            INIT_72 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_73 => X"000000000000000000000000000000000000002d000000000000003800000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_75 => X"0000000900000000000000000000000000000000000000000000003b00000000",
            INIT_76 => X"0000000500000000000000090000000000000000000000000000000300000000",
            INIT_77 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000001800000000000000020000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000002000000000000000500000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"000000000000000000000009000000000000000d000000000000001000000000",
            INIT_7E => X"0000000000000000000000050000000000000011000000000000001000000000",
            INIT_7F => X"0000000000000000000000000000000000000039000000000000002000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE31;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32 : if BRAM_NAME = "samplegold_layersamples_instance32" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000004a00000000000000150000000000000008000000000000000000000000",
            INIT_01 => X"0000000000000000000000150000000000000003000000000000003600000000",
            INIT_02 => X"0000000000000000000000000000000000000004000000000000001400000000",
            INIT_03 => X"0000000000000000000000000000000000000026000000000000002000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000003000000000000000190000000000000007000000000000001200000000",
            INIT_06 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_07 => X"000000000000000000000003000000000000001e000000000000000300000000",
            INIT_08 => X"00000033000000000000000c0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000014000000000000004f00000000",
            INIT_0A => X"000000230000000000000012000000000000003a000000000000000000000000",
            INIT_0B => X"00000030000000000000000a0000000000000024000000000000003c00000000",
            INIT_0C => X"00000050000000000000004f0000000000000047000000000000002a00000000",
            INIT_0D => X"000000300000000000000024000000000000004e000000000000004100000000",
            INIT_0E => X"000000430000000000000045000000000000002a000000000000004b00000000",
            INIT_0F => X"00000024000000000000002f0000000000000009000000000000001a00000000",
            INIT_10 => X"00000045000000000000004b000000000000003e000000000000004e00000000",
            INIT_11 => X"00000052000000000000004d000000000000002d000000000000006200000000",
            INIT_12 => X"00000011000000000000003a0000000000000049000000000000004600000000",
            INIT_13 => X"0000004c000000000000003e000000000000002e000000000000000900000000",
            INIT_14 => X"000000850000000000000052000000000000004b000000000000003200000000",
            INIT_15 => X"0000003c00000000000000370000000000000070000000000000005f00000000",
            INIT_16 => X"0000003a0000000000000008000000000000002c000000000000004500000000",
            INIT_17 => X"00000034000000000000002f0000000000000028000000000000005b00000000",
            INIT_18 => X"0000007900000000000000a50000000000000065000000000000003b00000000",
            INIT_19 => X"0000006f000000000000006c0000000000000037000000000000007200000000",
            INIT_1A => X"00000037000000000000005e0000000000000031000000000000003000000000",
            INIT_1B => X"0000006b0000000000000054000000000000004e000000000000001800000000",
            INIT_1C => X"0000005f0000000000000088000000000000008d000000000000006d00000000",
            INIT_1D => X"0000004700000000000000980000000000000069000000000000003100000000",
            INIT_1E => X"0000004f000000000000003e0000000000000057000000000000004100000000",
            INIT_1F => X"0000004e0000000000000053000000000000005a000000000000005700000000",
            INIT_20 => X"00000034000000000000004f000000000000008f000000000000008600000000",
            INIT_21 => X"00000055000000000000008f000000000000007e000000000000005200000000",
            INIT_22 => X"000000510000000000000046000000000000003e000000000000004700000000",
            INIT_23 => X"00000070000000000000004d000000000000004e000000000000005100000000",
            INIT_24 => X"00000060000000000000004a000000000000005d000000000000007c00000000",
            INIT_25 => X"0000002d000000000000006a0000000000000093000000000000006c00000000",
            INIT_26 => X"000000470000000000000052000000000000005f000000000000005300000000",
            INIT_27 => X"00000075000000000000005c0000000000000078000000000000004c00000000",
            INIT_28 => X"00000072000000000000005f0000000000000056000000000000004700000000",
            INIT_29 => X"0000005200000000000000650000000000000083000000000000007d00000000",
            INIT_2A => X"0000006b000000000000006e000000000000005c000000000000006700000000",
            INIT_2B => X"00000042000000000000005d000000000000007d000000000000006000000000",
            INIT_2C => X"0000006300000000000000550000000000000067000000000000006e00000000",
            INIT_2D => X"00000071000000000000006a0000000000000084000000000000006d00000000",
            INIT_2E => X"0000006700000000000000630000000000000075000000000000007900000000",
            INIT_2F => X"000000620000000000000054000000000000003e000000000000005100000000",
            INIT_30 => X"00000057000000000000005d000000000000004a000000000000005100000000",
            INIT_31 => X"0000008200000000000000880000000000000080000000000000005a00000000",
            INIT_32 => X"0000004d00000000000000620000000000000066000000000000007a00000000",
            INIT_33 => X"0000006400000000000000680000000000000070000000000000005500000000",
            INIT_34 => X"0000006b0000000000000076000000000000005c000000000000005700000000",
            INIT_35 => X"0000006e00000000000000860000000000000086000000000000007800000000",
            INIT_36 => X"000000590000000000000051000000000000005f000000000000006700000000",
            INIT_37 => X"0000009c00000000000000b6000000000000007d000000000000008500000000",
            INIT_38 => X"00000082000000000000007e0000000000000069000000000000007200000000",
            INIT_39 => X"000000770000000000000076000000000000007d000000000000006d00000000",
            INIT_3A => X"0000007c000000000000003c0000000000000047000000000000005c00000000",
            INIT_3B => X"000000a7000000000000009b0000000000000037000000000000004800000000",
            INIT_3C => X"000000660000000000000077000000000000006b000000000000007600000000",
            INIT_3D => X"0000005e00000000000000750000000000000075000000000000004b00000000",
            INIT_3E => X"0000004f0000000000000067000000000000003b000000000000003b00000000",
            INIT_3F => X"000000b3000000000000009f000000000000002b000000000000001400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006800000000000000790000000000000076000000000000008300000000",
            INIT_41 => X"000000340000000000000060000000000000006f000000000000007000000000",
            INIT_42 => X"0000000000000000000000000000000000000068000000000000003a00000000",
            INIT_43 => X"00000000000000000000001d0000000000000000000000000000000000000000",
            INIT_44 => X"0000000600000000000000140000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000290000000000000000000000000000001200000000",
            INIT_46 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000030000000000000006000000000000001c000000000000000000000000",
            INIT_48 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000001700000000000000000000000000000000000000000000003800000000",
            INIT_4B => X"0000001800000000000000000000000000000000000000000000001200000000",
            INIT_4C => X"0000000000000000000000000000000000000045000000000000000000000000",
            INIT_4D => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_4F => X"0000000000000000000000280000000000000024000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"00000000000000000000000a000000000000003c000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_54 => X"0000000000000000000000000000000000000002000000000000000600000000",
            INIT_55 => X"0000000000000000000000000000000000000026000000000000004200000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000002700000000000000000000000000000015000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000300000000000000000000000000000000000000000000000700000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_5C => X"00000008000000000000000c0000000000000000000000000000000100000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_5F => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_60 => X"000000000000000000000000000000000000004f000000000000000000000000",
            INIT_61 => X"0000000000000000000000220000000000000006000000000000002000000000",
            INIT_62 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000002c00000000000000230000000000000009000000000000000000000000",
            INIT_64 => X"0000002100000000000000230000000000000009000000000000000000000000",
            INIT_65 => X"0000000000000000000000280000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000007000000000000000200000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000003300000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_6A => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000c00000000000000020000000000000000000000000000000000000000",
            INIT_6F => X"00000001000000000000004d0000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000080000000000000057000000000000000700000000",
            INIT_72 => X"0000001700000000000000110000000000000000000000000000000000000000",
            INIT_73 => X"00000000000000000000006d0000000000000018000000000000001800000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000045000000000000002300000000",
            INIT_77 => X"0000000000000000000000380000000000000000000000000000001a00000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000350000000000000013000000000000002400000000",
            INIT_7A => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"00000000000000000000001b0000000000000019000000000000000000000000",
            INIT_7C => X"0000000a00000000000000180000000000000006000000000000002e00000000",
            INIT_7D => X"0000000000000000000000340000000000000000000000000000001100000000",
            INIT_7E => X"000000010000000000000007000000000000000e000000000000002500000000",
            INIT_7F => X"0000002900000000000000000000000000000018000000000000000600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE32;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33 : if BRAM_NAME = "samplegold_layersamples_instance33" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001300000000000000000000000000000025000000000000001200000000",
            INIT_01 => X"0000001e00000000000000000000000000000042000000000000000000000000",
            INIT_02 => X"000000110000000000000012000000000000000f000000000000000100000000",
            INIT_03 => X"0000001400000000000000200000000000000000000000000000001100000000",
            INIT_04 => X"000000120000000000000000000000000000001d000000000000000900000000",
            INIT_05 => X"00000000000000000000000c0000000000000000000000000000003c00000000",
            INIT_06 => X"000000020000000000000000000000000000002b000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000001c000000000000000e00000000",
            INIT_08 => X"0000002c00000000000000190000000000000000000000000000003500000000",
            INIT_09 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_0A => X"0000002100000000000000000000000000000000000000000000003d00000000",
            INIT_0B => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000100000000000000000000000000000000e00000000",
            INIT_0D => X"0000004400000000000000000000000000000000000000000000000d00000000",
            INIT_0E => X"0000000000000000000000180000000000000000000000000000000900000000",
            INIT_0F => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_10 => X"000000170000000000000000000000000000001d000000000000000000000000",
            INIT_11 => X"00000028000000000000002d0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_15 => X"00000006000000000000001e0000000000000028000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000c0000000000000000000000000000000d000000000000000000000000",
            INIT_19 => X"00000014000000000000000e0000000000000012000000000000001100000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000800000000000000100000000000000000000000000000000000000000",
            INIT_1D => X"0000001c000000000000000f0000000000000020000000000000000a00000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000001f0000000000000000000000000000001800000000",
            INIT_21 => X"0000001f0000000000000003000000000000000f000000000000001a00000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"00000018000000000000000a0000000000000000000000000000000000000000",
            INIT_24 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000080000000000000012000000000000000100000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000001f000000000000000f0000000000000015000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_29 => X"0000001600000000000000000000000000000000000000000000002100000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000003100000000000000000000000000000010000000000000001a00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000002e00000000",
            INIT_2D => X"0000000000000000000000170000000000000000000000000000000500000000",
            INIT_2E => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000003900000000000000000000000000000000000000000000000d00000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000002500000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000003100000000000000060000000000000000000000000000000000000000",
            INIT_33 => X"00000031000000000000004a000000000000000a000000000000002600000000",
            INIT_34 => X"00000039000000000000002b0000000000000062000000000000000000000000",
            INIT_35 => X"0000006a000000000000000b0000000000000030000000000000003a00000000",
            INIT_36 => X"0000002000000000000000270000000000000045000000000000000000000000",
            INIT_37 => X"000000000000000000000030000000000000001e000000000000001c00000000",
            INIT_38 => X"00000027000000000000004c000000000000001d000000000000004d00000000",
            INIT_39 => X"000000000000000000000084000000000000000a000000000000004100000000",
            INIT_3A => X"00000022000000000000001d0000000000000027000000000000006000000000",
            INIT_3B => X"0000005800000000000000000000000000000015000000000000002200000000",
            INIT_3C => X"000000000000000000000032000000000000002f000000000000005200000000",
            INIT_3D => X"000000350000000000000005000000000000007b000000000000004700000000",
            INIT_3E => X"0000001800000000000000700000000000000000000000000000002c00000000",
            INIT_3F => X"0000002d00000000000000750000000000000019000000000000000f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000006b00000000000000000000000000000070000000000000000000000000",
            INIT_41 => X"00000000000000000000002e0000000000000014000000000000007600000000",
            INIT_42 => X"0000000a00000000000000000000000000000088000000000000000800000000",
            INIT_43 => X"0000006000000000000000000000000000000038000000000000006400000000",
            INIT_44 => X"0000003f0000000000000044000000000000005e000000000000004200000000",
            INIT_45 => X"0000000000000000000000000000000000000029000000000000002500000000",
            INIT_46 => X"000000670000000000000000000000000000002d000000000000008300000000",
            INIT_47 => X"0000002d000000000000005a0000000000000003000000000000002c00000000",
            INIT_48 => X"000000140000000000000073000000000000000c000000000000002900000000",
            INIT_49 => X"0000006300000000000000000000000000000000000000000000003200000000",
            INIT_4A => X"00000026000000000000000e0000000000000020000000000000004200000000",
            INIT_4B => X"0000002400000000000000150000000000000029000000000000001800000000",
            INIT_4C => X"0000004700000000000000050000000000000033000000000000001e00000000",
            INIT_4D => X"00000041000000000000004f0000000000000008000000000000000000000000",
            INIT_4E => X"0000003500000000000000000000000000000026000000000000002d00000000",
            INIT_4F => X"0000002200000000000000230000000000000019000000000000002200000000",
            INIT_50 => X"00000000000000000000002f0000000000000005000000000000002e00000000",
            INIT_51 => X"00000024000000000000001b0000000000000044000000000000002f00000000",
            INIT_52 => X"00000014000000000000002d000000000000000b000000000000003b00000000",
            INIT_53 => X"0000002c0000000000000009000000000000001a000000000000002500000000",
            INIT_54 => X"000000340000000000000000000000000000000a000000000000000000000000",
            INIT_55 => X"00000028000000000000004a000000000000000c000000000000000e00000000",
            INIT_56 => X"00000013000000000000002d0000000000000022000000000000002f00000000",
            INIT_57 => X"0000000000000000000000100000000000000011000000000000001700000000",
            INIT_58 => X"0000004f00000000000000000000000000000043000000000000001d00000000",
            INIT_59 => X"00000026000000000000003f0000000000000046000000000000000d00000000",
            INIT_5A => X"000000020000000000000012000000000000001c000000000000005d00000000",
            INIT_5B => X"000000200000000000000007000000000000000d000000000000001800000000",
            INIT_5C => X"0000000e00000000000000620000000000000030000000000000005100000000",
            INIT_5D => X"0000004900000000000000420000000000000011000000000000005100000000",
            INIT_5E => X"0000002f0000000000000000000000000000000f000000000000001f00000000",
            INIT_5F => X"00000028000000000000003f0000000000000003000000000000001200000000",
            INIT_60 => X"00000029000000000000001f000000000000004e000000000000003f00000000",
            INIT_61 => X"000000000000000000000031000000000000004f000000000000002600000000",
            INIT_62 => X"00000000000000000000001b0000000000000013000000000000002a00000000",
            INIT_63 => X"0000000c00000000000000380000000000000027000000000000000100000000",
            INIT_64 => X"000000200000000000000036000000000000006f000000000000004800000000",
            INIT_65 => X"000000540000000000000012000000000000003e000000000000003b00000000",
            INIT_66 => X"000000000000000000000000000000000000001e000000000000002900000000",
            INIT_67 => X"000000290000000000000000000000000000003a000000000000006300000000",
            INIT_68 => X"0000002b0000000000000033000000000000007a000000000000007800000000",
            INIT_69 => X"0000002a0000000000000019000000000000003a000000000000003200000000",
            INIT_6A => X"0000003600000000000000020000000000000000000000000000001b00000000",
            INIT_6B => X"0000001700000000000000150000000000000008000000000000009e00000000",
            INIT_6C => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"000000000000000000000000000000000000000f000000000000000200000000",
            INIT_70 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000034000000000000000300000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000031000000000000002a00000000",
            INIT_75 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_76 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000001b00000000000000180000000000000000000000000000000000000000",
            INIT_78 => X"0000000200000000000000010000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000001f00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_7C => X"0000000000000000000000140000000000000013000000000000003500000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000300000000000000000000000000000000000000000000001800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE33;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34 : if BRAM_NAME = "samplegold_layersamples_instance34" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"00000042000000000000002f0000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000000f000000000000002a00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000016000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_35 => X"00000000000000000000000d0000000000000000000000000000000500000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_37 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_38 => X"0000000300000000000000070000000000000007000000000000000900000000",
            INIT_39 => X"0000000d00000000000000000000000000000017000000000000000000000000",
            INIT_3A => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000001a000000000000000c0000000000000017000000000000001300000000",
            INIT_3C => X"00000017000000000000000d0000000000000010000000000000000b00000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_3E => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000020000000000000001a0000000000000012000000000000000f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000002a000000000000000c000000000000001e000000000000001e00000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"00000018000000000000000c0000000000000000000000000000000000000000",
            INIT_43 => X"0000001f000000000000002a000000000000001c000000000000001900000000",
            INIT_44 => X"00000003000000000000001a0000000000000023000000000000001600000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000001600000000000000320000000000000021000000000000002100000000",
            INIT_48 => X"0000000000000000000000000000000000000016000000000000002300000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000003000000000000000040000000000000000000000000000000000000000",
            INIT_4B => X"0000001c000000000000001d0000000000000023000000000000002500000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_4D => X"000000000000000000000000000000000000000e000000000000001c00000000",
            INIT_4E => X"00000022000000000000002a000000000000001d000000000000000000000000",
            INIT_4F => X"0000001b00000000000000240000000000000028000000000000001d00000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000000000000000000000f000000000000001400000000",
            INIT_52 => X"0000001c0000000000000000000000000000002b000000000000001a00000000",
            INIT_53 => X"00000000000000000000001c0000000000000023000000000000002700000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"000000000000000000000000000000000000001a000000000000000800000000",
            INIT_56 => X"0000001a00000000000000230000000000000000000000000000000000000000",
            INIT_57 => X"000000000000000000000000000000000000000c000000000000002500000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"000000070000000000000009000000000000001c000000000000000d00000000",
            INIT_5A => X"0000000000000000000000160000000000000013000000000000000000000000",
            INIT_5B => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000054000000000000002c000000000000002c000000000000003400000000",
            INIT_5D => X"0000003a00000000000000180000000000000037000000000000000300000000",
            INIT_5E => X"0000007a00000000000000000000000000000046000000000000001f00000000",
            INIT_5F => X"000000360000000000000026000000000000001d000000000000000e00000000",
            INIT_60 => X"0000001a00000000000000510000000000000029000000000000004000000000",
            INIT_61 => X"0000002c00000000000000310000000000000013000000000000001f00000000",
            INIT_62 => X"00000019000000000000005d0000000000000000000000000000004600000000",
            INIT_63 => X"0000002400000000000000120000000000000034000000000000004000000000",
            INIT_64 => X"00000031000000000000000a0000000000000040000000000000002e00000000",
            INIT_65 => X"0000000700000000000000510000000000000011000000000000004d00000000",
            INIT_66 => X"00000034000000000000002f0000000000000046000000000000000000000000",
            INIT_67 => X"0000002c00000000000000460000000000000003000000000000004100000000",
            INIT_68 => X"00000040000000000000005e000000000000002e000000000000001800000000",
            INIT_69 => X"0000001b00000000000000200000000000000025000000000000000900000000",
            INIT_6A => X"00000045000000000000005e0000000000000026000000000000002c00000000",
            INIT_6B => X"0000000000000000000000450000000000000048000000000000000000000000",
            INIT_6C => X"0000004000000000000000020000000000000063000000000000003600000000",
            INIT_6D => X"00000034000000000000001d0000000000000047000000000000002a00000000",
            INIT_6E => X"0000000000000000000000480000000000000073000000000000002300000000",
            INIT_6F => X"000000170000000000000031000000000000004f000000000000001700000000",
            INIT_70 => X"0000002e00000000000000370000000000000012000000000000001800000000",
            INIT_71 => X"00000015000000000000004b0000000000000007000000000000003000000000",
            INIT_72 => X"0000000b0000000000000010000000000000003f000000000000007800000000",
            INIT_73 => X"0000000e000000000000000d000000000000002a000000000000002900000000",
            INIT_74 => X"000000000000000000000003000000000000000f000000000000001e00000000",
            INIT_75 => X"0000005f0000000000000023000000000000002b000000000000001500000000",
            INIT_76 => X"0000001e000000000000001a000000000000000d000000000000003300000000",
            INIT_77 => X"0000000600000000000000000000000000000037000000000000000000000000",
            INIT_78 => X"00000000000000000000001a0000000000000011000000000000000a00000000",
            INIT_79 => X"000000180000000000000062000000000000001d000000000000003000000000",
            INIT_7A => X"0000000a000000000000001d000000000000002a000000000000002d00000000",
            INIT_7B => X"0000000e00000000000000000000000000000006000000000000000100000000",
            INIT_7C => X"00000015000000000000000f0000000000000009000000000000000100000000",
            INIT_7D => X"00000028000000000000002d000000000000003b000000000000002800000000",
            INIT_7E => X"0000000000000000000000150000000000000011000000000000003900000000",
            INIT_7F => X"0000000f00000000000000030000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE34;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35 : if BRAM_NAME = "samplegold_layersamples_instance35" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002500000000000000290000000000000016000000000000000600000000",
            INIT_01 => X"000000440000000000000000000000000000004c000000000000000a00000000",
            INIT_02 => X"00000000000000000000001e0000000000000036000000000000001200000000",
            INIT_03 => X"0000000000000000000000130000000000000002000000000000000900000000",
            INIT_04 => X"0000003100000000000000140000000000000023000000000000000a00000000",
            INIT_05 => X"0000003300000000000000650000000000000029000000000000000300000000",
            INIT_06 => X"0000000000000000000000000000000000000014000000000000003000000000",
            INIT_07 => X"0000001100000000000000000000000000000013000000000000000000000000",
            INIT_08 => X"0000002000000000000000350000000000000012000000000000002a00000000",
            INIT_09 => X"0000004d000000000000005c000000000000002f000000000000000000000000",
            INIT_0A => X"00000000000000000000002b0000000000000014000000000000000c00000000",
            INIT_0B => X"0000002e00000000000000160000000000000007000000000000000000000000",
            INIT_0C => X"0000002500000000000000450000000000000043000000000000001600000000",
            INIT_0D => X"000000500000000000000061000000000000001a000000000000000000000000",
            INIT_0E => X"000000000000000000000016000000000000002a000000000000003600000000",
            INIT_0F => X"0000000f00000000000000430000000000000025000000000000000000000000",
            INIT_10 => X"0000001800000000000000370000000000000055000000000000000d00000000",
            INIT_11 => X"0000005c0000000000000051000000000000001a000000000000000000000000",
            INIT_12 => X"0000000a00000000000000010000000000000035000000000000004600000000",
            INIT_13 => X"0000000f0000000000000031000000000000003b000000000000000700000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000010000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_34 => X"00000010000000000000001f0000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_39 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_3A => X"0000000700000000000000000000000000000035000000000000000000000000",
            INIT_3B => X"0000000000000000000000180000000000000000000000000000000d00000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000008000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000001b00000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE35;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36 : if BRAM_NAME = "samplegold_layersamples_instance36" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000f00000000000000080000000000000000000000000000000200000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000500000000000000010000000000000008000000000000000600000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"00000004000000000000000e0000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000050000000000000003000000000000000900000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000400000000000000000000000000000008000000000000000c00000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000500000000000000000000000000000007000000000000000000000000",
            INIT_16 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_17 => X"0000000b00000000000000000000000000000015000000000000000300000000",
            INIT_18 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000080000000000000000000000000000000300000000",
            INIT_1A => X"0000000700000000000000000000000000000004000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000006000000000000002700000000",
            INIT_1C => X"0000000000000000000000000000000000000009000000000000000600000000",
            INIT_1D => X"0000000000000000000000000000000000000013000000000000001b00000000",
            INIT_1E => X"0000000200000000000000040000000000000003000000000000000500000000",
            INIT_1F => X"0000000e00000000000000010000000000000000000000000000002000000000",
            INIT_20 => X"0000000b00000000000000100000000000000006000000000000000300000000",
            INIT_21 => X"0000000200000000000000000000000000000000000000000000000400000000",
            INIT_22 => X"0000001c000000000000000b0000000000000000000000000000000a00000000",
            INIT_23 => X"0000000800000000000000030000000000000000000000000000000c00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000001600000000000000110000000000000000000000000000000000000000",
            INIT_26 => X"0000000c00000000000000250000000000000001000000000000000000000000",
            INIT_27 => X"000000000000000000000009000000000000000f000000000000000000000000",
            INIT_28 => X"0000000200000000000000000000000000000000000000000000000f00000000",
            INIT_29 => X"000000000000000000000020000000000000000c000000000000000300000000",
            INIT_2A => X"0000000000000000000000030000000000000019000000000000000800000000",
            INIT_2B => X"0000001100000000000000000000000000000001000000000000000c00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000300000000000000000000000000000021000000000000000c00000000",
            INIT_2E => X"0000000000000000000000050000000000000003000000000000001400000000",
            INIT_2F => X"0000000000000000000000000000000000000012000000000000000f00000000",
            INIT_30 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000e000000000000000f0000000000000000000000000000001100000000",
            INIT_32 => X"0000000000000000000000000000000000000002000000000000000f00000000",
            INIT_33 => X"0000000100000000000000010000000000000004000000000000000f00000000",
            INIT_34 => X"00000000000000000000000b0000000000000003000000000000000000000000",
            INIT_35 => X"000000020000000000000013000000000000000a000000000000001500000000",
            INIT_36 => X"00000016000000000000000c0000000000000000000000000000000700000000",
            INIT_37 => X"000000070000000000000008000000000000000b000000000000000100000000",
            INIT_38 => X"00000000000000000000000f0000000000000006000000000000000f00000000",
            INIT_39 => X"00000013000000000000000a000000000000001a000000000000000d00000000",
            INIT_3A => X"000000030000000000000009000000000000000f000000000000000a00000000",
            INIT_3B => X"0000000c000000000000000c000000000000000b000000000000000300000000",
            INIT_3C => X"0000002c000000000000000f0000000000000000000000000000000800000000",
            INIT_3D => X"00000012000000000000000a0000000000000010000000000000000000000000",
            INIT_3E => X"0000003300000000000000000000000000000011000000000000000900000000",
            INIT_3F => X"000000010000000000000010000000000000000b000000000000000900000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000260000000000000014000000000000002b000000000000000000000000",
            INIT_41 => X"0000000a00000000000000070000000000000009000000000000000300000000",
            INIT_42 => X"0000001200000000000000260000000000000002000000000000001400000000",
            INIT_43 => X"0000001f000000000000000b000000000000000d000000000000000000000000",
            INIT_44 => X"000000060000000000000005000000000000003a000000000000000c00000000",
            INIT_45 => X"00000015000000000000000c0000000000000007000000000000000600000000",
            INIT_46 => X"000000000000000000000026000000000000000c000000000000000000000000",
            INIT_47 => X"0000000f000000000000000f0000000000000012000000000000001c00000000",
            INIT_48 => X"00000000000000000000000d000000000000000a000000000000002800000000",
            INIT_49 => X"00000011000000000000001a000000000000000b000000000000001100000000",
            INIT_4A => X"0000002f000000000000000a000000000000000e000000000000000200000000",
            INIT_4B => X"0000000f000000000000000c0000000000000000000000000000001100000000",
            INIT_4C => X"0000000b0000000000000003000000000000000e000000000000000500000000",
            INIT_4D => X"0000002800000000000000100000000000000018000000000000001300000000",
            INIT_4E => X"00000001000000000000005c000000000000000b000000000000000000000000",
            INIT_4F => X"000000130000000000000000000000000000000e000000000000001100000000",
            INIT_50 => X"0000000000000000000000160000000000000013000000000000000000000000",
            INIT_51 => X"00000000000000000000003f0000000000000036000000000000004b00000000",
            INIT_52 => X"0000000b00000000000000000000000000000045000000000000002a00000000",
            INIT_53 => X"0000002b00000000000000000000000000000000000000000000000400000000",
            INIT_54 => X"0000002f00000000000000190000000000000000000000000000002800000000",
            INIT_55 => X"0000004f00000000000000110000000000000000000000000000002f00000000",
            INIT_56 => X"0000000e00000000000000030000000000000000000000000000003200000000",
            INIT_57 => X"0000001300000000000000340000000000000000000000000000002400000000",
            INIT_58 => X"0000001500000000000000200000000000000031000000000000000000000000",
            INIT_59 => X"00000041000000000000006c000000000000002f000000000000002d00000000",
            INIT_5A => X"0000002700000000000000380000000000000000000000000000000000000000",
            INIT_5B => X"0000001800000000000000390000000000000029000000000000000000000000",
            INIT_5C => X"000000270000000000000025000000000000005c000000000000000000000000",
            INIT_5D => X"000000000000000000000022000000000000006b000000000000003e00000000",
            INIT_5E => X"00000000000000000000002c0000000000000079000000000000000000000000",
            INIT_5F => X"00000011000000000000000000000000000000a7000000000000002d00000000",
            INIT_60 => X"0000001e00000000000000550000000000000000000000000000006200000000",
            INIT_61 => X"0000000000000000000000000000000000000020000000000000001100000000",
            INIT_62 => X"000000370000000000000000000000000000003700000000000000a500000000",
            INIT_63 => X"0000001600000000000000010000000000000000000000000000008f00000000",
            INIT_64 => X"0000001400000000000000210000000000000051000000000000000000000000",
            INIT_65 => X"0000009000000000000000000000000000000000000000000000000700000000",
            INIT_66 => X"00000034000000000000000e0000000000000010000000000000002300000000",
            INIT_67 => X"0000003900000000000000070000000000000005000000000000002900000000",
            INIT_68 => X"0000000000000000000000140000000000000009000000000000001800000000",
            INIT_69 => X"0000000d00000000000000180000000000000000000000000000000000000000",
            INIT_6A => X"0000004200000000000000030000000000000016000000000000001600000000",
            INIT_6B => X"0000002400000000000000320000000000000004000000000000002e00000000",
            INIT_6C => X"0000000000000000000000000000000000000011000000000000001000000000",
            INIT_6D => X"00000000000000000000002d0000000000000000000000000000000000000000",
            INIT_6E => X"0000000700000000000000360000000000000003000000000000003e00000000",
            INIT_6F => X"0000001e00000000000000100000000000000037000000000000000000000000",
            INIT_70 => X"0000000300000000000000120000000000000001000000000000001100000000",
            INIT_71 => X"000000230000000000000009000000000000000f000000000000002400000000",
            INIT_72 => X"0000001c000000000000001b0000000000000018000000000000000e00000000",
            INIT_73 => X"0000000a0000000000000015000000000000001b000000000000002000000000",
            INIT_74 => X"000000000000000000000027000000000000001b000000000000000800000000",
            INIT_75 => X"000000190000000000000005000000000000005f000000000000001800000000",
            INIT_76 => X"0000000b0000000000000009000000000000000c000000000000000b00000000",
            INIT_77 => X"0000000e00000000000000000000000000000000000000000000000300000000",
            INIT_78 => X"0000001100000000000000060000000000000014000000000000000b00000000",
            INIT_79 => X"0000001400000000000000100000000000000008000000000000000000000000",
            INIT_7A => X"0000001c00000000000000180000000000000019000000000000001c00000000",
            INIT_7B => X"0000000800000000000000000000000000000000000000000000000900000000",
            INIT_7C => X"0000000000000000000000050000000000000003000000000000000b00000000",
            INIT_7D => X"0000000a00000000000000100000000000000006000000000000001100000000",
            INIT_7E => X"0000004900000000000000180000000000000008000000000000001300000000",
            INIT_7F => X"0000000000000000000000000000000000000022000000000000004800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE36;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37 : if BRAM_NAME = "samplegold_layersamples_instance37" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_01 => X"0000000000000000000000010000000000000003000000000000000e00000000",
            INIT_02 => X"0000001100000000000000000000000000000000000000000000000700000000",
            INIT_03 => X"00000001000000000000000b0000000000000000000000000000001400000000",
            INIT_04 => X"00000004000000000000000b000000000000000c000000000000000000000000",
            INIT_05 => X"0000002e0000000000000003000000000000000f000000000000000a00000000",
            INIT_06 => X"0000000000000000000000020000000000000000000000000000000d00000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"00000000000000000000000d0000000000000020000000000000000900000000",
            INIT_09 => X"000000000000000000000000000000000000002a000000000000001f00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_0B => X"00000000000000000000002e0000000000000000000000000000000000000000",
            INIT_0C => X"0000001000000000000000190000000000000004000000000000000000000000",
            INIT_0D => X"0000003a00000000000000660000000000000040000000000000000000000000",
            INIT_0E => X"0000000600000000000000030000000000000000000000000000000100000000",
            INIT_0F => X"0000000000000000000000050000000000000009000000000000000000000000",
            INIT_10 => X"000000250000000000000012000000000000001b000000000000000000000000",
            INIT_11 => X"0000002700000000000000080000000000000001000000000000000f00000000",
            INIT_12 => X"00000016000000000000002f0000000000000000000000000000000000000000",
            INIT_13 => X"000000000000000000000011000000000000001e000000000000001900000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000030000000000000016000000000000000b000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000003000000000000001200000000",
            INIT_18 => X"00000018000000000000003c0000000000000000000000000000000000000000",
            INIT_19 => X"00000003000000000000002a000000000000000f000000000000000000000000",
            INIT_1A => X"0000000000000000000000100000000000000028000000000000001500000000",
            INIT_1B => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_1E => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_1F => X"00000045000000000000004f000000000000002d000000000000004800000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"00000000000000000000000b0000000000000000000000000000001500000000",
            INIT_23 => X"00000037000000000000000f0000000000000000000000000000002700000000",
            INIT_24 => X"00000027000000000000002f0000000000000036000000000000003a00000000",
            INIT_25 => X"0000000100000000000000000000000000000000000000000000001500000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"00000021000000000000000c000000000000000b000000000000000f00000000",
            INIT_28 => X"00000044000000000000004f0000000000000034000000000000003200000000",
            INIT_29 => X"0000003300000000000000030000000000000000000000000000003b00000000",
            INIT_2A => X"0000001a00000000000000250000000000000023000000000000000700000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2C => X"0000001100000000000000170000000000000011000000000000001600000000",
            INIT_2D => X"0000008900000000000000780000000000000074000000000000002000000000",
            INIT_2E => X"0000008c0000000000000093000000000000008f000000000000008b00000000",
            INIT_2F => X"0000004b000000000000004a0000000000000069000000000000007400000000",
            INIT_30 => X"0000004f0000000000000052000000000000004b000000000000005100000000",
            INIT_31 => X"0000008d000000000000008a0000000000000089000000000000008000000000",
            INIT_32 => X"0000009500000000000000a1000000000000009a000000000000009600000000",
            INIT_33 => X"0000005400000000000000450000000000000059000000000000008a00000000",
            INIT_34 => X"0000008500000000000000530000000000000062000000000000005600000000",
            INIT_35 => X"000000960000000000000095000000000000008f000000000000007500000000",
            INIT_36 => X"00000091000000000000009d00000000000000a600000000000000a000000000",
            INIT_37 => X"00000066000000000000006c0000000000000061000000000000006e00000000",
            INIT_38 => X"000000740000000000000064000000000000005d000000000000005e00000000",
            INIT_39 => X"000000a6000000000000009a0000000000000090000000000000008d00000000",
            INIT_3A => X"0000008e0000000000000090000000000000009900000000000000a500000000",
            INIT_3B => X"0000006000000000000000600000000000000087000000000000008700000000",
            INIT_3C => X"0000008b0000000000000077000000000000005e000000000000006000000000",
            INIT_3D => X"00000080000000000000009d000000000000009d000000000000009200000000",
            INIT_3E => X"000000830000000000000088000000000000008e000000000000007d00000000",
            INIT_3F => X"0000005c000000000000005b0000000000000051000000000000007f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000910000000000000089000000000000007b000000000000002900000000",
            INIT_41 => X"0000006600000000000000660000000000000061000000000000009300000000",
            INIT_42 => X"0000005a00000000000000780000000000000062000000000000005e00000000",
            INIT_43 => X"0000004a00000000000000590000000000000055000000000000004300000000",
            INIT_44 => X"00000068000000000000007b000000000000007a000000000000005a00000000",
            INIT_45 => X"0000004e00000000000000540000000000000063000000000000007600000000",
            INIT_46 => X"0000003600000000000000460000000000000064000000000000005600000000",
            INIT_47 => X"0000004b00000000000000660000000000000059000000000000005100000000",
            INIT_48 => X"00000073000000000000005b0000000000000067000000000000007700000000",
            INIT_49 => X"000000520000000000000054000000000000005f000000000000008600000000",
            INIT_4A => X"0000004700000000000000240000000000000045000000000000006e00000000",
            INIT_4B => X"0000006d000000000000004d000000000000007d000000000000006400000000",
            INIT_4C => X"00000099000000000000005b000000000000005c000000000000007600000000",
            INIT_4D => X"00000056000000000000006a0000000000000066000000000000007100000000",
            INIT_4E => X"0000006700000000000000420000000000000026000000000000003300000000",
            INIT_4F => X"0000008a00000000000000560000000000000056000000000000008200000000",
            INIT_50 => X"0000005c0000000000000077000000000000005c000000000000002200000000",
            INIT_51 => X"0000004100000000000000360000000000000045000000000000008900000000",
            INIT_52 => X"0000008900000000000000630000000000000033000000000000002f00000000",
            INIT_53 => X"0000003c0000000000000064000000000000005c000000000000005e00000000",
            INIT_54 => X"00000068000000000000006e0000000000000051000000000000004500000000",
            INIT_55 => X"00000043000000000000002f0000000000000032000000000000004100000000",
            INIT_56 => X"0000007700000000000000780000000000000057000000000000003900000000",
            INIT_57 => X"0000004f00000000000000650000000000000067000000000000005000000000",
            INIT_58 => X"000000230000000000000039000000000000005d000000000000005c00000000",
            INIT_59 => X"00000057000000000000002c0000000000000021000000000000001a00000000",
            INIT_5A => X"0000007500000000000000760000000000000084000000000000003f00000000",
            INIT_5B => X"00000067000000000000006d000000000000007f000000000000005800000000",
            INIT_5C => X"00000026000000000000002d0000000000000045000000000000006e00000000",
            INIT_5D => X"00000055000000000000003c0000000000000037000000000000001a00000000",
            INIT_5E => X"00000069000000000000007e0000000000000067000000000000008300000000",
            INIT_5F => X"0000008200000000000000710000000000000066000000000000006800000000",
            INIT_60 => X"000000520000000000000050000000000000005a000000000000006000000000",
            INIT_61 => X"00000070000000000000004f000000000000005d000000000000005600000000",
            INIT_62 => X"0000006d0000000000000076000000000000007d000000000000007e00000000",
            INIT_63 => X"0000007900000000000000790000000000000087000000000000007f00000000",
            INIT_64 => X"0000007a00000000000000760000000000000076000000000000007300000000",
            INIT_65 => X"0000003300000000000000040000000000000062000000000000007700000000",
            INIT_66 => X"0000003200000000000000290000000000000039000000000000002a00000000",
            INIT_67 => X"0000002300000000000000030000000000000033000000000000002c00000000",
            INIT_68 => X"00000039000000000000002c0000000000000020000000000000002b00000000",
            INIT_69 => X"0000003100000000000000140000000000000026000000000000001300000000",
            INIT_6A => X"0000002d00000000000000330000000000000034000000000000002e00000000",
            INIT_6B => X"000000380000000000000017000000000000000e000000000000003b00000000",
            INIT_6C => X"0000002c00000000000000200000000000000035000000000000003400000000",
            INIT_6D => X"00000034000000000000002e000000000000002d000000000000000300000000",
            INIT_6E => X"0000004100000000000000280000000000000030000000000000003300000000",
            INIT_6F => X"0000002100000000000000390000000000000005000000000000003100000000",
            INIT_70 => X"00000008000000000000002d0000000000000033000000000000003500000000",
            INIT_71 => X"0000002f0000000000000039000000000000002b000000000000002700000000",
            INIT_72 => X"00000040000000000000002f0000000000000032000000000000003500000000",
            INIT_73 => X"0000002a00000000000000100000000000000027000000000000003300000000",
            INIT_74 => X"0000003300000000000000230000000000000033000000000000003d00000000",
            INIT_75 => X"000000290000000000000033000000000000002d000000000000002b00000000",
            INIT_76 => X"0000004e000000000000001d000000000000002f000000000000002900000000",
            INIT_77 => X"0000002c00000000000000360000000000000000000000000000003700000000",
            INIT_78 => X"0000003a0000000000000018000000000000007f000000000000002f00000000",
            INIT_79 => X"00000000000000000000003d0000000000000022000000000000002a00000000",
            INIT_7A => X"00000020000000000000003d0000000000000004000000000000001c00000000",
            INIT_7B => X"00000036000000000000002b0000000000000036000000000000000000000000",
            INIT_7C => X"0000001200000000000000150000000000000048000000000000006b00000000",
            INIT_7D => X"0000000000000000000000080000000000000021000000000000003400000000",
            INIT_7E => X"000000030000000000000000000000000000001e000000000000002c00000000",
            INIT_7F => X"00000015000000000000002c000000000000002d000000000000002c00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE37;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38 : if BRAM_NAME = "samplegold_layersamples_instance38" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000003400000000000000230000000000000012000000000000007100000000",
            INIT_01 => X"0000001000000000000000260000000000000022000000000000001100000000",
            INIT_02 => X"0000003300000000000000000000000000000000000000000000000800000000",
            INIT_03 => X"0000005c000000000000002d0000000000000008000000000000003400000000",
            INIT_04 => X"000000340000000000000023000000000000000a000000000000001c00000000",
            INIT_05 => X"0000001500000000000000220000000000000024000000000000000700000000",
            INIT_06 => X"0000004700000000000000500000000000000009000000000000000000000000",
            INIT_07 => X"00000015000000000000006b0000000000000020000000000000000000000000",
            INIT_08 => X"0000000000000000000000310000000000000068000000000000000000000000",
            INIT_09 => X"0000001d000000000000000e0000000000000000000000000000004900000000",
            INIT_0A => X"000000000000000000000060000000000000004a000000000000001900000000",
            INIT_0B => X"00000000000000000000000b0000000000000056000000000000002500000000",
            INIT_0C => X"00000051000000000000002c000000000000002d000000000000002d00000000",
            INIT_0D => X"0000002d000000000000001d0000000000000013000000000000000800000000",
            INIT_0E => X"0000002f00000000000000000000000000000073000000000000003d00000000",
            INIT_0F => X"0000000e000000000000000c0000000000000025000000000000003d00000000",
            INIT_10 => X"0000000900000000000000000000000000000031000000000000003300000000",
            INIT_11 => X"000000490000000000000026000000000000000d000000000000001800000000",
            INIT_12 => X"0000003800000000000000440000000000000020000000000000004c00000000",
            INIT_13 => X"00000019000000000000000d0000000000000038000000000000002b00000000",
            INIT_14 => X"0000000d000000000000000b0000000000000017000000000000004400000000",
            INIT_15 => X"000000290000000000000033000000000000001c000000000000000b00000000",
            INIT_16 => X"0000001d0000000000000057000000000000002b000000000000003e00000000",
            INIT_17 => X"0000004a00000000000000350000000000000011000000000000003400000000",
            INIT_18 => X"000000230000000000000023000000000000002e000000000000002000000000",
            INIT_19 => X"000000160000000000000032000000000000001d000000000000003000000000",
            INIT_1A => X"0000004000000000000000320000000000000044000000000000003c00000000",
            INIT_1B => X"0000003600000000000000340000000000000035000000000000002a00000000",
            INIT_1C => X"0000003f00000000000000410000000000000037000000000000002f00000000",
            INIT_1D => X"0000002300000000000000400000000000000020000000000000002f00000000",
            INIT_1E => X"00000038000000000000002f0000000000000036000000000000000100000000",
            INIT_1F => X"0000003000000000000000360000000000000043000000000000003c00000000",
            INIT_20 => X"000000260000000000000029000000000000002c000000000000002a00000000",
            INIT_21 => X"0000002200000000000000140000000000000028000000000000002100000000",
            INIT_22 => X"000000330000000000000036000000000000002f000000000000003200000000",
            INIT_23 => X"0000002c00000000000000480000000000000041000000000000003f00000000",
            INIT_24 => X"0000002f000000000000002c0000000000000030000000000000002c00000000",
            INIT_25 => X"000000270000000000000019000000000000001a000000000000002d00000000",
            INIT_26 => X"0000003e000000000000003a000000000000002e000000000000003200000000",
            INIT_27 => X"00000018000000000000001d000000000000003e000000000000003d00000000",
            INIT_28 => X"0000002b00000000000000390000000000000036000000000000002d00000000",
            INIT_29 => X"0000002c000000000000002b0000000000000016000000000000001a00000000",
            INIT_2A => X"0000004000000000000000420000000000000043000000000000002b00000000",
            INIT_2B => X"000000360000000000000039000000000000003d000000000000003a00000000",
            INIT_2C => X"0000002300000000000000300000000000000031000000000000003c00000000",
            INIT_2D => X"0000002c000000000000002e0000000000000021000000000000001800000000",
            INIT_2E => X"0000002a000000000000001a0000000000000026000000000000003800000000",
            INIT_2F => X"0000002a000000000000002f0000000000000032000000000000004000000000",
            INIT_30 => X"0000002200000000000000230000000000000030000000000000003100000000",
            INIT_31 => X"0000000d00000000000000310000000000000022000000000000001500000000",
            INIT_32 => X"00000023000000000000002c0000000000000014000000000000000000000000",
            INIT_33 => X"0000002f0000000000000024000000000000003b000000000000002c00000000",
            INIT_34 => X"0000000f00000000000000210000000000000000000000000000002e00000000",
            INIT_35 => X"0000001e0000000000000000000000000000000e000000000000001600000000",
            INIT_36 => X"0000001e00000000000000000000000000000000000000000000000600000000",
            INIT_37 => X"0000002e00000000000000280000000000000019000000000000002800000000",
            INIT_38 => X"0000001900000000000000120000000000000012000000000000003000000000",
            INIT_39 => X"0000000400000000000000110000000000000000000000000000000000000000",
            INIT_3A => X"0000001e00000000000000050000000000000000000000000000000000000000",
            INIT_3B => X"0000003800000000000000200000000000000011000000000000001900000000",
            INIT_3C => X"0000000600000000000000170000000000000003000000000000000f00000000",
            INIT_3D => X"000000300000000000000037000000000000001b000000000000002000000000",
            INIT_3E => X"0000001400000000000000380000000000000051000000000000003700000000",
            INIT_3F => X"0000001a00000000000000450000000000000017000000000000000f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c00000000000000240000000000000025000000000000000000000000",
            INIT_41 => X"0000003e000000000000002f0000000000000013000000000000003800000000",
            INIT_42 => X"00000009000000000000001b000000000000001d000000000000001b00000000",
            INIT_43 => X"0000000d000000000000002a0000000000000036000000000000000000000000",
            INIT_44 => X"00000048000000000000003f000000000000001c000000000000004100000000",
            INIT_45 => X"0000002b00000000000000320000000000000058000000000000004b00000000",
            INIT_46 => X"0000000b0000000000000018000000000000001d000000000000003000000000",
            INIT_47 => X"00000000000000000000001f000000000000002a000000000000004700000000",
            INIT_48 => X"0000003f000000000000001c000000000000001a000000000000002800000000",
            INIT_49 => X"0000001e00000000000000200000000000000025000000000000002f00000000",
            INIT_4A => X"00000036000000000000002a000000000000002b000000000000002c00000000",
            INIT_4B => X"0000000e00000000000000270000000000000021000000000000003f00000000",
            INIT_4C => X"0000001b000000000000002e0000000000000035000000000000003400000000",
            INIT_4D => X"00000017000000000000000f0000000000000013000000000000001500000000",
            INIT_4E => X"00000039000000000000003b000000000000001f000000000000003100000000",
            INIT_4F => X"0000002900000000000000350000000000000030000000000000003600000000",
            INIT_50 => X"0000001f000000000000002a0000000000000041000000000000003000000000",
            INIT_51 => X"0000001800000000000000180000000000000013000000000000002000000000",
            INIT_52 => X"0000003b0000000000000027000000000000003e000000000000003200000000",
            INIT_53 => X"0000003e000000000000002d0000000000000023000000000000002d00000000",
            INIT_54 => X"00000036000000000000003e000000000000003d000000000000004300000000",
            INIT_55 => X"0000002800000000000000340000000000000032000000000000003400000000",
            INIT_56 => X"0000001100000000000000180000000000000000000000000000000000000000",
            INIT_57 => X"000000040000000000000017000000000000000d000000000000000f00000000",
            INIT_58 => X"00000000000000000000000a0000000000000013000000000000001200000000",
            INIT_59 => X"0000001100000000000000120000000000000004000000000000000000000000",
            INIT_5A => X"0000000d0000000000000006000000000000000b000000000000001900000000",
            INIT_5B => X"00000002000000000000000a0000000000000010000000000000000a00000000",
            INIT_5C => X"00000014000000000000001f000000000000000b000000000000000100000000",
            INIT_5D => X"000000080000000000000017000000000000000c000000000000000d00000000",
            INIT_5E => X"00000010000000000000000d0000000000000013000000000000000700000000",
            INIT_5F => X"0000000000000000000000150000000000000015000000000000000b00000000",
            INIT_60 => X"0000001e00000000000000170000000000000008000000000000000000000000",
            INIT_61 => X"00000012000000000000000f0000000000000012000000000000000b00000000",
            INIT_62 => X"00000026000000000000001d0000000000000017000000000000001100000000",
            INIT_63 => X"0000000000000000000000190000000000000024000000000000001e00000000",
            INIT_64 => X"0000000f0000000000000001000000000000000f000000000000000900000000",
            INIT_65 => X"00000005000000000000000d0000000000000007000000000000002200000000",
            INIT_66 => X"000000000000000000000010000000000000001e000000000000001100000000",
            INIT_67 => X"0000002b000000000000001f0000000000000025000000000000000b00000000",
            INIT_68 => X"000000040000000000000013000000000000001e000000000000001500000000",
            INIT_69 => X"0000001c00000000000000120000000000000000000000000000000000000000",
            INIT_6A => X"00000037000000000000004f0000000000000001000000000000000000000000",
            INIT_6B => X"000000150000000000000026000000000000001a000000000000000d00000000",
            INIT_6C => X"0000002300000000000000000000000000000010000000000000001300000000",
            INIT_6D => X"000000070000000000000000000000000000000d000000000000001700000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_6F => X"000000020000000000000000000000000000000c000000000000001000000000",
            INIT_70 => X"0000001b00000000000000070000000000000003000000000000001400000000",
            INIT_71 => X"0000000900000000000000100000000000000000000000000000002000000000",
            INIT_72 => X"0000000900000000000000070000000000000012000000000000001000000000",
            INIT_73 => X"0000000a00000000000000000000000000000007000000000000001f00000000",
            INIT_74 => X"00000022000000000000000c0000000000000000000000000000001900000000",
            INIT_75 => X"000000470000000000000030000000000000000c000000000000001800000000",
            INIT_76 => X"0000001500000000000000670000000000000063000000000000004900000000",
            INIT_77 => X"0000000d000000000000000b0000000000000000000000000000000000000000",
            INIT_78 => X"0000006600000000000000250000000000000011000000000000000000000000",
            INIT_79 => X"0000000d000000000000000c0000000000000042000000000000002d00000000",
            INIT_7A => X"0000000600000000000000000000000000000000000000000000001b00000000",
            INIT_7B => X"00000018000000000000001c0000000000000000000000000000000000000000",
            INIT_7C => X"0000002a00000000000000000000000000000030000000000000002300000000",
            INIT_7D => X"0000001a00000000000000620000000000000030000000000000003600000000",
            INIT_7E => X"0000001a0000000000000000000000000000001f000000000000002000000000",
            INIT_7F => X"000000170000000000000007000000000000002f000000000000002100000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE38;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39 : if BRAM_NAME = "samplegold_layersamples_instance39" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_01 => X"0000000b00000000000000040000000000000000000000000000001100000000",
            INIT_02 => X"0000002c0000000000000021000000000000000a000000000000000600000000",
            INIT_03 => X"0000003e00000000000000000000000000000018000000000000001400000000",
            INIT_04 => X"0000000000000000000000030000000000000023000000000000002300000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000001f00000000000000030000000000000000000000000000000000000000",
            INIT_07 => X"0000002d00000000000000090000000000000030000000000000002300000000",
            INIT_08 => X"0000000000000000000000170000000000000010000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000000000000a0000000000000021000000000000000000000000",
            INIT_0B => X"0000000a0000000000000000000000000000000d000000000000001800000000",
            INIT_0C => X"0000001500000000000000190000000000000031000000000000002100000000",
            INIT_0D => X"0000000f000000000000000e0000000000000010000000000000000e00000000",
            INIT_0E => X"000000150000000000000003000000000000001a000000000000000300000000",
            INIT_0F => X"0000000200000000000000060000000000000011000000000000001200000000",
            INIT_10 => X"000000050000000000000003000000000000000b000000000000000000000000",
            INIT_11 => X"0000000a00000000000000070000000000000000000000000000000000000000",
            INIT_12 => X"0000001900000000000000140000000000000035000000000000003800000000",
            INIT_13 => X"0000000000000000000000000000000000000010000000000000001700000000",
            INIT_14 => X"0000000a00000000000000060000000000000000000000000000000000000000",
            INIT_15 => X"0000003c00000000000000080000000000000008000000000000000b00000000",
            INIT_16 => X"000000240000000000000022000000000000001e000000000000003b00000000",
            INIT_17 => X"0000000d0000000000000008000000000000000f000000000000001900000000",
            INIT_18 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"00000036000000000000003e0000000000000008000000000000000d00000000",
            INIT_1A => X"0000001a000000000000002c0000000000000027000000000000002b00000000",
            INIT_1B => X"0000001b000000000000001a000000000000000d000000000000001d00000000",
            INIT_1C => X"0000000200000000000000040000000000000008000000000000000800000000",
            INIT_1D => X"0000002d00000000000000360000000000000033000000000000000e00000000",
            INIT_1E => X"000000330000000000000027000000000000002c000000000000002600000000",
            INIT_1F => X"0000001f000000000000001e0000000000000015000000000000002900000000",
            INIT_20 => X"00000011000000000000000e000000000000000c000000000000001f00000000",
            INIT_21 => X"00000038000000000000003a000000000000002d000000000000002800000000",
            INIT_22 => X"000000560000000000000051000000000000004f000000000000002c00000000",
            INIT_23 => X"0000001600000000000000230000000000000026000000000000003700000000",
            INIT_24 => X"00000007000000000000000e0000000000000005000000000000000900000000",
            INIT_25 => X"0000003900000000000000490000000000000057000000000000004d00000000",
            INIT_26 => X"0000003100000000000000380000000000000058000000000000005a00000000",
            INIT_27 => X"000000000000000000000007000000000000002a000000000000003b00000000",
            INIT_28 => X"000000350000000000000007000000000000000a000000000000000200000000",
            INIT_29 => X"00000069000000000000005f000000000000004c000000000000005800000000",
            INIT_2A => X"00000069000000000000006e0000000000000065000000000000003800000000",
            INIT_2B => X"000000180000000000000007000000000000000d000000000000003c00000000",
            INIT_2C => X"0000005f00000000000000300000000000000012000000000000000300000000",
            INIT_2D => X"0000004f00000000000000600000000000000073000000000000003700000000",
            INIT_2E => X"000000410000000000000055000000000000005a000000000000004e00000000",
            INIT_2F => X"0000001d00000000000000340000000000000000000000000000000000000000",
            INIT_30 => X"0000002f00000000000000780000000000000036000000000000001300000000",
            INIT_31 => X"0000002f00000000000000480000000000000053000000000000005f00000000",
            INIT_32 => X"0000000000000000000000000000000000000003000000000000000800000000",
            INIT_33 => X"00000020000000000000003f0000000000000041000000000000000000000000",
            INIT_34 => X"00000000000000000000002e000000000000006b000000000000002f00000000",
            INIT_35 => X"0000002b00000000000000260000000000000026000000000000002400000000",
            INIT_36 => X"0000000000000000000000090000000000000007000000000000000000000000",
            INIT_37 => X"0000001d00000000000000250000000000000064000000000000003e00000000",
            INIT_38 => X"0000000000000000000000000000000000000026000000000000004a00000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000001100000000000000070000000000000000000000000000000000000000",
            INIT_3B => X"0000002200000000000000290000000000000015000000000000005500000000",
            INIT_3C => X"0000001400000000000000170000000000000027000000000000005200000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000001c00000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"00000011000000000000002b0000000000000028000000000000001f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000011000000000000001d0000000000000011000000000000003000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_42 => X"0000001e00000000000000150000000000000000000000000000000000000000",
            INIT_43 => X"000000160000000000000013000000000000001e000000000000001500000000",
            INIT_44 => X"0000000f000000000000001f0000000000000016000000000000001a00000000",
            INIT_45 => X"0000001200000000000000150000000000000009000000000000000c00000000",
            INIT_46 => X"0000000000000000000000000000000000000007000000000000000c00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000100000000000000070000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000100000000000000000000000000000000000000000000000300000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000020000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000400000000000000000000000000000010000000000000000000000000",
            INIT_5B => X"0000001c00000000000000000000000000000002000000000000003500000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_5F => X"0000000d00000000000000180000000000000000000000000000000000000000",
            INIT_60 => X"0000000400000000000000040000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000170000000000000007000000000000000000000000",
            INIT_64 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_65 => X"000000000000000000000003000000000000002f000000000000000000000000",
            INIT_66 => X"0000005a00000000000000210000000000000039000000000000003000000000",
            INIT_67 => X"0000000000000000000000000000000000000012000000000000005e00000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_69 => X"0000001c000000000000000f0000000000000000000000000000005700000000",
            INIT_6A => X"000000000000000000000018000000000000002f000000000000000000000000",
            INIT_6B => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000002600000000000000170000000000000000000000000000000100000000",
            INIT_6D => X"0000003f00000000000000210000000000000059000000000000001400000000",
            INIT_6E => X"0000000000000000000000210000000000000021000000000000003500000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"00000021000000000000001c0000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000001f000000000000000a000000000000000c00000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_74 => X"0000000200000000000000000000000000000000000000000000001200000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000a00000000000000000000000000000010000000000000002700000000",
            INIT_78 => X"0000000000000000000000000000000000000003000000000000000c00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE39;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40 : if BRAM_NAME = "samplegold_layersamples_instance40" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000022000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"000000000000000000000000000000000000000f000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000c00000000000000000000000000000000000000000000000300000000",
            INIT_21 => X"0000000000000000000000200000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"00000010000000000000000d0000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"000000000000000000000019000000000000001b000000000000000000000000",
            INIT_26 => X"0000000800000000000000000000000000000000000000000000000400000000",
            INIT_27 => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000001900000000000000090000000000000009000000000000000000000000",
            INIT_2B => X"000000000000000000000000000000000000000a000000000000000f00000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000e00000000000000060000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000002200000000000000150000000000000048000000000000000000000000",
            INIT_38 => X"0000001e000000000000000b000000000000001a000000000000001400000000",
            INIT_39 => X"0000001000000000000000160000000000000015000000000000000000000000",
            INIT_3A => X"0000001f0000000000000000000000000000002a000000000000001600000000",
            INIT_3B => X"0000001d000000000000001d0000000000000014000000000000001100000000",
            INIT_3C => X"00000000000000000000001c0000000000000010000000000000001b00000000",
            INIT_3D => X"0000002000000000000000130000000000000025000000000000000500000000",
            INIT_3E => X"0000002c0000000000000000000000000000000d000000000000000d00000000",
            INIT_3F => X"00000015000000000000001e000000000000001c000000000000002000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000e0000000000000020000000000000000d00000000",
            INIT_41 => X"0000000f0000000000000019000000000000000a000000000000003400000000",
            INIT_42 => X"0000001a00000000000000290000000000000000000000000000001700000000",
            INIT_43 => X"0000000a0000000000000015000000000000001c000000000000002600000000",
            INIT_44 => X"0000000a0000000000000010000000000000001e000000000000001100000000",
            INIT_45 => X"000000160000000000000020000000000000000b000000000000000000000000",
            INIT_46 => X"0000001f0000000000000020000000000000002b000000000000000e00000000",
            INIT_47 => X"0000001d000000000000000c0000000000000018000000000000001f00000000",
            INIT_48 => X"0000000000000000000000170000000000000026000000000000000400000000",
            INIT_49 => X"0000005900000000000000170000000000000016000000000000002600000000",
            INIT_4A => X"0000000c000000000000001b000000000000002f000000000000000c00000000",
            INIT_4B => X"0000000000000000000000100000000000000007000000000000003800000000",
            INIT_4C => X"0000002a00000000000000000000000000000005000000000000002e00000000",
            INIT_4D => X"0000003200000000000000860000000000000020000000000000001800000000",
            INIT_4E => X"0000003100000000000000230000000000000010000000000000001300000000",
            INIT_4F => X"0000002e000000000000003c0000000000000000000000000000000000000000",
            INIT_50 => X"0000002100000000000000240000000000000000000000000000000000000000",
            INIT_51 => X"0000000900000000000000680000000000000006000000000000001900000000",
            INIT_52 => X"0000001400000000000000090000000000000041000000000000001100000000",
            INIT_53 => X"0000000000000000000000100000000000000016000000000000002c00000000",
            INIT_54 => X"0000000000000000000000360000000000000027000000000000000000000000",
            INIT_55 => X"000000000000000000000011000000000000005c000000000000000300000000",
            INIT_56 => X"0000001400000000000000000000000000000017000000000000004700000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_58 => X"000000000000000000000000000000000000004e000000000000004900000000",
            INIT_59 => X"0000005200000000000000000000000000000018000000000000005a00000000",
            INIT_5A => X"0000000000000000000000420000000000000000000000000000003400000000",
            INIT_5B => X"0000004300000000000000150000000000000005000000000000000000000000",
            INIT_5C => X"0000003800000000000000000000000000000000000000000000006900000000",
            INIT_5D => X"0000000e000000000000003e0000000000000000000000000000001000000000",
            INIT_5E => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_5F => X"0000006700000000000000350000000000000014000000000000001200000000",
            INIT_60 => X"0000001300000000000000250000000000000000000000000000000000000000",
            INIT_61 => X"0000002a000000000000001b0000000000000000000000000000000000000000",
            INIT_62 => X"0000000e000000000000000b0000000000000000000000000000000000000000",
            INIT_63 => X"0000001100000000000000330000000000000031000000000000002b00000000",
            INIT_64 => X"0000001b00000000000000180000000000000009000000000000001900000000",
            INIT_65 => X"000000000000000000000017000000000000000c000000000000000000000000",
            INIT_66 => X"00000027000000000000000e000000000000000f000000000000000100000000",
            INIT_67 => X"00000008000000000000003c000000000000000e000000000000003c00000000",
            INIT_68 => X"00000000000000000000001c0000000000000000000000000000002100000000",
            INIT_69 => X"0000000c0000000000000000000000000000002b000000000000001d00000000",
            INIT_6A => X"00000016000000000000002e0000000000000011000000000000000c00000000",
            INIT_6B => X"0000002e00000000000000070000000000000003000000000000002e00000000",
            INIT_6C => X"00000018000000000000000d0000000000000019000000000000000000000000",
            INIT_6D => X"00000005000000000000000b0000000000000003000000000000001300000000",
            INIT_6E => X"00000002000000000000000a000000000000001c000000000000001d00000000",
            INIT_6F => X"00000000000000000000001c0000000000000000000000000000001f00000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"000000000000000000000000000000000000001d000000000000001400000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE40;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41 : if BRAM_NAME = "samplegold_layersamples_instance41" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000002f00000000000000060000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000c000000000000000a0000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000002c000000000000000e0000000000000019000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000001f00000000000000200000000000000019000000000000000700000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000002600000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000002500000000000000180000000000000008000000000000000000000000",
            INIT_23 => X"000000000000000000000000000000000000000c000000000000001e00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000002800000000000000240000000000000000000000000000000000000000",
            INIT_28 => X"0000003500000000000000360000000000000034000000000000003100000000",
            INIT_29 => X"0000000100000000000000180000000000000022000000000000002b00000000",
            INIT_2A => X"0000000d0000000000000001000000000000000a000000000000000700000000",
            INIT_2B => X"0000002e0000000000000039000000000000002e000000000000000a00000000",
            INIT_2C => X"0000003d0000000000000039000000000000003a000000000000003600000000",
            INIT_2D => X"000000010000000000000001000000000000002a000000000000003500000000",
            INIT_2E => X"00000009000000000000001c0000000000000017000000000000000b00000000",
            INIT_2F => X"000000380000000000000036000000000000002b000000000000003600000000",
            INIT_30 => X"000000330000000000000041000000000000003f000000000000003c00000000",
            INIT_31 => X"0000001e00000000000000180000000000000022000000000000003700000000",
            INIT_32 => X"0000001f00000000000000170000000000000014000000000000001e00000000",
            INIT_33 => X"0000004100000000000000360000000000000036000000000000003200000000",
            INIT_34 => X"0000003500000000000000390000000000000043000000000000004500000000",
            INIT_35 => X"000000120000000000000025000000000000002e000000000000003700000000",
            INIT_36 => X"0000002900000000000000180000000000000017000000000000001100000000",
            INIT_37 => X"00000043000000000000003c000000000000003c000000000000003900000000",
            INIT_38 => X"0000002e00000000000000320000000000000034000000000000003100000000",
            INIT_39 => X"00000014000000000000000b000000000000002e000000000000002d00000000",
            INIT_3A => X"0000003100000000000000340000000000000000000000000000001600000000",
            INIT_3B => X"0000003900000000000000250000000000000038000000000000003f00000000",
            INIT_3C => X"0000002a00000000000000200000000000000024000000000000002500000000",
            INIT_3D => X"00000013000000000000000c0000000000000000000000000000000c00000000",
            INIT_3E => X"000000390000000000000040000000000000001d000000000000000d00000000",
            INIT_3F => X"0000002100000000000000200000000000000042000000000000001f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000220000000000000028000000000000001d00000000",
            INIT_41 => X"000000250000000000000011000000000000000a000000000000000000000000",
            INIT_42 => X"0000002d0000000000000027000000000000003a000000000000001300000000",
            INIT_43 => X"0000003000000000000000360000000000000041000000000000003800000000",
            INIT_44 => X"000000000000000000000003000000000000002e000000000000002e00000000",
            INIT_45 => X"00000021000000000000002e0000000000000016000000000000001000000000",
            INIT_46 => X"0000001b0000000000000038000000000000002b000000000000003400000000",
            INIT_47 => X"0000002400000000000000280000000000000033000000000000004500000000",
            INIT_48 => X"0000001500000000000000000000000000000000000000000000000f00000000",
            INIT_49 => X"0000002e000000000000001a0000000000000035000000000000001e00000000",
            INIT_4A => X"0000002e00000000000000300000000000000000000000000000004000000000",
            INIT_4B => X"0000000000000000000000000000000000000044000000000000002d00000000",
            INIT_4C => X"0000003300000000000000120000000000000000000000000000000300000000",
            INIT_4D => X"0000001b000000000000002e0000000000000023000000000000003c00000000",
            INIT_4E => X"0000002100000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_50 => X"0000002b000000000000002e000000000000000e000000000000000000000000",
            INIT_51 => X"0000002100000000000000200000000000000018000000000000003600000000",
            INIT_52 => X"000000000000000000000021000000000000001e000000000000000b00000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"00000032000000000000002e0000000000000012000000000000000d00000000",
            INIT_55 => X"00000032000000000000002c0000000000000014000000000000002e00000000",
            INIT_56 => X"0000000000000000000000030000000000000021000000000000002000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"00000034000000000000001f0000000000000036000000000000001800000000",
            INIT_59 => X"0000002b00000000000000210000000000000018000000000000002200000000",
            INIT_5A => X"0000000f00000000000000180000000000000017000000000000003200000000",
            INIT_5B => X"0000001400000000000000170000000000000014000000000000001600000000",
            INIT_5C => X"0000002e000000000000002f0000000000000036000000000000002400000000",
            INIT_5D => X"0000002a00000000000000340000000000000038000000000000002900000000",
            INIT_5E => X"0000002b0000000000000028000000000000001e000000000000002b00000000",
            INIT_5F => X"0000002500000000000000150000000000000029000000000000002c00000000",
            INIT_60 => X"0000000d0000000000000004000000000000000d000000000000001700000000",
            INIT_61 => X"000000230000000000000008000000000000000c000000000000001000000000",
            INIT_62 => X"00000004000000000000000f0000000000000002000000000000000c00000000",
            INIT_63 => X"0000001800000000000000090000000000000011000000000000000000000000",
            INIT_64 => X"0000000b0000000000000007000000000000000a000000000000000900000000",
            INIT_65 => X"0000002500000000000000210000000000000005000000000000001600000000",
            INIT_66 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000c0000000000000000000000000000002b000000000000000300000000",
            INIT_68 => X"00000012000000000000000d0000000000000007000000000000000600000000",
            INIT_69 => X"000000020000000000000023000000000000000a000000000000000800000000",
            INIT_6A => X"0000000200000000000000000000000000000002000000000000001400000000",
            INIT_6B => X"00000000000000000000000a000000000000000d000000000000001300000000",
            INIT_6C => X"0000000d000000000000000b0000000000000004000000000000000c00000000",
            INIT_6D => X"0000002800000000000000100000000000000000000000000000000100000000",
            INIT_6E => X"0000000500000000000000000000000000000000000000000000000600000000",
            INIT_6F => X"00000005000000000000000a0000000000000008000000000000000000000000",
            INIT_70 => X"0000002200000000000000050000000000000007000000000000001000000000",
            INIT_71 => X"00000000000000000000003b0000000000000000000000000000000000000000",
            INIT_72 => X"0000001300000000000000000000000000000000000000000000000500000000",
            INIT_73 => X"0000000000000000000000160000000000000011000000000000000000000000",
            INIT_74 => X"00000000000000000000000c0000000000000011000000000000002e00000000",
            INIT_75 => X"000000070000000000000000000000000000002c000000000000001600000000",
            INIT_76 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000200000000000000180000000000000000000000000000000f00000000",
            INIT_78 => X"0000002d00000000000000110000000000000006000000000000000f00000000",
            INIT_79 => X"0000000700000000000000070000000000000007000000000000002100000000",
            INIT_7A => X"00000004000000000000000c0000000000000000000000000000001600000000",
            INIT_7B => X"000000000000000000000013000000000000000c000000000000000000000000",
            INIT_7C => X"0000002900000000000000380000000000000005000000000000000600000000",
            INIT_7D => X"0000000300000000000000320000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000280000000000000005000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000025000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE41;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42 : if BRAM_NAME = "samplegold_layersamples_instance42" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000130000000000000025000000000000000e00000000",
            INIT_01 => X"0000000000000000000000090000000000000048000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000062000000000000000000000000",
            INIT_03 => X"0000001200000000000000400000000000000000000000000000001800000000",
            INIT_04 => X"000000000000000000000000000000000000001c000000000000000b00000000",
            INIT_05 => X"000000060000000000000000000000000000000a000000000000005b00000000",
            INIT_06 => X"0000000000000000000000010000000000000010000000000000004600000000",
            INIT_07 => X"00000010000000000000001e0000000000000012000000000000000000000000",
            INIT_08 => X"0000003500000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000002800000000000000070000000000000000000000000000002a00000000",
            INIT_0B => X"00000013000000000000001b0000000000000017000000000000002400000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000250000000000000000000000000000000b000000000000000000000000",
            INIT_0E => X"0000001e000000000000001a0000000000000000000000000000000f00000000",
            INIT_0F => X"0000000d000000000000000f0000000000000024000000000000001e00000000",
            INIT_10 => X"0000000000000000000000050000000000000003000000000000000000000000",
            INIT_11 => X"0000000000000000000000090000000000000000000000000000000a00000000",
            INIT_12 => X"0000000e00000000000000000000000000000007000000000000000000000000",
            INIT_13 => X"0000000c00000000000000120000000000000005000000000000000700000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_17 => X"00000000000000000000000f0000000000000004000000000000000000000000",
            INIT_18 => X"00000013000000000000000c000000000000000b000000000000000000000000",
            INIT_19 => X"00000011000000000000000b0000000000000010000000000000001600000000",
            INIT_1A => X"000000030000000000000006000000000000001b000000000000000000000000",
            INIT_1B => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000400000000000000070000000000000008000000000000000900000000",
            INIT_1D => X"0000000000000000000000030000000000000000000000000000000100000000",
            INIT_1E => X"0000000400000000000000000000000000000004000000000000000000000000",
            INIT_1F => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000000000000000000012000000000000001e000000000000000300000000",
            INIT_31 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000004200000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000040000000000000000000000000000000d00000000",
            INIT_3F => X"0000004000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_48 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000001f00000000000000340000000000000025000000000000000800000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"00000007000000000000001b0000000000000007000000000000000900000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"00000000000000000000000b000000000000000a000000000000000400000000",
            INIT_74 => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000700000000000000020000000000000000000000000000002000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_78 => X"00000001000000000000003a0000000000000035000000000000003b00000000",
            INIT_79 => X"000000000000000000000000000000000000002b000000000000000700000000",
            INIT_7A => X"0000000300000000000000000000000000000000000000000000000200000000",
            INIT_7B => X"0000000100000000000000000000000000000000000000000000000500000000",
            INIT_7C => X"00000005000000000000000e0000000000000028000000000000000000000000",
            INIT_7D => X"0000000d00000000000000030000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000030000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE42;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43 : if BRAM_NAME = "samplegold_layersamples_instance43" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000003000000000000000e0000000000000027000000000000000000000000",
            INIT_01 => X"0000001d000000000000001a0000000000000000000000000000000000000000",
            INIT_02 => X"0000005900000000000000580000000000000057000000000000003f00000000",
            INIT_03 => X"0000000000000000000000110000000000000018000000000000002e00000000",
            INIT_04 => X"000000000000000000000007000000000000000d000000000000002c00000000",
            INIT_05 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000100000000000000070000000000000006000000000000001900000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000004000000000000000e0000000000000000000000000000000100000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000009000000000000000100000000",
            INIT_14 => X"0000000400000000000000020000000000000004000000000000000500000000",
            INIT_15 => X"000000020000000000000005000000000000000b000000000000000500000000",
            INIT_16 => X"00000005000000000000000a0000000000000000000000000000000400000000",
            INIT_17 => X"0000000800000000000000070000000000000000000000000000000000000000",
            INIT_18 => X"0000000a00000000000000090000000000000006000000000000000700000000",
            INIT_19 => X"0000002100000000000000180000000000000007000000000000000000000000",
            INIT_1A => X"000000000000000000000006000000000000000a000000000000000a00000000",
            INIT_1B => X"0000000500000000000000080000000000000009000000000000000000000000",
            INIT_1C => X"0000002c000000000000001f0000000000000009000000000000000400000000",
            INIT_1D => X"0000001500000000000000000000000000000005000000000000001200000000",
            INIT_1E => X"0000000200000000000000000000000000000005000000000000000000000000",
            INIT_1F => X"0000000500000000000000050000000000000008000000000000000800000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_21 => X"00000000000000000000004c0000000000000039000000000000000000000000",
            INIT_22 => X"0000000800000000000000000000000000000001000000000000000800000000",
            INIT_23 => X"0000000300000000000000190000000000000012000000000000000600000000",
            INIT_24 => X"0000004800000000000000190000000000000000000000000000001200000000",
            INIT_25 => X"0000000000000000000000000000000000000035000000000000005a00000000",
            INIT_26 => X"0000000c00000000000000090000000000000021000000000000000600000000",
            INIT_27 => X"000000010000000000000000000000000000000d000000000000000e00000000",
            INIT_28 => X"0000002c000000000000002b0000000000000048000000000000002b00000000",
            INIT_29 => X"00000044000000000000002c0000000000000000000000000000001900000000",
            INIT_2A => X"00000000000000000000004b000000000000000c000000000000002c00000000",
            INIT_2B => X"0000003900000000000000130000000000000000000000000000001700000000",
            INIT_2C => X"00000013000000000000001d0000000000000032000000000000003400000000",
            INIT_2D => X"0000001700000000000000240000000000000033000000000000001400000000",
            INIT_2E => X"000000060000000000000000000000000000000c000000000000003100000000",
            INIT_2F => X"0000002f00000000000000520000000000000017000000000000000000000000",
            INIT_30 => X"0000003700000000000000180000000000000000000000000000001100000000",
            INIT_31 => X"0000001400000000000000000000000000000013000000000000001700000000",
            INIT_32 => X"0000000b00000000000000000000000000000015000000000000001500000000",
            INIT_33 => X"0000000000000000000000300000000000000047000000000000002900000000",
            INIT_34 => X"00000021000000000000002d0000000000000007000000000000000b00000000",
            INIT_35 => X"0000001300000000000000100000000000000000000000000000000000000000",
            INIT_36 => X"0000003400000000000000310000000000000001000000000000001a00000000",
            INIT_37 => X"0000001900000000000000000000000000000030000000000000004a00000000",
            INIT_38 => X"00000000000000000000001d0000000000000011000000000000000c00000000",
            INIT_39 => X"0000000a0000000000000017000000000000000f000000000000000200000000",
            INIT_3A => X"000000020000000000000006000000000000000b000000000000000000000000",
            INIT_3B => X"0000000000000000000000160000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000f000000000000000e0000000000000006000000000000000c00000000",
            INIT_3E => X"000000060000000000000009000000000000000a000000000000000900000000",
            INIT_3F => X"0000000000000000000000000000000000000018000000000000000200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000003200000000000000030000000000000003000000000000000d00000000",
            INIT_44 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_46 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_47 => X"0000000000000000000000260000000000000022000000000000000000000000",
            INIT_48 => X"00000003000000000000000e0000000000000006000000000000000900000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_4A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"000000150000000000000000000000000000000d000000000000003c00000000",
            INIT_4C => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000520000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000090000000000000007000000000000000200000000",
            INIT_50 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000003000000000000000300000000",
            INIT_52 => X"000000190000000000000004000000000000003f000000000000002700000000",
            INIT_53 => X"0000000100000000000000000000000000000003000000000000000a00000000",
            INIT_54 => X"0000000000000000000000000000000000000004000000000000000400000000",
            INIT_55 => X"0000006100000000000000530000000000000045000000000000000a00000000",
            INIT_56 => X"0000002f000000000000000000000000000000a4000000000000003800000000",
            INIT_57 => X"0000000f00000000000000040000000000000000000000000000000a00000000",
            INIT_58 => X"00000049000000000000001b0000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000020000000000000004400000000",
            INIT_5A => X"000000150000000000000013000000000000002400000000000000fb00000000",
            INIT_5B => X"0000001a00000000000000000000000000000007000000000000000100000000",
            INIT_5C => X"00000000000000000000002f0000000000000006000000000000003a00000000",
            INIT_5D => X"000000fd000000000000004e0000000000000000000000000000000000000000",
            INIT_5E => X"0000000700000000000000000000000000000000000000000000006c00000000",
            INIT_5F => X"0000005c0000000000000013000000000000001d000000000000000000000000",
            INIT_60 => X"0000005700000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000ad0000000000000096000000000000005700000000",
            INIT_62 => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_63 => X"000000000000000000000050000000000000000900000000000000b700000000",
            INIT_64 => X"00000098000000000000004c0000000000000034000000000000000000000000",
            INIT_65 => X"0000004c000000000000002f000000000000007a000000000000004100000000",
            INIT_66 => X"000000a400000000000000360000000000000000000000000000007400000000",
            INIT_67 => X"0000000000000000000000000000000000000024000000000000004000000000",
            INIT_68 => X"00000000000000000000007100000000000000c2000000000000004100000000",
            INIT_69 => X"000000920000000000000080000000000000007f000000000000000000000000",
            INIT_6A => X"00000064000000000000003e0000000000000010000000000000000000000000",
            INIT_6B => X"0000005100000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"00000000000000000000002c000000000000000d000000000000010c00000000",
            INIT_6D => X"00000000000000000000001300000000000000b4000000000000002d00000000",
            INIT_6E => X"00000000000000000000004a0000000000000022000000000000000e00000000",
            INIT_6F => X"000000f500000000000000480000000000000000000000000000000b00000000",
            INIT_70 => X"000000000000000000000011000000000000004e000000000000000000000000",
            INIT_71 => X"0000000f00000000000000010000000000000000000000000000008f00000000",
            INIT_72 => X"0000003800000000000000150000000000000041000000000000003b00000000",
            INIT_73 => X"000000000000000000000090000000000000004e000000000000004200000000",
            INIT_74 => X"0000002200000000000000050000000000000041000000000000004500000000",
            INIT_75 => X"0000000d000000000000001b000000000000000e000000000000000100000000",
            INIT_76 => X"00000014000000000000000f000000000000000f000000000000002700000000",
            INIT_77 => X"0000004100000000000000000000000000000016000000000000001600000000",
            INIT_78 => X"0000000000000000000000050000000000000007000000000000003400000000",
            INIT_79 => X"0000000000000000000000000000000000000010000000000000003a00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"00000000000000000000001e000000000000000c000000000000000800000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE43;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44 : if BRAM_NAME = "samplegold_layersamples_instance44" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000000000000e000000000000000d00000000",
            INIT_01 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"000000110000000000000011000000000000000b000000000000000700000000",
            INIT_03 => X"00000027000000000000001a0000000000000000000000000000003200000000",
            INIT_04 => X"0000000700000000000000040000000000000000000000000000000e00000000",
            INIT_05 => X"0000001d000000000000000f000000000000000d000000000000000c00000000",
            INIT_06 => X"0000000000000000000000240000000000000026000000000000002800000000",
            INIT_07 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_08 => X"000000090000000000000006000000000000000a000000000000000900000000",
            INIT_09 => X"0000000e00000000000000060000000000000020000000000000000900000000",
            INIT_0A => X"00000029000000000000004b0000000000000080000000000000004200000000",
            INIT_0B => X"0000000a00000000000000000000000000000003000000000000000900000000",
            INIT_0C => X"0000000c0000000000000007000000000000000a000000000000000c00000000",
            INIT_0D => X"0000000000000000000000460000000000000082000000000000003c00000000",
            INIT_0E => X"0000000000000000000000440000000000000064000000000000000000000000",
            INIT_0F => X"00000009000000000000000c0000000000000000000000000000000400000000",
            INIT_10 => X"0000000000000000000000380000000000000004000000000000000a00000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"00000000000000000000002e000000000000004f000000000000002500000000",
            INIT_13 => X"00000022000000000000000a0000000000000005000000000000000000000000",
            INIT_14 => X"00000003000000000000000d0000000000000000000000000000004500000000",
            INIT_15 => X"0000001100000000000000fa00000000000000f3000000000000007300000000",
            INIT_16 => X"00000061000000000000000c0000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000120000000000000018000000000000000600000000",
            INIT_18 => X"0000006b00000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"00000015000000000000003b00000000000000a8000000000000002f00000000",
            INIT_1B => X"000000000000000000000000000000000000003000000000000000ab00000000",
            INIT_1C => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_1D => X"0000008600000000000000600000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000200000000000000000000000000000001800000000",
            INIT_1F => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000004c00000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_23 => X"0000000f0000000000000024000000000000001b000000000000000000000000",
            INIT_24 => X"0000000400000000000000090000000000000000000000000000000c00000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000001600000000000000000000000000000000000000000000000100000000",
            INIT_27 => X"00000000000000000000004d0000000000000078000000000000005f00000000",
            INIT_28 => X"000000080000000000000033000000000000000f000000000000000000000000",
            INIT_29 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000b000000000000000e0000000000000000000000000000000000000000",
            INIT_2E => X"000000260000000000000023000000000000004a000000000000001200000000",
            INIT_2F => X"00000000000000000000000a0000000000000011000000000000001f00000000",
            INIT_30 => X"0000000800000000000000070000000000000000000000000000000000000000",
            INIT_31 => X"00000145000000000000013c000000000000012f000000000000000c00000000",
            INIT_32 => X"0000011900000000000001270000000000000141000000000000014b00000000",
            INIT_33 => X"000000ba00000000000000bb00000000000000f0000000000000010c00000000",
            INIT_34 => X"0000008a000000000000003e000000000000005c000000000000009c00000000",
            INIT_35 => X"0000011700000000000001200000000000000126000000000000013400000000",
            INIT_36 => X"000000db00000000000000e400000000000000ec000000000000010200000000",
            INIT_37 => X"00000084000000000000009d00000000000000b900000000000000ca00000000",
            INIT_38 => X"000000e3000000000000009c0000000000000047000000000000002d00000000",
            INIT_39 => X"000000cc00000000000000d800000000000000de00000000000000df00000000",
            INIT_3A => X"000000bc00000000000000c100000000000000c500000000000000c400000000",
            INIT_3B => X"000000460000000000000029000000000000006d00000000000000b200000000",
            INIT_3C => X"000000b900000000000000b300000000000000a3000000000000007900000000",
            INIT_3D => X"000000c300000000000000c000000000000000bd00000000000000bb00000000",
            INIT_3E => X"000000a800000000000000bc00000000000000c200000000000000bf00000000",
            INIT_3F => X"000000a5000000000000007e0000000000000017000000000000004700000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000bf00000000000000bd00000000000000af00000000000000a900000000",
            INIT_41 => X"000000a300000000000000b900000000000000bd00000000000000bf00000000",
            INIT_42 => X"00000029000000000000008c000000000000008d00000000000000a100000000",
            INIT_43 => X"000000a100000000000000a2000000000000008a000000000000003100000000",
            INIT_44 => X"000000bd00000000000000bf00000000000000be00000000000000ba00000000",
            INIT_45 => X"0000003c000000000000004f000000000000006e00000000000000a700000000",
            INIT_46 => X"0000005500000000000000000000000000000000000000000000002e00000000",
            INIT_47 => X"000000c00000000000000093000000000000006f000000000000001900000000",
            INIT_48 => X"0000007c00000000000000a200000000000000be00000000000000c000000000",
            INIT_49 => X"00000017000000000000001c0000000000000022000000000000003800000000",
            INIT_4A => X"0000002700000000000000330000000000000000000000000000000000000000",
            INIT_4B => X"000000be00000000000000be000000000000005f000000000000001f00000000",
            INIT_4C => X"0000001e00000000000000310000000000000070000000000000008500000000",
            INIT_4D => X"0000000300000000000000000000000000000000000000000000000b00000000",
            INIT_4E => X"0000000000000000000000170000000000000035000000000000000000000000",
            INIT_4F => X"0000005c000000000000009000000000000000bd000000000000001100000000",
            INIT_50 => X"0000000000000000000000000000000000000011000000000000000600000000",
            INIT_51 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000070000000000000013000000000000004500000000",
            INIT_53 => X"0000000000000000000000340000000000000042000000000000009800000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000001300000000",
            INIT_55 => X"000000000000000000000000000000000000001b000000000000000000000000",
            INIT_56 => X"0000007500000000000000220000000000000000000000000000000000000000",
            INIT_57 => X"0000000700000000000000090000000000000000000000000000000800000000",
            INIT_58 => X"0000002a00000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_5A => X"00000001000000000000006b0000000000000019000000000000000a00000000",
            INIT_5B => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_5C => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_5D => X"0000001f00000000000000000000000000000000000000000000000900000000",
            INIT_5E => X"000000000000000000000000000000000000004e000000000000001100000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000d0000000000000000000000000000002b000000000000000000000000",
            INIT_61 => X"0000001900000000000000110000000000000000000000000000000f00000000",
            INIT_62 => X"0000000000000000000000000000000000000010000000000000004c00000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000001700000000000000020000000000000000000000000000000000000000",
            INIT_65 => X"00000045000000000000000a0000000000000006000000000000000100000000",
            INIT_66 => X"0000000000000000000000020000000000000000000000000000001800000000",
            INIT_67 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000700000000000000070000000000000006000000000000000000000000",
            INIT_69 => X"0000007800000000000000820000000000000002000000000000000600000000",
            INIT_6A => X"0000007500000000000000770000000000000083000000000000008800000000",
            INIT_6B => X"0000004a000000000000006e0000000000000066000000000000007900000000",
            INIT_6C => X"0000004100000000000000150000000000000046000000000000005100000000",
            INIT_6D => X"0000007300000000000000780000000000000087000000000000004400000000",
            INIT_6E => X"00000070000000000000006d0000000000000077000000000000007a00000000",
            INIT_6F => X"00000055000000000000005a0000000000000061000000000000006200000000",
            INIT_70 => X"0000004e000000000000004b0000000000000008000000000000002f00000000",
            INIT_71 => X"0000006b000000000000006e0000000000000062000000000000006500000000",
            INIT_72 => X"0000006000000000000000650000000000000066000000000000006a00000000",
            INIT_73 => X"00000001000000000000003b000000000000005f000000000000005d00000000",
            INIT_74 => X"000000630000000000000042000000000000004f000000000000002800000000",
            INIT_75 => X"0000006a00000000000000630000000000000065000000000000006900000000",
            INIT_76 => X"0000005d0000000000000060000000000000006b000000000000006700000000",
            INIT_77 => X"00000049000000000000003a0000000000000000000000000000005000000000",
            INIT_78 => X"0000006b00000000000000650000000000000051000000000000004900000000",
            INIT_79 => X"00000066000000000000006f0000000000000066000000000000006a00000000",
            INIT_7A => X"0000002400000000000000570000000000000059000000000000005300000000",
            INIT_7B => X"0000005700000000000000420000000000000029000000000000000000000000",
            INIT_7C => X"00000065000000000000006a0000000000000069000000000000005300000000",
            INIT_7D => X"0000004a0000000000000063000000000000006a000000000000006400000000",
            INIT_7E => X"0000000000000000000000000000000000000012000000000000002100000000",
            INIT_7F => X"000000500000000000000028000000000000003f000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE44;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45 : if BRAM_NAME = "samplegold_layersamples_instance45" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000064000000000000005f0000000000000069000000000000006b00000000",
            INIT_01 => X"0000000000000000000000000000000000000023000000000000005f00000000",
            INIT_02 => X"0000000000000000000000360000000000000072000000000000000e00000000",
            INIT_03 => X"0000006c000000000000003d0000000000000022000000000000000200000000",
            INIT_04 => X"00000005000000000000003e0000000000000063000000000000006300000000",
            INIT_05 => X"0000003b00000000000000120000000000000000000000000000002f00000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000004400000000",
            INIT_07 => X"0000006500000000000000680000000000000036000000000000001f00000000",
            INIT_08 => X"0000001700000000000000000000000000000020000000000000002200000000",
            INIT_09 => X"000000000000000000000000000000000000003e000000000000005b00000000",
            INIT_0A => X"0000004c000000000000003c0000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000007c0000000000000073000000000000001800000000",
            INIT_0C => X"0000007300000000000000310000000000000000000000000000001f00000000",
            INIT_0D => X"0000000c00000000000000000000000000000000000000000000000600000000",
            INIT_0E => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000018000000000000009500000000",
            INIT_10 => X"0000000000000000000000720000000000000030000000000000000000000000",
            INIT_11 => X"0000006900000000000000210000000000000000000000000000000000000000",
            INIT_12 => X"0000005d00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000001e00000000000000000000000000000000000000000000001500000000",
            INIT_14 => X"0000000000000000000000000000000000000056000000000000003300000000",
            INIT_15 => X"00000006000000000000005d0000000000000000000000000000001200000000",
            INIT_16 => X"0000001800000000000000500000000000000015000000000000000000000000",
            INIT_17 => X"0000000b000000000000003b0000000000000000000000000000000600000000",
            INIT_18 => X"0000002b00000000000000000000000000000000000000000000002f00000000",
            INIT_19 => X"00000000000000000000002f0000000000000017000000000000000000000000",
            INIT_1A => X"000000000000000000000029000000000000003e000000000000002600000000",
            INIT_1B => X"0000000300000000000000080000000000000017000000000000000000000000",
            INIT_1C => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_1D => X"0000001b00000000000000020000000000000014000000000000000000000000",
            INIT_1E => X"000000000000000000000006000000000000000b000000000000003500000000",
            INIT_1F => X"0000000600000000000000070000000000000008000000000000000800000000",
            INIT_20 => X"0000000000000000000000000000000000000034000000000000000700000000",
            INIT_21 => X"000000ac000000000000001a0000000000000011000000000000001000000000",
            INIT_22 => X"000000cc00000000000000cd00000000000000c400000000000000bf00000000",
            INIT_23 => X"000000a700000000000000b100000000000000b600000000000000bf00000000",
            INIT_24 => X"00000041000000000000007a0000000000000088000000000000008b00000000",
            INIT_25 => X"000000b100000000000000c40000000000000068000000000000003200000000",
            INIT_26 => X"000000a800000000000000b800000000000000c100000000000000ba00000000",
            INIT_27 => X"00000086000000000000008f000000000000009b00000000000000a100000000",
            INIT_28 => X"0000002600000000000000320000000000000053000000000000007200000000",
            INIT_29 => X"000000a400000000000000aa000000000000009c000000000000007200000000",
            INIT_2A => X"000000910000000000000090000000000000009a00000000000000a200000000",
            INIT_2B => X"0000003600000000000000820000000000000083000000000000008800000000",
            INIT_2C => X"0000007100000000000000400000000000000027000000000000001800000000",
            INIT_2D => X"0000008b000000000000008b000000000000008d000000000000008900000000",
            INIT_2E => X"0000007a0000000000000081000000000000008d000000000000008c00000000",
            INIT_2F => X"000000180000000000000039000000000000006f000000000000007400000000",
            INIT_30 => X"000000820000000000000082000000000000007a000000000000005500000000",
            INIT_31 => X"0000008d000000000000008f000000000000008f000000000000008f00000000",
            INIT_32 => X"0000004600000000000000680000000000000060000000000000007900000000",
            INIT_33 => X"0000004e00000000000000000000000000000000000000000000001800000000",
            INIT_34 => X"00000090000000000000008e0000000000000078000000000000007300000000",
            INIT_35 => X"000000420000000000000086000000000000008d000000000000008d00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"00000034000000000000001f0000000000000000000000000000000000000000",
            INIT_38 => X"0000008f000000000000008f0000000000000090000000000000006d00000000",
            INIT_39 => X"000000260000000000000031000000000000003e000000000000008600000000",
            INIT_3A => X"0000000000000000000000000000000000000034000000000000003100000000",
            INIT_3B => X"0000004200000000000000250000000000000000000000000000000000000000",
            INIT_3C => X"0000002b00000000000000680000000000000091000000000000008f00000000",
            INIT_3D => X"0000000000000000000000050000000000000003000000000000001200000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000009000000000000000000000000000000019000000000000000a00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000005000000000000000f000000000000002e000000000000008200000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_42 => X"00000015000000000000001f0000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000950000000000000000000000000000000000000000",
            INIT_44 => X"0000000900000000000000120000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000110000000000000068000000000000000000000000",
            INIT_48 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_49 => X"00000012000000000000002d0000000000000000000000000000000000000000",
            INIT_4A => X"0000002f00000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000007600000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_4E => X"0000005900000000000000190000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000001600000000000000440000000000000021000000000000001800000000",
            INIT_53 => X"000000200000000000000008000000000000000a000000000000000000000000",
            INIT_54 => X"00000000000000000000002e0000000000000027000000000000002200000000",
            INIT_55 => X"0000002200000000000000210000000000000011000000000000000c00000000",
            INIT_56 => X"00000000000000000000001e0000000000000035000000000000001700000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000c000000000000000b000000000000000b000000000000000200000000",
            INIT_59 => X"0000000a00000000000000100000000000000012000000000000001c00000000",
            INIT_5A => X"00000055000000000000004c000000000000003f000000000000002600000000",
            INIT_5B => X"0000004a000000000000004c0000000000000051000000000000005900000000",
            INIT_5C => X"00000030000000000000002b0000000000000042000000000000004000000000",
            INIT_5D => X"0000004c000000000000001a000000000000001b000000000000002f00000000",
            INIT_5E => X"0000004f0000000000000053000000000000004f000000000000004500000000",
            INIT_5F => X"00000032000000000000003b000000000000003f000000000000004600000000",
            INIT_60 => X"0000000a000000000000001a0000000000000014000000000000002900000000",
            INIT_61 => X"000000530000000000000057000000000000001c000000000000000000000000",
            INIT_62 => X"0000002c00000000000000340000000000000041000000000000004700000000",
            INIT_63 => X"0000001f00000000000000230000000000000024000000000000002b00000000",
            INIT_64 => X"0000000100000000000000000000000000000025000000000000002c00000000",
            INIT_65 => X"00000029000000000000002a000000000000002b000000000000002500000000",
            INIT_66 => X"0000001c00000000000000280000000000000026000000000000002800000000",
            INIT_67 => X"00000029000000000000001e0000000000000015000000000000001200000000",
            INIT_68 => X"0000002b00000000000000270000000000000010000000000000000000000000",
            INIT_69 => X"0000002e000000000000002d000000000000002b000000000000002500000000",
            INIT_6A => X"0000001300000000000000280000000000000030000000000000002c00000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000002a00000000000000270000000000000026000000000000001a00000000",
            INIT_6D => X"00000020000000000000002c000000000000002b000000000000002c00000000",
            INIT_6E => X"0000008a0000000000000054000000000000000a000000000000000000000000",
            INIT_6F => X"0000002e00000000000000000000000000000000000000000000009700000000",
            INIT_70 => X"0000002d000000000000002b0000000000000023000000000000000f00000000",
            INIT_71 => X"0000003a00000000000000270000000000000025000000000000003200000000",
            INIT_72 => X"0000000000000000000000130000000000000024000000000000002900000000",
            INIT_73 => X"0000003200000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000001e000000000000002e000000000000002e000000000000002200000000",
            INIT_75 => X"0000000000000000000000070000000000000006000000000000000a00000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"000000000000000000000000000000000000000e000000000000006b00000000",
            INIT_78 => X"0000002100000000000000010000000000000016000000000000003100000000",
            INIT_79 => X"0000000000000000000000000000000000000003000000000000002500000000",
            INIT_7A => X"0000000600000000000000000000000000000013000000000000001f00000000",
            INIT_7B => X"0000001d00000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001400000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000300000000000000000000000000000000000000000000000f00000000",
            INIT_7E => X"000000000000000000000000000000000000008c000000000000006d00000000",
            INIT_7F => X"00000086000000000000002f0000000000000022000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE45;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46 : if BRAM_NAME = "samplegold_layersamples_instance46" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000060000000000000000000000000000002300000000",
            INIT_01 => X"0000003100000000000000300000000000000000000000000000000000000000",
            INIT_02 => X"00000037000000000000002e0000000000000053000000000000000100000000",
            INIT_03 => X"0000000000000000000000000000000000000029000000000000005600000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_05 => X"0000000000000000000000000000000000000030000000000000000000000000",
            INIT_06 => X"000000010000000000000027000000000000000f000000000000000600000000",
            INIT_07 => X"0000000000000000000000000000000000000003000000000000001d00000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_0A => X"0000000900000000000000070000000000000035000000000000002c00000000",
            INIT_0B => X"0000004f0000000000000047000000000000003e000000000000001f00000000",
            INIT_0C => X"0000007a0000000000000090000000000000008b000000000000007e00000000",
            INIT_0D => X"000000120000000000000005000000000000000e000000000000000000000000",
            INIT_0E => X"0000000000000000000000130000000000000000000000000000001000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000001000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"000000000000000000000000000000000000000e000000000000003300000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000001c0000000000000007000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000002000000000000001200000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000001e000000000000000b0000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000006300000000000000490000000000000000000000000000000000000000",
            INIT_27 => X"00000002000000000000009d00000000000000ab000000000000008600000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000002d00000000000000410000000000000064000000000000003600000000",
            INIT_2B => X"00000000000000000000007800000000000000d9000000000000004000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_2D => X"00000024000000000000002c0000000000000000000000000000000000000000",
            INIT_2E => X"00000076000000000000002f000000000000001f000000000000003000000000",
            INIT_2F => X"00000000000000000000001600000000000000ba00000000000000e800000000",
            INIT_30 => X"0000000500000000000000000000000000000000000000000000001f00000000",
            INIT_31 => X"0000004500000000000000200000000000000036000000000000004900000000",
            INIT_32 => X"000000e1000000000000010200000000000000ee00000000000000bf00000000",
            INIT_33 => X"0000007e00000000000000220000000000000016000000000000005100000000",
            INIT_34 => X"00000027000000000000003e000000000000003c000000000000000000000000",
            INIT_35 => X"000000df00000000000000530000000000000009000000000000000c00000000",
            INIT_36 => X"0000009800000000000000f100000000000000d600000000000000e600000000",
            INIT_37 => X"000000000000000000000091000000000000009f000000000000007900000000",
            INIT_38 => X"00000000000000000000001c0000000000000087000000000000009800000000",
            INIT_39 => X"000000c500000000000000d60000000000000056000000000000000a00000000",
            INIT_3A => X"000000c700000000000000ce0000000000000037000000000000005f00000000",
            INIT_3B => X"000000290000000000000000000000000000005200000000000000a500000000",
            INIT_3C => X"0000004000000000000000000000000000000016000000000000007700000000",
            INIT_3D => X"00000017000000000000009300000000000000d8000000000000009800000000",
            INIT_3E => X"0000005b00000000000000a8000000000000002c000000000000001200000000",
            INIT_3F => X"00000075000000000000002e0000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000009e00000000000000670000000000000034000000000000002200000000",
            INIT_41 => X"00000023000000000000002e000000000000007e00000000000000d700000000",
            INIT_42 => X"0000000000000000000000320000000000000075000000000000000000000000",
            INIT_43 => X"0000003b0000000000000054000000000000001c000000000000000000000000",
            INIT_44 => X"000000a2000000000000009d000000000000008d000000000000005600000000",
            INIT_45 => X"0000000000000000000000430000000000000031000000000000007200000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000e00000000",
            INIT_47 => X"0000000000000000000000080000000000000019000000000000000300000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_49 => X"0000000000000000000000000000000000000029000000000000001600000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000001500000000000000160000000000000011000000000000000000000000",
            INIT_4C => X"0000002600000000000000170000000000000011000000000000000f00000000",
            INIT_4D => X"0000000100000000000000390000000000000000000000000000000c00000000",
            INIT_4E => X"0000001800000000000000050000000000000008000000000000000000000000",
            INIT_4F => X"0000000a000000000000000e0000000000000012000000000000001600000000",
            INIT_50 => X"0000000000000000000000000000000000000003000000000000000700000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_52 => X"0000000d000000000000000d0000000000000028000000000000002600000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_54 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000048000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"00000000000000000000001f000000000000003b000000000000000000000000",
            INIT_60 => X"0000000300000000000000000000000000000000000000000000005d00000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"000000740000000000000060000000000000004f000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000002d00000000",
            INIT_64 => X"000000000000000000000009000000000000000e000000000000003100000000",
            INIT_65 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"00000000000000000000006e0000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000180000000000000039000000000000000c000000000000003d00000000",
            INIT_6A => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_6B => X"000000000000000000000000000000000000003e000000000000002d00000000",
            INIT_6C => X"0000003900000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"000000000000000000000000000000000000002a000000000000000500000000",
            INIT_6E => X"0000000000000000000000810000000000000000000000000000000000000000",
            INIT_6F => X"0000004200000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001e00000000000000020000000000000077000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_72 => X"0000000000000000000000750000000000000059000000000000007a00000000",
            INIT_73 => X"00000014000000000000007a000000000000004c000000000000002900000000",
            INIT_74 => X"0000000000000000000000250000000000000000000000000000000000000000",
            INIT_75 => X"0000005d00000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000002b0000000000000001000000000000000000000000",
            INIT_77 => X"0000000000000000000000090000000000000000000000000000006100000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"00000000000000000000003b0000000000000000000000000000000000000000",
            INIT_7A => X"0000004000000000000000180000000000000025000000000000000000000000",
            INIT_7B => X"0000003900000000000000020000000000000000000000000000000500000000",
            INIT_7C => X"0000009d00000000000000930000000000000069000000000000003800000000",
            INIT_7D => X"000000190000000000000000000000000000004800000000000000a500000000",
            INIT_7E => X"000000000000000000000007000000000000003f000000000000002100000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE46;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47 : if BRAM_NAME = "samplegold_layersamples_instance47" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000b0000000000000020000000000000001e000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000180000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000001c000000000000000d0000000000000000000000000000000000000000",
            INIT_1B => X"0000004600000000000000690000000000000023000000000000001d00000000",
            INIT_1C => X"000000000000000000000013000000000000000b000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000001200000000000000020000000000000011000000000000000000000000",
            INIT_1F => X"00000000000000000000001f000000000000003b000000000000001100000000",
            INIT_20 => X"00000000000000000000000d000000000000001b000000000000000000000000",
            INIT_21 => X"00000001000000000000001d0000000000000000000000000000000000000000",
            INIT_22 => X"0000001c000000000000003c0000000000000046000000000000002e00000000",
            INIT_23 => X"0000000e00000000000000000000000000000002000000000000001a00000000",
            INIT_24 => X"0000000d00000000000000000000000000000014000000000000001d00000000",
            INIT_25 => X"0000003500000000000000000000000000000030000000000000000000000000",
            INIT_26 => X"0000001600000000000000280000000000000037000000000000007600000000",
            INIT_27 => X"0000001800000000000000140000000000000000000000000000002700000000",
            INIT_28 => X"00000000000000000000002c0000000000000004000000000000000a00000000",
            INIT_29 => X"000000780000000000000036000000000000000d000000000000001400000000",
            INIT_2A => X"0000005500000000000000050000000000000006000000000000002e00000000",
            INIT_2B => X"0000000000000000000000110000000000000016000000000000008100000000",
            INIT_2C => X"00000000000000000000001f0000000000000028000000000000000000000000",
            INIT_2D => X"000000220000000000000069000000000000004b000000000000002500000000",
            INIT_2E => X"00000069000000000000000b0000000000000024000000000000000000000000",
            INIT_2F => X"0000000000000000000000080000000000000000000000000000003500000000",
            INIT_30 => X"0000004200000000000000000000000000000031000000000000002600000000",
            INIT_31 => X"00000000000000000000002b0000000000000053000000000000002600000000",
            INIT_32 => X"0000005200000000000000260000000000000000000000000000003100000000",
            INIT_33 => X"0000002000000000000000000000000000000015000000000000000000000000",
            INIT_34 => X"0000005100000000000000540000000000000025000000000000002d00000000",
            INIT_35 => X"0000004600000000000000000000000000000049000000000000004f00000000",
            INIT_36 => X"0000001200000000000000310000000000000006000000000000001000000000",
            INIT_37 => X"0000001c000000000000000b0000000000000000000000000000001900000000",
            INIT_38 => X"0000001a000000000000001c000000000000001d000000000000001000000000",
            INIT_39 => X"0000001700000000000000390000000000000013000000000000001800000000",
            INIT_3A => X"0000001a00000000000000150000000000000014000000000000000200000000",
            INIT_3B => X"0000000b00000000000000190000000000000013000000000000002b00000000",
            INIT_3C => X"00000000000000000000000c0000000000000002000000000000000000000000",
            INIT_3D => X"0000000500000000000000000000000000000000000000000000000800000000",
            INIT_3E => X"0000000600000000000000080000000000000014000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000500000000000000000000000000000007000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000014000000000000000700000000",
            INIT_42 => X"0000000000000000000000040000000000000007000000000000003d00000000",
            INIT_43 => X"0000000400000000000000030000000000000000000000000000000000000000",
            INIT_44 => X"0000000f000000000000000c0000000000000009000000000000000700000000",
            INIT_45 => X"0000003400000000000000090000000000000000000000000000003000000000",
            INIT_46 => X"0000000600000000000000060000000000000004000000000000000500000000",
            INIT_47 => X"0000000e000000000000000a000000000000000a000000000000000300000000",
            INIT_48 => X"0000000000000000000000150000000000000012000000000000001100000000",
            INIT_49 => X"00000000000000000000000a0000000000000019000000000000002000000000",
            INIT_4A => X"0000000300000000000000040000000000000006000000000000000b00000000",
            INIT_4B => X"0000000e000000000000001c0000000000000017000000000000000c00000000",
            INIT_4C => X"0000002b00000000000000000000000000000004000000000000001a00000000",
            INIT_4D => X"0000000900000000000000080000000000000004000000000000000d00000000",
            INIT_4E => X"0000001200000000000000040000000000000004000000000000000400000000",
            INIT_4F => X"0000002c0000000000000033000000000000004c000000000000002a00000000",
            INIT_50 => X"000000250000000000000000000000000000003c000000000000000000000000",
            INIT_51 => X"0000000200000000000000050000000000000005000000000000000800000000",
            INIT_52 => X"0000000e0000000000000034000000000000000b000000000000000000000000",
            INIT_53 => X"0000006000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000001c00000000000000000000000000000000000000000000006c00000000",
            INIT_55 => X"0000001600000000000000000000000000000003000000000000000700000000",
            INIT_56 => X"0000000000000000000000250000000000000000000000000000001900000000",
            INIT_57 => X"0000001f000000000000009c000000000000005f000000000000002e00000000",
            INIT_58 => X"00000051000000000000001b0000000000000000000000000000000000000000",
            INIT_59 => X"000000090000000000000003000000000000000e000000000000000100000000",
            INIT_5A => X"000000950000000000000041000000000000001f000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000006000000000000002200000000",
            INIT_5C => X"0000000c00000000000000430000000000000051000000000000002200000000",
            INIT_5D => X"0000000000000000000000230000000000000000000000000000008000000000",
            INIT_5E => X"0000001000000000000000370000000000000086000000000000003600000000",
            INIT_5F => X"000000390000000000000000000000000000000b000000000000000000000000",
            INIT_60 => X"0000000e00000000000000450000000000000000000000000000001500000000",
            INIT_61 => X"0000004700000000000000000000000000000007000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000020000000000000009300000000",
            INIT_63 => X"0000000000000000000000000000000000000061000000000000002b00000000",
            INIT_64 => X"00000025000000000000000e000000000000001a000000000000000000000000",
            INIT_65 => X"0000007c00000000000000600000000000000028000000000000000000000000",
            INIT_66 => X"00000000000000000000001e0000000000000000000000000000001700000000",
            INIT_67 => X"0000000200000000000000000000000000000020000000000000006700000000",
            INIT_68 => X"000000000000000000000032000000000000001e000000000000001200000000",
            INIT_69 => X"00000009000000000000006a000000000000003a000000000000005a00000000",
            INIT_6A => X"0000001c00000000000000000000000000000039000000000000000000000000",
            INIT_6B => X"0000001600000000000000220000000000000000000000000000005300000000",
            INIT_6C => X"000000300000000000000000000000000000001e000000000000002200000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_6E => X"0000002100000000000000000000000000000000000000000000004d00000000",
            INIT_6F => X"0000000300000000000000130000000000000022000000000000000000000000",
            INIT_70 => X"0000001c00000000000000190000000000000012000000000000000900000000",
            INIT_71 => X"0000003d00000000000000100000000000000012000000000000001800000000",
            INIT_72 => X"0000001c000000000000001a0000000000000000000000000000000400000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE47;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48 : if BRAM_NAME = "samplegold_layersamples_instance48" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000002b000000000000002b0000000000000019000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000002700000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"00000000000000000000003b0000000000000015000000000000000000000000",
            INIT_08 => X"00000002000000000000002a0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000f00000000000000020000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000006e00000000000000d1000000000000006d000000000000000000000000",
            INIT_10 => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000005100000000",
            INIT_12 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_14 => X"0000001000000000000000680000000000000031000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000045000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000002a00000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"000000000000000000000000000000000000001f000000000000003000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00000004000000000000001f0000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000000000000000000004e0000000000000050000000000000001100000000",
            INIT_22 => X"0000001900000000000000110000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_28 => X"000000250000000000000038000000000000001d000000000000000000000000",
            INIT_29 => X"0000000f0000000000000012000000000000001e000000000000002400000000",
            INIT_2A => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000008400000000000000800000000000000013000000000000000f00000000",
            INIT_2C => X"0000007400000000000000850000000000000089000000000000008900000000",
            INIT_2D => X"0000003c000000000000005a0000000000000064000000000000006d00000000",
            INIT_2E => X"00000000000000000000000e0000000000000028000000000000003800000000",
            INIT_2F => X"000000760000000000000076000000000000007b000000000000001f00000000",
            INIT_30 => X"0000005200000000000000550000000000000061000000000000006c00000000",
            INIT_31 => X"0000002d00000000000000360000000000000043000000000000004b00000000",
            INIT_32 => X"0000002c00000000000000000000000000000000000000000000002100000000",
            INIT_33 => X"0000004900000000000000490000000000000050000000000000005600000000",
            INIT_34 => X"0000003f00000000000000420000000000000041000000000000004300000000",
            INIT_35 => X"0000000000000000000000240000000000000037000000000000003c00000000",
            INIT_36 => X"000000330000000000000036000000000000001c000000000000000000000000",
            INIT_37 => X"0000003f000000000000003c000000000000003d000000000000003900000000",
            INIT_38 => X"0000004000000000000000440000000000000042000000000000004200000000",
            INIT_39 => X"000000180000000000000000000000000000000c000000000000003a00000000",
            INIT_3A => X"0000003d0000000000000036000000000000002e000000000000003200000000",
            INIT_3B => X"00000041000000000000003e000000000000003f000000000000003f00000000",
            INIT_3C => X"00000038000000000000002e0000000000000038000000000000003f00000000",
            INIT_3D => X"0000002b00000000000000270000000000000000000000000000000000000000",
            INIT_3E => X"0000003f000000000000003f000000000000003c000000000000002c00000000",
            INIT_3F => X"0000002400000000000000200000000000000033000000000000003e00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000d000000000000000d0000000000000038000000000000003500000000",
            INIT_41 => X"0000002500000000000000260000000000000000000000000000001900000000",
            INIT_42 => X"0000002e00000000000000400000000000000040000000000000004000000000",
            INIT_43 => X"0000000000000000000000000000000000000019000000000000002800000000",
            INIT_44 => X"0000002400000000000000150000000000000000000000000000000000000000",
            INIT_45 => X"0000003f00000000000000080000000000000000000000000000000000000000",
            INIT_46 => X"0000000c00000000000000280000000000000021000000000000003f00000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"00000000000000000000002a0000000000000020000000000000001a00000000",
            INIT_49 => X"00000028000000000000003f0000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_4B => X"0000001b000000000000002e000000000000001d000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000003500000000",
            INIT_4D => X"0000001c00000000000000250000000000000024000000000000001400000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"000000000000000000000021000000000000000a000000000000001500000000",
            INIT_50 => X"00000017000000000000000f000000000000001a000000000000001500000000",
            INIT_51 => X"0000000000000000000000000000000000000011000000000000001c00000000",
            INIT_52 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000003000000000",
            INIT_54 => X"0000001a00000000000000000000000000000009000000000000000c00000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000002200000000000000100000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000040000000000000000000000000000000500000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000100000000000000003000000000000000200000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_66 => X"0000002900000000000000000000000000000003000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000190000000000000027000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000600000000000000000000000000000016000000000000001b00000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"00000000000000000000003e0000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000b0000000000000014000000000000002f000000000000002400000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"00000000000000000000000b0000000000000012000000000000000000000000",
            INIT_79 => X"0000000f0000000000000000000000000000008a000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000a00000000000000050000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_7D => X"0000000300000000000000000000000000000044000000000000006000000000",
            INIT_7E => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000190000000000000000000000000000001f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE48;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49 : if BRAM_NAME = "samplegold_layersamples_instance49" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000005d00000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000002000000000000001d00000000",
            INIT_02 => X"0000003300000000000000000000000000000025000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_04 => X"00000000000000000000003f000000000000001a000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000320000000000000000000000000000007800000000",
            INIT_07 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000800000000000000100000000000000001000000000000000000000000",
            INIT_09 => X"0000001e00000000000000000000000000000000000000000000001f00000000",
            INIT_0A => X"0000000000000000000000000000000000000019000000000000002800000000",
            INIT_0B => X"0000000900000000000000130000000000000040000000000000000000000000",
            INIT_0C => X"0000003900000000000000190000000000000008000000000000000000000000",
            INIT_0D => X"0000004200000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_0F => X"0000000000000000000000200000000000000004000000000000007800000000",
            INIT_10 => X"0000000000000000000000030000000000000059000000000000000000000000",
            INIT_11 => X"00000000000000000000002c0000000000000000000000000000000000000000",
            INIT_12 => X"0000006d00000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000000000001e0000000000000030000000000000000000000000",
            INIT_14 => X"000000000000000000000000000000000000000a000000000000003c00000000",
            INIT_15 => X"000000000000000000000000000000000000000c000000000000000d00000000",
            INIT_16 => X"00000000000000000000000b0000000000000000000000000000000000000000",
            INIT_17 => X"0000001000000000000000140000000000000031000000000000001200000000",
            INIT_18 => X"0000001100000000000000130000000000000000000000000000001200000000",
            INIT_19 => X"00000020000000000000001c000000000000001e000000000000002c00000000",
            INIT_1A => X"0000001200000000000000030000000000000020000000000000001e00000000",
            INIT_1B => X"00000013000000000000001c000000000000001d000000000000002100000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"00000000000000000000000b0000000000000010000000000000000100000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000001700000000000000140000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000080000000000000025000000000000001c00000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000001d0000000000000021000000000000001f000000000000000000000000",
            INIT_29 => X"0000000000000000000000110000000000000015000000000000001400000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000001400000000000000040000000000000005000000000000000700000000",
            INIT_2D => X"00000017000000000000001c000000000000001e000000000000002000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000c00000000000000000000000000000007000000000000000000000000",
            INIT_30 => X"0000001b00000000000000220000000000000013000000000000000000000000",
            INIT_31 => X"000000020000000000000021000000000000001f000000000000001b00000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000150000000000000014000000000000001f000000000000001100000000",
            INIT_35 => X"00000000000000000000000d0000000000000018000000000000001f00000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"000000210000000000000013000000000000000a000000000000000a00000000",
            INIT_39 => X"00000000000000000000000a000000000000001d000000000000001c00000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000022000000000000001c000000000000001b000000000000001400000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000001300000000000000180000000000000000000000000000000c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001900000000000000220000000000000016000000000000001600000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_42 => X"0000002c0000000000000007000000000000002b000000000000001100000000",
            INIT_43 => X"00000011000000000000000b0000000000000010000000000000001400000000",
            INIT_44 => X"0000000400000000000000180000000000000029000000000000001600000000",
            INIT_45 => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_46 => X"00000010000000000000001c000000000000000c000000000000000000000000",
            INIT_47 => X"0000000900000000000000200000000000000017000000000000000000000000",
            INIT_48 => X"0000000100000000000000000000000000000011000000000000001400000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000001300000000000000000000000000000007000000000000000300000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_4D => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"00000017000000000000001c0000000000000012000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_52 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_53 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"00000020000000000000000c0000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE49;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50 : if BRAM_NAME = "samplegold_layersamples_instance50" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000002000000000000000800000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000300000000000000000000000000000001000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000500000000000000080000000000000005000000000000000200000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000001a00000000000000150000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000120000000000000015000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000008000000000000000d000000000000000e00000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"000000000000000000000000000000000000000e000000000000001400000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000001c00000000000000120000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000000000000000000000000001a000000000000002100000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000001d00000000000000330000000000000038000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"000000000000000000000000000000000000001f000000000000002c00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000005000000000000000300000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000030000000000000001000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000001500000000000000260000000000000011000000000000002200000000",
            INIT_46 => X"0000001f000000000000001b000000000000001e000000000000000c00000000",
            INIT_47 => X"00000017000000000000001e000000000000001c000000000000001d00000000",
            INIT_48 => X"00000025000000000000001f0000000000000010000000000000000a00000000",
            INIT_49 => X"000000000000000000000016000000000000000e000000000000001800000000",
            INIT_4A => X"0000001100000000000000110000000000000009000000000000000e00000000",
            INIT_4B => X"0000000d00000000000000080000000000000008000000000000000900000000",
            INIT_4C => X"0000002f000000000000001f000000000000001d000000000000001800000000",
            INIT_4D => X"0000000000000000000000000000000000000005000000000000000500000000",
            INIT_4E => X"00000017000000000000000d0000000000000000000000000000000000000000",
            INIT_4F => X"000000250000000000000027000000000000001d000000000000001a00000000",
            INIT_50 => X"00000000000000000000002b0000000000000010000000000000001600000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000001d00000000000000080000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000150000000000000020000000000000001500000000",
            INIT_54 => X"0000000000000000000000240000000000000066000000000000000800000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000002e00000000000000210000000000000011000000000000001400000000",
            INIT_58 => X"0000000000000000000000000000000000000023000000000000007b00000000",
            INIT_59 => X"0000000000000000000000000000000000000001000000000000000200000000",
            INIT_5A => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000003a0000000000000032000000000000002f000000000000002000000000",
            INIT_5C => X"0000001000000000000000000000000000000000000000000000006000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000002f000000000000000d0000000000000000000000000000000000000000",
            INIT_5F => X"00000031000000000000003b000000000000001d000000000000001d00000000",
            INIT_60 => X"00000000000000000000000d0000000000000000000000000000005300000000",
            INIT_61 => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_62 => X"0000001500000000000000110000000000000000000000000000000000000000",
            INIT_63 => X"0000003c000000000000003e000000000000001e000000000000000800000000",
            INIT_64 => X"000000000000000000000008000000000000000d000000000000005200000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_66 => X"00000038000000000000001b0000000000000029000000000000000400000000",
            INIT_67 => X"00000069000000000000001f00000000000000a3000000000000006500000000",
            INIT_68 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_69 => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"00000097000000000000007b0000000000000051000000000000000d00000000",
            INIT_6B => X"00000000000000000000001d0000000000000014000000000000003300000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000001800000000000000050000000000000000000000000000000000000000",
            INIT_6E => X"0000003800000000000000510000000000000061000000000000007d00000000",
            INIT_6F => X"0000001900000000000000000000000000000000000000000000002d00000000",
            INIT_70 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"00000034000000000000002c0000000000000000000000000000000300000000",
            INIT_72 => X"00000033000000000000001c0000000000000021000000000000002900000000",
            INIT_73 => X"0000000000000000000000160000000000000000000000000000001800000000",
            INIT_74 => X"00000012000000000000000c000000000000000a000000000000000000000000",
            INIT_75 => X"0000001500000000000000140000000000000004000000000000000000000000",
            INIT_76 => X"0000000e000000000000000a0000000000000027000000000000002500000000",
            INIT_77 => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_78 => X"00000003000000000000000c0000000000000001000000000000000000000000",
            INIT_79 => X"0000000b000000000000001e0000000000000027000000000000000000000000",
            INIT_7A => X"0000001100000000000000020000000000000000000000000000000b00000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_7C => X"000000070000000000000000000000000000000b000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE50;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51 : if BRAM_NAME = "samplegold_layersamples_instance51" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000000d0000000000000003000000000000000000000000",
            INIT_01 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_03 => X"00000035000000000000002a0000000000000015000000000000000300000000",
            INIT_04 => X"000000000000000000000000000000000000002a000000000000003600000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000003200000000000000180000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000050000000000000018000000000000002100000000",
            INIT_08 => X"0000001b00000000000000030000000000000000000000000000000000000000",
            INIT_09 => X"0000000f00000000000000050000000000000000000000000000001b00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_0B => X"0000000b00000000000000070000000000000000000000000000000000000000",
            INIT_0C => X"00000007000000000000004f0000000000000064000000000000004e00000000",
            INIT_0D => X"0000001400000000000000270000000000000007000000000000000500000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_0F => X"0000001b0000000000000021000000000000001b000000000000000600000000",
            INIT_10 => X"0000001a00000000000000120000000000000000000000000000000300000000",
            INIT_11 => X"0000000700000000000000000000000000000000000000000000002500000000",
            INIT_12 => X"0000000000000000000000000000000000000005000000000000000800000000",
            INIT_13 => X"0000000000000000000000000000000000000005000000000000000200000000",
            INIT_14 => X"000000000000000000000000000000000000003b000000000000000000000000",
            INIT_15 => X"00000010000000000000000d0000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_17 => X"0000000f00000000000000110000000000000000000000000000000000000000",
            INIT_18 => X"0000001f00000000000000480000000000000054000000000000000000000000",
            INIT_19 => X"00000005000000000000000b000000000000000d000000000000000f00000000",
            INIT_1A => X"0000000b00000000000000000000000000000000000000000000000400000000",
            INIT_1B => X"0000006b000000000000005e0000000000000025000000000000001400000000",
            INIT_1C => X"0000001b0000000000000015000000000000003f000000000000003100000000",
            INIT_1D => X"0000000b000000000000000f0000000000000000000000000000000000000000",
            INIT_1E => X"0000007b00000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000005800000000",
            INIT_20 => X"0000000500000000000000050000000000000000000000000000000000000000",
            INIT_21 => X"000000000000000000000008000000000000000b000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_27 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000001200000000000000000000000000000000000000000000000d00000000",
            INIT_29 => X"0000001000000000000000000000000000000000000000000000000b00000000",
            INIT_2A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000023000000000000001300000000",
            INIT_2C => X"00000000000000000000001d000000000000000a000000000000001300000000",
            INIT_2D => X"0000000000000000000000000000000000000001000000000000000800000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_2F => X"000000000000000000000000000000000000000f000000000000000400000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000a000000000000000c0000000000000008000000000000000000000000",
            INIT_36 => X"000000250000000000000025000000000000001b000000000000001000000000",
            INIT_37 => X"0000000f00000000000000120000000000000010000000000000001100000000",
            INIT_38 => X"0000000e000000000000000b000000000000000d000000000000000e00000000",
            INIT_39 => X"000000110000000000000011000000000000000c000000000000000800000000",
            INIT_3A => X"0000003300000000000000330000000000000035000000000000002d00000000",
            INIT_3B => X"0000001b000000000000001b0000000000000013000000000000001f00000000",
            INIT_3C => X"0000000a000000000000001d000000000000001a000000000000001a00000000",
            INIT_3D => X"000000330000000000000015000000000000001e000000000000000a00000000",
            INIT_3E => X"000000320000000000000051000000000000004c000000000000004100000000",
            INIT_3F => X"0000002a000000000000002b0000000000000025000000000000002100000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000000d0000000000000029000000000000002700000000",
            INIT_41 => X"000000420000000000000033000000000000002d000000000000001b00000000",
            INIT_42 => X"0000003b000000000000005f000000000000005e000000000000004f00000000",
            INIT_43 => X"000000290000000000000029000000000000003a000000000000002d00000000",
            INIT_44 => X"00000037000000000000000e000000000000000b000000000000003000000000",
            INIT_45 => X"0000003f00000000000000280000000000000039000000000000002e00000000",
            INIT_46 => X"00000052000000000000005f0000000000000062000000000000005a00000000",
            INIT_47 => X"0000004700000000000000430000000000000039000000000000004700000000",
            INIT_48 => X"000000320000000000000027000000000000001b000000000000001700000000",
            INIT_49 => X"0000004b0000000000000042000000000000002e000000000000002a00000000",
            INIT_4A => X"0000004e00000000000000670000000000000061000000000000005200000000",
            INIT_4B => X"00000016000000000000004e0000000000000051000000000000004f00000000",
            INIT_4C => X"00000038000000000000003d0000000000000015000000000000001800000000",
            INIT_4D => X"0000004400000000000000470000000000000043000000000000002800000000",
            INIT_4E => X"000000560000000000000051000000000000005d000000000000005000000000",
            INIT_4F => X"000000190000000000000013000000000000003c000000000000004400000000",
            INIT_50 => X"000000300000000000000037000000000000001d000000000000002c00000000",
            INIT_51 => X"000000450000000000000040000000000000004f000000000000004c00000000",
            INIT_52 => X"0000003900000000000000470000000000000059000000000000005500000000",
            INIT_53 => X"0000001b00000000000000150000000000000018000000000000003600000000",
            INIT_54 => X"0000003a00000000000000550000000000000033000000000000004900000000",
            INIT_55 => X"0000004c000000000000003d000000000000003d000000000000005800000000",
            INIT_56 => X"0000005200000000000000490000000000000041000000000000005500000000",
            INIT_57 => X"00000037000000000000002d0000000000000021000000000000001900000000",
            INIT_58 => X"0000005700000000000000380000000000000048000000000000002e00000000",
            INIT_59 => X"000000530000000000000046000000000000003a000000000000003e00000000",
            INIT_5A => X"0000001a00000000000000500000000000000053000000000000004900000000",
            INIT_5B => X"0000003e00000000000000340000000000000044000000000000002d00000000",
            INIT_5C => X"0000004400000000000000420000000000000048000000000000003f00000000",
            INIT_5D => X"000000520000000000000051000000000000004b000000000000004500000000",
            INIT_5E => X"00000015000000000000001e000000000000005a000000000000004c00000000",
            INIT_5F => X"0000003b000000000000003c0000000000000020000000000000002200000000",
            INIT_60 => X"0000003b00000000000000370000000000000040000000000000002e00000000",
            INIT_61 => X"0000004f0000000000000060000000000000004c000000000000003d00000000",
            INIT_62 => X"000000170000000000000014000000000000001a000000000000005d00000000",
            INIT_63 => X"0000003800000000000000340000000000000029000000000000002500000000",
            INIT_64 => X"00000034000000000000002a000000000000002f000000000000003900000000",
            INIT_65 => X"0000004f00000000000000620000000000000060000000000000004500000000",
            INIT_66 => X"0000004000000000000000350000000000000026000000000000001c00000000",
            INIT_67 => X"00000049000000000000003c0000000000000040000000000000003f00000000",
            INIT_68 => X"0000003b000000000000002b000000000000003e000000000000004300000000",
            INIT_69 => X"00000035000000000000005a0000000000000060000000000000005b00000000",
            INIT_6A => X"0000004f00000000000000530000000000000047000000000000003e00000000",
            INIT_6B => X"0000005b000000000000005a0000000000000051000000000000004900000000",
            INIT_6C => X"00000058000000000000004e0000000000000048000000000000005100000000",
            INIT_6D => X"000000000000000000000000000000000000005f000000000000006300000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000b00000000000000010000000000000000000000000000000000000000",
            INIT_71 => X"0000000500000000000000000000000000000000000000000000000500000000",
            INIT_72 => X"0000000000000000000000020000000000000000000000000000000500000000",
            INIT_73 => X"0000000600000000000000030000000000000000000000000000000000000000",
            INIT_74 => X"00000009000000000000000f000000000000000d000000000000000a00000000",
            INIT_75 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000600000000000000050000000000000003000000000000000a00000000",
            INIT_78 => X"0000000000000000000000060000000000000007000000000000000800000000",
            INIT_79 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_7B => X"0000000d00000000000000000000000000000000000000000000000800000000",
            INIT_7C => X"0000000e0000000000000010000000000000000c000000000000000600000000",
            INIT_7D => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000001300000000000000110000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE51;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52 : if BRAM_NAME = "samplegold_layersamples_instance52" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000006000000000000001500000000",
            INIT_01 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"000000120000000000000019000000000000001a000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000010000000000000001800000000",
            INIT_06 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000100000000000000030000000000000018000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_09 => X"0000000000000000000000020000000000000000000000000000002400000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000f00000000000000070000000000000010000000000000000900000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_0E => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000080000000000000014000000000000000600000000",
            INIT_10 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000002200000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000017000000000000000e000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"000000070000000000000000000000000000000a000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000002c00000000",
            INIT_1B => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_1C => X"0000000900000000000000000000000000000000000000000000000700000000",
            INIT_1D => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"00000001000000000000000c0000000000000008000000000000002000000000",
            INIT_1F => X"0000000f00000000000000130000000000000014000000000000000100000000",
            INIT_20 => X"0000000000000000000000060000000000000001000000000000000400000000",
            INIT_21 => X"0000002a000000000000001c0000000000000000000000000000000000000000",
            INIT_22 => X"0000001a00000000000000160000000000000009000000000000000300000000",
            INIT_23 => X"00000012000000000000000e0000000000000022000000000000003400000000",
            INIT_24 => X"00000012000000000000001a0000000000000017000000000000001e00000000",
            INIT_25 => X"0000000000000000000000270000000000000026000000000000000900000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000004000000000000000400000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000c00000000000000010000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000003000000000000000500000000",
            INIT_34 => X"0000000000000000000000080000000000000000000000000000000300000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000007000000000000000700000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000001200000000000000060000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000001300000000000000130000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000060000000000000008000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"000000000000000000000000000000000000002b000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000001600000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000003300000000",
            INIT_4C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_4E => X"0000002600000000000000100000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"000000000000000000000020000000000000001d000000000000000c00000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000022000000000000002400000000",
            INIT_57 => X"00000013000000000000002b000000000000001d000000000000000000000000",
            INIT_58 => X"0000000000000000000000080000000000000003000000000000000600000000",
            INIT_59 => X"0000002e00000000000000010000000000000000000000000000000000000000",
            INIT_5A => X"0000002e0000000000000027000000000000000a000000000000002e00000000",
            INIT_5B => X"00000011000000000000001d000000000000002c000000000000002b00000000",
            INIT_5C => X"0000001a0000000000000021000000000000002f000000000000002900000000",
            INIT_5D => X"0000003b00000000000000360000000000000028000000000000001e00000000",
            INIT_5E => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000003000000000000000a00000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000007000000000000001200000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000e00000000000000050000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"00000009000000000000000d000000000000000c000000000000000800000000",
            INIT_75 => X"0000001e00000000000000030000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_77 => X"0000001800000000000000020000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000270000000000000008000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE52;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53 : if BRAM_NAME = "samplegold_layersamples_instance53" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001a0000000000000035000000000000003d000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000002100000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000001e0000000000000003000000000000000e000000000000000200000000",
            INIT_04 => X"0000002500000000000000180000000000000013000000000000001b00000000",
            INIT_05 => X"000000000000000000000000000000000000001a000000000000000600000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000210000000000000043000000000000006a000000000000000200000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000013000000000000001d00000000",
            INIT_0C => X"00000000000000000000000b0000000000000000000000000000001200000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000120000000000000003000000000000000000000000",
            INIT_0F => X"0000001300000000000000250000000000000017000000000000000000000000",
            INIT_10 => X"0000000200000000000000020000000000000000000000000000000100000000",
            INIT_11 => X"0000000500000000000000000000000000000019000000000000000800000000",
            INIT_12 => X"0000002200000000000000200000000000000011000000000000001300000000",
            INIT_13 => X"0000000b000000000000000a000000000000000a000000000000000f00000000",
            INIT_14 => X"000000010000000000000007000000000000000e000000000000000300000000",
            INIT_15 => X"0000001100000000000000120000000000000014000000000000000300000000",
            INIT_16 => X"000000460000000000000044000000000000004a000000000000001500000000",
            INIT_17 => X"0000003c00000000000000420000000000000040000000000000004900000000",
            INIT_18 => X"00000024000000000000002a000000000000002f000000000000003b00000000",
            INIT_19 => X"000000020000000000000008000000000000000f000000000000001900000000",
            INIT_1A => X"0000003000000000000000400000000000000042000000000000004800000000",
            INIT_1B => X"0000002a00000000000000380000000000000035000000000000003100000000",
            INIT_1C => X"0000001300000000000000190000000000000022000000000000002a00000000",
            INIT_1D => X"0000004300000000000000140000000000000012000000000000001100000000",
            INIT_1E => X"00000021000000000000001f0000000000000033000000000000004200000000",
            INIT_1F => X"00000028000000000000001c0000000000000017000000000000001600000000",
            INIT_20 => X"0000003100000000000000340000000000000035000000000000003300000000",
            INIT_21 => X"0000003a00000000000000390000000000000025000000000000003100000000",
            INIT_22 => X"0000001100000000000000120000000000000000000000000000002200000000",
            INIT_23 => X"0000004200000000000000190000000000000011000000000000000c00000000",
            INIT_24 => X"000000240000000000000032000000000000003b000000000000004300000000",
            INIT_25 => X"0000005900000000000000550000000000000045000000000000001600000000",
            INIT_26 => X"0000002d000000000000002c000000000000000d000000000000000600000000",
            INIT_27 => X"0000002a00000000000000170000000000000016000000000000001600000000",
            INIT_28 => X"0000001900000000000000200000000000000033000000000000003a00000000",
            INIT_29 => X"0000000b0000000000000088000000000000008f000000000000008100000000",
            INIT_2A => X"0000002d000000000000003c0000000000000027000000000000001300000000",
            INIT_2B => X"0000002b00000000000000110000000000000011000000000000002200000000",
            INIT_2C => X"0000008f000000000000002c0000000000000030000000000000003500000000",
            INIT_2D => X"0000001c00000000000000220000000000000086000000000000008b00000000",
            INIT_2E => X"0000003200000000000000280000000000000038000000000000003800000000",
            INIT_2F => X"00000034000000000000001c0000000000000018000000000000002400000000",
            INIT_30 => X"00000080000000000000007e0000000000000034000000000000003c00000000",
            INIT_31 => X"0000000e00000000000000270000000000000073000000000000008100000000",
            INIT_32 => X"0000003b0000000000000041000000000000001f000000000000002000000000",
            INIT_33 => X"0000002b00000000000000310000000000000016000000000000001d00000000",
            INIT_34 => X"0000009b00000000000000910000000000000083000000000000002300000000",
            INIT_35 => X"0000004800000000000000500000000000000087000000000000006500000000",
            INIT_36 => X"0000002900000000000000440000000000000043000000000000001d00000000",
            INIT_37 => X"00000017000000000000002a0000000000000029000000000000001d00000000",
            INIT_38 => X"000000c600000000000000e000000000000000ce00000000000000b300000000",
            INIT_39 => X"0000002f00000000000000490000000000000085000000000000009300000000",
            INIT_3A => X"0000002300000000000000360000000000000044000000000000003c00000000",
            INIT_3B => X"0000010100000000000000000000000000000016000000000000002300000000",
            INIT_3C => X"000000620000000000000089000000000000009400000000000000fb00000000",
            INIT_3D => X"0000003700000000000000340000000000000042000000000000005b00000000",
            INIT_3E => X"0000001a00000000000000240000000000000033000000000000004000000000",
            INIT_3F => X"000000cb00000000000000e80000000000000000000000000000001400000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001900000000000000220000000000000056000000000000008200000000",
            INIT_41 => X"000000330000000000000023000000000000000c000000000000003300000000",
            INIT_42 => X"000000170000000000000011000000000000002d000000000000003700000000",
            INIT_43 => X"0000005c00000000000000650000000000000075000000000000000600000000",
            INIT_44 => X"000000230000000000000010000000000000003b000000000000004d00000000",
            INIT_45 => X"0000004f0000000000000038000000000000001b000000000000002e00000000",
            INIT_46 => X"0000001a0000000000000004000000000000001e000000000000003f00000000",
            INIT_47 => X"0000002f000000000000003d000000000000003e000000000000004500000000",
            INIT_48 => X"000000190000000000000007000000000000001e000000000000001c00000000",
            INIT_49 => X"00000037000000000000004b0000000000000022000000000000000c00000000",
            INIT_4A => X"0000002e00000000000000010000000000000002000000000000002600000000",
            INIT_4B => X"000000000000000000000000000000000000000c000000000000001e00000000",
            INIT_4C => X"0000000000000000000000020000000000000010000000000000001300000000",
            INIT_4D => X"00000003000000000000000d0000000000000000000000000000000000000000",
            INIT_4E => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000030000000000000007000000000000000000000000",
            INIT_50 => X"0000000100000000000000000000000000000000000000000000000500000000",
            INIT_51 => X"0000000000000000000000000000000000000004000000000000000400000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"00000000000000000000000c0000000000000000000000000000000900000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000220000000000000000000000000000000400000000",
            INIT_57 => X"0000000000000000000000090000000000000000000000000000000400000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"00000000000000000000000c0000000000000007000000000000000000000000",
            INIT_5A => X"00000000000000000000000d0000000000000000000000000000000000000000",
            INIT_5B => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000060000000000000000000000000000000100000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000010000000000000009000000000000000000000000",
            INIT_5F => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000001100000000000000000000000000000000000000000000001500000000",
            INIT_63 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000007000000000000000a00000000",
            INIT_66 => X"000000000000000000000002000000000000000b000000000000001900000000",
            INIT_67 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_68 => X"00000000000000000000001d0000000000000008000000000000000500000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_6F => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000002d00000000000000000000000000000000000000000000002500000000",
            INIT_71 => X"0000000000000000000000030000000000000018000000000000000400000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_73 => X"0000000000000000000000130000000000000005000000000000000000000000",
            INIT_74 => X"00000046000000000000007b000000000000001b000000000000000000000000",
            INIT_75 => X"00000012000000000000001a000000000000002c000000000000002e00000000",
            INIT_76 => X"0000000000000000000000090000000000000002000000000000000000000000",
            INIT_77 => X"0000007300000000000000020000000000000000000000000000000000000000",
            INIT_78 => X"0000002500000000000000000000000000000002000000000000005e00000000",
            INIT_79 => X"0000000a000000000000001a0000000000000000000000000000000f00000000",
            INIT_7A => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"00000019000000000000001f0000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_7E => X"0000000700000000000000000000000000000002000000000000000000000000",
            INIT_7F => X"0000001600000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE53;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54 : if BRAM_NAME = "samplegold_layersamples_instance54" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000011000000000000002a00000000",
            INIT_01 => X"0000001500000000000000230000000000000009000000000000000800000000",
            INIT_02 => X"0000000a00000000000000070000000000000010000000000000000300000000",
            INIT_03 => X"0000000000000000000000090000000000000025000000000000001e00000000",
            INIT_04 => X"0000000400000000000000010000000000000000000000000000000000000000",
            INIT_05 => X"00000014000000000000000d0000000000000000000000000000000100000000",
            INIT_06 => X"0000001000000000000000070000000000000003000000000000000700000000",
            INIT_07 => X"00000006000000000000000e0000000000000016000000000000000d00000000",
            INIT_08 => X"00000009000000000000000d0000000000000003000000000000000000000000",
            INIT_09 => X"0000000d000000000000000b000000000000000c000000000000000900000000",
            INIT_0A => X"0000000b0000000000000010000000000000000a000000000000001100000000",
            INIT_0B => X"000000000000000000000000000000000000000a000000000000001200000000",
            INIT_0C => X"0000000700000000000000090000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000001000000000000000300000000",
            INIT_0E => X"00000004000000000000000e0000000000000012000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"000000030000000000000000000000000000000f000000000000000e00000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000800000000000000090000000000000000000000000000000000000000",
            INIT_1A => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"00000000000000000000000a000000000000000e000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000003000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000009000000000000000d00000000",
            INIT_22 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"000000000000000000000000000000000000000f000000000000000e00000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000000000000000000002000000000000000b000000000000001000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000200000000000000070000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000001700000000000000250000000000000018000000000000001c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000019000000000000001a0000000000000027000000000000002800000000",
            INIT_41 => X"000000100000000000000014000000000000001a000000000000001600000000",
            INIT_42 => X"0000001b0000000000000013000000000000001b000000000000001400000000",
            INIT_43 => X"0000002d00000000000000130000000000000026000000000000001700000000",
            INIT_44 => X"000000170000000000000029000000000000002b000000000000003d00000000",
            INIT_45 => X"000000240000000000000020000000000000001c000000000000001b00000000",
            INIT_46 => X"0000001a000000000000001c000000000000001c000000000000002600000000",
            INIT_47 => X"0000003d000000000000002a000000000000002b000000000000000f00000000",
            INIT_48 => X"00000033000000000000003a000000000000003f000000000000004000000000",
            INIT_49 => X"0000001200000000000000180000000000000023000000000000002600000000",
            INIT_4A => X"000000030000000000000021000000000000001e000000000000000b00000000",
            INIT_4B => X"000000440000000000000042000000000000003a000000000000002b00000000",
            INIT_4C => X"0000003200000000000000360000000000000040000000000000004700000000",
            INIT_4D => X"0000001600000000000000110000000000000015000000000000001600000000",
            INIT_4E => X"000000000000000000000015000000000000003e000000000000003600000000",
            INIT_4F => X"0000003200000000000000470000000000000058000000000000003f00000000",
            INIT_50 => X"0000003200000000000000480000000000000044000000000000004300000000",
            INIT_51 => X"0000002e000000000000001e0000000000000019000000000000002700000000",
            INIT_52 => X"0000003300000000000000000000000000000000000000000000002100000000",
            INIT_53 => X"0000004400000000000000310000000000000033000000000000006400000000",
            INIT_54 => X"0000003500000000000000460000000000000042000000000000003d00000000",
            INIT_55 => X"0000001200000000000000190000000000000011000000000000001b00000000",
            INIT_56 => X"0000004700000000000000340000000000000000000000000000000800000000",
            INIT_57 => X"000000350000000000000048000000000000003f000000000000002a00000000",
            INIT_58 => X"0000002300000000000000330000000000000051000000000000003700000000",
            INIT_59 => X"0000001e00000000000000260000000000000024000000000000000200000000",
            INIT_5A => X"0000002b00000000000000450000000000000000000000000000000400000000",
            INIT_5B => X"000000340000000000000030000000000000004d000000000000004700000000",
            INIT_5C => X"000000150000000000000024000000000000003b000000000000004500000000",
            INIT_5D => X"0000001600000000000000230000000000000030000000000000002e00000000",
            INIT_5E => X"0000002a00000000000000330000000000000013000000000000002800000000",
            INIT_5F => X"0000003a00000000000000390000000000000033000000000000004900000000",
            INIT_60 => X"000000430000000000000005000000000000002a000000000000004800000000",
            INIT_61 => X"000000260000000000000000000000000000000e000000000000003e00000000",
            INIT_62 => X"000000490000000000000019000000000000003c000000000000000000000000",
            INIT_63 => X"0000003f0000000000000032000000000000003d000000000000003f00000000",
            INIT_64 => X"000000010000000000000018000000000000000d000000000000000b00000000",
            INIT_65 => X"00000018000000000000002a0000000000000003000000000000000000000000",
            INIT_66 => X"0000003e00000000000000440000000000000024000000000000003700000000",
            INIT_67 => X"000000220000000000000031000000000000002e000000000000003000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000a00000000",
            INIT_69 => X"000000470000000000000035000000000000000a000000000000000c00000000",
            INIT_6A => X"000000410000000000000041000000000000003f000000000000001500000000",
            INIT_6B => X"000000010000000000000033000000000000001a000000000000002f00000000",
            INIT_6C => X"0000001d00000000000000100000000000000012000000000000000500000000",
            INIT_6D => X"0000001d000000000000003e0000000000000027000000000000000b00000000",
            INIT_6E => X"0000003000000000000000400000000000000058000000000000004600000000",
            INIT_6F => X"00000018000000000000001e0000000000000028000000000000001d00000000",
            INIT_70 => X"0000000c0000000000000009000000000000001d000000000000002600000000",
            INIT_71 => X"0000002d00000000000000260000000000000024000000000000001e00000000",
            INIT_72 => X"00000023000000000000002d0000000000000032000000000000003f00000000",
            INIT_73 => X"0000000800000000000000130000000000000026000000000000001600000000",
            INIT_74 => X"0000002900000000000000260000000000000011000000000000000d00000000",
            INIT_75 => X"000000210000000000000017000000000000000e000000000000001f00000000",
            INIT_76 => X"0000001c00000000000000110000000000000022000000000000002c00000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000001600000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000001900000000000000090000000000000000000000000000000000000000",
            INIT_7E => X"000000000000000000000011000000000000001d000000000000002300000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE54;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55 : if BRAM_NAME = "samplegold_layersamples_instance55" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000001000000000000000a00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000a0000000000000034000000000000002d000000000000000000000000",
            INIT_07 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"000000000000000000000000000000000000000c000000000000000900000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000002d000000000000001b0000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000002300000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000001200000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000002400000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000002200000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000100000000000000040000000000000002000000000000000200000000",
            INIT_41 => X"0000000800000000000000040000000000000001000000000000000000000000",
            INIT_42 => X"0000001800000000000000110000000000000010000000000000000b00000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000700000000000000040000000000000001000000000000000000000000",
            INIT_45 => X"0000001200000000000000160000000000000006000000000000000000000000",
            INIT_46 => X"0000000900000000000000060000000000000009000000000000000900000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_49 => X"000000020000000000000005000000000000000a000000000000000c00000000",
            INIT_4A => X"0000001800000000000000000000000000000017000000000000000800000000",
            INIT_4B => X"000000010000000000000000000000000000000b000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000100000000",
            INIT_4D => X"00000010000000000000000d0000000000000000000000000000000000000000",
            INIT_4E => X"0000002900000000000000230000000000000022000000000000001700000000",
            INIT_4F => X"000000000000000000000000000000000000000b000000000000000700000000",
            INIT_50 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"00000036000000000000003c0000000000000026000000000000000d00000000",
            INIT_52 => X"0000000200000000000000240000000000000014000000000000003000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_54 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_55 => X"00000000000000000000001b000000000000003b000000000000003400000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_58 => X"00000024000000000000000a0000000000000006000000000000000000000000",
            INIT_59 => X"0000000000000000000000060000000000000000000000000000000900000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000600000000000000070000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000012000000000000000700000000",
            INIT_5D => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000d000000000000000c0000000000000000000000000000000400000000",
            INIT_60 => X"0000000500000000000000000000000000000000000000000000000700000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000c000000000000000a000000000000000a000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_65 => X"0000000900000000000000080000000000000009000000000000000000000000",
            INIT_66 => X"0000000100000000000000000000000000000000000000000000000600000000",
            INIT_67 => X"00000018000000000000000b0000000000000008000000000000000600000000",
            INIT_68 => X"0000001c0000000000000014000000000000000c000000000000001c00000000",
            INIT_69 => X"0000001f0000000000000018000000000000002a000000000000002100000000",
            INIT_6A => X"0000001e0000000000000020000000000000001e000000000000001f00000000",
            INIT_6B => X"0000001d0000000000000019000000000000001c000000000000001600000000",
            INIT_6C => X"0000002e000000000000002f0000000000000018000000000000001500000000",
            INIT_6D => X"0000001900000000000000220000000000000036000000000000003100000000",
            INIT_6E => X"00000018000000000000001a000000000000001a000000000000001d00000000",
            INIT_6F => X"000000290000000000000019000000000000001a000000000000001c00000000",
            INIT_70 => X"0000004600000000000000410000000000000039000000000000001300000000",
            INIT_71 => X"0000001d000000000000001c0000000000000020000000000000003e00000000",
            INIT_72 => X"0000001900000000000000180000000000000019000000000000001c00000000",
            INIT_73 => X"0000003200000000000000260000000000000017000000000000001a00000000",
            INIT_74 => X"0000004500000000000000440000000000000046000000000000004100000000",
            INIT_75 => X"0000002b000000000000001e0000000000000020000000000000004200000000",
            INIT_76 => X"0000000a00000000000000170000000000000017000000000000000e00000000",
            INIT_77 => X"0000004700000000000000400000000000000045000000000000000d00000000",
            INIT_78 => X"0000004d00000000000000580000000000000041000000000000002500000000",
            INIT_79 => X"000000140000000000000031000000000000003a000000000000004a00000000",
            INIT_7A => X"0000000900000000000000070000000000000016000000000000001200000000",
            INIT_7B => X"0000002900000000000000340000000000000041000000000000003600000000",
            INIT_7C => X"000000510000000000000046000000000000004d000000000000004d00000000",
            INIT_7D => X"0000000c0000000000000018000000000000003c000000000000005400000000",
            INIT_7E => X"0000000b00000000000000060000000000000006000000000000001500000000",
            INIT_7F => X"00000045000000000000001d0000000000000028000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE55;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56 : if BRAM_NAME = "samplegold_layersamples_instance56" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000055000000000000004d000000000000003c000000000000004400000000",
            INIT_01 => X"0000001c000000000000000e0000000000000033000000000000004100000000",
            INIT_02 => X"0000000800000000000000170000000000000002000000000000000600000000",
            INIT_03 => X"0000003b00000000000000440000000000000020000000000000004a00000000",
            INIT_04 => X"0000005300000000000000570000000000000050000000000000003c00000000",
            INIT_05 => X"0000000300000000000000130000000000000023000000000000003900000000",
            INIT_06 => X"0000001900000000000000410000000000000000000000000000000000000000",
            INIT_07 => X"0000003f00000000000000510000000000000012000000000000004000000000",
            INIT_08 => X"0000003f000000000000005c0000000000000052000000000000004900000000",
            INIT_09 => X"000000000000000000000000000000000000001f000000000000003200000000",
            INIT_0A => X"00000039000000000000001d000000000000002b000000000000000e00000000",
            INIT_0B => X"000000440000000000000043000000000000004e000000000000001f00000000",
            INIT_0C => X"00000036000000000000004b0000000000000060000000000000004b00000000",
            INIT_0D => X"0000004c00000000000000090000000000000000000000000000000d00000000",
            INIT_0E => X"000000390000000000000037000000000000002e000000000000002300000000",
            INIT_0F => X"000000450000000000000043000000000000003f000000000000002e00000000",
            INIT_10 => X"0000002500000000000000190000000000000045000000000000005300000000",
            INIT_11 => X"00000029000000000000000b0000000000000004000000000000000f00000000",
            INIT_12 => X"0000004900000000000000230000000000000042000000000000005300000000",
            INIT_13 => X"0000004d00000000000000380000000000000035000000000000002e00000000",
            INIT_14 => X"0000000d00000000000000260000000000000009000000000000003f00000000",
            INIT_15 => X"00000022000000000000000f000000000000000a000000000000000f00000000",
            INIT_16 => X"0000003b00000000000000360000000000000029000000000000003800000000",
            INIT_17 => X"00000040000000000000004b0000000000000040000000000000002c00000000",
            INIT_18 => X"00000012000000000000000f0000000000000008000000000000001d00000000",
            INIT_19 => X"0000000e000000000000000a000000000000001d000000000000002000000000",
            INIT_1A => X"0000003000000000000000340000000000000030000000000000002800000000",
            INIT_1B => X"0000001c00000000000000450000000000000041000000000000002600000000",
            INIT_1C => X"0000000f0000000000000016000000000000001e000000000000001000000000",
            INIT_1D => X"00000022000000000000000d0000000000000008000000000000001700000000",
            INIT_1E => X"000000230000000000000020000000000000001d000000000000001f00000000",
            INIT_1F => X"0000001200000000000000150000000000000023000000000000002200000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000040000000000000002000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000004000000000000000100000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000002000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE56;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57 : if BRAM_NAME = "samplegold_layersamples_instance57" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000002600000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000200000000000000070000000000000003000000000000000900000000",
            INIT_12 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_13 => X"00000006000000000000000a0000000000000013000000000000002300000000",
            INIT_14 => X"0000000d00000000000000170000000000000002000000000000000300000000",
            INIT_15 => X"0000000b00000000000000120000000000000019000000000000001000000000",
            INIT_16 => X"000000390000000000000000000000000000000e000000000000000b00000000",
            INIT_17 => X"0000000a000000000000000c000000000000000c000000000000000f00000000",
            INIT_18 => X"0000001c00000000000000170000000000000007000000000000000200000000",
            INIT_19 => X"00000011000000000000000a0000000000000006000000000000002f00000000",
            INIT_1A => X"000000120000000000000025000000000000000c000000000000000000000000",
            INIT_1B => X"00000007000000000000000f0000000000000014000000000000001100000000",
            INIT_1C => X"000000280000000000000001000000000000002d000000000000002700000000",
            INIT_1D => X"00000014000000000000000a0000000000000015000000000000001700000000",
            INIT_1E => X"0000002200000000000000290000000000000014000000000000002e00000000",
            INIT_1F => X"000000180000000000000001000000000000000f000000000000000c00000000",
            INIT_20 => X"0000002100000000000000300000000000000000000000000000000d00000000",
            INIT_21 => X"0000002300000000000000150000000000000000000000000000001500000000",
            INIT_22 => X"0000000000000000000000170000000000000021000000000000001b00000000",
            INIT_23 => X"00000002000000000000000e0000000000000007000000000000000b00000000",
            INIT_24 => X"00000009000000000000001d0000000000000024000000000000000400000000",
            INIT_25 => X"0000001b0000000000000028000000000000001d000000000000000e00000000",
            INIT_26 => X"0000000000000000000000000000000000000010000000000000002300000000",
            INIT_27 => X"0000000e00000000000000000000000000000009000000000000000200000000",
            INIT_28 => X"0000001f00000000000000140000000000000024000000000000001400000000",
            INIT_29 => X"000000210000000000000023000000000000001a000000000000001600000000",
            INIT_2A => X"0000000000000000000000000000000000000008000000000000001500000000",
            INIT_2B => X"00000019000000000000002a0000000000000000000000000000000a00000000",
            INIT_2C => X"0000000e00000000000000200000000000000018000000000000001600000000",
            INIT_2D => X"000000090000000000000010000000000000000d000000000000001c00000000",
            INIT_2E => X"0000000a00000000000000000000000000000008000000000000000900000000",
            INIT_2F => X"00000022000000000000001b0000000000000030000000000000001800000000",
            INIT_30 => X"0000000800000000000000210000000000000008000000000000002400000000",
            INIT_31 => X"00000000000000000000001b0000000000000000000000000000000f00000000",
            INIT_32 => X"0000001a000000000000000d0000000000000000000000000000000f00000000",
            INIT_33 => X"0000001c000000000000001f000000000000001d000000000000001400000000",
            INIT_34 => X"00000001000000000000001d0000000000000013000000000000001600000000",
            INIT_35 => X"0000000c000000000000000c0000000000000015000000000000000a00000000",
            INIT_36 => X"0000001d000000000000001a0000000000000003000000000000000500000000",
            INIT_37 => X"0000002100000000000000210000000000000008000000000000001c00000000",
            INIT_38 => X"0000001500000000000000070000000000000004000000000000000d00000000",
            INIT_39 => X"00000007000000000000000c0000000000000006000000000000001200000000",
            INIT_3A => X"0000001a000000000000001f0000000000000023000000000000000000000000",
            INIT_3B => X"00000013000000000000001a000000000000001d000000000000000c00000000",
            INIT_3C => X"00000014000000000000000e0000000000000018000000000000000000000000",
            INIT_3D => X"0000000000000000000000010000000000000002000000000000000b00000000",
            INIT_3E => X"0000001c0000000000000009000000000000001c000000000000001300000000",
            INIT_3F => X"000000000000000000000005000000000000000f000000000000001b00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000005000000000000000d000000000000000a000000000000000f00000000",
            INIT_41 => X"0000000a00000000000000000000000000000000000000000000000900000000",
            INIT_42 => X"0000000a0000000000000027000000000000000c000000000000001c00000000",
            INIT_43 => X"0000000d00000000000000000000000000000003000000000000000600000000",
            INIT_44 => X"0000001000000000000000110000000000000003000000000000000a00000000",
            INIT_45 => X"0000001e00000000000000080000000000000000000000000000000000000000",
            INIT_46 => X"000000030000000000000000000000000000000e000000000000001200000000",
            INIT_47 => X"0000000c0000000000000008000000000000000d000000000000000000000000",
            INIT_48 => X"0000001400000000000000080000000000000011000000000000000500000000",
            INIT_49 => X"0000002800000000000000250000000000000006000000000000000000000000",
            INIT_4A => X"000000370000000000000010000000000000001e000000000000000e00000000",
            INIT_4B => X"0000002000000000000000190000000000000000000000000000005800000000",
            INIT_4C => X"0000000000000000000000110000000000000023000000000000001d00000000",
            INIT_4D => X"00000037000000000000002f0000000000000003000000000000000000000000",
            INIT_4E => X"00000079000000000000003a000000000000001a000000000000002000000000",
            INIT_4F => X"00000027000000000000002e000000000000002e000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000011000000000000002c00000000",
            INIT_51 => X"0000002c00000000000000860000000000000016000000000000000100000000",
            INIT_52 => X"00000000000000000000000b000000000000003d000000000000001700000000",
            INIT_53 => X"0000003500000000000000310000000000000035000000000000001c00000000",
            INIT_54 => X"0000004b00000000000000000000000000000000000000000000003500000000",
            INIT_55 => X"00000042000000000000004b0000000000000062000000000000000200000000",
            INIT_56 => X"00000000000000000000003c0000000000000000000000000000001700000000",
            INIT_57 => X"0000004a000000000000001d0000000000000063000000000000004900000000",
            INIT_58 => X"00000000000000000000005d0000000000000031000000000000000100000000",
            INIT_59 => X"0000001b000000000000006a000000000000005e000000000000003c00000000",
            INIT_5A => X"0000004600000000000000090000000000000016000000000000000000000000",
            INIT_5B => X"0000002300000000000000350000000000000009000000000000006800000000",
            INIT_5C => X"000000440000000000000014000000000000003f000000000000003e00000000",
            INIT_5D => X"000000020000000000000027000000000000003a000000000000006500000000",
            INIT_5E => X"0000006400000000000000440000000000000000000000000000001600000000",
            INIT_5F => X"0000005000000000000000220000000000000033000000000000001f00000000",
            INIT_60 => X"0000006300000000000000180000000000000031000000000000001e00000000",
            INIT_61 => X"00000014000000000000001b000000000000004f000000000000001000000000",
            INIT_62 => X"0000003a000000000000004f0000000000000037000000000000000200000000",
            INIT_63 => X"0000000000000000000000710000000000000023000000000000004100000000",
            INIT_64 => X"0000004d00000000000000480000000000000041000000000000005400000000",
            INIT_65 => X"000000110000000000000045000000000000001f000000000000001f00000000",
            INIT_66 => X"0000005a00000000000000250000000000000059000000000000001400000000",
            INIT_67 => X"0000003f000000000000000a000000000000003c000000000000001400000000",
            INIT_68 => X"000000000000000000000078000000000000004a000000000000003e00000000",
            INIT_69 => X"000000000000000000000034000000000000003a000000000000003300000000",
            INIT_6A => X"0000002200000000000000490000000000000000000000000000003800000000",
            INIT_6B => X"00000044000000000000002b000000000000003c000000000000003200000000",
            INIT_6C => X"00000013000000000000004b000000000000004f000000000000004600000000",
            INIT_6D => X"00000034000000000000000e000000000000001f000000000000005000000000",
            INIT_6E => X"00000013000000000000004f0000000000000036000000000000000a00000000",
            INIT_6F => X"0000001400000000000000650000000000000037000000000000003600000000",
            INIT_70 => X"00000018000000000000005f000000000000005c000000000000003200000000",
            INIT_71 => X"0000002d00000000000000400000000000000028000000000000001600000000",
            INIT_72 => X"000000420000000000000000000000000000005c000000000000003200000000",
            INIT_73 => X"0000003400000000000000260000000000000050000000000000005600000000",
            INIT_74 => X"0000002e00000000000000000000000000000061000000000000004d00000000",
            INIT_75 => X"0000003900000000000000360000000000000042000000000000002800000000",
            INIT_76 => X"0000007d000000000000003f0000000000000000000000000000004500000000",
            INIT_77 => X"0000005000000000000000390000000000000025000000000000001000000000",
            INIT_78 => X"000000330000000000000029000000000000000b000000000000004400000000",
            INIT_79 => X"00000040000000000000003f000000000000002c000000000000002700000000",
            INIT_7A => X"0000002900000000000000670000000000000030000000000000000000000000",
            INIT_7B => X"0000002100000000000000400000000000000032000000000000004600000000",
            INIT_7C => X"0000000000000000000000390000000000000022000000000000001200000000",
            INIT_7D => X"0000000000000000000000300000000000000036000000000000002100000000",
            INIT_7E => X"000000520000000000000057000000000000004c000000000000001c00000000",
            INIT_7F => X"0000001900000000000000000000000000000045000000000000002700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE57;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58 : if BRAM_NAME = "samplegold_layersamples_instance58" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001e00000000000000160000000000000028000000000000001f00000000",
            INIT_01 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"00000014000000000000000d0000000000000000000000000000000400000000",
            INIT_03 => X"000000290000000000000000000000000000002b000000000000002c00000000",
            INIT_04 => X"000000010000000000000014000000000000001a000000000000001f00000000",
            INIT_05 => X"0000002500000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000200000000000000090000000000000000000000000000001300000000",
            INIT_07 => X"00000015000000000000001a0000000000000050000000000000000700000000",
            INIT_08 => X"000000000000000000000003000000000000000b000000000000001000000000",
            INIT_09 => X"0000000e000000000000000a0000000000000018000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000001700000000000000050000000000000000000000000000003a00000000",
            INIT_0C => X"0000008d000000000000007d0000000000000097000000000000001f00000000",
            INIT_0D => X"0000004e00000000000000120000000000000000000000000000000000000000",
            INIT_0E => X"00000000000000000000000a0000000000000008000000000000002100000000",
            INIT_0F => X"000000000000000000000001000000000000001f000000000000000e00000000",
            INIT_10 => X"000000000000000000000012000000000000005c000000000000003400000000",
            INIT_11 => X"0000000000000000000000010000000000000000000000000000000600000000",
            INIT_12 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000800000000000000000000000000000000000000000000000b00000000",
            INIT_14 => X"00000012000000000000000a0000000000000000000000000000000500000000",
            INIT_15 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_17 => X"0000000000000000000000000000000000000005000000000000000e00000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000b00000000000000180000000000000009000000000000000700000000",
            INIT_1A => X"0000001400000000000000000000000000000001000000000000000700000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_1C => X"0000000000000000000000000000000000000015000000000000000800000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000002400000000000000120000000000000000000000000000000200000000",
            INIT_20 => X"000000080000000000000031000000000000003a000000000000000800000000",
            INIT_21 => X"00000012000000000000000a0000000000000000000000000000000000000000",
            INIT_22 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"00000000000000000000000e0000000000000006000000000000001c00000000",
            INIT_24 => X"0000004c00000000000000180000000000000000000000000000000000000000",
            INIT_25 => X"0000002200000000000000000000000000000000000000000000001b00000000",
            INIT_26 => X"0000000200000000000000000000000000000000000000000000001000000000",
            INIT_27 => X"000000000000000000000018000000000000000e000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000090000000000000016000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000001600000000000000000000000000000000000000000000000600000000",
            INIT_2D => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000005400000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000001100000000000000030000000000000000000000000000000000000000",
            INIT_39 => X"0000005500000000000000070000000000000006000000000000000000000000",
            INIT_3A => X"00000067000000000000005d0000000000000053000000000000005c00000000",
            INIT_3B => X"000000070000000000000058000000000000004e000000000000005900000000",
            INIT_3C => X"00000074000000000000006f000000000000006e000000000000005400000000",
            INIT_3D => X"0000003f0000000000000040000000000000000d000000000000000800000000",
            INIT_3E => X"00000041000000000000003d0000000000000045000000000000001d00000000",
            INIT_3F => X"00000049000000000000000f0000000000000047000000000000004f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000c000000000000006c0000000000000066000000000000005e00000000",
            INIT_41 => X"0000000e000000000000004f0000000000000018000000000000000d00000000",
            INIT_42 => X"0000003e000000000000003e0000000000000038000000000000003900000000",
            INIT_43 => X"0000003f00000000000000320000000000000026000000000000001700000000",
            INIT_44 => X"0000000100000000000000380000000000000046000000000000004000000000",
            INIT_45 => X"0000002000000000000000070000000000000055000000000000002a00000000",
            INIT_46 => X"0000001500000000000000280000000000000038000000000000003100000000",
            INIT_47 => X"0000003c000000000000002d000000000000001d000000000000002200000000",
            INIT_48 => X"00000037000000000000002c000000000000003a000000000000002700000000",
            INIT_49 => X"00000031000000000000001d0000000000000014000000000000004f00000000",
            INIT_4A => X"0000001800000000000000140000000000000020000000000000003900000000",
            INIT_4B => X"0000003a000000000000004d0000000000000036000000000000002700000000",
            INIT_4C => X"00000045000000000000003e0000000000000035000000000000003c00000000",
            INIT_4D => X"0000002600000000000000310000000000000022000000000000001f00000000",
            INIT_4E => X"00000021000000000000001d0000000000000014000000000000001e00000000",
            INIT_4F => X"000000460000000000000047000000000000004c000000000000003200000000",
            INIT_50 => X"000000310000000000000037000000000000005b000000000000003e00000000",
            INIT_51 => X"00000021000000000000000f0000000000000034000000000000001b00000000",
            INIT_52 => X"000000310000000000000021000000000000001a000000000000001400000000",
            INIT_53 => X"0000003e000000000000004a000000000000003e000000000000003300000000",
            INIT_54 => X"0000002000000000000000320000000000000020000000000000006600000000",
            INIT_55 => X"0000002c00000000000000140000000000000036000000000000001800000000",
            INIT_56 => X"00000041000000000000001b0000000000000035000000000000002f00000000",
            INIT_57 => X"0000003f000000000000003a000000000000004c000000000000002a00000000",
            INIT_58 => X"00000028000000000000001b000000000000001a000000000000003200000000",
            INIT_59 => X"00000039000000000000003b000000000000002d000000000000003300000000",
            INIT_5A => X"00000026000000000000003b000000000000003d000000000000004f00000000",
            INIT_5B => X"0000003000000000000000300000000000000037000000000000003d00000000",
            INIT_5C => X"0000001a00000000000000150000000000000029000000000000002b00000000",
            INIT_5D => X"0000004300000000000000480000000000000038000000000000004a00000000",
            INIT_5E => X"0000003400000000000000420000000000000049000000000000003b00000000",
            INIT_5F => X"0000002f0000000000000032000000000000001b000000000000004300000000",
            INIT_60 => X"0000002e00000000000000290000000000000024000000000000003e00000000",
            INIT_61 => X"0000003c000000000000003c0000000000000031000000000000005300000000",
            INIT_62 => X"0000004100000000000000360000000000000046000000000000004300000000",
            INIT_63 => X"0000003800000000000000370000000000000029000000000000001d00000000",
            INIT_64 => X"00000049000000000000003d0000000000000033000000000000003000000000",
            INIT_65 => X"000000450000000000000034000000000000003c000000000000003500000000",
            INIT_66 => X"000000250000000000000043000000000000003a000000000000003c00000000",
            INIT_67 => X"00000039000000000000003e000000000000004d000000000000002600000000",
            INIT_68 => X"0000003600000000000000460000000000000046000000000000004100000000",
            INIT_69 => X"000000400000000000000032000000000000003e000000000000003b00000000",
            INIT_6A => X"0000001f000000000000002c0000000000000049000000000000003e00000000",
            INIT_6B => X"0000004900000000000000480000000000000046000000000000003900000000",
            INIT_6C => X"0000003b00000000000000390000000000000038000000000000004c00000000",
            INIT_6D => X"0000003b00000000000000390000000000000031000000000000003f00000000",
            INIT_6E => X"0000002e00000000000000100000000000000038000000000000003f00000000",
            INIT_6F => X"0000004b0000000000000041000000000000004c000000000000004600000000",
            INIT_70 => X"00000038000000000000003a0000000000000036000000000000003400000000",
            INIT_71 => X"0000007e000000000000000e0000000000000035000000000000003d00000000",
            INIT_72 => X"000000240000000000000012000000000000000c000000000000003100000000",
            INIT_73 => X"000000000000000000000000000000000000001b000000000000001500000000",
            INIT_74 => X"00000017000000000000001a000000000000001d000000000000006500000000",
            INIT_75 => X"0000004900000000000000500000000000000011000000000000001400000000",
            INIT_76 => X"0000001b00000000000000050000000000000006000000000000002600000000",
            INIT_77 => X"0000006c00000000000000000000000000000003000000000000001600000000",
            INIT_78 => X"0000001200000000000000120000000000000009000000000000000400000000",
            INIT_79 => X"0000002b00000000000000670000000000000024000000000000001200000000",
            INIT_7A => X"00000026000000000000000b0000000000000000000000000000002700000000",
            INIT_7B => X"0000000b0000000000000023000000000000001a000000000000000400000000",
            INIT_7C => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_7D => X"0000003200000000000000000000000000000043000000000000004200000000",
            INIT_7E => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000260000000000000000000000000000004a00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE58;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59 : if BRAM_NAME = "samplegold_layersamples_instance59" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001900000000000000000000000000000008000000000000000000000000",
            INIT_01 => X"00000007000000000000003c0000000000000000000000000000000000000000",
            INIT_02 => X"0000003400000000000000190000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000016000000000000001b00000000",
            INIT_04 => X"0000000000000000000000020000000000000000000000000000000c00000000",
            INIT_05 => X"000000000000000000000002000000000000001f000000000000000000000000",
            INIT_06 => X"000000190000000000000029000000000000000d000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000002300000000",
            INIT_08 => X"0000000c00000000000000000000000000000001000000000000000000000000",
            INIT_09 => X"0000002800000000000000000000000000000016000000000000000000000000",
            INIT_0A => X"00000020000000000000001b0000000000000010000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"00000000000000000000004b0000000000000000000000000000000600000000",
            INIT_0D => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000f000000000000002b0000000000000000000000000000001200000000",
            INIT_0F => X"0000000900000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000030000000000000000b00000000",
            INIT_11 => X"00000000000000000000003e0000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000410000000000000000000000000000000500000000",
            INIT_13 => X"0000000700000000000000000000000000000000000000000000002700000000",
            INIT_14 => X"0000000000000000000000020000000000000005000000000000000000000000",
            INIT_15 => X"0000000000000000000000240000000000000000000000000000000000000000",
            INIT_16 => X"0000001b0000000000000006000000000000001e000000000000001600000000",
            INIT_17 => X"0000000000000000000000150000000000000000000000000000000000000000",
            INIT_18 => X"0000000d000000000000001d0000000000000000000000000000000200000000",
            INIT_19 => X"0000001b00000000000000130000000000000000000000000000000000000000",
            INIT_1A => X"00000000000000000000000f0000000000000000000000000000001100000000",
            INIT_1B => X"0000000000000000000000010000000000000025000000000000000000000000",
            INIT_1C => X"000000000000000000000008000000000000000f000000000000000000000000",
            INIT_1D => X"00000013000000000000000a000000000000002f000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000002f00000000000000000000000000000000000000000000001500000000",
            INIT_20 => X"0000000000000000000000000000000000000005000000000000001c00000000",
            INIT_21 => X"0000000d000000000000000c000000000000000b000000000000002100000000",
            INIT_22 => X"0000001600000000000000000000000000000000000000000000000700000000",
            INIT_23 => X"0000000000000000000000220000000000000000000000000000000500000000",
            INIT_24 => X"0000001b000000000000000a0000000000000000000000000000000600000000",
            INIT_25 => X"0000001500000000000000270000000000000000000000000000000f00000000",
            INIT_26 => X"00000013000000000000000f0000000000000000000000000000000000000000",
            INIT_27 => X"0000001100000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000001300000000000000130000000000000027000000000000000000000000",
            INIT_29 => X"0000000d0000000000000012000000000000001d000000000000000600000000",
            INIT_2A => X"0000000000000000000000050000000000000000000000000000000100000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"00000004000000000000000f0000000000000000000000000000000000000000",
            INIT_2E => X"000000000000000000000000000000000000000c000000000000000900000000",
            INIT_2F => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"00000000000000000000000b0000000000000011000000000000000000000000",
            INIT_32 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000000d000000000000000500000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000a00000000000000030000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"000000000000000000000000000000000000000c000000000000000700000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"00000013000000000000000b0000000000000000000000000000000000000000",
            INIT_63 => X"0000000200000000000000060000000000000012000000000000000300000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000030000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000160000000000000016000000000000000000000000",
            INIT_67 => X"0000000e00000000000000070000000000000021000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000001000000000",
            INIT_69 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"00000001000000000000003b000000000000002b000000000000000f00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000013000000000000001700000000",
            INIT_6F => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000c00000000000000150000000000000002000000000000000000000000",
            INIT_71 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000001600000000000000110000000000000008000000000000000000000000",
            INIT_73 => X"0000000000000000000000060000000000000000000000000000000300000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000300000000000000000000000000000007000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000010000000000000001700000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_7A => X"000000000000000000000000000000000000000f000000000000000200000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000001000000000000000100000000000000005000000000000000000000000",
            INIT_7D => X"000000100000000000000001000000000000000b000000000000000900000000",
            INIT_7E => X"00000011000000000000000b0000000000000014000000000000000000000000",
            INIT_7F => X"0000000000000000000000120000000000000029000000000000005f00000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE59;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60 : if BRAM_NAME = "samplegold_layersamples_instance60" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_02 => X"0000000000000000000000090000000000000009000000000000000900000000",
            INIT_03 => X"00000000000000000000001a0000000000000039000000000000001500000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000000000000000000001b000000000000001f00000000",
            INIT_06 => X"00000000000000000000000d000000000000001c000000000000000000000000",
            INIT_07 => X"000000000000000000000000000000000000000b000000000000000700000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000180000000000000019000000000000000f000000000000000300000000",
            INIT_0A => X"0000000c00000000000000010000000000000000000000000000000e00000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_0C => X"00000000000000000000002b0000000000000010000000000000000c00000000",
            INIT_0D => X"000000000000000000000016000000000000000b000000000000000300000000",
            INIT_0E => X"00000001000000000000000a000000000000000b000000000000001000000000",
            INIT_0F => X"0000000000000000000000000000000000000009000000000000000000000000",
            INIT_10 => X"00000018000000000000000f0000000000000017000000000000001000000000",
            INIT_11 => X"0000001100000000000000070000000000000018000000000000002100000000",
            INIT_12 => X"000000050000000000000000000000000000001b000000000000002200000000",
            INIT_13 => X"0000000800000000000000020000000000000000000000000000000400000000",
            INIT_14 => X"0000001e00000000000000170000000000000016000000000000000000000000",
            INIT_15 => X"0000000d00000000000000050000000000000003000000000000001300000000",
            INIT_16 => X"0000000000000000000000170000000000000006000000000000000000000000",
            INIT_17 => X"0000000d0000000000000004000000000000000a000000000000000700000000",
            INIT_18 => X"0000000000000000000000190000000000000021000000000000003100000000",
            INIT_19 => X"0000000100000000000000000000000000000005000000000000000900000000",
            INIT_1A => X"00000062000000000000000e0000000000000000000000000000001000000000",
            INIT_1B => X"0000005e00000000000000620000000000000061000000000000006500000000",
            INIT_1C => X"0000004c00000000000000230000000000000062000000000000006400000000",
            INIT_1D => X"0000006b000000000000006e000000000000006e000000000000007500000000",
            INIT_1E => X"0000006b000000000000005f0000000000000000000000000000000000000000",
            INIT_1F => X"0000007f000000000000007d000000000000006c000000000000008800000000",
            INIT_20 => X"0000009d000000000000005c0000000000000055000000000000008800000000",
            INIT_21 => X"0000000000000000000000810000000000000087000000000000009100000000",
            INIT_22 => X"000000ae000000000000005f0000000000000049000000000000000000000000",
            INIT_23 => X"000000800000000000000076000000000000005d000000000000008700000000",
            INIT_24 => X"000000b600000000000000b8000000000000008b000000000000007000000000",
            INIT_25 => X"0000000a000000000000000000000000000000a600000000000000b100000000",
            INIT_26 => X"000000ab00000000000000b00000000000000076000000000000005700000000",
            INIT_27 => X"0000006e0000000000000053000000000000004f000000000000006200000000",
            INIT_28 => X"000000c300000000000000ca00000000000000c000000000000000b100000000",
            INIT_29 => X"000000a10000000000000073000000000000008e00000000000000c300000000",
            INIT_2A => X"000000a200000000000000b40000000000000090000000000000007100000000",
            INIT_2B => X"000000aa00000000000000710000000000000060000000000000006d00000000",
            INIT_2C => X"000000a700000000000000b400000000000000da00000000000000cb00000000",
            INIT_2D => X"0000007d00000000000000ac00000000000000a200000000000000a800000000",
            INIT_2E => X"00000069000000000000009600000000000000aa000000000000009800000000",
            INIT_2F => X"000000d800000000000000980000000000000072000000000000006900000000",
            INIT_30 => X"000000a9000000000000009800000000000000bb00000000000000e300000000",
            INIT_31 => X"0000008a0000000000000091000000000000008800000000000000a000000000",
            INIT_32 => X"00000087000000000000007b0000000000000090000000000000009700000000",
            INIT_33 => X"000000e500000000000000cb0000000000000099000000000000008b00000000",
            INIT_34 => X"000000a300000000000000a900000000000000a300000000000000da00000000",
            INIT_35 => X"0000009f00000000000000a80000000000000095000000000000007000000000",
            INIT_36 => X"000000840000000000000094000000000000007200000000000000a300000000",
            INIT_37 => X"000000e100000000000000e000000000000000ae000000000000009700000000",
            INIT_38 => X"00000093000000000000009100000000000000a700000000000000ca00000000",
            INIT_39 => X"0000009c00000000000000b200000000000000c2000000000000008700000000",
            INIT_3A => X"0000008d00000000000000750000000000000066000000000000008d00000000",
            INIT_3B => X"000000bb00000000000000b70000000000000080000000000000004700000000",
            INIT_3C => X"000000a700000000000000af000000000000009600000000000000b800000000",
            INIT_3D => X"000000a600000000000000cd00000000000000cb00000000000000b400000000",
            INIT_3E => X"0000006b000000000000007a000000000000007d000000000000006200000000",
            INIT_3F => X"000000c40000000000000076000000000000006e000000000000005c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000b300000000000000af00000000000000ba00000000000000a600000000",
            INIT_41 => X"000000b100000000000000b200000000000000a8000000000000009e00000000",
            INIT_42 => X"0000007c000000000000006d000000000000006b000000000000007a00000000",
            INIT_43 => X"000000ae00000000000000c00000000000000065000000000000007200000000",
            INIT_44 => X"0000009d00000000000000be00000000000000ca00000000000000b200000000",
            INIT_45 => X"0000006e000000000000009d00000000000000a0000000000000009600000000",
            INIT_46 => X"0000007100000000000000890000000000000078000000000000006000000000",
            INIT_47 => X"000000ad00000000000000a900000000000000b7000000000000005d00000000",
            INIT_48 => X"0000009e000000000000006300000000000000ae00000000000000c800000000",
            INIT_49 => X"000000670000000000000063000000000000008d000000000000009900000000",
            INIT_4A => X"0000006000000000000000720000000000000076000000000000006d00000000",
            INIT_4B => X"000000cc000000000000009c000000000000009500000000000000ae00000000",
            INIT_4C => X"0000007a0000000000000083000000000000006900000000000000af00000000",
            INIT_4D => X"0000005f000000000000005d0000000000000050000000000000006b00000000",
            INIT_4E => X"0000009f000000000000006d0000000000000055000000000000005600000000",
            INIT_4F => X"000000b500000000000000c70000000000000083000000000000009000000000",
            INIT_50 => X"0000004f00000000000000640000000000000073000000000000009b00000000",
            INIT_51 => X"00000052000000000000005e0000000000000056000000000000004300000000",
            INIT_52 => X"0000000000000000000000000000000000000067000000000000005300000000",
            INIT_53 => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_54 => X"0000002d00000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_5B => X"0000002c000000000000002c0000000000000010000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000210000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000001100000000",
            INIT_62 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000018000000000000000000000000",
            INIT_64 => X"0000001300000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_66 => X"0000001700000000000000060000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000360000000000000000000000000000000000000000",
            INIT_6A => X"00000000000000000000000a0000000000000000000000000000000b00000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_6E => X"0000000000000000000000130000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000430000000000000010000000000000000700000000",
            INIT_70 => X"0000000000000000000000070000000000000000000000000000001500000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"00000000000000000000000a0000000000000000000000000000000000000000",
            INIT_73 => X"0000002d00000000000000430000000000000001000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"00000000000000000000001e000000000000000c000000000000000000000000",
            INIT_76 => X"0000002000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000011000000000000000000000000",
            INIT_79 => X"0000000600000000000000000000000000000018000000000000000000000000",
            INIT_7A => X"000000000000000000000000000000000000002d000000000000000000000000",
            INIT_7B => X"0000000000000000000000090000000000000007000000000000000000000000",
            INIT_7C => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000400000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000040000000000000000000000000000000f00000000",
            INIT_7F => X"0000000700000000000000010000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE60;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61 : if BRAM_NAME = "samplegold_layersamples_instance61" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002100000000000000290000000000000000000000000000000000000000",
            INIT_01 => X"0000000d0000000000000018000000000000000e000000000000000000000000",
            INIT_02 => X"0000000000000000000000220000000000000003000000000000000000000000",
            INIT_03 => X"00000000000000000000000e0000000000000007000000000000000000000000",
            INIT_04 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"000000000000000000000008000000000000001a000000000000001100000000",
            INIT_06 => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_07 => X"0000000000000000000000140000000000000000000000000000001900000000",
            INIT_08 => X"0000000600000000000000250000000000000014000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000001c00000000",
            INIT_0A => X"0000001300000000000000030000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000004900000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"000000000000000000000000000000000000002e000000000000000000000000",
            INIT_0E => X"0000003800000000000000140000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000003a00000000",
            INIT_12 => X"0000002700000000000000220000000000000012000000000000000000000000",
            INIT_13 => X"000000030000000000000000000000000000001d000000000000000000000000",
            INIT_14 => X"0000001700000000000000000000000000000000000000000000000e00000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000019000000000000001a000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000002b00000000",
            INIT_18 => X"000000130000000000000000000000000000002c000000000000000500000000",
            INIT_19 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_1A => X"0000003000000000000000000000000000000000000000000000000100000000",
            INIT_1B => X"0000000d00000000000000000000000000000000000000000000000900000000",
            INIT_1C => X"00000000000000000000000f000000000000000a000000000000002400000000",
            INIT_1D => X"0000000000000000000000000000000000000008000000000000000000000000",
            INIT_1E => X"0000000500000000000000130000000000000000000000000000000000000000",
            INIT_1F => X"0000001d00000000000000070000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000018000000000000001200000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000150000000000000003000000000000000000000000",
            INIT_23 => X"0000001200000000000000160000000000000000000000000000001000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000001400000000",
            INIT_25 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000005000000000000000000000000",
            INIT_27 => X"0000001600000000000000000000000000000005000000000000000700000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_29 => X"0000000000000000000000100000000000000000000000000000000000000000",
            INIT_2A => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000002b00000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_2D => X"0000000e000000000000000d0000000000000000000000000000000000000000",
            INIT_2E => X"0000000100000000000000000000000000000000000000000000000500000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000d00000000000000000000000000000000000000000000000900000000",
            INIT_31 => X"0000001700000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000c00000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"00000000000000000000001e0000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000040000000000000014000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000001000000000000000500000000",
            INIT_3A => X"0000000000000000000000000000000000000004000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000008000000000000001300000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000c00000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000001800000000",
            INIT_41 => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000f0000000000000044000000000000007b000000000000001400000000",
            INIT_44 => X"00000026000000000000001c0000000000000024000000000000001b00000000",
            INIT_45 => X"0000003600000000000000620000000000000000000000000000000100000000",
            INIT_46 => X"00000016000000000000001b0000000000000023000000000000002100000000",
            INIT_47 => X"0000001d00000000000000160000000000000062000000000000005300000000",
            INIT_48 => X"00000015000000000000002c0000000000000024000000000000001000000000",
            INIT_49 => X"000000190000000000000024000000000000009c000000000000000000000000",
            INIT_4A => X"0000002e00000000000000140000000000000017000000000000001c00000000",
            INIT_4B => X"0000000000000000000000390000000000000028000000000000008000000000",
            INIT_4C => X"0000001300000000000000020000000000000026000000000000000600000000",
            INIT_4D => X"00000021000000000000001a0000000000000027000000000000006100000000",
            INIT_4E => X"00000091000000000000004f0000000000000005000000000000001b00000000",
            INIT_4F => X"0000000200000000000000000000000000000047000000000000000000000000",
            INIT_50 => X"000000270000000000000053000000000000001c000000000000000000000000",
            INIT_51 => X"00000029000000000000000c000000000000001a000000000000004800000000",
            INIT_52 => X"0000000000000000000000290000000000000056000000000000000600000000",
            INIT_53 => X"0000000000000000000000000000000000000012000000000000005700000000",
            INIT_54 => X"0000005300000000000000370000000000000039000000000000002000000000",
            INIT_55 => X"0000001b000000000000003e0000000000000000000000000000001a00000000",
            INIT_56 => X"0000003e0000000000000000000000000000001a000000000000002900000000",
            INIT_57 => X"0000002800000000000000000000000000000000000000000000001100000000",
            INIT_58 => X"0000001d00000000000000560000000000000033000000000000003900000000",
            INIT_59 => X"0000001d000000000000001c000000000000002a000000000000000000000000",
            INIT_5A => X"00000015000000000000000f000000000000002d000000000000000000000000",
            INIT_5B => X"0000002d0000000000000010000000000000001e000000000000000000000000",
            INIT_5C => X"0000001100000000000000240000000000000058000000000000003000000000",
            INIT_5D => X"0000000000000000000000210000000000000012000000000000000c00000000",
            INIT_5E => X"0000000000000000000000190000000000000007000000000000005f00000000",
            INIT_5F => X"0000001c000000000000001d0000000000000021000000000000001b00000000",
            INIT_60 => X"000000240000000000000014000000000000003d000000000000003400000000",
            INIT_61 => X"000000420000000000000004000000000000001f000000000000000000000000",
            INIT_62 => X"000000000000000000000008000000000000001e000000000000001200000000",
            INIT_63 => X"0000000400000000000000220000000000000001000000000000003b00000000",
            INIT_64 => X"0000000c000000000000004f000000000000000a000000000000004800000000",
            INIT_65 => X"0000002000000000000000150000000000000028000000000000002400000000",
            INIT_66 => X"000000090000000000000000000000000000000d000000000000001400000000",
            INIT_67 => X"0000002500000000000000190000000000000000000000000000003100000000",
            INIT_68 => X"00000007000000000000001c0000000000000032000000000000001a00000000",
            INIT_69 => X"00000000000000000000001d0000000000000018000000000000003300000000",
            INIT_6A => X"0000000000000000000000000000000000000018000000000000003200000000",
            INIT_6B => X"000000000000000000000023000000000000002c000000000000000f00000000",
            INIT_6C => X"0000004c00000000000000000000000000000022000000000000001700000000",
            INIT_6D => X"000000310000000000000000000000000000000d000000000000001600000000",
            INIT_6E => X"000000430000000000000000000000000000000c000000000000001700000000",
            INIT_6F => X"0000000200000000000000070000000000000026000000000000001300000000",
            INIT_70 => X"000000190000000000000042000000000000000d000000000000001c00000000",
            INIT_71 => X"0000000f00000000000000300000000000000000000000000000000000000000",
            INIT_72 => X"0000000e00000000000000330000000000000000000000000000000000000000",
            INIT_73 => X"000000130000000000000011000000000000000b000000000000001500000000",
            INIT_74 => X"0000000000000000000000290000000000000041000000000000000f00000000",
            INIT_75 => X"00000000000000000000000c000000000000000b000000000000002700000000",
            INIT_76 => X"000000000000000000000015000000000000002a000000000000000000000000",
            INIT_77 => X"0000001d000000000000000c0000000000000020000000000000002f00000000",
            INIT_78 => X"000000060000000000000005000000000000003b000000000000002f00000000",
            INIT_79 => X"0000002e00000000000000000000000000000014000000000000000000000000",
            INIT_7A => X"0000002c000000000000000b000000000000001f000000000000001b00000000",
            INIT_7B => X"0000000000000000000000000000000000000002000000000000001b00000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000200000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE61;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62 : if BRAM_NAME = "samplegold_layersamples_instance62" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"00000000000000000000000e0000000000000000000000000000000000000000",
            INIT_02 => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"00000073000000000000005e0000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000003700000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000900000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000020000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"000000250000000000000025000000000000002c000000000000002a00000000",
            INIT_35 => X"0000001b000000000000002b0000000000000029000000000000003000000000",
            INIT_36 => X"0000003b000000000000003c0000000000000036000000000000000000000000",
            INIT_37 => X"0000001d00000000000000000000000000000000000000000000003d00000000",
            INIT_38 => X"0000001e00000000000000230000000000000018000000000000001600000000",
            INIT_39 => X"0000000200000000000000160000000000000032000000000000002900000000",
            INIT_3A => X"0000003c000000000000003a0000000000000039000000000000003300000000",
            INIT_3B => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"00000012000000000000000d0000000000000028000000000000001500000000",
            INIT_3D => X"0000002100000000000000250000000000000000000000000000001b00000000",
            INIT_3E => X"0000000b00000000000000340000000000000031000000000000002e00000000",
            INIT_3F => X"00000012000000000000002e000000000000001f000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000050000000000000019000000000000001c000000000000001c00000000",
            INIT_41 => X"00000036000000000000001e0000000000000024000000000000000200000000",
            INIT_42 => X"000000220000000000000020000000000000001e000000000000003900000000",
            INIT_43 => X"0000001b000000000000000f0000000000000021000000000000002800000000",
            INIT_44 => X"000000010000000000000003000000000000001b000000000000002400000000",
            INIT_45 => X"0000003000000000000000300000000000000031000000000000001300000000",
            INIT_46 => X"0000002b00000000000000230000000000000027000000000000002000000000",
            INIT_47 => X"000000240000000000000020000000000000001d000000000000001d00000000",
            INIT_48 => X"0000001300000000000000060000000000000010000000000000000200000000",
            INIT_49 => X"0000002200000000000000320000000000000033000000000000002600000000",
            INIT_4A => X"0000002300000000000000300000000000000023000000000000002b00000000",
            INIT_4B => X"0000000000000000000000210000000000000004000000000000002000000000",
            INIT_4C => X"0000002b000000000000000c000000000000000f000000000000002100000000",
            INIT_4D => X"0000002b00000000000000290000000000000033000000000000003200000000",
            INIT_4E => X"0000002a000000000000001e0000000000000038000000000000002300000000",
            INIT_4F => X"0000000a0000000000000025000000000000000c000000000000002300000000",
            INIT_50 => X"0000002800000000000000180000000000000026000000000000001200000000",
            INIT_51 => X"00000017000000000000002f000000000000001b000000000000003c00000000",
            INIT_52 => X"0000002a000000000000001c000000000000002e000000000000002400000000",
            INIT_53 => X"0000001600000000000000090000000000000022000000000000002200000000",
            INIT_54 => X"0000001b000000000000000f0000000000000020000000000000002400000000",
            INIT_55 => X"0000002b000000000000001f000000000000002a000000000000001600000000",
            INIT_56 => X"0000001b00000000000000240000000000000023000000000000002600000000",
            INIT_57 => X"0000002c0000000000000016000000000000002a000000000000001c00000000",
            INIT_58 => X"0000002200000000000000280000000000000016000000000000001b00000000",
            INIT_59 => X"0000002b0000000000000018000000000000002a000000000000002800000000",
            INIT_5A => X"0000001d00000000000000170000000000000030000000000000002700000000",
            INIT_5B => X"0000002000000000000000080000000000000036000000000000002300000000",
            INIT_5C => X"00000027000000000000001b000000000000001d000000000000002400000000",
            INIT_5D => X"00000036000000000000002a0000000000000018000000000000002a00000000",
            INIT_5E => X"0000002c0000000000000026000000000000002a000000000000002100000000",
            INIT_5F => X"0000001f000000000000001e0000000000000013000000000000001e00000000",
            INIT_60 => X"0000002500000000000000260000000000000018000000000000002100000000",
            INIT_61 => X"00000006000000000000003a0000000000000027000000000000001900000000",
            INIT_62 => X"0000001600000000000000260000000000000027000000000000002700000000",
            INIT_63 => X"00000010000000000000001d0000000000000015000000000000001500000000",
            INIT_64 => X"0000001100000000000000230000000000000026000000000000001900000000",
            INIT_65 => X"000000320000000000000023000000000000002b000000000000002200000000",
            INIT_66 => X"000000140000000000000006000000000000001b000000000000002100000000",
            INIT_67 => X"00000016000000000000000b0000000000000011000000000000001200000000",
            INIT_68 => X"0000001b0000000000000010000000000000001b000000000000001900000000",
            INIT_69 => X"00000019000000000000001e000000000000002f000000000000002300000000",
            INIT_6A => X"00000013000000000000000f0000000000000001000000000000001700000000",
            INIT_6B => X"0000001600000000000000150000000000000015000000000000000f00000000",
            INIT_6C => X"00000010000000000000000d0000000000000000000000000000000000000000",
            INIT_6D => X"0000001800000000000000060000000000000010000000000000000000000000",
            INIT_6E => X"0000000600000000000000030000000000000000000000000000004b00000000",
            INIT_6F => X"000000000000000000000014000000000000000b000000000000000a00000000",
            INIT_70 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000002f000000000000000c0000000000000000000000000000000000000000",
            INIT_72 => X"00000008000000000000000c0000000000000007000000000000000000000000",
            INIT_73 => X"0000000000000000000000090000000000000015000000000000000800000000",
            INIT_74 => X"0000000e000000000000002e0000000000000000000000000000000100000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000b00000000000000020000000000000002000000000000000000000000",
            INIT_77 => X"0000002d00000000000000000000000000000000000000000000005100000000",
            INIT_78 => X"00000023000000000000001c0000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000001f00000000000000000000000000000019000000000000000000000000",
            INIT_7B => X"0000000000000000000000350000000000000011000000000000000900000000",
            INIT_7C => X"0000000000000000000000250000000000000009000000000000000000000000",
            INIT_7D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"00000009000000000000000f0000000000000007000000000000003400000000",
            INIT_7F => X"0000000000000000000000000000000000000019000000000000001300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE62;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63 : if BRAM_NAME = "samplegold_layersamples_instance63" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000010000000000000007000000000000001200000000",
            INIT_01 => X"0000003500000000000000080000000000000000000000000000000000000000",
            INIT_02 => X"00000029000000000000000a000000000000001b000000000000002700000000",
            INIT_03 => X"0000001a0000000000000000000000000000000e000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_05 => X"0000002f00000000000000100000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000240000000000000003000000000000002600000000",
            INIT_07 => X"0000001500000000000000000000000000000002000000000000001300000000",
            INIT_08 => X"0000000000000000000000090000000000000006000000000000000000000000",
            INIT_09 => X"0000003600000000000000000000000000000016000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_0B => X"000000000000000000000021000000000000000f000000000000000000000000",
            INIT_0C => X"0000000000000000000000210000000000000001000000000000000700000000",
            INIT_0D => X"0000001500000000000000240000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000000000000000000002a0000000000000002000000000000000000000000",
            INIT_10 => X"0000001400000000000000000000000000000000000000000000001d00000000",
            INIT_11 => X"00000000000000000000002a0000000000000011000000000000000300000000",
            INIT_12 => X"0000000000000000000000240000000000000000000000000000000200000000",
            INIT_13 => X"00000000000000000000002a0000000000000001000000000000000000000000",
            INIT_14 => X"0000000d000000000000000f0000000000000000000000000000000000000000",
            INIT_15 => X"000000000000000000000000000000000000002a000000000000001100000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_17 => X"0000000600000000000000000000000000000022000000000000000a00000000",
            INIT_18 => X"0000001900000000000000110000000000000011000000000000000000000000",
            INIT_19 => X"0000002100000000000000000000000000000000000000000000002900000000",
            INIT_1A => X"0000000e00000000000000010000000000000000000000000000000000000000",
            INIT_1B => X"0000000800000000000000050000000000000000000000000000001400000000",
            INIT_1C => X"0000002f000000000000001e000000000000000c000000000000000000000000",
            INIT_1D => X"0000000000000000000000140000000000000000000000000000000000000000",
            INIT_1E => X"0000000900000000000000110000000000000005000000000000001600000000",
            INIT_1F => X"0000000000000000000000140000000000000005000000000000000100000000",
            INIT_20 => X"000000150000000000000020000000000000001a000000000000000000000000",
            INIT_21 => X"0000001900000000000000180000000000000005000000000000000000000000",
            INIT_22 => X"000000060000000000000000000000000000001e000000000000000000000000",
            INIT_23 => X"000000000000000000000008000000000000000c000000000000000300000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"00000025000000000000001e0000000000000019000000000000001200000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000001b00000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000001800000000000000010000000000000000000000000000000900000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000001e00000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000000000000000000008000000000000001c000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000001d0000000000000024000000000000001a000000000000000d00000000",
            INIT_6D => X"0000000a00000000000000160000000000000018000000000000001d00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"000000280000000000000016000000000000001f000000000000003500000000",
            INIT_71 => X"0000002800000000000000290000000000000028000000000000003000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000e0000000000000015000000000000001a000000000000001200000000",
            INIT_75 => X"00000018000000000000000d0000000000000009000000000000000d00000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_77 => X"0000002100000000000000220000000000000000000000000000000000000000",
            INIT_78 => X"00000033000000000000002a0000000000000010000000000000001800000000",
            INIT_79 => X"000000290000000000000045000000000000002f000000000000001f00000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"000000000000000000000000000000000000000a000000000000001700000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_7F => X"00000012000000000000002a0000000000000017000000000000002700000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE63;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64 : if BRAM_NAME = "samplegold_layersamples_instance64" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d000000000000002c0000000000000027000000000000002900000000",
            INIT_01 => X"000000000000000000000015000000000000001e000000000000001600000000",
            INIT_02 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000002f00000000000000000000000000000000000000000000001700000000",
            INIT_04 => X"0000000300000000000000060000000000000014000000000000000900000000",
            INIT_05 => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_06 => X"0000000900000000000000000000000000000000000000000000000b00000000",
            INIT_07 => X"00000005000000000000000f000000000000001a000000000000003100000000",
            INIT_08 => X"00000032000000000000000b0000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000004000000000000001a00000000",
            INIT_0A => X"0000000600000000000000000000000000000000000000000000000300000000",
            INIT_0B => X"000000000000000000000000000000000000000d000000000000000b00000000",
            INIT_0C => X"0000000a000000000000000c0000000000000001000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000500000000",
            INIT_0F => X"0000000400000000000000260000000000000035000000000000000000000000",
            INIT_10 => X"0000000a0000000000000016000000000000000a000000000000000000000000",
            INIT_11 => X"0000000a000000000000000a0000000000000000000000000000000400000000",
            INIT_12 => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"00000000000000000000000e0000000000000018000000000000000d00000000",
            INIT_14 => X"000000220000000000000022000000000000000c000000000000000c00000000",
            INIT_15 => X"00000028000000000000001d0000000000000012000000000000002500000000",
            INIT_16 => X"0000001c0000000000000027000000000000002b000000000000002300000000",
            INIT_17 => X"000000190000000000000016000000000000001e000000000000001900000000",
            INIT_18 => X"00000023000000000000002b000000000000002b000000000000000900000000",
            INIT_19 => X"0000002b000000000000002c000000000000001f000000000000000b00000000",
            INIT_1A => X"0000000f000000000000000f0000000000000022000000000000002100000000",
            INIT_1B => X"000000150000000000000004000000000000001c000000000000002400000000",
            INIT_1C => X"0000000c000000000000001f000000000000002e000000000000002d00000000",
            INIT_1D => X"0000004a00000000000000510000000000000050000000000000004800000000",
            INIT_1E => X"00000027000000000000002b000000000000003e000000000000004800000000",
            INIT_1F => X"0000002d000000000000000f0000000000000000000000000000001b00000000",
            INIT_20 => X"00000060000000000000000e0000000000000028000000000000002800000000",
            INIT_21 => X"0000004d000000000000004d0000000000000042000000000000004a00000000",
            INIT_22 => X"00000019000000000000002c0000000000000034000000000000005400000000",
            INIT_23 => X"00000027000000000000002c0000000000000008000000000000001100000000",
            INIT_24 => X"0000004d000000000000004f0000000000000018000000000000001b00000000",
            INIT_25 => X"0000004e00000000000000510000000000000050000000000000003a00000000",
            INIT_26 => X"00000018000000000000002b0000000000000044000000000000003e00000000",
            INIT_27 => X"0000002200000000000000200000000000000032000000000000002f00000000",
            INIT_28 => X"0000004c0000000000000046000000000000003f000000000000002000000000",
            INIT_29 => X"000000400000000000000047000000000000003d000000000000004200000000",
            INIT_2A => X"0000002e000000000000002c0000000000000043000000000000003500000000",
            INIT_2B => X"0000002200000000000000240000000000000015000000000000003400000000",
            INIT_2C => X"0000003e000000000000003e000000000000004d000000000000004a00000000",
            INIT_2D => X"0000003500000000000000250000000000000037000000000000004a00000000",
            INIT_2E => X"00000021000000000000002c000000000000002c000000000000003100000000",
            INIT_2F => X"00000034000000000000001b0000000000000031000000000000000b00000000",
            INIT_30 => X"0000002200000000000000330000000000000040000000000000002f00000000",
            INIT_31 => X"0000002f000000000000001e0000000000000028000000000000002000000000",
            INIT_32 => X"0000000a000000000000002a0000000000000047000000000000004300000000",
            INIT_33 => X"0000003800000000000000380000000000000003000000000000003300000000",
            INIT_34 => X"000000470000000000000040000000000000001f000000000000002a00000000",
            INIT_35 => X"0000004300000000000000510000000000000033000000000000002300000000",
            INIT_36 => X"0000001a00000000000000070000000000000023000000000000004800000000",
            INIT_37 => X"0000002b000000000000001d0000000000000029000000000000000d00000000",
            INIT_38 => X"0000002b000000000000003d000000000000001f000000000000004500000000",
            INIT_39 => X"0000005700000000000000200000000000000032000000000000002e00000000",
            INIT_3A => X"0000001300000000000000230000000000000000000000000000002f00000000",
            INIT_3B => X"0000002400000000000000370000000000000025000000000000001900000000",
            INIT_3C => X"0000003e00000000000000320000000000000032000000000000002f00000000",
            INIT_3D => X"00000034000000000000004e000000000000003c000000000000003000000000",
            INIT_3E => X"0000000d00000000000000310000000000000020000000000000000000000000",
            INIT_3F => X"0000003e00000000000000000000000000000026000000000000001500000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000340000000000000027000000000000001300000000",
            INIT_41 => X"00000020000000000000003c0000000000000053000000000000001e00000000",
            INIT_42 => X"0000000d00000000000000140000000000000029000000000000003d00000000",
            INIT_43 => X"0000004e00000000000000200000000000000011000000000000000b00000000",
            INIT_44 => X"00000020000000000000000a000000000000000e000000000000002c00000000",
            INIT_45 => X"0000002700000000000000320000000000000045000000000000005b00000000",
            INIT_46 => X"0000000f00000000000000050000000000000025000000000000002000000000",
            INIT_47 => X"00000033000000000000002d0000000000000022000000000000001900000000",
            INIT_48 => X"00000053000000000000002d0000000000000006000000000000000800000000",
            INIT_49 => X"0000001b000000000000002b000000000000003a000000000000003e00000000",
            INIT_4A => X"0000001900000000000000140000000000000010000000000000002000000000",
            INIT_4B => X"000000140000000000000032000000000000002a000000000000002000000000",
            INIT_4C => X"0000004600000000000000620000000000000025000000000000000b00000000",
            INIT_4D => X"0000003d00000000000000600000000000000055000000000000003a00000000",
            INIT_4E => X"00000034000000000000002b0000000000000033000000000000003a00000000",
            INIT_4F => X"000000520000000000000039000000000000004a000000000000004c00000000",
            INIT_50 => X"0000004d00000000000000500000000000000040000000000000003500000000",
            INIT_51 => X"00000049000000000000005a0000000000000099000000000000007400000000",
            INIT_52 => X"00000038000000000000004f0000000000000056000000000000004600000000",
            INIT_53 => X"0000005d0000000000000044000000000000002f000000000000003600000000",
            INIT_54 => X"0000007500000000000000520000000000000053000000000000001600000000",
            INIT_55 => X"000000460000000000000045000000000000002500000000000000c700000000",
            INIT_56 => X"000000000000000000000032000000000000004b000000000000005b00000000",
            INIT_57 => X"00000000000000000000005e000000000000005d000000000000003500000000",
            INIT_58 => X"000000da00000000000000560000000000000063000000000000005200000000",
            INIT_59 => X"0000006c00000000000000930000000000000056000000000000001200000000",
            INIT_5A => X"00000010000000000000004d0000000000000055000000000000006a00000000",
            INIT_5B => X"0000004d000000000000002d0000000000000065000000000000004c00000000",
            INIT_5C => X"0000002d00000000000000ab0000000000000086000000000000006c00000000",
            INIT_5D => X"0000005e000000000000005e000000000000007c000000000000004b00000000",
            INIT_5E => X"0000003500000000000000100000000000000073000000000000005500000000",
            INIT_5F => X"0000008300000000000000310000000000000030000000000000006700000000",
            INIT_60 => X"00000045000000000000001800000000000000b5000000000000007100000000",
            INIT_61 => X"000000480000000000000059000000000000005d000000000000006800000000",
            INIT_62 => X"000000540000000000000001000000000000001f000000000000005100000000",
            INIT_63 => X"0000004a00000000000000800000000000000036000000000000005100000000",
            INIT_64 => X"0000007d000000000000005c000000000000003a000000000000006e00000000",
            INIT_65 => X"0000005e0000000000000069000000000000004b000000000000005e00000000",
            INIT_66 => X"0000004300000000000000310000000000000025000000000000001f00000000",
            INIT_67 => X"0000008d00000000000000000000000000000080000000000000005f00000000",
            INIT_68 => X"00000063000000000000003c000000000000004e000000000000005700000000",
            INIT_69 => X"0000003a000000000000004d0000000000000036000000000000004700000000",
            INIT_6A => X"000000620000000000000000000000000000001e000000000000000600000000",
            INIT_6B => X"0000001e0000000000000083000000000000000e000000000000008700000000",
            INIT_6C => X"0000001900000000000000520000000000000049000000000000004100000000",
            INIT_6D => X"0000000800000000000000230000000000000061000000000000000c00000000",
            INIT_6E => X"000000af00000000000000690000000000000000000000000000005600000000",
            INIT_6F => X"0000004900000000000000180000000000000055000000000000002500000000",
            INIT_70 => X"0000003a00000000000000690000000000000004000000000000001e00000000",
            INIT_71 => X"00000067000000000000004f0000000000000046000000000000005c00000000",
            INIT_72 => X"0000003100000000000000bd0000000000000055000000000000000000000000",
            INIT_73 => X"00000006000000000000000b0000000000000031000000000000004400000000",
            INIT_74 => X"00000039000000000000004e0000000000000000000000000000007100000000",
            INIT_75 => X"00000000000000000000002b000000000000005a000000000000000500000000",
            INIT_76 => X"0000003c000000000000000200000000000000d1000000000000006800000000",
            INIT_77 => X"0000006900000000000000090000000000000019000000000000006900000000",
            INIT_78 => X"0000004a0000000000000041000000000000004e000000000000000000000000",
            INIT_79 => X"0000005700000000000000000000000000000027000000000000008500000000",
            INIT_7A => X"00000060000000000000005e0000000000000029000000000000009300000000",
            INIT_7B => X"000000000000000000000010000000000000001c000000000000004b00000000",
            INIT_7C => X"0000005600000000000000ba0000000000000060000000000000000000000000",
            INIT_7D => X"0000007a00000000000000500000000000000000000000000000000000000000",
            INIT_7E => X"0000006800000000000000460000000000000066000000000000008000000000",
            INIT_7F => X"00000006000000000000000a000000000000000d000000000000001500000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE64;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65 : if BRAM_NAME = "samplegold_layersamples_instance65" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000003f00000000000000bf000000000000002800000000",
            INIT_01 => X"0000008000000000000000610000000000000066000000000000000000000000",
            INIT_02 => X"000000200000000000000046000000000000003d000000000000006300000000",
            INIT_03 => X"00000022000000000000001e0000000000000019000000000000001d00000000",
            INIT_04 => X"0000000000000000000000000000000000000042000000000000007700000000",
            INIT_05 => X"0000000000000000000000170000000000000021000000000000001c00000000",
            INIT_06 => X"000000610000000000000036000000000000001d000000000000000000000000",
            INIT_07 => X"0000000000000000000000040000000000000007000000000000003000000000",
            INIT_08 => X"0000000d0000000000000013000000000000002e000000000000002600000000",
            INIT_09 => X"0000000000000000000000000000000000000002000000000000000d00000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_0D => X"0000003200000000000000000000000000000001000000000000000000000000",
            INIT_0E => X"00000000000000000000000e000000000000003d000000000000003a00000000",
            INIT_0F => X"000000000000000000000000000000000000000a000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000700000000000000000000000000000012000000000000000000000000",
            INIT_12 => X"00000002000000000000001d0000000000000006000000000000000000000000",
            INIT_13 => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000700000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"00000000000000000000006a0000000000000021000000000000000c00000000",
            INIT_18 => X"0000000000000000000000020000000000000006000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000004a0000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000002000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"000000000000000000000009000000000000000d000000000000001f00000000",
            INIT_24 => X"0000003a00000000000000060000000000000005000000000000000000000000",
            INIT_25 => X"000000bd00000000000000ab00000000000000b500000000000000b800000000",
            INIT_26 => X"000000000000000000000000000000000000002e00000000000000a000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_2C => X"000000040000000000000000000000000000001c000000000000002e00000000",
            INIT_2D => X"0000001f0000000000000000000000000000001e000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_2F => X"000000000000000000000000000000000000001f000000000000004300000000",
            INIT_30 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"00000000000000000000006b0000000000000053000000000000000000000000",
            INIT_33 => X"000000000000000000000000000000000000001a000000000000000a00000000",
            INIT_34 => X"0000003a000000000000005b0000000000000062000000000000000000000000",
            INIT_35 => X"00000006000000000000001d0000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000001a00000000000000140000000000000013000000000000000400000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_3B => X"000000000000000000000004000000000000000f000000000000001100000000",
            INIT_3C => X"00000000000000000000000c0000000000000000000000000000000000000000",
            INIT_3D => X"000000270000000000000022000000000000001d000000000000001b00000000",
            INIT_3E => X"00000006000000000000000d000000000000001b000000000000003200000000",
            INIT_3F => X"00000029000000000000001b0000000000000014000000000000000c00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000022000000000000002a0000000000000020000000000000001b00000000",
            INIT_41 => X"0000002800000000000000250000000000000017000000000000001600000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000001f000000000000001f0000000000000004000000000000000000000000",
            INIT_44 => X"000000170000000000000022000000000000003a000000000000002400000000",
            INIT_45 => X"000000000000000000000031000000000000001d000000000000001700000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"00000039000000000000001b0000000000000000000000000000000000000000",
            INIT_48 => X"0000001e00000000000000170000000000000024000000000000003c00000000",
            INIT_49 => X"000000000000000000000000000000000000001c000000000000001600000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000003d000000000000001b000000000000000c000000000000000000000000",
            INIT_4C => X"00000022000000000000001f0000000000000015000000000000003400000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"000000240000000000000020000000000000000b000000000000000000000000",
            INIT_50 => X"00000003000000000000000a0000000000000029000000000000001100000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000001d00000000000000170000000000000016000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000021000000000000002d00000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000003800000000000000330000000000000004000000000000000000000000",
            INIT_58 => X"000000000000000000000000000000000000002f000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"000000140000000000000027000000000000002c000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000001a00000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000f0000000000000002000000000000003a000000000000001f00000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000001800000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000400000000000000000000000000000007000000000000002700000000",
            INIT_64 => X"0000000000000000000000190000000000000000000000000000000000000000",
            INIT_65 => X"0000000f00000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000003300000000000000040000000000000000000000000000000000000000",
            INIT_67 => X"00000004000000000000000d0000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"000000000000000000000004000000000000000b000000000000000000000000",
            INIT_6A => X"0000000500000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000009000000000000001800000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_70 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000a00000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000d00000000000000020000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000007000000000000000500000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000001400000000000000120000000000000000000000000000000000000000",
            INIT_7B => X"000000000000000000000008000000000000000f000000000000000a00000000",
            INIT_7C => X"0000000800000000000000000000000000000000000000000000000900000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"00000000000000000000000e000000000000000c000000000000002200000000",
            INIT_7F => X"00000002000000000000003e0000000000000019000000000000000600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE65;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66 : if BRAM_NAME = "samplegold_layersamples_instance66" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000000000000000000001a0000000000000000000000000000000000000000",
            INIT_01 => X"0000004a00000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_03 => X"00000000000000000000002d0000000000000000000000000000000d00000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"00000016000000000000002a0000000000000000000000000000000000000000",
            INIT_06 => X"0000000c000000000000000c000000000000000a000000000000000000000000",
            INIT_07 => X"00000000000000000000000b000000000000003c000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000017000000000000000500000000",
            INIT_09 => X"000000070000000000000011000000000000002b000000000000000000000000",
            INIT_0A => X"0000000f00000000000000130000000000000004000000000000000800000000",
            INIT_0B => X"0000000000000000000000000000000000000039000000000000001b00000000",
            INIT_0C => X"0000000000000000000000080000000000000000000000000000001900000000",
            INIT_0D => X"000000050000000000000000000000000000000f000000000000001900000000",
            INIT_0E => X"0000002d00000000000000000000000000000006000000000000001f00000000",
            INIT_0F => X"0000000100000000000000030000000000000024000000000000002a00000000",
            INIT_10 => X"000000060000000000000000000000000000004a000000000000000000000000",
            INIT_11 => X"0000000e00000000000000040000000000000012000000000000000000000000",
            INIT_12 => X"0000002e0000000000000016000000000000000c000000000000000f00000000",
            INIT_13 => X"0000000000000000000000000000000000000050000000000000003300000000",
            INIT_14 => X"0000001f000000000000002a0000000000000000000000000000003500000000",
            INIT_15 => X"00000027000000000000001c0000000000000000000000000000000500000000",
            INIT_16 => X"0000000f000000000000002f0000000000000009000000000000000000000000",
            INIT_17 => X"0000002300000000000000000000000000000000000000000000005b00000000",
            INIT_18 => X"0000001f00000000000000000000000000000025000000000000000000000000",
            INIT_19 => X"00000000000000000000001c0000000000000000000000000000004f00000000",
            INIT_1A => X"0000008100000000000000000000000000000013000000000000000a00000000",
            INIT_1B => X"00000000000000000000000a0000000000000000000000000000000100000000",
            INIT_1C => X"00000000000000000000002b0000000000000029000000000000000d00000000",
            INIT_1D => X"00000029000000000000000a0000000000000000000000000000003900000000",
            INIT_1E => X"0000000000000000000000630000000000000020000000000000000000000000",
            INIT_1F => X"0000000000000000000000090000000000000034000000000000000000000000",
            INIT_20 => X"0000006500000000000000000000000000000035000000000000001900000000",
            INIT_21 => X"0000000000000000000000190000000000000008000000000000000000000000",
            INIT_22 => X"0000000000000000000000060000000000000085000000000000001800000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000001d00000000",
            INIT_24 => X"0000006a000000000000002d000000000000001a000000000000001100000000",
            INIT_25 => X"0000002900000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000011000000000000007a00000000",
            INIT_27 => X"0000001200000000000000000000000000000007000000000000000000000000",
            INIT_28 => X"00000023000000000000002e000000000000002d000000000000001f00000000",
            INIT_29 => X"00000065000000000000003e0000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"00000014000000000000000e0000000000000000000000000000000900000000",
            INIT_2C => X"0000000000000000000000270000000000000020000000000000001b00000000",
            INIT_2D => X"0000000000000000000000720000000000000032000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000012000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000d0000000000000003000000000000001b000000000000001400000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000d00000000",
            INIT_4C => X"00000000000000000000002a0000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000030000000000000000000000000000000700000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"00000000000000000000000e0000000000000007000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000007000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000090000000000000001000000000000000000000000",
            INIT_58 => X"0000002200000000000000150000000000000007000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000012000000000000001200000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"00000001000000000000000a000000000000000c000000000000000000000000",
            INIT_5D => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_61 => X"00000000000000000000000f0000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000001000000000000000000000000",
            INIT_66 => X"0000000e00000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000005000000000000001200000000",
            INIT_68 => X"0000000300000000000000000000000000000005000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"000000410000000000000046000000000000000f000000000000000000000000",
            INIT_6B => X"000000660000000000000063000000000000004a000000000000004100000000",
            INIT_6C => X"0000000800000000000000000000000000000017000000000000003e00000000",
            INIT_6D => X"0000000300000000000000020000000000000000000000000000000600000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000001700000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000001300000000000000070000000000000000000000000000000b00000000",
            INIT_71 => X"0000000600000000000000040000000000000001000000000000000c00000000",
            INIT_72 => X"00000012000000000000002e0000000000000011000000000000003100000000",
            INIT_73 => X"0000000000000000000000020000000000000002000000000000001400000000",
            INIT_74 => X"0000000400000000000000000000000000000001000000000000001b00000000",
            INIT_75 => X"0000003d00000000000000410000000000000009000000000000000500000000",
            INIT_76 => X"0000001200000000000000310000000000000014000000000000000900000000",
            INIT_77 => X"0000000600000000000000090000000000000013000000000000001600000000",
            INIT_78 => X"0000001600000000000000000000000000000000000000000000000100000000",
            INIT_79 => X"00000013000000000000000c000000000000000b000000000000002400000000",
            INIT_7A => X"0000001b000000000000001f0000000000000008000000000000000400000000",
            INIT_7B => X"0000000000000000000000010000000000000029000000000000000200000000",
            INIT_7C => X"0000003300000000000000090000000000000001000000000000000200000000",
            INIT_7D => X"000000140000000000000000000000000000000b000000000000002100000000",
            INIT_7E => X"0000004000000000000000240000000000000013000000000000002800000000",
            INIT_7F => X"00000053000000000000003e0000000000000026000000000000002600000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE66;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67 : if BRAM_NAME = "samplegold_layersamples_instance67" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000e00000000000000370000000000000028000000000000000e00000000",
            INIT_01 => X"0000000000000000000000000000000000000016000000000000001a00000000",
            INIT_02 => X"0000002200000000000000290000000000000036000000000000000b00000000",
            INIT_03 => X"0000000a000000000000000e0000000000000029000000000000004100000000",
            INIT_04 => X"000000510000000000000000000000000000001b000000000000000800000000",
            INIT_05 => X"00000000000000000000001a0000000000000034000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"000000070000000000000018000000000000000f000000000000000000000000",
            INIT_08 => X"0000001e00000000000000080000000000000035000000000000001d00000000",
            INIT_09 => X"0000001f00000000000000300000000000000007000000000000000a00000000",
            INIT_0A => X"00000034000000000000001b0000000000000027000000000000001400000000",
            INIT_0B => X"00000022000000000000000e0000000000000000000000000000001c00000000",
            INIT_0C => X"0000001000000000000000000000000000000004000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"00000023000000000000002d000000000000001c000000000000000000000000",
            INIT_10 => X"0000002f00000000000000010000000000000000000000000000000000000000",
            INIT_11 => X"0000000a000000000000003e000000000000002a000000000000003900000000",
            INIT_12 => X"0000000000000000000000220000000000000036000000000000003600000000",
            INIT_13 => X"0000000e00000000000000000000000000000000000000000000000f00000000",
            INIT_14 => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_15 => X"0000000e00000000000000020000000000000000000000000000000000000000",
            INIT_16 => X"0000000600000000000000000000000000000000000000000000001300000000",
            INIT_17 => X"0000000e000000000000001f0000000000000009000000000000001f00000000",
            INIT_18 => X"0000000a00000000000000000000000000000000000000000000000300000000",
            INIT_19 => X"0000000b00000000000000260000000000000029000000000000001b00000000",
            INIT_1A => X"0000000900000000000000170000000000000000000000000000000000000000",
            INIT_1B => X"00000009000000000000000b000000000000001d000000000000000400000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000029000000000000001100000000",
            INIT_1E => X"000000d600000000000000cb00000000000000d5000000000000000000000000",
            INIT_1F => X"000000a900000000000000a200000000000000b000000000000000a800000000",
            INIT_20 => X"000000d700000000000000e200000000000000cf00000000000000af00000000",
            INIT_21 => X"000000b000000000000000b300000000000000c700000000000000e000000000",
            INIT_22 => X"000000a500000000000000ee00000000000000f000000000000000f200000000",
            INIT_23 => X"000000ca00000000000000b200000000000000b500000000000000a800000000",
            INIT_24 => X"000000da00000000000000d800000000000000d700000000000000e100000000",
            INIT_25 => X"000000fb00000000000000cd00000000000000c300000000000000e100000000",
            INIT_26 => X"0000008c000000000000008a00000000000000ef00000000000000fc00000000",
            INIT_27 => X"0000008c0000000000000088000000000000008d000000000000008e00000000",
            INIT_28 => X"000000ce00000000000000de00000000000000bb000000000000008d00000000",
            INIT_29 => X"000000f800000000000000fa00000000000000b700000000000000b100000000",
            INIT_2A => X"000000d200000000000000ab00000000000000ae00000000000000dd00000000",
            INIT_2B => X"000000b900000000000000be00000000000000c900000000000000c000000000",
            INIT_2C => X"000000ae00000000000000d500000000000000de000000000000009b00000000",
            INIT_2D => X"000000cb00000000000000f700000000000000f8000000000000008d00000000",
            INIT_2E => X"000000c400000000000000ad00000000000000a100000000000000a800000000",
            INIT_2F => X"000000c900000000000000c100000000000000be00000000000000b500000000",
            INIT_30 => X"000000ab00000000000000d900000000000000e100000000000000bf00000000",
            INIT_31 => X"0000007800000000000000b000000000000000ef00000000000000eb00000000",
            INIT_32 => X"0000009600000000000000930000000000000098000000000000007800000000",
            INIT_33 => X"000000ac00000000000000b1000000000000009e000000000000009800000000",
            INIT_34 => X"000000c600000000000000fb00000000000000fc00000000000000e800000000",
            INIT_35 => X"0000006a0000000000000085000000000000009700000000000000c100000000",
            INIT_36 => X"0000008400000000000000760000000000000099000000000000008a00000000",
            INIT_37 => X"000000cc000000000000008e0000000000000078000000000000009700000000",
            INIT_38 => X"0000007b00000000000000b200000000000000ff00000000000000f200000000",
            INIT_39 => X"0000006900000000000000880000000000000081000000000000008700000000",
            INIT_3A => X"000000550000000000000056000000000000005b000000000000006600000000",
            INIT_3B => X"00000092000000000000007a0000000000000052000000000000004d00000000",
            INIT_3C => X"0000006f000000000000006200000000000000aa00000000000000e900000000",
            INIT_3D => X"0000007b00000000000000750000000000000070000000000000006c00000000",
            INIT_3E => X"0000005000000000000000410000000000000038000000000000005500000000",
            INIT_3F => X"000000c100000000000000880000000000000054000000000000003000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000300000000000000072000000000000006400000000000000c200000000",
            INIT_41 => X"0000007e0000000000000053000000000000004f000000000000005200000000",
            INIT_42 => X"0000009a00000000000000a0000000000000009b000000000000009d00000000",
            INIT_43 => X"000000c90000000000000098000000000000007700000000000000ad00000000",
            INIT_44 => X"0000001d000000000000003d0000000000000039000000000000006f00000000",
            INIT_45 => X"0000006e0000000000000035000000000000004f000000000000004000000000",
            INIT_46 => X"0000005700000000000000700000000000000064000000000000006300000000",
            INIT_47 => X"0000006000000000000000cb000000000000007b000000000000007400000000",
            INIT_48 => X"00000014000000000000001d0000000000000056000000000000005d00000000",
            INIT_49 => X"000000810000000000000047000000000000004b000000000000004b00000000",
            INIT_4A => X"0000005d0000000000000050000000000000008c000000000000007a00000000",
            INIT_4B => X"0000003e000000000000007c00000000000000c2000000000000007d00000000",
            INIT_4C => X"00000008000000000000000d0000000000000047000000000000008600000000",
            INIT_4D => X"0000009c0000000000000085000000000000001c000000000000000f00000000",
            INIT_4E => X"00000069000000000000002e000000000000001d000000000000008300000000",
            INIT_4F => X"0000007d000000000000008900000000000000bd00000000000000bb00000000",
            INIT_50 => X"0000001100000000000000050000000000000025000000000000005b00000000",
            INIT_51 => X"0000009000000000000000ac0000000000000073000000000000002b00000000",
            INIT_52 => X"000000be000000000000007b000000000000002c000000000000001600000000",
            INIT_53 => X"000000500000000000000058000000000000009200000000000000ad00000000",
            INIT_54 => X"0000002b00000000000000200000000000000018000000000000003100000000",
            INIT_55 => X"0000000c00000000000000790000000000000067000000000000004600000000",
            INIT_56 => X"0000000000000000000000000000000000000083000000000000002d00000000",
            INIT_57 => X"000000000000000000000000000000000000001e000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"000000540000000000000031000000000000003d000000000000005200000000",
            INIT_5C => X"00000008000000000000001c0000000000000047000000000000006900000000",
            INIT_5D => X"0000000000000000000000110000000000000000000000000000000000000000",
            INIT_5E => X"0000003a00000000000000010000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_61 => X"000000000000000000000002000000000000001c000000000000001600000000",
            INIT_62 => X"00000000000000000000003d0000000000000005000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000019000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000029000000000000000000000000",
            INIT_65 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_66 => X"0000002300000000000000000000000000000031000000000000005d00000000",
            INIT_67 => X"0000000400000000000000030000000000000000000000000000001600000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_6A => X"0000001800000000000000000000000000000019000000000000003e00000000",
            INIT_6B => X"0000001b000000000000000c000000000000001c000000000000001a00000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000300000000",
            INIT_6D => X"00000000000000000000002c0000000000000036000000000000000a00000000",
            INIT_6E => X"000000000000000000000000000000000000000e000000000000000000000000",
            INIT_6F => X"00000024000000000000001e0000000000000004000000000000000000000000",
            INIT_70 => X"0000001300000000000000000000000000000029000000000000004700000000",
            INIT_71 => X"00000021000000000000001d0000000000000000000000000000006500000000",
            INIT_72 => X"000000380000000000000032000000000000001e000000000000000e00000000",
            INIT_73 => X"00000014000000000000003a0000000000000031000000000000002400000000",
            INIT_74 => X"0000001300000000000000000000000000000000000000000000001c00000000",
            INIT_75 => X"000000000000000000000000000000000000006e000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000001300000000000000540000000000000000000000000000000000000000",
            INIT_79 => X"000000370000000000000017000000000000001c000000000000000e00000000",
            INIT_7A => X"000000460000000000000039000000000000003a000000000000000900000000",
            INIT_7B => X"00000000000000000000003d0000000000000025000000000000003600000000",
            INIT_7C => X"000000000000000000000003000000000000001e000000000000000000000000",
            INIT_7D => X"0000004800000000000000000000000000000000000000000000002000000000",
            INIT_7E => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_7F => X"0000000f00000000000000000000000000000000000000000000004300000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE67;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68 : if BRAM_NAME = "samplegold_layersamples_instance68" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001000000000000000000000000000000000000000000000006f00000000",
            INIT_01 => X"0000001400000000000000140000000000000053000000000000001f00000000",
            INIT_02 => X"0000003700000000000000380000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000004800000000",
            INIT_04 => X"0000001000000000000000000000000000000002000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"00000000000000000000002b0000000000000000000000000000000000000000",
            INIT_07 => X"0000000900000000000000160000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000040000000000000000000000000000000900000000",
            INIT_09 => X"0000001d00000000000000430000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000008000000000000003b00000000",
            INIT_0B => X"0000002d00000000000000040000000000000000000000000000000e00000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000200000000",
            INIT_0D => X"00000003000000000000001a0000000000000005000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000f00000000",
            INIT_0F => X"0000000400000000000000000000000000000000000000000000000100000000",
            INIT_10 => X"0000000600000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_12 => X"0000000400000000000000040000000000000000000000000000000000000000",
            INIT_13 => X"0000003a00000000000000240000000000000000000000000000000000000000",
            INIT_14 => X"00000019000000000000002e000000000000002f000000000000003700000000",
            INIT_15 => X"000000000000000000000001000000000000000c000000000000000700000000",
            INIT_16 => X"00000000000000000000000b000000000000000a000000000000000a00000000",
            INIT_17 => X"000000440000000000000042000000000000004f000000000000000000000000",
            INIT_18 => X"0000003000000000000000430000000000000042000000000000003900000000",
            INIT_19 => X"0000001400000000000000000000000000000000000000000000000b00000000",
            INIT_1A => X"0000000000000000000000080000000000000006000000000000000a00000000",
            INIT_1B => X"0000004d000000000000002a0000000000000031000000000000006100000000",
            INIT_1C => X"0000002b000000000000002f0000000000000042000000000000004300000000",
            INIT_1D => X"0000000c00000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000005f0000000000000003000000000000000a000000000000000000000000",
            INIT_1F => X"0000005000000000000000540000000000000039000000000000005c00000000",
            INIT_20 => X"0000001000000000000000350000000000000033000000000000005100000000",
            INIT_21 => X"00000000000000000000001b0000000000000000000000000000000000000000",
            INIT_22 => X"0000005200000000000000610000000000000000000000000000000000000000",
            INIT_23 => X"0000005a00000000000000510000000000000052000000000000004500000000",
            INIT_24 => X"00000009000000000000003f0000000000000053000000000000005400000000",
            INIT_25 => X"0000001300000000000000000000000000000019000000000000000b00000000",
            INIT_26 => X"0000003d0000000000000045000000000000003e000000000000000200000000",
            INIT_27 => X"0000002500000000000000380000000000000048000000000000003b00000000",
            INIT_28 => X"00000015000000000000002e0000000000000042000000000000004600000000",
            INIT_29 => X"0000000000000000000000290000000000000000000000000000000000000000",
            INIT_2A => X"0000003200000000000000420000000000000039000000000000004300000000",
            INIT_2B => X"0000004700000000000000380000000000000048000000000000004300000000",
            INIT_2C => X"00000000000000000000004d000000000000005a000000000000006500000000",
            INIT_2D => X"000000420000000000000000000000000000002e000000000000000000000000",
            INIT_2E => X"0000000a00000000000000040000000000000022000000000000002c00000000",
            INIT_2F => X"0000002e00000000000000000000000000000000000000000000001100000000",
            INIT_30 => X"000000000000000000000000000000000000005b000000000000002d00000000",
            INIT_31 => X"0000002700000000000000480000000000000003000000000000002900000000",
            INIT_32 => X"0000004b0000000000000027000000000000005a000000000000004a00000000",
            INIT_33 => X"0000001f000000000000003c0000000000000040000000000000003800000000",
            INIT_34 => X"0000001700000000000000000000000000000009000000000000007c00000000",
            INIT_35 => X"0000003b000000000000003d0000000000000022000000000000001400000000",
            INIT_36 => X"00000038000000000000002c0000000000000058000000000000001600000000",
            INIT_37 => X"0000006200000000000000380000000000000020000000000000004500000000",
            INIT_38 => X"0000001400000000000000350000000000000000000000000000001500000000",
            INIT_39 => X"000000070000000000000056000000000000002e000000000000000000000000",
            INIT_3A => X"0000003000000000000000200000000000000014000000000000005d00000000",
            INIT_3B => X"0000002d00000000000000820000000000000040000000000000000000000000",
            INIT_3C => X"00000006000000000000001e0000000000000020000000000000000000000000",
            INIT_3D => X"000000330000000000000026000000000000001d000000000000000300000000",
            INIT_3E => X"0000000800000000000000000000000000000000000000000000004b00000000",
            INIT_3F => X"0000001b000000000000002d000000000000007b000000000000003300000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000250000000000000016000000000000000f00000000",
            INIT_41 => X"00000053000000000000002f0000000000000022000000000000001800000000",
            INIT_42 => X"00000046000000000000000a0000000000000000000000000000004300000000",
            INIT_43 => X"0000000c000000000000002b000000000000002f000000000000007400000000",
            INIT_44 => X"00000018000000000000000f0000000000000027000000000000001100000000",
            INIT_45 => X"000000450000000000000035000000000000002a000000000000001f00000000",
            INIT_46 => X"0000007d000000000000003e0000000000000006000000000000000800000000",
            INIT_47 => X"0000000000000000000000100000000000000020000000000000001700000000",
            INIT_48 => X"000000440000000000000025000000000000001c000000000000001500000000",
            INIT_49 => X"0000001e000000000000001b000000000000001d000000000000004200000000",
            INIT_4A => X"000000150000000000000008000000000000002d000000000000000500000000",
            INIT_4B => X"0000000000000000000000000000000000000002000000000000001700000000",
            INIT_4C => X"0000000e00000000000000000000000000000000000000000000000900000000",
            INIT_4D => X"0000001800000000000000310000000000000014000000000000001d00000000",
            INIT_4E => X"0000001300000000000000110000000000000039000000000000000100000000",
            INIT_4F => X"0000000a00000000000000130000000000000000000000000000000000000000",
            INIT_50 => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"000000000000000000000009000000000000002c000000000000004700000000",
            INIT_52 => X"00000000000000000000000a0000000000000010000000000000004300000000",
            INIT_53 => X"0000000000000000000000140000000000000055000000000000000000000000",
            INIT_54 => X"0000002200000000000000030000000000000000000000000000000000000000",
            INIT_55 => X"0000001f00000000000000040000000000000001000000000000003d00000000",
            INIT_56 => X"0000000000000000000000000000000000000002000000000000001400000000",
            INIT_57 => X"000000000000000000000000000000000000000d000000000000003100000000",
            INIT_58 => X"0000004800000000000000000000000000000000000000000000000300000000",
            INIT_59 => X"00000023000000000000001f0000000000000000000000000000002d00000000",
            INIT_5A => X"0000001500000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000004f00000000000000210000000000000000000000000000000700000000",
            INIT_5D => X"00000000000000000000001f0000000000000013000000000000001000000000",
            INIT_5E => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_5F => X"00000008000000000000000f0000000000000000000000000000000000000000",
            INIT_60 => X"00000014000000000000002e000000000000002a000000000000000000000000",
            INIT_61 => X"0000003200000000000000000000000000000002000000000000002600000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"00000060000000000000001a000000000000001e000000000000000e00000000",
            INIT_65 => X"0000000000000000000000540000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000060000000000000017000000000000002800000000",
            INIT_67 => X"000000260000000000000002000000000000003c000000000000003000000000",
            INIT_68 => X"0000000000000000000000640000000000000011000000000000005100000000",
            INIT_69 => X"0000002000000000000000000000000000000021000000000000000000000000",
            INIT_6A => X"00000000000000000000002a000000000000000c000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000077000000000000000000000000",
            INIT_6D => X"0000001100000000000000000000000000000000000000000000001900000000",
            INIT_6E => X"0000000000000000000000270000000000000000000000000000002300000000",
            INIT_6F => X"0000002600000000000000000000000000000026000000000000000000000000",
            INIT_70 => X"0000002000000000000000000000000000000000000000000000005a00000000",
            INIT_71 => X"0000002a00000000000000170000000000000000000000000000001a00000000",
            INIT_72 => X"0000001400000000000000000000000000000069000000000000000000000000",
            INIT_73 => X"0000006600000000000000120000000000000000000000000000002e00000000",
            INIT_74 => X"0000000a00000000000000270000000000000000000000000000000000000000",
            INIT_75 => X"0000001700000000000000110000000000000000000000000000000000000000",
            INIT_76 => X"00000000000000000000001d0000000000000094000000000000002000000000",
            INIT_77 => X"0000000d000000000000007a000000000000001f000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000003100000000000000210000000000000014000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000002000000000000003b00000000",
            INIT_7B => X"000000000000000000000000000000000000005b000000000000003f00000000",
            INIT_7C => X"0000000000000000000000050000000000000000000000000000000000000000",
            INIT_7D => X"0000001800000000000000160000000000000013000000000000000d00000000",
            INIT_7E => X"0000003100000000000000000000000000000000000000000000001c00000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000007900000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE68;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69 : if BRAM_NAME = "samplegold_layersamples_instance69" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000050000000000000007000000000000000600000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_11 => X"0000001a00000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_16 => X"0000000d00000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000006a000000000000007a0000000000000083000000000000002400000000",
            INIT_20 => X"0000000000000000000000000000000000000054000000000000008800000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000017000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000000000000000000000000000000000001a000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000002600000000000000200000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000060000000000000000000000000000000000000000",
            INIT_2E => X"0000000a00000000000000350000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000c000000000000000e0000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000020000000000000006000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000002c00000000000000270000000000000000000000000000000000000000",
            INIT_38 => X"0000001800000000000000170000000000000020000000000000002d00000000",
            INIT_39 => X"0000002b00000000000000340000000000000025000000000000001a00000000",
            INIT_3A => X"0000002a00000000000000260000000000000027000000000000002f00000000",
            INIT_3B => X"0000003a00000000000000310000000000000030000000000000001e00000000",
            INIT_3C => X"000000000000000000000002000000000000000f000000000000001c00000000",
            INIT_3D => X"0000001b000000000000000e0000000000000010000000000000000600000000",
            INIT_3E => X"0000001c000000000000002a000000000000002b000000000000002a00000000",
            INIT_3F => X"00000022000000000000002e0000000000000030000000000000002f00000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000002e00000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000002f00000000000000140000000000000028000000000000003600000000",
            INIT_43 => X"00000000000000000000001b000000000000001e000000000000003600000000",
            INIT_44 => X"0000000000000000000000000000000000000013000000000000000000000000",
            INIT_45 => X"00000022000000000000000f0000000000000015000000000000000000000000",
            INIT_46 => X"00000036000000000000002e0000000000000026000000000000003200000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000002200000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000002f000000000000002a000000000000000b000000000000000000000000",
            INIT_4A => X"0000000b000000000000003a0000000000000023000000000000002400000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000700000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"000000300000000000000030000000000000000d000000000000000000000000",
            INIT_4E => X"0000000000000000000000130000000000000025000000000000002900000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"00000031000000000000002a0000000000000008000000000000000c00000000",
            INIT_52 => X"00000000000000000000002f0000000000000000000000000000001200000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"00000009000000000000002c0000000000000007000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000001900000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000100000000000000060000000000000000000000000000000d00000000",
            INIT_59 => X"00000000000000000000000f0000000000000027000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"000000000000000000000000000000000000000d000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000010000000000000007000000000000002200000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000001e00000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000800000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000120000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_65 => X"000000000000000000000000000000000000000a000000000000000400000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"000000000000000000000000000000000000002a000000000000002300000000",
            INIT_68 => X"00000000000000000000000f000000000000000c000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000600000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_6C => X"0000000000000000000000060000000000000000000000000000000400000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"00000000000000000000001a0000000000000000000000000000000100000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000900000000000000000000000000000009000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000015000000000000001400000000",
            INIT_74 => X"000000000000000000000000000000000000002f000000000000000800000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000001f00000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000004a00000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"00000000000000000000001d000000000000000f000000000000000000000000",
            INIT_7B => X"0000003d00000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000010000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000190000000000000023000000000000000000000000",
            INIT_7F => X"0000000000000000000000040000000000000017000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE69;


    MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70 : if BRAM_NAME = "samplegold_layersamples_instance70" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_02 => X"0000000600000000000000000000000000000000000000000000000600000000",
            INIT_03 => X"0000000000000000000000000000000000000031000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000070000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0A => X"0000002600000000000000000000000000000020000000000000000000000000",
            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000100000000000000000000000000000000000000000000000000000000",
            INIT_0E => X"0000000000000000000000260000000000000000000000000000002a00000000",
            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_10 => X"00000000000000000000000f0000000000000019000000000000000000000000",
            INIT_11 => X"0000004900000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000000000000000000015000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"0000000a000000000000003f0000000000000000000000000000000000000000",
            INIT_16 => X"000000000000000000000000000000000000000e000000000000000300000000",
            INIT_17 => X"0000000000000000000000020000000000000000000000000000003500000000",
            INIT_18 => X"000000000000000000000000000000000000001c000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000051000000000000000000000000",
            INIT_1A => X"000000000000000000000000000000000000000b000000000000003200000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000001500000000",
            INIT_1D => X"0000000800000000000000000000000000000010000000000000000700000000",
            INIT_1E => X"000000000000000000000001000000000000000c000000000000002c00000000",
            INIT_1F => X"0000002600000000000000380000000000000005000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000002200000000000000000000000000000000000000000000000100000000",
            INIT_22 => X"0000000000000000000000000000000000000002000000000000000e00000000",
            INIT_23 => X"0000000000000000000000130000000000000028000000000000000000000000",
            INIT_24 => X"0000000300000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000c00000000000000090000000000000000000000000000001300000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000400000000",
            INIT_27 => X"0000000000000000000000000000000000000024000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_SAMPLEGOLD_LAYERSAMPLES_INSTANCE70;

MEM_EMPTY_36Kb : if BRAM_NAME(1 to 7) = "default" generate
    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
        BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
        DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
        DO_REG => 0,                     -- Optional output register (0 or 1)
        INIT => X"000000000000000000",   -- Initial values on output port
        INIT_FILE => "NONE",
        WRITE_WIDTH => 44, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH => 44, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        SRVAL => X"000000000000000000",  -- Set/Reset value for port output
        WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
    )
    port map (
        DO => bram_do,      -- Output data, width defined by READ_WIDTH parameter
        ADDR => bram_addr,  -- Input address, width defined by read/write port depth
        CLK => CLK,    -- 1-bit input clock
        DI => bram_di,      -- Input data port, width defined by WRITE_WIDTH parameter
        EN => EN,      -- 1-bit input RAM enable
        REGCE => '1', -- 1-bit input output register enable
        RST => RST,    -- 1-bit input reset
        WE => bram_wr_en       -- Input write enable, width defined by write port depth
    );
-- End of BRAM_SINGLE_MACRO_inst instantiation
end generate;


end a1;