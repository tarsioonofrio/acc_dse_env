library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 6, 12, 14, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 9, 2, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 5, 24, 16, 
    79, 28, 0, 0, 39, 68, 63, 60, 37, 27, 28, 34, 31, 33, 31, 
    38, 69, 16, 0, 41, 23, 26, 28, 27, 25, 27, 22, 32, 38, 22, 
    42, 40, 63, 34, 20, 26, 20, 26, 28, 28, 40, 48, 43, 30, 64, 
    36, 41, 50, 70, 41, 47, 42, 25, 16, 19, 30, 36, 14, 19, 36, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    9, 0, 0, 0, 16, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 0, 0, 35, 0, 23, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 42, 0, 0, 0, 0, 33, 3, 7, 0, 15, 0, 0, 0, 0, 
    0, 38, 0, 0, 0, 14, 26, 3, 2, 0, 14, 0, 0, 0, 0, 
    18, 23, 0, 7, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    35, 18, 31, 0, 0, 0, 0, 20, 0, 0, 9, 0, 0, 0, 0, 
    39, 12, 31, 0, 38, 0, 10, 43, 23, 0, 0, 0, 0, 0, 0, 
    20, 35, 13, 16, 68, 26, 11, 8, 10, 5, 10, 13, 16, 13, 16, 
    19, 4, 0, 58, 35, 11, 11, 8, 8, 7, 12, 12, 21, 22, 19, 
    28, 13, 0, 103, 19, 9, 11, 6, 10, 13, 18, 24, 22, 16, 42, 
    29, 22, 11, 32, 9, 10, 19, 15, 11, 15, 15, 11, 10, 34, 30, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 4, 0, 0, 
    17, 19, 0, 0, 0, 47, 1, 6, 0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 5, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 6, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 23, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 27, 35, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 29, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 
    67, 6, 0, 0, 64, 51, 34, 32, 4, 0, 0, 0, 0, 0, 0, 
    0, 49, 0, 4, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 41, 46, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 35, 
    0, 0, 0, 55, 13, 18, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    9, 2, 4, 6, 6, 0, 7, 8, 6, 8, 9, 5, 2, 6, 8, 
    5, 1, 2, 7, 2, 0, 10, 5, 8, 0, 0, 0, 0, 5, 9, 
    12, 6, 10, 6, 8, 0, 3, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 18, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 5, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 8, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 6, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 13, 20, 14, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 42, 26, 18, 8, 5, 0, 
    4, 19, 0, 0, 0, 2, 22, 13, 15, 39, 8, 17, 7, 2, 8, 
    16, 45, 0, 7, 49, 29, 19, 11, 11, 32, 28, 9, 20, 7, 6, 
    22, 42, 0, 0, 50, 19, 23, 14, 8, 72, 18, 2, 25, 15, 10, 
    20, 37, 0, 0, 34, 38, 40, 16, 11, 71, 12, 13, 20, 29, 9, 
    33, 42, 10, 3, 21, 68, 7, 16, 7, 39, 10, 9, 28, 20, 0, 
    41, 59, 11, 37, 12, 14, 8, 23, 25, 1, 28, 0, 14, 2, 0, 
    41, 48, 16, 54, 28, 14, 29, 41, 20, 14, 0, 17, 30, 5, 0, 
    74, 48, 17, 88, 35, 50, 72, 51, 24, 21, 42, 53, 53, 50, 41, 
    84, 64, 37, 88, 32, 26, 49, 48, 46, 53, 58, 61, 64, 61, 60, 
    59, 72, 60, 65, 14, 55, 55, 52, 51, 57, 63, 69, 66, 67, 75, 
    61, 64, 89, 42, 40, 58, 52, 56, 58, 63, 64, 66, 61, 83, 66, 
    59, 68, 59, 51, 44, 56, 55, 54, 61, 63, 59, 59, 78, 75, 50, 
    
    -- channel=5
    36, 37, 42, 43, 42, 34, 44, 48, 42, 22, 15, 21, 32, 36, 36, 
    44, 43, 44, 43, 44, 41, 39, 25, 3, 0, 0, 0, 0, 20, 33, 
    0, 22, 43, 45, 40, 0, 6, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 8, 36, 43, 26, 21, 1, 0, 0, 0, 0, 0, 0, 0, 3, 
    7, 0, 40, 42, 31, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 9, 31, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 29, 
    0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 19, 27, 
    0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 23, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 24, 23, 0, 0, 
    51, 0, 0, 0, 0, 0, 25, 13, 11, 0, 34, 0, 15, 7, 0, 
    62, 23, 5, 0, 75, 27, 29, 25, 7, 0, 24, 32, 14, 34, 0, 
    4, 15, 17, 0, 0, 0, 56, 27, 47, 0, 24, 21, 0, 23, 29, 
    18, 31, 0, 15, 0, 0, 14, 35, 38, 0, 31, 23, 2, 8, 22, 
    20, 50, 7, 28, 0, 0, 24, 0, 23, 0, 21, 17, 0, 0, 6, 
    34, 15, 38, 10, 0, 0, 3, 14, 1, 0, 0, 6, 0, 1, 0, 
    13, 4, 63, 0, 18, 0, 0, 53, 0, 0, 13, 0, 5, 0, 0, 
    0, 7, 48, 0, 129, 46, 0, 12, 43, 28, 19, 30, 11, 0, 0, 
    0, 0, 37, 0, 5, 0, 0, 0, 8, 8, 13, 11, 20, 13, 19, 
    25, 0, 0, 5, 24, 20, 18, 15, 15, 16, 20, 21, 16, 13, 30, 
    30, 17, 0, 42, 20, 14, 28, 15, 14, 17, 12, 7, 19, 14, 7, 
    36, 21, 3, 0, 1, 0, 1, 21, 23, 29, 21, 14, 22, 39, 45, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 9, 6, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 1, 4, 6, 0, 
    13, 0, 0, 0, 0, 0, 1, 7, 10, 0, 0, 7, 4, 9, 0, 
    27, 0, 0, 0, 0, 0, 0, 5, 14, 0, 9, 8, 4, 9, 6, 
    23, 10, 0, 0, 0, 0, 0, 0, 14, 0, 7, 11, 5, 3, 7, 
    15, 11, 5, 0, 0, 0, 13, 0, 0, 0, 0, 14, 5, 1, 0, 
    20, 14, 26, 0, 0, 0, 0, 3, 0, 0, 0, 7, 0, 0, 0, 
    6, 15, 24, 1, 16, 1, 0, 3, 18, 0, 3, 6, 0, 0, 0, 
    0, 8, 22, 0, 11, 30, 13, 16, 18, 15, 29, 31, 34, 18, 17, 
    50, 9, 12, 0, 34, 38, 41, 43, 48, 52, 57, 60, 63, 66, 66, 
    79, 47, 0, 19, 54, 55, 57, 55, 58, 61, 65, 70, 69, 66, 71, 
    84, 67, 39, 32, 49, 59, 59, 59, 58, 65, 72, 74, 72, 81, 81, 
    84, 75, 58, 55, 59, 60, 59, 57, 57, 64, 72, 68, 65, 88, 81, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 4, 1, 0, 
    20, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 3, 0, 10, 0, 
    5, 0, 0, 0, 0, 0, 9, 0, 22, 0, 3, 5, 0, 2, 3, 
    1, 28, 0, 0, 0, 0, 0, 0, 12, 0, 10, 8, 0, 0, 0, 
    6, 21, 0, 0, 0, 0, 3, 0, 0, 0, 3, 8, 0, 0, 0, 
    20, 8, 30, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    4, 3, 41, 0, 2, 0, 0, 12, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 33, 0, 56, 15, 0, 11, 28, 19, 23, 30, 32, 19, 23, 
    13, 7, 5, 0, 41, 44, 33, 33, 47, 43, 50, 51, 58, 57, 60, 
    76, 14, 0, 19, 50, 50, 49, 48, 50, 53, 58, 60, 59, 58, 65, 
    82, 64, 0, 59, 46, 47, 56, 49, 49, 55, 62, 63, 69, 68, 73, 
    81, 70, 58, 38, 47, 44, 46, 48, 50, 59, 62, 57, 53, 80, 84, 
    
    -- channel=9
    34, 40, 35, 38, 38, 34, 38, 42, 40, 34, 29, 26, 29, 36, 38, 
    33, 39, 36, 41, 31, 32, 47, 41, 35, 10, 15, 22, 18, 17, 33, 
    46, 7, 36, 41, 34, 46, 47, 30, 4, 0, 21, 15, 26, 3, 18, 
    62, 0, 34, 35, 48, 12, 27, 15, 7, 0, 42, 14, 25, 15, 0, 
    34, 0, 45, 0, 27, 17, 49, 34, 26, 0, 23, 35, 12, 25, 0, 
    19, 6, 49, 29, 3, 20, 48, 33, 47, 0, 46, 41, 3, 17, 12, 
    13, 40, 19, 67, 0, 0, 34, 29, 49, 0, 47, 30, 4, 0, 19, 
    12, 37, 10, 37, 0, 0, 61, 24, 30, 0, 33, 39, 0, 9, 24, 
    26, 8, 43, 0, 19, 12, 28, 23, 0, 39, 13, 46, 0, 6, 20, 
    18, 6, 59, 0, 32, 7, 0, 28, 15, 23, 38, 4, 0, 6, 34, 
    0, 9, 58, 0, 40, 6, 0, 22, 31, 20, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 74, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 24, 0, 0, 0, 19, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 32, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 1, 
    0, 9, 0, 0, 67, 0, 0, 0, 0, 68, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 46, 0, 0, 0, 0, 76, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 50, 0, 0, 0, 47, 0, 0, 0, 0, 0, 
    0, 2, 0, 7, 0, 26, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 22, 0, 0, 1, 0, 0, 0, 0, 0, 5, 0, 0, 
    38, 0, 0, 52, 0, 0, 31, 15, 0, 0, 0, 0, 0, 1, 0, 
    90, 44, 0, 57, 0, 0, 6, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 68, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    0, 0, 107, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 12, 
    0, 0, 3, 19, 0, 9, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 14, 0, 7, 0, 5, 0, 
    0, 50, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 20, 9, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 11, 14, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 0, 0, 4, 7, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 15, 13, 7, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 19, 13, 0, 
    0, 0, 0, 13, 0, 8, 13, 0, 0, 0, 0, 23, 43, 0, 0, 
    0, 0, 0, 44, 0, 0, 0, 0, 0, 11, 49, 56, 38, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 22, 31, 38, 38, 44, 39, 35, 
    47, 10, 23, 0, 0, 38, 34, 39, 41, 48, 53, 50, 32, 34, 56, 
    42, 52, 23, 0, 9, 41, 40, 39, 42, 43, 40, 33, 42, 56, 6, 
    35, 51, 41, 0, 24, 34, 28, 41, 46, 45, 36, 52, 65, 24, 39, 
    
    -- channel=12
    18, 14, 21, 20, 21, 16, 19, 20, 22, 15, 10, 13, 16, 15, 17, 
    23, 16, 19, 18, 21, 32, 18, 17, 0, 16, 12, 10, 10, 15, 19, 
    10, 12, 23, 19, 23, 0, 8, 0, 18, 9, 0, 0, 0, 8, 13, 
    0, 36, 18, 22, 23, 20, 9, 9, 5, 0, 0, 0, 0, 6, 6, 
    0, 8, 14, 26, 12, 13, 0, 6, 0, 24, 0, 1, 5, 0, 13, 
    2, 0, 15, 27, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 10, 
    12, 0, 6, 7, 0, 29, 0, 6, 0, 11, 0, 3, 6, 9, 4, 
    15, 0, 9, 7, 7, 0, 0, 0, 0, 4, 0, 0, 1, 0, 5, 
    0, 0, 8, 2, 30, 0, 0, 7, 7, 0, 0, 0, 3, 5, 18, 
    0, 0, 0, 0, 0, 19, 13, 0, 10, 0, 0, 0, 6, 18, 14, 
    0, 0, 0, 33, 9, 13, 7, 0, 0, 0, 11, 15, 6, 3, 8, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    
    -- channel=13
    40, 38, 38, 40, 41, 35, 43, 46, 40, 31, 22, 23, 27, 37, 39, 
    41, 41, 41, 42, 38, 18, 41, 29, 21, 6, 7, 15, 17, 26, 35, 
    22, 20, 42, 43, 44, 27, 21, 19, 9, 0, 1, 0, 12, 21, 24, 
    21, 14, 46, 38, 32, 12, 11, 5, 3, 0, 0, 7, 5, 17, 18, 
    0, 3, 42, 11, 0, 0, 2, 3, 6, 0, 5, 11, 2, 10, 17, 
    0, 0, 35, 23, 0, 0, 0, 9, 13, 0, 0, 3, 1, 1, 10, 
    0, 0, 25, 34, 0, 0, 0, 0, 11, 0, 0, 6, 2, 0, 12, 
    0, 0, 10, 22, 9, 0, 0, 0, 7, 0, 0, 11, 0, 3, 21, 
    0, 0, 0, 0, 8, 0, 13, 5, 0, 21, 13, 2, 5, 19, 35, 
    0, 0, 0, 0, 8, 0, 0, 0, 6, 0, 0, 3, 2, 18, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 22, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 12, 27, 0, 0, 0, 22, 16, 0, 
    36, 41, 0, 0, 0, 35, 15, 10, 0, 0, 0, 0, 0, 24, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 4, 0, 4, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 15, 
    0, 5, 0, 0, 63, 4, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 33, 0, 9, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 22, 24, 1, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 31, 34, 14, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 43, 31, 5, 0, 0, 1, 
    10, 0, 0, 0, 0, 0, 0, 36, 14, 0, 0, 0, 0, 22, 16, 
    67, 29, 0, 0, 46, 54, 31, 29, 13, 0, 0, 0, 0, 0, 0, 
    0, 48, 2, 11, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 46, 59, 1, 0, 0, 0, 0, 0, 0, 6, 0, 0, 28, 
    0, 0, 3, 45, 9, 17, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 6, 20, 0, 0, 0, 13, 0, 0, 4, 6, 0, 
    0, 25, 0, 0, 4, 10, 0, 0, 6, 49, 0, 0, 0, 6, 16, 
    0, 68, 0, 4, 0, 16, 0, 0, 0, 58, 0, 0, 0, 0, 51, 
    0, 26, 0, 53, 0, 0, 0, 0, 0, 86, 0, 0, 1, 0, 17, 
    0, 11, 0, 0, 68, 0, 0, 0, 0, 148, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 62, 46, 0, 0, 0, 118, 0, 0, 6, 14, 0, 
    0, 0, 0, 0, 32, 48, 0, 0, 0, 79, 0, 0, 20, 0, 0, 
    0, 0, 0, 26, 0, 7, 0, 0, 22, 0, 11, 0, 25, 29, 9, 
    0, 1, 0, 56, 0, 0, 35, 0, 0, 0, 0, 0, 28, 23, 0, 
    54, 0, 0, 138, 0, 0, 21, 0, 0, 0, 1, 4, 2, 0, 0, 
    46, 27, 0, 84, 0, 0, 2, 1, 0, 0, 0, 3, 4, 1, 0, 
    0, 45, 72, 0, 0, 0, 0, 0, 0, 2, 6, 4, 0, 0, 13, 
    0, 0, 93, 0, 0, 4, 0, 0, 2, 2, 0, 0, 0, 22, 0, 
    0, 0, 2, 0, 0, 12, 1, 0, 6, 0, 0, 6, 38, 0, 0, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 6, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 0, 0, 0, 0, 0, 
    7, 27, 0, 0, 27, 20, 0, 0, 0, 6, 0, 0, 5, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 6, 14, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 9, 3, 
    6, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 1, 0, 14, 1, 0, 0, 0, 17, 0, 0, 
    1, 0, 0, 49, 45, 55, 48, 0, 5, 6, 34, 61, 44, 9, 4, 
    15, 2, 9, 35, 0, 0, 0, 0, 20, 41, 50, 50, 55, 52, 51, 
    63, 20, 12, 0, 0, 46, 47, 43, 45, 54, 61, 66, 57, 56, 70, 
    60, 57, 34, 0, 27, 49, 48, 47, 51, 57, 57, 51, 53, 77, 49, 
    62, 62, 45, 0, 30, 38, 40, 49, 61, 59, 55, 55, 79, 73, 54, 
    
    -- channel=17
    26, 35, 27, 33, 31, 28, 31, 35, 36, 32, 23, 15, 18, 24, 29, 
    26, 32, 28, 37, 25, 36, 37, 39, 28, 0, 5, 6, 0, 6, 26, 
    50, 0, 31, 35, 31, 49, 38, 7, 0, 0, 18, 0, 17, 0, 8, 
    57, 0, 30, 28, 50, 0, 28, 3, 0, 0, 36, 7, 13, 2, 0, 
    24, 0, 36, 0, 37, 2, 40, 21, 16, 0, 16, 25, 0, 12, 0, 
    3, 11, 37, 30, 8, 0, 50, 19, 41, 0, 45, 24, 0, 3, 0, 
    0, 57, 4, 65, 0, 0, 50, 20, 43, 0, 42, 18, 0, 0, 8, 
    0, 35, 0, 34, 0, 7, 52, 17, 20, 0, 33, 28, 0, 4, 4, 
    23, 9, 34, 0, 14, 0, 16, 25, 0, 30, 18, 27, 0, 0, 16, 
    24, 9, 60, 0, 31, 0, 0, 37, 2, 21, 24, 0, 0, 1, 28, 
    0, 10, 55, 0, 51, 8, 0, 28, 22, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 105, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 78, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 91, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 39, 8, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 3, 0, 12, 0, 0, 0, 7, 0, 0, 0, 0, 
    41, 12, 9, 0, 74, 30, 9, 0, 0, 0, 11, 10, 0, 1, 0, 
    0, 0, 18, 0, 0, 0, 36, 5, 10, 0, 6, 0, 0, 0, 5, 
    16, 0, 0, 2, 0, 1, 0, 17, 2, 0, 10, 0, 0, 0, 0, 
    21, 17, 13, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 117, 38, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 9, 0, 0, 0, 13, 0, 0, 0, 0, 
    21, 16, 0, 0, 50, 35, 26, 3, 0, 0, 17, 6, 0, 0, 0, 
    25, 26, 4, 7, 16, 25, 40, 4, 0, 0, 36, 0, 0, 0, 0, 
    27, 41, 0, 0, 0, 22, 36, 19, 2, 1, 26, 1, 0, 0, 0, 
    44, 37, 4, 0, 0, 30, 30, 3, 0, 0, 21, 0, 0, 0, 0, 
    56, 42, 30, 4, 10, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    42, 40, 35, 5, 16, 0, 0, 31, 5, 0, 0, 0, 0, 0, 0, 
    24, 39, 30, 20, 78, 33, 30, 30, 13, 0, 0, 0, 0, 0, 0, 
    0, 21, 28, 57, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 75, 13, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 4, 23, 0, 
    
    -- channel=20
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 1, 0, 2, 25, 0, 0, 0, 5, 0, 0, 7, 2, 0, 
    0, 10, 0, 0, 1, 30, 0, 0, 0, 41, 0, 0, 0, 8, 11, 
    0, 61, 0, 6, 0, 6, 0, 0, 0, 48, 0, 0, 0, 0, 41, 
    0, 48, 0, 36, 10, 0, 0, 0, 0, 46, 0, 0, 1, 0, 18, 
    0, 14, 0, 0, 48, 0, 0, 0, 0, 118, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 64, 22, 0, 0, 0, 109, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 30, 60, 0, 0, 0, 72, 0, 0, 13, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 14, 0, 14, 0, 8, 11, 8, 
    0, 0, 0, 45, 0, 0, 10, 0, 0, 0, 0, 0, 29, 31, 0, 
    48, 0, 0, 105, 0, 0, 31, 0, 0, 0, 4, 7, 13, 13, 0, 
    56, 7, 0, 90, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 45, 23, 1, 0, 0, 0, 0, 0, 0, 3, 5, 0, 0, 5, 
    0, 0, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    0, 0, 0, 2, 0, 4, 0, 0, 0, 0, 0, 0, 23, 0, 0, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 
    0, 0, 0, 0, 0, 4, 22, 0, 0, 0, 29, 22, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 17, 13, 3, 0, 9, 7, 34, 0, 0, 
    80, 0, 5, 0, 10, 0, 21, 15, 7, 0, 28, 0, 18, 21, 0, 
    60, 0, 29, 0, 22, 16, 27, 27, 13, 0, 16, 43, 5, 37, 0, 
    20, 0, 33, 0, 0, 0, 33, 28, 58, 0, 25, 32, 0, 18, 33, 
    24, 18, 0, 34, 0, 0, 0, 25, 44, 0, 38, 34, 2, 0, 23, 
    15, 18, 27, 36, 0, 0, 19, 0, 18, 0, 12, 33, 0, 0, 2, 
    17, 0, 61, 0, 19, 0, 11, 13, 0, 30, 0, 17, 0, 0, 0, 
    0, 0, 65, 0, 22, 0, 0, 31, 7, 0, 18, 3, 0, 0, 2, 
    0, 0, 56, 0, 92, 39, 0, 0, 30, 37, 19, 12, 0, 0, 16, 
    0, 0, 9, 0, 28, 9, 0, 0, 4, 0, 0, 0, 0, 0, 3, 
    19, 0, 0, 0, 43, 1, 4, 1, 4, 1, 0, 0, 0, 0, 0, 
    17, 3, 0, 14, 12, 0, 16, 3, 0, 0, 0, 0, 3, 0, 0, 
    23, 0, 0, 0, 5, 0, 0, 0, 0, 7, 11, 0, 0, 18, 39, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 2, 23, 13, 0, 0, 0, 0, 12, 2, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 4, 13, 15, 0, 
    7, 0, 10, 0, 0, 0, 5, 3, 14, 0, 0, 8, 0, 5, 2, 
    24, 0, 16, 3, 0, 12, 0, 0, 6, 0, 17, 34, 0, 0, 0, 
    9, 0, 13, 8, 0, 0, 0, 0, 17, 0, 27, 3, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 50, 18, 7, 0, 9, 15, 0, 0, 5, 
    0, 0, 33, 0, 0, 26, 3, 0, 0, 8, 0, 55, 0, 0, 0, 
    0, 0, 26, 0, 7, 4, 0, 0, 0, 20, 52, 8, 0, 0, 0, 
    0, 0, 31, 0, 0, 0, 0, 14, 35, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 76, 57, 13, 12, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    2, 0, 0, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    
    -- channel=23
    23, 17, 21, 16, 19, 19, 20, 23, 17, 15, 22, 26, 20, 18, 17, 
    18, 19, 24, 15, 22, 0, 3, 12, 26, 10, 0, 0, 26, 27, 14, 
    4, 51, 22, 18, 24, 27, 0, 19, 15, 6, 0, 0, 0, 32, 20, 
    0, 33, 12, 22, 0, 24, 0, 0, 0, 37, 0, 0, 0, 0, 51, 
    0, 0, 0, 53, 0, 0, 0, 0, 0, 54, 0, 0, 0, 0, 45, 
    0, 0, 0, 31, 9, 0, 0, 0, 0, 50, 0, 0, 1, 0, 0, 
    0, 0, 11, 0, 35, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 0, 0, 0, 0, 23, 0, 0, 7, 0, 2, 
    0, 0, 0, 0, 0, 27, 0, 0, 5, 0, 0, 0, 24, 8, 6, 
    0, 0, 0, 5, 0, 22, 14, 0, 0, 0, 0, 13, 12, 14, 9, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 4, 2, 1, 0, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 4, 3, 1, 17, 1, 2, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 1, 3, 28, 0, 0, 0, 6, 14, 0, 0, 0, 0, 
    0, 0, 0, 2, 5, 0, 5, 0, 0, 16, 13, 5, 0, 0, 0, 
    0, 23, 0, 2, 33, 28, 25, 0, 0, 0, 17, 0, 0, 0, 0, 
    20, 41, 6, 21, 61, 35, 33, 2, 0, 22, 34, 0, 0, 0, 0, 
    15, 47, 0, 0, 24, 33, 50, 15, 0, 38, 21, 0, 0, 0, 0, 
    34, 38, 0, 0, 4, 61, 32, 19, 0, 37, 23, 0, 0, 9, 0, 
    47, 50, 12, 18, 7, 17, 6, 7, 0, 4, 17, 0, 0, 0, 1, 
    54, 53, 19, 21, 14, 0, 5, 25, 12, 11, 0, 0, 0, 7, 2, 
    47, 49, 21, 46, 36, 12, 42, 44, 5, 0, 0, 0, 0, 0, 0, 
    30, 39, 26, 86, 73, 5, 5, 1, 0, 0, 0, 0, 0, 4, 1, 
    0, 23, 32, 90, 5, 0, 0, 0, 0, 0, 0, 0, 6, 2, 2, 
    0, 0, 38, 51, 0, 0, 0, 0, 0, 0, 1, 3, 0, 5, 16, 
    2, 0, 2, 5, 0, 0, 0, 0, 0, 1, 0, 0, 7, 19, 0, 
    
    -- channel=25
    0, 3, 6, 7, 7, 5, 2, 2, 7, 0, 0, 0, 7, 4, 6, 
    8, 8, 7, 6, 10, 59, 8, 3, 0, 16, 29, 4, 0, 0, 10, 
    0, 0, 5, 5, 0, 0, 0, 0, 7, 31, 5, 18, 13, 0, 8, 
    26, 28, 2, 10, 13, 20, 35, 13, 9, 0, 8, 0, 0, 0, 0, 
    36, 49, 4, 27, 103, 44, 5, 6, 0, 9, 22, 13, 17, 22, 0, 
    0, 7, 0, 0, 0, 0, 30, 16, 23, 37, 0, 0, 3, 18, 22, 
    0, 2, 0, 11, 0, 21, 5, 19, 10, 22, 0, 2, 3, 17, 9, 
    0, 26, 3, 29, 13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 7, 0, 17, 0, 0, 0, 14, 16, 0, 0, 0, 0, 5, 14, 
    0, 0, 7, 16, 0, 0, 19, 51, 0, 0, 0, 0, 24, 21, 3, 
    10, 0, 0, 50, 103, 54, 26, 0, 7, 21, 27, 46, 22, 8, 7, 
    0, 0, 20, 41, 0, 0, 0, 0, 0, 3, 7, 3, 9, 2, 2, 
    3, 0, 0, 0, 0, 6, 2, 2, 4, 9, 15, 16, 3, 3, 26, 
    1, 2, 0, 0, 0, 6, 10, 1, 5, 7, 0, 0, 1, 14, 0, 
    2, 2, 0, 0, 0, 0, 0, 7, 19, 19, 1, 3, 34, 21, 4, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 40, 0, 0, 42, 14, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 13, 0, 0, 0, 0, 4, 0, 0, 17, 0, 0, 0, 0, 0, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    3, 30, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 3, 23, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 
    17, 13, 0, 57, 70, 49, 19, 0, 0, 0, 15, 28, 23, 4, 0, 
    16, 6, 22, 57, 0, 0, 0, 0, 8, 18, 28, 32, 42, 42, 36, 
    47, 12, 10, 19, 0, 29, 28, 25, 26, 34, 45, 52, 42, 37, 64, 
    48, 42, 14, 0, 3, 35, 35, 31, 29, 38, 38, 37, 39, 60, 31, 
    48, 47, 27, 10, 8, 14, 15, 28, 41, 50, 41, 40, 69, 75, 46, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 16, 10, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 6, 7, 0, 12, 3, 10, 3, 0, 
    32, 0, 0, 0, 0, 3, 11, 8, 8, 0, 10, 11, 4, 9, 0, 
    39, 14, 0, 0, 0, 5, 6, 12, 12, 0, 21, 18, 6, 13, 7, 
    40, 21, 0, 0, 0, 0, 10, 14, 16, 0, 27, 15, 9, 7, 9, 
    31, 32, 17, 0, 0, 0, 29, 10, 9, 0, 14, 17, 6, 4, 0, 
    37, 29, 34, 1, 0, 9, 7, 2, 5, 1, 0, 14, 1, 0, 0, 
    25, 30, 36, 15, 17, 6, 7, 13, 14, 0, 13, 7, 0, 0, 0, 
    13, 26, 37, 5, 40, 24, 13, 30, 31, 23, 23, 24, 33, 25, 23, 
    44, 33, 35, 8, 50, 52, 43, 44, 45, 44, 49, 53, 56, 59, 60, 
    71, 42, 27, 26, 65, 49, 50, 49, 51, 53, 59, 60, 61, 63, 67, 
    77, 61, 32, 49, 48, 53, 55, 50, 51, 56, 63, 65, 68, 65, 71, 
    76, 66, 54, 55, 52, 49, 52, 53, 51, 58, 62, 62, 60, 76, 77, 
    
    -- channel=28
    10, 4, 9, 11, 13, 4, 8, 10, 13, 9, 6, 3, 6, 13, 16, 
    14, 3, 7, 10, 8, 5, 19, 4, 2, 6, 20, 18, 8, 4, 13, 
    8, 0, 9, 10, 10, 0, 19, 15, 16, 0, 18, 23, 31, 12, 1, 
    36, 8, 10, 7, 13, 5, 12, 27, 24, 0, 25, 13, 25, 32, 0, 
    36, 2, 26, 0, 0, 17, 14, 28, 23, 0, 12, 33, 19, 33, 19, 
    34, 0, 27, 14, 0, 1, 14, 23, 37, 0, 24, 31, 10, 26, 33, 
    38, 8, 7, 17, 0, 0, 0, 23, 26, 0, 25, 31, 21, 14, 30, 
    28, 6, 36, 12, 0, 0, 26, 9, 19, 0, 20, 29, 8, 8, 24, 
    21, 0, 48, 0, 27, 0, 15, 17, 8, 22, 0, 28, 10, 10, 14, 
    1, 2, 36, 0, 14, 25, 6, 9, 27, 4, 25, 18, 6, 6, 15, 
    0, 2, 30, 0, 46, 28, 0, 0, 27, 33, 25, 25, 22, 9, 17, 
    0, 0, 13, 0, 14, 24, 10, 12, 23, 23, 25, 23, 25, 28, 29, 
    42, 0, 0, 0, 41, 25, 25, 27, 30, 30, 28, 28, 25, 23, 26, 
    39, 28, 0, 4, 32, 25, 33, 26, 24, 25, 28, 24, 32, 24, 25, 
    41, 27, 27, 4, 31, 20, 20, 27, 25, 30, 32, 30, 21, 34, 45, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 10, 10, 7, 7, 0, 0, 0, 3, 14, 9, 1, 0, 
    6, 0, 0, 26, 0, 0, 0, 0, 0, 7, 14, 14, 17, 18, 13, 
    22, 3, 0, 6, 0, 9, 10, 10, 11, 16, 20, 22, 18, 13, 23, 
    18, 18, 0, 0, 0, 12, 12, 12, 11, 16, 18, 15, 15, 26, 20, 
    19, 20, 13, 0, 4, 6, 5, 9, 17, 21, 17, 15, 28, 34, 16, 
    
    -- channel=30
    47, 43, 48, 47, 49, 40, 49, 57, 52, 36, 30, 33, 37, 41, 45, 
    49, 46, 48, 47, 48, 15, 40, 33, 33, 12, 0, 1, 16, 31, 38, 
    17, 42, 51, 52, 52, 24, 35, 24, 8, 0, 0, 0, 0, 11, 25, 
    0, 4, 41, 50, 34, 32, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 36, 37, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 12, 
    0, 0, 35, 45, 0, 9, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 22, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 8, 9, 2, 0, 0, 14, 0, 11, 3, 8, 21, 
    0, 0, 0, 0, 0, 12, 3, 0, 0, 0, 4, 0, 0, 8, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 76, 0, 0, 0, 13, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 0, 37, 0, 0, 0, 0, 19, 
    18, 24, 0, 0, 13, 0, 38, 0, 0, 0, 2, 0, 0, 0, 2, 
    0, 55, 0, 0, 74, 0, 0, 0, 7, 0, 10, 0, 17, 8, 0, 
    0, 36, 0, 0, 62, 0, 49, 0, 37, 39, 0, 0, 1, 0, 0, 
    0, 69, 0, 23, 43, 14, 31, 0, 11, 62, 0, 0, 0, 14, 0, 
    0, 43, 0, 27, 0, 42, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    0, 9, 0, 39, 0, 0, 0, 42, 0, 4, 20, 0, 0, 14, 0, 
    5, 0, 0, 27, 0, 0, 0, 73, 0, 0, 0, 0, 19, 20, 0, 
    82, 0, 0, 41, 30, 0, 0, 0, 0, 0, 8, 12, 0, 1, 0, 
    0, 0, 0, 71, 0, 0, 0, 0, 0, 0, 3, 2, 9, 2, 0, 
    0, 0, 0, 67, 0, 0, 0, 0, 0, 4, 6, 7, 0, 0, 8, 
    0, 0, 0, 78, 0, 0, 0, 0, 0, 1, 0, 1, 0, 14, 0, 
    0, 8, 0, 25, 0, 0, 0, 0, 6, 13, 0, 0, 16, 22, 0, 
    
    -- channel=33
    4, 8, 4, 6, 3, 2, 9, 7, 0, 0, 0, 0, 0, 0, 0, 
    1, 5, 7, 8, 4, 22, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 6, 5, 38, 0, 0, 0, 7, 20, 4, 0, 0, 2, 
    4, 0, 10, 2, 2, 0, 13, 0, 0, 11, 20, 1, 0, 0, 0, 
    13, 42, 12, 0, 53, 11, 28, 0, 0, 0, 25, 0, 0, 0, 0, 
    0, 57, 15, 0, 59, 16, 46, 12, 4, 0, 35, 0, 2, 0, 0, 
    0, 70, 6, 5, 26, 14, 72, 14, 19, 31, 29, 0, 0, 0, 1, 
    4, 61, 0, 12, 0, 68, 36, 21, 7, 34, 26, 3, 0, 13, 3, 
    33, 56, 0, 29, 0, 11, 10, 9, 2, 9, 16, 0, 0, 7, 10, 
    52, 53, 34, 17, 25, 0, 0, 48, 0, 11, 0, 0, 0, 13, 4, 
    56, 42, 37, 27, 56, 14, 32, 54, 13, 0, 0, 0, 0, 0, 0, 
    39, 40, 37, 85, 85, 0, 0, 0, 0, 0, 0, 0, 2, 7, 2, 
    4, 18, 7, 103, 5, 0, 0, 0, 0, 0, 0, 3, 12, 4, 8, 
    7, 0, 8, 95, 0, 0, 0, 0, 0, 0, 2, 10, 1, 4, 28, 
    10, 3, 0, 35, 0, 0, 4, 0, 2, 6, 6, 0, 8, 33, 8, 
    
    -- channel=34
    0, 0, 0, 1, 2, 4, 0, 0, 5, 0, 0, 0, 0, 0, 2, 
    7, 5, 0, 0, 5, 45, 0, 0, 0, 27, 28, 9, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 12, 18, 18, 0, 6, 0, 0, 0, 
    15, 32, 0, 8, 3, 27, 20, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 21, 0, 30, 44, 1, 0, 0, 0, 32, 25, 1, 9, 8, 0, 
    0, 0, 0, 0, 0, 0, 19, 14, 7, 31, 0, 0, 0, 5, 16, 
    10, 0, 0, 0, 0, 25, 0, 1, 0, 2, 0, 8, 10, 21, 0, 
    4, 16, 5, 18, 6, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 15, 15, 17, 0, 0, 0, 0, 14, 2, 
    0, 0, 0, 27, 0, 0, 27, 30, 0, 0, 0, 4, 10, 0, 0, 
    7, 0, 0, 56, 55, 20, 0, 0, 0, 8, 34, 24, 2, 0, 4, 
    0, 0, 9, 1, 0, 0, 0, 0, 1, 0, 0, 0, 7, 2, 2, 
    0, 0, 15, 0, 0, 2, 0, 0, 3, 7, 11, 8, 0, 0, 20, 
    0, 0, 0, 0, 0, 1, 7, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 0, 6, 31, 0, 0, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 3, 0, 0, 
    16, 3, 0, 0, 0, 18, 4, 0, 0, 0, 12, 0, 3, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 9, 21, 3, 17, 8, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 15, 0, 0, 0, 0, 0, 13, 
    23, 15, 0, 25, 36, 9, 0, 0, 0, 1, 16, 9, 8, 0, 0, 
    6, 21, 6, 0, 13, 0, 15, 0, 1, 12, 9, 4, 5, 1, 5, 
    11, 0, 1, 0, 2, 26, 24, 23, 7, 19, 13, 9, 11, 19, 0, 
    12, 11, 19, 2, 11, 22, 4, 4, 0, 0, 32, 20, 15, 0, 0, 
    21, 20, 8, 0, 13, 11, 0, 0, 20, 30, 17, 3, 0, 0, 0, 
    18, 14, 10, 0, 0, 0, 26, 29, 15, 0, 0, 0, 15, 18, 18, 
    62, 28, 0, 13, 64, 46, 37, 34, 30, 26, 28, 28, 26, 31, 31, 
    39, 56, 15, 44, 36, 23, 25, 24, 25, 26, 24, 26, 36, 34, 21, 
    38, 31, 59, 45, 31, 24, 21, 26, 26, 28, 36, 42, 33, 36, 62, 
    37, 34, 40, 39, 38, 43, 41, 26, 21, 20, 32, 29, 17, 31, 31, 
    
    -- channel=36
    28, 32, 31, 29, 29, 30, 33, 34, 29, 24, 19, 26, 26, 24, 25, 
    32, 35, 34, 30, 33, 46, 8, 25, 14, 21, 3, 6, 19, 31, 28, 
    15, 43, 33, 32, 35, 46, 0, 1, 5, 35, 0, 0, 0, 16, 40, 
    0, 54, 31, 35, 24, 22, 13, 0, 0, 36, 0, 0, 0, 0, 52, 
    0, 38, 0, 32, 21, 0, 0, 0, 0, 31, 0, 0, 8, 0, 14, 
    0, 14, 0, 3, 51, 0, 0, 0, 0, 78, 0, 0, 12, 0, 0, 
    0, 2, 3, 10, 59, 19, 5, 0, 0, 77, 0, 0, 3, 10, 0, 
    0, 0, 0, 15, 26, 46, 0, 0, 0, 54, 0, 0, 12, 7, 0, 
    0, 0, 0, 28, 0, 0, 0, 9, 13, 6, 23, 0, 14, 27, 29, 
    0, 0, 0, 29, 0, 0, 4, 9, 0, 0, 0, 2, 32, 42, 15, 
    43, 0, 0, 55, 0, 0, 9, 0, 0, 0, 0, 0, 0, 5, 0, 
    20, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 34, 10, 0, 0, 0, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 7, 0, 9, 0, 0, 
    14, 25, 0, 0, 0, 0, 29, 14, 0, 0, 0, 0, 0, 0, 0, 
    13, 61, 3, 13, 83, 68, 0, 0, 0, 0, 16, 16, 4, 9, 0, 
    0, 0, 0, 0, 0, 0, 4, 9, 12, 45, 0, 0, 0, 3, 20, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 21, 0, 0, 0, 8, 11, 
    0, 0, 17, 1, 22, 12, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 4, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 0, 2, 0, 0, 0, 41, 7, 0, 0, 0, 18, 22, 0, 
    0, 0, 0, 48, 87, 89, 34, 0, 0, 0, 19, 45, 18, 0, 0, 
    0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 14, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 12, 2, 0, 30, 26, 0, 
    
    -- channel=38
    32, 30, 28, 27, 28, 27, 31, 35, 26, 22, 21, 24, 18, 23, 23, 
    27, 29, 30, 28, 27, 0, 9, 21, 18, 0, 0, 0, 23, 23, 21, 
    23, 39, 31, 30, 37, 62, 0, 9, 0, 0, 0, 0, 0, 27, 23, 
    0, 27, 27, 28, 13, 5, 0, 0, 0, 32, 0, 4, 0, 0, 41, 
    0, 0, 3, 13, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 34, 
    0, 0, 0, 45, 40, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 43, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 11, 0, 3, 0, 44, 0, 0, 3, 10, 5, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 11, 25, 0, 21, 11, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 0, 0, 18, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=39
    5, 4, 6, 0, 0, 5, 5, 4, 0, 0, 7, 15, 7, 0, 0, 
    4, 5, 7, 0, 6, 0, 0, 1, 2, 6, 0, 0, 16, 18, 0, 
    0, 43, 5, 1, 6, 22, 0, 0, 2, 25, 0, 0, 0, 17, 21, 
    0, 44, 0, 8, 0, 8, 0, 0, 0, 50, 0, 0, 0, 0, 54, 
    0, 4, 0, 36, 0, 0, 0, 0, 0, 58, 0, 0, 0, 0, 26, 
    0, 1, 0, 3, 63, 0, 0, 0, 0, 98, 0, 0, 6, 0, 0, 
    0, 0, 4, 0, 55, 20, 0, 0, 0, 82, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 36, 0, 0, 0, 52, 0, 0, 13, 2, 0, 
    0, 0, 0, 17, 0, 17, 0, 0, 12, 0, 13, 0, 19, 13, 2, 
    0, 0, 0, 27, 0, 1, 17, 0, 0, 1, 0, 1, 27, 23, 0, 
    33, 0, 0, 69, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 21, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 41, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    6, 6, 0, 2, 4, 0, 5, 9, 8, 16, 21, 12, 3, 4, 8, 
    0, 0, 0, 6, 0, 0, 9, 14, 47, 0, 0, 0, 7, 5, 3, 
    32, 14, 3, 6, 3, 44, 48, 32, 0, 0, 0, 0, 6, 1, 0, 
    28, 0, 5, 0, 11, 0, 0, 0, 0, 0, 18, 6, 20, 5, 0, 
    8, 0, 16, 0, 0, 0, 14, 3, 16, 0, 0, 4, 0, 0, 0, 
    16, 0, 19, 18, 9, 12, 0, 0, 11, 0, 22, 37, 0, 0, 0, 
    0, 14, 21, 37, 0, 0, 10, 0, 25, 0, 40, 6, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 54, 27, 16, 0, 22, 25, 0, 0, 2, 
    0, 0, 27, 0, 0, 39, 21, 0, 0, 28, 11, 61, 0, 0, 0, 
    0, 0, 36, 0, 9, 0, 0, 0, 0, 27, 55, 5, 0, 0, 15, 
    0, 0, 48, 0, 0, 0, 0, 23, 28, 11, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 117, 78, 28, 27, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 88, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 43, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=41
    39, 39, 41, 40, 42, 39, 42, 49, 46, 37, 31, 33, 34, 32, 34, 
    44, 43, 43, 42, 44, 28, 32, 37, 34, 20, 0, 0, 16, 35, 33, 
    19, 53, 43, 46, 44, 35, 22, 19, 0, 0, 0, 0, 0, 10, 31, 
    0, 15, 41, 48, 33, 36, 0, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 23, 51, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 1, 0, 0, 1, 2, 0, 0, 0, 4, 16, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 16, 31, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    4, 0, 0, 0, 0, 0, 0, 0, 0, 2, 11, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 13, 13, 0, 
    0, 42, 0, 0, 2, 48, 0, 18, 3, 0, 0, 0, 0, 27, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 61, 0, 14, 0, 0, 42, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 30, 
    10, 0, 0, 28, 80, 37, 0, 0, 0, 38, 0, 0, 10, 0, 0, 
    1, 0, 22, 0, 46, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 30, 19, 0, 24, 0, 35, 0, 0, 20, 10, 4, 
    0, 0, 0, 0, 0, 69, 2, 0, 6, 0, 39, 15, 33, 6, 0, 
    0, 1, 0, 11, 0, 16, 12, 0, 0, 31, 5, 17, 0, 0, 0, 
    5, 0, 0, 14, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    81, 31, 0, 0, 0, 46, 43, 42, 13, 5, 0, 4, 0, 0, 0, 
    0, 71, 52, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 106, 0, 0, 1, 0, 0, 4, 0, 4, 13, 2, 0, 12, 
    0, 0, 11, 40, 13, 30, 25, 1, 0, 0, 0, 6, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 41, 16, 0, 0, 0, 30, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 10, 10, 22, 0, 0, 
    52, 7, 0, 0, 12, 0, 32, 17, 6, 0, 15, 0, 0, 7, 0, 
    42, 26, 14, 0, 65, 49, 17, 23, 0, 0, 22, 34, 10, 27, 0, 
    3, 0, 13, 0, 0, 0, 36, 23, 45, 0, 11, 2, 0, 15, 32, 
    18, 7, 0, 17, 0, 0, 0, 21, 20, 0, 7, 22, 3, 7, 19, 
    20, 12, 21, 19, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    20, 0, 38, 0, 26, 0, 0, 20, 0, 13, 0, 0, 0, 0, 11, 
    0, 0, 36, 0, 2, 0, 0, 44, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 117, 66, 0, 0, 0, 22, 24, 33, 7, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 2, 
    12, 0, 0, 0, 0, 2, 0, 0, 1, 5, 7, 11, 0, 0, 12, 
    5, 0, 0, 0, 0, 0, 14, 1, 0, 0, 0, 0, 0, 4, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 9, 18, 8, 0, 14, 28, 15, 
    
    -- channel=44
    0, 0, 4, 0, 2, 5, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    3, 6, 8, 0, 12, 35, 0, 0, 0, 14, 11, 0, 0, 0, 0, 
    0, 0, 2, 0, 6, 0, 0, 0, 15, 53, 0, 0, 0, 0, 2, 
    0, 65, 0, 11, 0, 26, 12, 0, 0, 43, 0, 0, 0, 0, 29, 
    0, 55, 0, 77, 44, 44, 0, 0, 0, 75, 7, 0, 4, 0, 15, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 136, 0, 0, 6, 0, 2, 
    0, 0, 0, 0, 43, 44, 0, 0, 0, 105, 0, 0, 8, 21, 0, 
    0, 0, 2, 0, 60, 42, 0, 0, 0, 57, 0, 0, 13, 0, 0, 
    0, 4, 0, 13, 1, 0, 0, 0, 23, 0, 0, 0, 0, 9, 19, 
    0, 0, 0, 59, 0, 2, 35, 9, 0, 0, 0, 0, 32, 30, 0, 
    27, 1, 0, 130, 0, 31, 44, 0, 0, 0, 22, 39, 26, 10, 0, 
    6, 0, 0, 101, 0, 0, 0, 0, 0, 0, 1, 5, 6, 4, 0, 
    0, 13, 47, 0, 0, 0, 0, 0, 0, 7, 14, 14, 0, 1, 20, 
    0, 2, 61, 0, 0, 7, 0, 0, 3, 5, 0, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 11, 0, 5, 48, 0, 0, 
    
    -- channel=45
    0, 2, 6, 6, 6, 2, 6, 4, 1, 0, 0, 0, 5, 7, 4, 
    7, 5, 4, 7, 3, 32, 17, 1, 0, 0, 14, 0, 0, 0, 7, 
    0, 0, 6, 4, 1, 0, 0, 0, 0, 0, 9, 10, 18, 0, 0, 
    24, 6, 5, 1, 9, 0, 20, 20, 13, 0, 20, 0, 0, 6, 0, 
    35, 24, 25, 0, 61, 59, 14, 18, 0, 0, 7, 30, 5, 22, 0, 
    14, 0, 33, 9, 0, 0, 28, 11, 28, 0, 24, 5, 0, 13, 27, 
    25, 6, 0, 15, 0, 6, 0, 31, 9, 0, 8, 12, 0, 1, 21, 
    31, 1, 21, 13, 0, 0, 16, 0, 1, 0, 5, 0, 0, 0, 6, 
    24, 0, 42, 0, 33, 0, 0, 3, 0, 3, 0, 0, 0, 0, 15, 
    0, 0, 29, 0, 0, 19, 0, 26, 12, 0, 0, 0, 4, 11, 1, 
    0, 0, 10, 0, 106, 53, 20, 0, 21, 13, 1, 26, 1, 0, 0, 
    0, 0, 13, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 2, 13, 7, 
    
    -- channel=46
    55, 58, 58, 58, 57, 52, 63, 73, 58, 32, 21, 29, 37, 48, 48, 
    57, 65, 62, 61, 57, 27, 40, 34, 19, 0, 0, 0, 0, 25, 40, 
    10, 35, 63, 66, 66, 44, 10, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 52, 59, 32, 8, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 33, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 29, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 32, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=47
    0, 0, 3, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 3, 3, 0, 6, 58, 5, 0, 0, 5, 21, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 23, 0, 9, 0, 0, 2, 
    2, 48, 3, 4, 2, 9, 26, 5, 0, 0, 0, 0, 0, 0, 0, 
    17, 58, 4, 26, 92, 42, 0, 0, 0, 20, 16, 4, 9, 10, 0, 
    0, 3, 2, 0, 0, 0, 17, 5, 7, 60, 0, 0, 0, 5, 22, 
    0, 0, 0, 0, 0, 26, 0, 6, 0, 21, 0, 0, 0, 15, 8, 
    0, 6, 10, 17, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 1, 0, 0, 4, 18, 0, 0, 0, 0, 8, 19, 
    0, 0, 0, 9, 0, 0, 15, 37, 0, 0, 0, 0, 25, 23, 0, 
    0, 0, 0, 74, 95, 60, 13, 0, 0, 0, 24, 42, 13, 0, 0, 
    0, 0, 11, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 5, 10, 0, 0, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 34, 7, 0, 
    
    -- channel=48
    69, 71, 71, 72, 70, 68, 76, 80, 71, 55, 44, 50, 59, 66, 65, 
    70, 80, 76, 74, 72, 71, 65, 57, 41, 29, 22, 25, 31, 50, 61, 
    36, 50, 75, 77, 75, 64, 36, 30, 23, 25, 16, 14, 17, 24, 54, 
    30, 34, 73, 74, 59, 45, 40, 14, 11, 20, 20, 19, 14, 13, 43, 
    11, 35, 58, 51, 50, 30, 28, 17, 13, 17, 32, 21, 20, 18, 18, 
    0, 15, 54, 42, 28, 20, 36, 29, 24, 21, 11, 9, 18, 14, 17, 
    0, 18, 37, 67, 41, 26, 27, 17, 24, 22, 13, 15, 14, 18, 21, 
    0, 22, 6, 49, 38, 26, 2, 13, 23, 34, 15, 17, 13, 19, 39, 
    0, 7, 0, 20, 17, 19, 28, 24, 19, 38, 27, 7, 17, 42, 60, 
    6, 5, 6, 15, 15, 2, 17, 36, 7, 11, 4, 11, 22, 53, 53, 
    10, 8, 9, 17, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    4, 0, 3, 0, 0, 2, 1, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 3, 6, 0, 8, 1, 0, 0, 0, 3, 0, 0, 7, 10, 0, 
    0, 33, 2, 0, 5, 19, 0, 0, 3, 46, 0, 0, 0, 17, 16, 
    0, 64, 0, 5, 0, 15, 0, 0, 0, 71, 0, 0, 0, 0, 60, 
    0, 37, 0, 66, 0, 0, 0, 0, 0, 82, 0, 0, 0, 0, 29, 
    0, 10, 0, 0, 48, 0, 0, 0, 0, 138, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 64, 29, 0, 0, 0, 118, 0, 0, 4, 9, 0, 
    0, 0, 0, 0, 48, 57, 0, 0, 0, 79, 0, 0, 20, 6, 0, 
    0, 4, 0, 20, 0, 16, 0, 0, 29, 0, 2, 0, 20, 24, 13, 
    0, 4, 0, 56, 0, 7, 35, 0, 0, 0, 0, 0, 34, 32, 0, 
    43, 0, 0, 124, 0, 0, 38, 0, 0, 0, 0, 5, 13, 9, 0, 
    66, 31, 0, 88, 0, 0, 0, 0, 0, 0, 0, 5, 1, 2, 0, 
    0, 59, 71, 0, 0, 0, 0, 0, 0, 0, 6, 5, 0, 2, 10, 
    0, 1, 111, 0, 0, 7, 0, 0, 3, 3, 0, 0, 0, 15, 0, 
    0, 0, 3, 0, 0, 10, 3, 0, 7, 0, 0, 6, 33, 0, 0, 
    
    -- channel=50
    94, 98, 98, 98, 96, 93, 102, 107, 99, 84, 75, 78, 84, 86, 86, 
    97, 103, 102, 101, 100, 86, 88, 88, 73, 47, 28, 29, 45, 76, 84, 
    65, 88, 102, 104, 102, 79, 62, 40, 34, 24, 18, 20, 18, 38, 75, 
    27, 40, 95, 101, 83, 67, 44, 25, 19, 31, 28, 25, 21, 19, 57, 
    23, 28, 81, 88, 60, 37, 31, 22, 15, 29, 31, 25, 21, 20, 25, 
    6, 23, 80, 62, 42, 46, 37, 29, 14, 29, 23, 23, 22, 20, 19, 
    12, 9, 66, 84, 42, 43, 38, 31, 23, 20, 24, 17, 15, 21, 24, 
    12, 17, 21, 61, 50, 41, 22, 25, 34, 31, 29, 17, 19, 26, 52, 
    8, 8, 4, 31, 33, 29, 34, 22, 33, 31, 36, 21, 20, 49, 74, 
    20, 10, 10, 7, 26, 21, 30, 26, 10, 39, 21, 17, 28, 66, 81, 
    14, 16, 9, 18, 18, 10, 7, 12, 11, 1, 0, 0, 0, 0, 0, 
    0, 4, 23, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    63, 65, 65, 65, 64, 62, 68, 68, 65, 58, 49, 50, 52, 53, 51, 
    63, 65, 69, 67, 69, 75, 65, 60, 46, 41, 33, 28, 34, 49, 51, 
    45, 57, 65, 67, 68, 76, 47, 29, 25, 48, 43, 37, 27, 29, 50, 
    25, 41, 66, 70, 60, 52, 50, 28, 25, 56, 43, 36, 22, 12, 45, 
    46, 65, 63, 84, 87, 62, 52, 28, 18, 43, 59, 32, 29, 17, 18, 
    45, 72, 62, 46, 85, 71, 65, 44, 17, 67, 58, 30, 36, 27, 14, 
    48, 63, 59, 48, 62, 73, 85, 49, 34, 72, 54, 29, 27, 37, 29, 
    58, 69, 46, 50, 60, 95, 51, 51, 33, 67, 55, 30, 35, 37, 41, 
    68, 78, 30, 62, 38, 50, 47, 40, 49, 43, 50, 18, 18, 45, 60, 
    76, 77, 44, 57, 52, 28, 53, 62, 34, 46, 18, 11, 30, 60, 62, 
    78, 74, 45, 87, 75, 53, 65, 67, 35, 14, 12, 15, 24, 38, 32, 
    51, 68, 68, 112, 73, 22, 21, 21, 17, 14, 14, 14, 16, 20, 16, 
    10, 39, 71, 94, 25, 16, 14, 13, 11, 11, 15, 18, 20, 20, 23, 
    11, 12, 54, 63, 19, 18, 14, 13, 14, 15, 13, 17, 13, 19, 16, 
    9, 11, 14, 32, 8, 13, 18, 15, 19, 19, 14, 14, 30, 27, 7, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 
    0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 2, 5, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 7, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 6, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 13, 4, 0, 7, 0, 0, 6, 22, 2, 
    0, 0, 0, 14, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 5, 10, 0, 0, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 15, 0, 28, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 60, 26, 0, 0, 8, 8, 29, 0, 0, 
    91, 0, 0, 0, 3, 0, 0, 7, 0, 0, 55, 0, 44, 23, 0, 
    80, 0, 39, 0, 0, 0, 43, 36, 28, 0, 0, 45, 0, 36, 0, 
    54, 0, 59, 0, 0, 12, 33, 28, 59, 0, 58, 83, 0, 16, 5, 
    43, 20, 18, 63, 0, 0, 7, 30, 75, 0, 90, 40, 0, 0, 17, 
    14, 27, 5, 24, 0, 0, 106, 22, 54, 0, 51, 60, 0, 0, 26, 
    25, 0, 95, 0, 0, 8, 34, 0, 0, 19, 0, 97, 0, 0, 0, 
    2, 0, 116, 0, 43, 0, 0, 0, 0, 25, 84, 5, 0, 0, 6, 
    0, 0, 113, 0, 50, 0, 0, 23, 80, 31, 0, 0, 0, 0, 1, 
    0, 0, 20, 0, 151, 107, 6, 11, 19, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 187, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 130, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    31, 0, 0, 35, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 
    
    -- channel=54
    78, 83, 82, 83, 84, 80, 85, 92, 89, 75, 65, 66, 69, 72, 73, 
    82, 88, 87, 86, 86, 77, 76, 79, 65, 43, 24, 26, 39, 61, 70, 
    61, 70, 86, 89, 87, 80, 54, 39, 25, 20, 9, 12, 13, 28, 60, 
    24, 33, 78, 90, 79, 62, 37, 16, 10, 22, 19, 17, 11, 9, 45, 
    11, 19, 63, 82, 51, 30, 23, 13, 9, 20, 24, 14, 14, 11, 20, 
    0, 14, 56, 56, 37, 30, 27, 21, 9, 23, 16, 13, 15, 12, 8, 
    0, 8, 44, 71, 43, 34, 32, 20, 15, 21, 14, 9, 9, 12, 10, 
    0, 12, 14, 48, 44, 34, 14, 18, 17, 29, 18, 10, 12, 13, 34, 
    1, 4, 0, 22, 22, 23, 24, 19, 22, 33, 28, 14, 10, 32, 58, 
    12, 5, 0, 8, 11, 15, 25, 20, 4, 27, 14, 10, 14, 53, 69, 
    11, 10, 1, 14, 5, 1, 4, 6, 0, 2, 0, 0, 0, 0, 3, 
    0, 0, 6, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    49, 42, 45, 45, 50, 39, 50, 55, 47, 33, 25, 27, 30, 42, 42, 
    49, 45, 47, 47, 44, 9, 47, 29, 23, 3, 0, 19, 28, 28, 36, 
    21, 28, 50, 50, 55, 50, 24, 29, 4, 0, 0, 0, 6, 30, 24, 
    0, 30, 51, 46, 32, 19, 0, 0, 0, 5, 0, 9, 0, 14, 28, 
    0, 0, 47, 19, 0, 3, 0, 0, 6, 10, 0, 0, 0, 0, 40, 
    0, 0, 37, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 28, 23, 12, 0, 0, 0, 0, 0, 0, 0, 8, 0, 4, 
    0, 0, 20, 7, 17, 0, 0, 4, 0, 17, 0, 8, 0, 6, 27, 
    0, 0, 0, 0, 18, 25, 11, 0, 0, 49, 3, 7, 16, 18, 35, 
    0, 0, 0, 0, 0, 8, 0, 0, 22, 0, 0, 0, 0, 22, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 3, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    6, 13, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    9, 12, 0, 20, 0, 0, 2, 0, 0, 0, 5, 5, 0, 0, 0, 
    21, 2, 0, 15, 0, 0, 27, 25, 15, 7, 11, 27, 32, 21, 13, 
    61, 44, 12, 9, 9, 39, 40, 40, 42, 48, 54, 59, 60, 59, 58, 
    68, 56, 42, 0, 29, 51, 52, 50, 50, 54, 62, 59, 64, 72, 67, 
    73, 66, 59, 26, 44, 54, 49, 48, 58, 59, 68, 70, 73, 70, 77, 
    70, 73, 65, 44, 49, 57, 62, 58, 57, 55, 57, 66, 68, 62, 68, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 19, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 16, 0, 0, 0, 3, 2, 0, 0, 27, 0, 0, 0, 0, 0, 
    6, 4, 0, 0, 0, 20, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    11, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 15, 0, 14, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    21, 13, 0, 34, 16, 17, 30, 4, 0, 0, 0, 9, 12, 0, 0, 
    24, 11, 0, 51, 6, 0, 3, 0, 0, 5, 12, 15, 18, 20, 17, 
    22, 22, 10, 35, 0, 12, 13, 10, 9, 13, 18, 23, 22, 18, 26, 
    18, 21, 35, 0, 0, 14, 13, 13, 14, 18, 21, 19, 16, 32, 27, 
    21, 23, 23, 0, 3, 10, 8, 9, 19, 21, 19, 15, 30, 36, 11, 
    
    -- channel=58
    3, 4, 10, 11, 9, 7, 10, 13, 11, 0, 0, 0, 0, 4, 2, 
    13, 16, 13, 10, 13, 38, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 8, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 18, 33, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    0, 2, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 2, 1, 5, 
    0, 0, 0, 2, 0, 6, 2, 0, 7, 0, 7, 0, 0, 0, 4, 
    0, 0, 0, 3, 0, 0, 29, 4, 0, 0, 1, 14, 19, 0, 1, 
    57, 0, 0, 0, 5, 0, 7, 0, 1, 0, 38, 0, 26, 5, 0, 
    62, 0, 16, 0, 23, 0, 25, 18, 10, 0, 6, 22, 1, 30, 0, 
    0, 0, 30, 0, 0, 0, 46, 20, 44, 0, 19, 37, 0, 16, 11, 
    0, 21, 3, 40, 0, 0, 11, 26, 47, 0, 46, 18, 0, 0, 10, 
    0, 44, 0, 35, 0, 0, 42, 0, 34, 0, 32, 24, 0, 0, 19, 
    10, 0, 30, 0, 0, 0, 18, 1, 0, 5, 0, 38, 0, 0, 0, 
    7, 0, 70, 0, 11, 0, 0, 28, 0, 0, 41, 3, 0, 0, 3, 
    0, 0, 64, 0, 85, 0, 0, 11, 45, 24, 0, 0, 0, 0, 0, 
    0, 0, 23, 0, 41, 31, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 73, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 83, 16, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 15, 23, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 32, 8, 0, 0, 0, 0, 10, 0, 
    3, 21, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 12, 0, 0, 25, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 0, 0, 25, 31, 
    0, 0, 0, 0, 0, 26, 31, 27, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=61
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 
    0, 0, 0, 0, 0, 0, 24, 0, 10, 0, 5, 7, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 29, 10, 0, 0, 8, 7, 28, 0, 0, 
    63, 0, 4, 0, 8, 0, 0, 11, 2, 0, 35, 0, 20, 16, 0, 
    55, 0, 39, 0, 0, 9, 33, 26, 14, 0, 2, 39, 0, 26, 0, 
    40, 0, 49, 0, 0, 3, 26, 22, 44, 0, 45, 47, 0, 13, 17, 
    37, 20, 8, 36, 0, 0, 0, 27, 44, 0, 54, 28, 0, 0, 18, 
    24, 17, 27, 22, 0, 0, 63, 4, 22, 0, 25, 34, 0, 0, 11, 
    26, 0, 71, 0, 15, 0, 12, 0, 0, 27, 0, 45, 0, 0, 0, 
    0, 0, 73, 0, 27, 2, 0, 6, 9, 0, 42, 0, 0, 0, 8, 
    0, 0, 68, 0, 67, 13, 0, 7, 50, 30, 0, 0, 0, 0, 4, 
    0, 0, 15, 0, 81, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 52, 13, 0, 4, 0, 0, 0, 0, 0, 0, 0, 8, 
    21, 0, 0, 0, 3, 0, 0, 0, 0, 0, 1, 0, 0, 3, 36, 
    
    -- channel=62
    0, 0, 2, 5, 4, 0, 2, 3, 3, 0, 0, 0, 4, 7, 8, 
    6, 3, 0, 5, 0, 41, 17, 0, 0, 0, 24, 8, 0, 0, 8, 
    0, 0, 3, 6, 0, 0, 17, 0, 0, 0, 11, 15, 26, 0, 0, 
    63, 0, 5, 0, 18, 0, 26, 14, 11, 0, 42, 0, 19, 14, 0, 
    58, 3, 28, 0, 56, 24, 30, 35, 12, 0, 16, 40, 10, 38, 0, 
    8, 0, 43, 0, 0, 0, 59, 24, 60, 0, 32, 30, 0, 20, 32, 
    21, 25, 0, 42, 0, 0, 0, 40, 38, 0, 36, 32, 0, 0, 26, 
    23, 30, 8, 36, 0, 0, 33, 0, 24, 0, 24, 26, 0, 0, 13, 
    30, 0, 63, 0, 23, 0, 4, 18, 0, 15, 0, 15, 0, 0, 3, 
    1, 0, 73, 0, 9, 0, 0, 42, 0, 0, 16, 0, 0, 0, 4, 
    0, 0, 54, 0, 133, 35, 0, 0, 36, 30, 7, 13, 0, 0, 0, 
    0, 0, 14, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    9, 0, 0, 31, 12, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 8, 2, 0, 0, 17, 28, 
    
    -- channel=63
    30, 33, 29, 30, 29, 29, 33, 38, 34, 31, 33, 31, 28, 29, 29, 
    28, 32, 30, 32, 27, 0, 31, 34, 47, 5, 0, 2, 15, 23, 24, 
    33, 29, 31, 35, 31, 37, 45, 28, 2, 0, 0, 0, 0, 9, 15, 
    9, 0, 27, 30, 27, 12, 0, 0, 0, 0, 12, 9, 13, 7, 1, 
    2, 0, 28, 4, 0, 0, 12, 8, 7, 0, 0, 6, 0, 0, 3, 
    15, 0, 35, 42, 12, 33, 0, 1, 0, 0, 12, 27, 0, 0, 0, 
    12, 0, 30, 44, 0, 0, 0, 3, 10, 0, 21, 5, 0, 0, 0, 
    3, 0, 0, 6, 0, 0, 30, 17, 13, 0, 15, 14, 0, 0, 18, 
    0, 0, 17, 0, 6, 30, 18, 0, 0, 10, 12, 41, 2, 0, 3, 
    0, 0, 11, 0, 7, 8, 0, 0, 0, 27, 31, 8, 0, 0, 28, 
    0, 0, 15, 0, 0, 0, 0, 2, 11, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 39, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 24, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 30, 18, 22, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    91, 79, 18, 0, 0, 0, 0, 0, 0, 0, 21, 52, 65, 47, 0, 
    0, 0, 0, 17, 14, 47, 61, 49, 33, 0, 0, 0, 0, 0, 0, 
    95, 98, 46, 0, 0, 9, 28, 1, 0, 1, 24, 43, 35, 45, 48, 
    33, 0, 19, 28, 4, 0, 0, 0, 50, 42, 20, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 21, 0, 0, 2, 4, 16, 41, 62, 50, 
    38, 77, 83, 83, 76, 64, 54, 43, 41, 30, 47, 39, 23, 19, 17, 
    62, 65, 71, 87, 94, 98, 97, 91, 79, 72, 58, 44, 26, 0, 0, 
    1, 7, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 13, 25, 10, 0, 0, 48, 0, 0, 0, 19, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    35, 35, 35, 35, 35, 36, 35, 36, 34, 36, 38, 35, 36, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 49, 39, 32, 35, 35, 35, 
    37, 36, 36, 35, 34, 37, 35, 42, 40, 43, 24, 39, 35, 35, 36, 
    33, 35, 35, 35, 36, 50, 29, 41, 25, 23, 11, 5, 37, 37, 37, 
    26, 21, 44, 35, 35, 45, 24, 38, 31, 40, 50, 49, 39, 28, 40, 
    18, 16, 32, 27, 45, 42, 56, 55, 49, 52, 23, 14, 21, 0, 36, 
    34, 23, 32, 26, 50, 1, 0, 0, 0, 41, 50, 50, 50, 51, 31, 
    0, 0, 0, 5, 33, 16, 5, 30, 32, 23, 6, 0, 0, 3, 2, 
    0, 45, 19, 23, 38, 50, 50, 55, 35, 39, 50, 48, 46, 40, 31, 
    28, 45, 44, 44, 42, 38, 42, 22, 25, 19, 23, 20, 10, 9, 11, 
    0, 0, 0, 0, 3, 11, 26, 26, 29, 21, 13, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 3, 3, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 9, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    84, 72, 0, 0, 0, 0, 0, 0, 0, 0, 24, 57, 72, 31, 0, 
    0, 0, 0, 19, 13, 88, 95, 74, 31, 0, 0, 0, 0, 0, 0, 
    100, 91, 41, 0, 0, 0, 0, 0, 0, 0, 42, 67, 58, 60, 41, 
    2, 0, 0, 6, 0, 0, 0, 0, 40, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 22, 2, 0, 8, 3, 26, 51, 63, 34, 
    41, 79, 76, 71, 56, 39, 20, 3, 11, 0, 24, 15, 0, 0, 0, 
    60, 47, 67, 92, 109, 114, 107, 97, 79, 67, 46, 22, 0, 0, 0, 
    9, 11, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 36, 20, 2, 0, 56, 21, 0, 17, 53, 23, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 12, 34, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=67
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 8, 0, 3, 9, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 8, 4, 7, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 10, 7, 8, 5, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=68
    59, 60, 60, 60, 60, 60, 60, 60, 59, 60, 63, 60, 60, 60, 61, 
    59, 60, 60, 60, 60, 60, 60, 59, 60, 51, 61, 65, 60, 60, 61, 
    59, 60, 60, 60, 61, 60, 61, 55, 52, 50, 65, 67, 60, 60, 61, 
    69, 64, 62, 60, 61, 52, 62, 49, 58, 58, 60, 78, 62, 62, 62, 
    41, 49, 68, 58, 60, 54, 66, 60, 66, 64, 56, 46, 44, 60, 62, 
    66, 72, 67, 50, 57, 45, 53, 55, 59, 55, 56, 61, 52, 80, 65, 
    43, 50, 58, 58, 57, 13, 42, 57, 81, 63, 54, 45, 51, 49, 58, 
    42, 63, 29, 59, 52, 54, 74, 53, 44, 43, 41, 48, 54, 62, 68, 
    94, 72, 66, 78, 76, 61, 65, 52, 65, 64, 68, 60, 55, 46, 44, 
    80, 56, 64, 65, 66, 65, 64, 60, 65, 52, 57, 47, 53, 51, 51, 
    14, 28, 29, 27, 27, 35, 49, 50, 48, 45, 45, 47, 52, 48, 46, 
    0, 28, 17, 8, 6, 17, 55, 41, 45, 47, 50, 56, 43, 32, 44, 
    0, 6, 10, 1, 1, 5, 64, 26, 26, 20, 15, 17, 32, 40, 52, 
    0, 3, 7, 5, 3, 4, 28, 36, 18, 24, 33, 38, 29, 39, 52, 
    0, 0, 1, 1, 3, 4, 11, 27, 30, 32, 24, 23, 33, 40, 53, 
    
    -- channel=69
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 2, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 17, 3, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 6, 32, 17, 11, 17, 0, 0, 0, 0, 
    4, 10, 3, 2, 3, 1, 0, 5, 25, 12, 0, 0, 0, 0, 0, 
    
    -- channel=70
    12, 11, 11, 11, 10, 10, 10, 12, 10, 10, 12, 11, 11, 11, 10, 
    11, 10, 10, 10, 9, 10, 9, 11, 8, 8, 0, 0, 10, 10, 9, 
    8, 7, 10, 10, 10, 11, 6, 7, 0, 11, 0, 0, 10, 8, 10, 
    7, 12, 8, 9, 10, 21, 0, 30, 32, 44, 41, 0, 9, 9, 9, 
    0, 0, 0, 4, 7, 29, 6, 20, 15, 17, 0, 0, 0, 0, 5, 
    66, 58, 10, 0, 0, 0, 0, 0, 0, 28, 42, 53, 71, 0, 1, 
    0, 0, 0, 15, 38, 38, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 0, 0, 11, 75, 58, 16, 0, 0, 10, 18, 16, 32, 5, 
    0, 40, 58, 33, 10, 5, 0, 28, 28, 9, 17, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 1, 0, 13, 0, 7, 6, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 17, 2, 
    11, 0, 41, 34, 12, 0, 50, 69, 44, 45, 45, 38, 14, 10, 3, 
    23, 0, 0, 0, 4, 1, 0, 22, 29, 16, 0, 0, 6, 3, 0, 
    52, 4, 0, 5, 4, 3, 0, 13, 0, 5, 20, 8, 2, 0, 0, 
    37, 16, 10, 10, 10, 10, 0, 4, 25, 8, 2, 0, 0, 0, 0, 
    
    -- channel=71
    10, 9, 9, 9, 9, 9, 9, 9, 8, 11, 11, 9, 9, 9, 9, 
    10, 9, 9, 9, 9, 9, 9, 8, 11, 18, 5, 7, 9, 9, 9, 
    8, 8, 8, 9, 9, 11, 10, 17, 21, 28, 20, 2, 9, 9, 9, 
    13, 13, 10, 8, 8, 12, 6, 20, 23, 31, 26, 22, 13, 12, 11, 
    26, 20, 2, 6, 9, 12, 9, 12, 16, 27, 30, 26, 23, 6, 12, 
    29, 20, 18, 11, 11, 26, 15, 13, 8, 19, 28, 28, 26, 16, 14, 
    26, 13, 18, 7, 25, 41, 25, 20, 21, 22, 22, 20, 16, 19, 11, 
    13, 24, 23, 4, 15, 24, 25, 32, 17, 16, 23, 22, 22, 23, 30, 
    5, 25, 15, 13, 16, 19, 23, 27, 32, 38, 32, 38, 30, 28, 25, 
    28, 32, 37, 36, 35, 36, 38, 38, 38, 40, 43, 39, 38, 32, 23, 
    31, 23, 36, 34, 32, 34, 42, 39, 39, 38, 38, 34, 30, 30, 17, 
    13, 16, 14, 19, 16, 17, 4, 47, 42, 37, 30, 33, 15, 8, 5, 
    20, 7, 0, 4, 9, 8, 0, 0, 0, 0, 0, 0, 0, 5, 9, 
    20, 8, 5, 6, 7, 7, 0, 0, 0, 0, 0, 0, 4, 8, 12, 
    19, 9, 10, 10, 8, 9, 0, 0, 0, 0, 0, 6, 6, 10, 13, 
    
    -- channel=72
    2, 1, 1, 1, 1, 1, 1, 0, 0, 2, 3, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 1, 3, 19, 0, 0, 1, 1, 1, 
    0, 0, 0, 1, 0, 3, 0, 13, 9, 23, 0, 0, 1, 0, 1, 
    6, 7, 1, 0, 0, 16, 0, 17, 19, 29, 27, 0, 6, 4, 2, 
    6, 0, 0, 0, 0, 11, 0, 5, 6, 16, 17, 12, 5, 0, 3, 
    23, 18, 5, 0, 2, 0, 0, 0, 0, 24, 26, 23, 37, 0, 2, 
    13, 0, 0, 3, 31, 46, 21, 15, 0, 5, 3, 1, 0, 3, 0, 
    0, 26, 4, 0, 9, 28, 14, 19, 8, 18, 27, 23, 16, 20, 11, 
    0, 16, 18, 4, 6, 15, 10, 24, 20, 18, 23, 25, 16, 13, 17, 
    0, 20, 23, 26, 28, 31, 42, 37, 32, 39, 33, 35, 29, 20, 12, 
    7, 10, 16, 12, 4, 4, 21, 23, 29, 30, 29, 25, 23, 19, 2, 
    6, 0, 12, 14, 4, 0, 19, 49, 39, 34, 23, 15, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=73
    14, 13, 13, 13, 12, 13, 12, 14, 13, 13, 12, 12, 13, 13, 12, 
    14, 13, 13, 13, 13, 13, 12, 13, 16, 34, 0, 3, 13, 13, 12, 
    13, 13, 13, 14, 12, 17, 9, 27, 18, 24, 0, 0, 13, 12, 12, 
    2, 9, 9, 13, 14, 35, 0, 32, 0, 6, 0, 0, 8, 9, 10, 
    8, 0, 0, 12, 13, 25, 0, 15, 4, 16, 15, 14, 15, 0, 4, 
    0, 0, 7, 15, 16, 22, 3, 1, 0, 17, 5, 0, 18, 0, 0, 
    10, 0, 0, 0, 29, 43, 0, 0, 0, 13, 17, 19, 9, 17, 0, 
    0, 0, 12, 0, 7, 3, 0, 21, 17, 20, 17, 1, 0, 0, 0, 
    0, 12, 0, 0, 0, 14, 7, 17, 0, 0, 0, 8, 0, 4, 8, 
    0, 8, 4, 4, 4, 5, 12, 4, 2, 9, 3, 8, 0, 0, 0, 
    14, 0, 16, 10, 7, 1, 4, 3, 5, 8, 1, 0, 0, 0, 0, 
    13, 0, 14, 19, 10, 0, 0, 8, 0, 0, 0, 0, 4, 12, 0, 
    28, 0, 12, 22, 9, 3, 0, 57, 55, 56, 44, 28, 5, 0, 0, 
    50, 5, 4, 10, 5, 4, 0, 86, 92, 44, 8, 0, 4, 0, 0, 
    43, 7, 2, 2, 3, 1, 0, 30, 11, 0, 7, 2, 0, 0, 0, 
    
    -- channel=74
    2, 5, 5, 5, 6, 6, 6, 4, 5, 4, 7, 6, 5, 5, 6, 
    4, 5, 5, 5, 5, 5, 6, 4, 0, 0, 36, 16, 4, 5, 5, 
    9, 9, 6, 4, 5, 2, 12, 0, 17, 0, 48, 51, 5, 6, 6, 
    7, 3, 8, 6, 6, 0, 27, 0, 0, 0, 0, 18, 7, 7, 7, 
    45, 65, 47, 12, 8, 0, 9, 0, 2, 0, 23, 39, 42, 76, 15, 
    0, 0, 18, 22, 26, 48, 83, 76, 66, 0, 0, 0, 0, 15, 20, 
    52, 80, 43, 11, 0, 0, 0, 0, 5, 20, 37, 46, 54, 49, 68, 
    44, 0, 0, 48, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 
    46, 5, 0, 2, 26, 18, 33, 0, 6, 25, 29, 24, 47, 48, 19, 
    85, 51, 54, 48, 41, 28, 6, 0, 7, 0, 10, 0, 0, 5, 13, 
    0, 12, 2, 27, 45, 57, 54, 52, 35, 22, 14, 8, 0, 0, 6, 
    0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 114, 2, 0, 0, 16, 4, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 3, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 14, 
    
    -- channel=75
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 29, 40, 0, 0, 0, 0, 0, 0, 0, 
    55, 29, 0, 0, 0, 0, 9, 0, 0, 0, 0, 3, 8, 4, 0, 
    121, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 4, 0, 
    10, 25, 3, 1, 0, 0, 0, 0, 0, 0, 11, 23, 36, 22, 3, 
    39, 55, 37, 49, 57, 64, 109, 79, 77, 79, 78, 45, 0, 0, 3, 
    38, 54, 26, 30, 55, 58, 35, 0, 0, 0, 0, 0, 8, 0, 0, 
    8, 59, 57, 54, 59, 59, 72, 0, 0, 0, 30, 8, 0, 0, 0, 
    7, 59, 61, 64, 65, 65, 69, 16, 39, 26, 0, 0, 0, 0, 0, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 8, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 15, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 1, 21, 0, 
    0, 0, 0, 7, 0, 0, 0, 17, 21, 0, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 0, 17, 23, 0, 0, 0, 0, 4, 9, 10, 12, 
    60, 0, 15, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 2, 14, 10, 1, 4, 8, 7, 0, 0, 8, 
    3, 7, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 10, 6, 12, 
    0, 4, 2, 2, 4, 4, 3, 0, 0, 0, 18, 15, 4, 9, 4, 
    0, 12, 11, 9, 9, 10, 12, 0, 20, 18, 6, 5, 8, 9, 7, 
    
    -- channel=77
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 8, 12, 5, 0, 9, 4, 0, 0, 0, 0, 0, 0, 
    24, 14, 11, 14, 15, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 17, 14, 15, 16, 16, 3, 0, 0, 0, 2, 0, 0, 0, 0, 
    22, 22, 20, 19, 19, 18, 14, 9, 10, 4, 0, 0, 0, 0, 0, 
    
    -- channel=78
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 19, 22, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    72, 67, 17, 0, 0, 0, 0, 0, 0, 0, 27, 53, 68, 38, 0, 
    0, 0, 0, 21, 26, 78, 98, 80, 38, 0, 0, 0, 0, 0, 0, 
    93, 80, 50, 0, 0, 0, 0, 0, 0, 6, 44, 66, 63, 56, 45, 
    0, 0, 0, 4, 0, 0, 0, 0, 36, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 33, 22, 0, 15, 20, 33, 53, 57, 35, 
    32, 77, 72, 70, 56, 43, 24, 7, 13, 6, 21, 18, 3, 5, 0, 
    39, 36, 47, 71, 86, 90, 92, 87, 73, 61, 43, 22, 0, 0, 0, 
    9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 33, 18, 4, 0, 47, 21, 0, 11, 42, 22, 0, 0, 0, 
    0, 0, 2, 2, 0, 0, 24, 37, 42, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 32, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 39, 0, 0, 0, 
    5, 31, 44, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 52, 1, 
    0, 2, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 57, 3, 
    0, 36, 17, 20, 0, 0, 26, 58, 62, 0, 0, 0, 0, 0, 31, 
    62, 39, 0, 63, 11, 0, 13, 0, 0, 0, 0, 4, 16, 13, 13, 
    172, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 2, 17, 
    0, 33, 1, 12, 17, 23, 10, 5, 0, 0, 0, 9, 28, 10, 20, 
    0, 47, 0, 0, 0, 17, 84, 0, 10, 18, 31, 17, 0, 7, 31, 
    0, 14, 11, 0, 0, 4, 133, 0, 0, 0, 0, 16, 19, 21, 34, 
    0, 0, 5, 0, 1, 2, 57, 6, 0, 19, 28, 20, 5, 23, 30, 
    0, 0, 1, 0, 3, 5, 24, 23, 26, 35, 5, 1, 13, 18, 26, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 28, 32, 22, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 9, 6, 0, 0, 0, 0, 0, 
    72, 72, 13, 0, 0, 0, 0, 0, 0, 0, 20, 44, 39, 45, 0, 
    0, 0, 0, 10, 9, 0, 6, 14, 32, 0, 0, 0, 0, 0, 0, 
    19, 58, 0, 0, 0, 48, 80, 16, 0, 0, 0, 4, 18, 30, 38, 
    84, 31, 55, 48, 22, 0, 0, 6, 42, 36, 33, 23, 6, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 3, 9, 7, 4, 24, 24, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 23, 26, 18, 
    5, 26, 29, 26, 17, 21, 67, 65, 49, 52, 57, 61, 31, 0, 14, 
    13, 6, 0, 0, 5, 12, 8, 0, 0, 0, 0, 0, 0, 16, 18, 
    1, 11, 8, 7, 11, 11, 0, 0, 0, 0, 8, 25, 1, 7, 10, 
    0, 16, 17, 16, 15, 17, 6, 0, 12, 27, 4, 0, 6, 11, 13, 
    
    -- channel=81
    27, 25, 25, 25, 25, 26, 25, 26, 25, 28, 24, 25, 26, 25, 25, 
    26, 26, 26, 26, 25, 26, 25, 26, 31, 54, 6, 15, 26, 25, 25, 
    25, 25, 25, 26, 24, 31, 21, 46, 30, 30, 0, 0, 26, 26, 25, 
    16, 21, 24, 26, 26, 55, 7, 42, 7, 12, 0, 0, 25, 25, 25, 
    11, 0, 4, 24, 26, 37, 14, 28, 17, 34, 38, 29, 26, 0, 22, 
    0, 0, 23, 25, 31, 42, 19, 17, 1, 32, 13, 6, 21, 0, 17, 
    8, 0, 4, 0, 51, 24, 0, 0, 0, 34, 36, 33, 21, 29, 0, 
    0, 0, 0, 0, 11, 8, 0, 40, 18, 10, 4, 0, 0, 0, 0, 
    0, 24, 0, 4, 12, 33, 32, 32, 7, 12, 8, 24, 10, 8, 6, 
    0, 5, 2, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 18, 13, 20, 12, 0, 0, 0, 0, 
    40, 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 2, 0, 0, 0, 
    
    -- channel=82
    6, 5, 5, 5, 4, 4, 4, 5, 4, 3, 4, 4, 4, 5, 4, 
    5, 4, 4, 4, 3, 4, 3, 6, 3, 0, 0, 0, 5, 4, 4, 
    0, 1, 3, 5, 5, 4, 0, 0, 0, 0, 0, 0, 4, 3, 4, 
    3, 6, 2, 4, 5, 5, 0, 14, 20, 30, 34, 0, 3, 3, 3, 
    0, 0, 0, 0, 1, 16, 3, 11, 8, 1, 0, 0, 0, 0, 0, 
    47, 47, 0, 0, 0, 0, 0, 0, 0, 8, 33, 45, 56, 0, 0, 
    0, 0, 0, 4, 12, 15, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 65, 51, 0, 0, 0, 0, 7, 7, 23, 0, 
    0, 9, 49, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 45, 16, 16, 21, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 7, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 
    
    -- channel=83
    72, 71, 71, 71, 71, 71, 71, 72, 71, 71, 71, 70, 71, 71, 71, 
    72, 71, 71, 72, 71, 71, 71, 71, 71, 68, 48, 64, 72, 71, 72, 
    70, 70, 72, 72, 72, 74, 68, 71, 49, 41, 36, 51, 71, 71, 72, 
    67, 70, 69, 72, 74, 75, 57, 66, 56, 57, 54, 58, 69, 70, 71, 
    14, 14, 49, 68, 72, 67, 66, 69, 71, 73, 59, 40, 31, 27, 68, 
    54, 62, 65, 52, 56, 40, 29, 36, 44, 63, 56, 58, 59, 55, 65, 
    7, 3, 28, 45, 63, 21, 0, 15, 49, 65, 55, 43, 34, 39, 33, 
    0, 32, 11, 25, 43, 58, 63, 62, 32, 28, 24, 21, 24, 36, 46, 
    0, 51, 55, 61, 65, 62, 56, 47, 44, 41, 41, 39, 26, 19, 19, 
    18, 22, 24, 28, 30, 31, 33, 26, 25, 21, 14, 6, 6, 6, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 1, 18, 17, 7, 13, 
    0, 0, 0, 0, 0, 0, 0, 34, 40, 33, 12, 0, 1, 8, 22, 
    0, 0, 0, 0, 0, 0, 0, 21, 14, 0, 0, 2, 4, 10, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 5, 16, 31, 
    
    -- channel=84
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 39, 0, 0, 0, 
    0, 2, 23, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 7, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 
    0, 2, 0, 0, 0, 0, 8, 35, 51, 0, 0, 0, 0, 0, 4, 
    22, 36, 0, 42, 0, 0, 20, 0, 0, 0, 0, 0, 10, 10, 17, 
    126, 11, 0, 14, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 10, 
    0, 38, 0, 0, 0, 8, 49, 0, 5, 6, 17, 17, 0, 0, 16, 
    0, 7, 5, 0, 0, 0, 118, 0, 0, 0, 0, 0, 3, 15, 27, 
    0, 0, 4, 0, 0, 0, 56, 1, 0, 0, 13, 24, 3, 15, 23, 
    0, 0, 1, 1, 2, 3, 25, 19, 8, 35, 5, 0, 9, 13, 20, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 15, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 16, 44, 0, 0, 
    0, 0, 0, 0, 15, 71, 3, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 29, 0, 2, 0, 0, 20, 16, 7, 7, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 19, 35, 21, 0, 0, 80, 47, 37, 22, 3, 0, 0, 0, 
    53, 0, 0, 9, 15, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    85, 15, 9, 15, 14, 13, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    67, 32, 24, 24, 22, 21, 5, 0, 14, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 23, 27, 0, 0, 
    0, 0, 0, 0, 0, 46, 32, 18, 0, 0, 0, 0, 0, 0, 0, 
    50, 29, 0, 0, 0, 38, 0, 0, 0, 0, 10, 33, 14, 25, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 16, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 19, 27, 10, 
    0, 42, 31, 32, 23, 12, 9, 0, 0, 6, 7, 14, 0, 0, 0, 
    46, 21, 48, 59, 62, 61, 62, 60, 51, 52, 33, 13, 0, 0, 0, 
    31, 0, 5, 15, 19, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 12, 29, 35, 19, 12, 0, 40, 29, 43, 64, 25, 0, 0, 0, 
    41, 11, 12, 17, 12, 11, 0, 56, 87, 21, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 31, 20, 34, 40, 42, 23, 21, 5, 5, 4, 2, 0, 0, 0, 
    8, 45, 0, 0, 19, 36, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 41, 42, 26, 26, 30, 115, 4, 5, 6, 27, 29, 0, 0, 0, 
    0, 27, 33, 30, 29, 29, 92, 76, 84, 61, 11, 0, 0, 0, 0, 
    0, 11, 15, 18, 21, 21, 43, 51, 19, 9, 0, 0, 0, 0, 0, 
    
    -- channel=88
    83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 82, 83, 83, 83, 
    83, 83, 83, 83, 83, 83, 83, 82, 82, 78, 72, 81, 83, 83, 83, 
    83, 84, 84, 83, 84, 85, 81, 82, 67, 51, 62, 76, 83, 83, 84, 
    77, 78, 81, 84, 85, 83, 78, 70, 56, 51, 46, 71, 80, 81, 82, 
    49, 54, 77, 83, 84, 73, 78, 77, 80, 81, 77, 67, 63, 65, 82, 
    43, 54, 80, 73, 79, 72, 70, 73, 74, 69, 50, 47, 40, 66, 82, 
    42, 45, 58, 53, 62, 0, 0, 16, 62, 86, 82, 73, 67, 69, 67, 
    0, 30, 23, 59, 58, 40, 53, 68, 55, 39, 24, 18, 22, 31, 51, 
    11, 61, 45, 62, 78, 78, 80, 54, 50, 53, 54, 53, 50, 47, 40, 
    51, 49, 53, 52, 52, 49, 42, 34, 37, 24, 29, 15, 14, 17, 25, 
    0, 0, 0, 0, 4, 11, 19, 18, 17, 10, 2, 0, 4, 14, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 29, 20, 23, 
    0, 0, 0, 0, 0, 0, 18, 69, 70, 63, 41, 13, 6, 16, 35, 
    0, 0, 0, 0, 0, 0, 0, 34, 22, 0, 0, 4, 13, 23, 43, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 9, 15, 27, 45, 
    
    -- channel=89
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 2, 0, 0, 0, 0, 0, 4, 28, 37, 42, 12, 0, 1, 0, 
    0, 0, 0, 0, 0, 10, 12, 8, 12, 0, 0, 0, 0, 0, 0, 
    80, 79, 12, 0, 0, 0, 0, 0, 0, 8, 35, 58, 59, 32, 0, 
    0, 0, 0, 20, 19, 0, 0, 18, 14, 0, 0, 0, 0, 0, 0, 
    0, 52, 0, 0, 0, 72, 88, 0, 0, 0, 0, 7, 21, 40, 19, 
    61, 46, 71, 54, 15, 0, 0, 0, 30, 2, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 
    0, 0, 30, 21, 3, 0, 82, 59, 35, 37, 48, 42, 5, 0, 17, 
    10, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 21, 21, 
    14, 5, 1, 1, 4, 5, 0, 0, 0, 0, 38, 35, 10, 8, 9, 
    3, 23, 19, 16, 16, 18, 0, 1, 43, 44, 15, 5, 13, 16, 15, 
    
    -- channel=90
    29, 30, 30, 30, 30, 29, 30, 29, 28, 29, 31, 30, 29, 30, 30, 
    29, 30, 30, 29, 29, 29, 29, 29, 27, 8, 9, 28, 30, 30, 30, 
    24, 26, 29, 30, 30, 29, 27, 17, 0, 9, 10, 18, 29, 29, 30, 
    36, 35, 32, 29, 30, 20, 20, 30, 48, 62, 67, 58, 33, 32, 32, 
    0, 0, 15, 23, 27, 35, 40, 35, 42, 34, 7, 0, 0, 0, 31, 
    75, 77, 48, 0, 0, 0, 0, 0, 0, 34, 58, 72, 68, 60, 34, 
    0, 0, 0, 24, 41, 0, 22, 54, 61, 23, 0, 0, 0, 0, 0, 
    0, 54, 1, 3, 27, 70, 89, 31, 0, 0, 16, 33, 44, 58, 46, 
    56, 62, 59, 56, 37, 17, 7, 8, 34, 19, 20, 8, 0, 0, 0, 
    8, 0, 0, 0, 0, 5, 17, 20, 19, 12, 11, 5, 15, 10, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 27, 15, 
    0, 0, 0, 0, 0, 0, 46, 74, 56, 54, 59, 53, 7, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 4, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 11, 23, 
    
    -- channel=91
    35, 34, 34, 34, 34, 34, 35, 34, 33, 35, 35, 34, 34, 34, 34, 
    35, 35, 35, 35, 35, 35, 35, 35, 34, 38, 32, 32, 35, 35, 35, 
    35, 34, 34, 35, 34, 35, 36, 38, 42, 45, 31, 31, 35, 35, 35, 
    38, 39, 36, 34, 34, 35, 29, 43, 42, 48, 44, 34, 40, 38, 37, 
    42, 37, 27, 33, 34, 40, 31, 37, 37, 42, 44, 44, 39, 34, 38, 
    40, 34, 35, 31, 29, 37, 32, 33, 38, 47, 47, 43, 42, 22, 39, 
    37, 34, 31, 31, 41, 54, 36, 33, 23, 37, 37, 37, 32, 36, 34, 
    24, 16, 35, 17, 39, 39, 32, 41, 39, 40, 41, 35, 34, 34, 32, 
    0, 40, 31, 26, 34, 41, 39, 45, 40, 42, 41, 43, 39, 43, 42, 
    21, 42, 45, 47, 47, 49, 52, 49, 44, 45, 44, 44, 36, 33, 31, 
    23, 20, 26, 25, 23, 27, 35, 36, 38, 38, 35, 33, 34, 28, 22, 
    7, 2, 10, 8, 4, 2, 11, 37, 33, 28, 24, 17, 14, 20, 16, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 12, 18, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 16, 24, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 14, 20, 26, 
    
    -- channel=92
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 11, 19, 20, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    18, 12, 0, 0, 0, 0, 0, 0, 0, 4, 18, 19, 28, 0, 0, 
    0, 0, 0, 0, 8, 53, 19, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 16, 20, 0, 0, 27, 17, 14, 0, 4, 18, 17, 16, 13, 8, 
    0, 0, 12, 0, 0, 0, 0, 4, 6, 1, 0, 2, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 14, 4, 11, 11, 9, 4, 
    20, 8, 9, 3, 0, 0, 0, 0, 0, 1, 6, 7, 8, 14, 7, 
    34, 8, 27, 38, 33, 23, 9, 49, 33, 28, 22, 13, 5, 10, 6, 
    47, 26, 8, 22, 30, 28, 0, 0, 0, 0, 0, 0, 8, 8, 4, 
    56, 30, 25, 27, 29, 29, 0, 0, 0, 0, 6, 9, 14, 9, 1, 
    53, 41, 38, 37, 34, 35, 21, 0, 5, 8, 13, 17, 12, 11, 4, 
    
    -- channel=93
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 21, 9, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 16, 0, 
    0, 0, 0, 0, 8, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 
    0, 28, 0, 0, 0, 4, 26, 3, 0, 0, 0, 0, 2, 7, 7, 
    16, 17, 7, 11, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 24, 28, 19, 16, 18, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 9, 8, 12, 9, 7, 0, 0, 0, 0, 3, 14, 0, 0, 0, 
    0, 7, 7, 9, 8, 7, 15, 26, 43, 38, 4, 0, 0, 0, 0, 
    8, 9, 7, 7, 7, 6, 9, 23, 13, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=96
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 3, 7, 3, 0, 0, 0, 
    0, 0, 30, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 16, 0, 0, 0, 0, 0, 0, 10, 2, 5, 18, 22, 0, 
    0, 0, 0, 0, 36, 0, 4, 31, 18, 0, 0, 0, 0, 0, 0, 
    0, 74, 0, 14, 12, 10, 18, 0, 0, 0, 0, 12, 9, 24, 0, 
    21, 36, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 0, 
    0, 0, 9, 0, 0, 0, 86, 25, 29, 27, 27, 22, 0, 0, 2, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 2, 8, 
    0, 1, 1, 0, 0, 2, 0, 18, 0, 0, 17, 12, 0, 0, 5, 
    0, 3, 7, 5, 7, 6, 0, 21, 15, 16, 5, 0, 0, 0, 4, 
    
    -- channel=97
    81, 81, 81, 81, 81, 82, 82, 82, 81, 81, 81, 82, 82, 81, 82, 
    81, 82, 82, 82, 81, 81, 81, 81, 80, 81, 70, 78, 81, 81, 82, 
    81, 81, 82, 82, 81, 83, 79, 82, 66, 60, 59, 73, 82, 82, 83, 
    75, 78, 83, 82, 82, 89, 72, 77, 57, 57, 46, 64, 83, 82, 83, 
    39, 44, 79, 80, 82, 87, 76, 82, 76, 80, 82, 68, 58, 58, 85, 
    50, 53, 87, 66, 77, 71, 69, 73, 74, 82, 59, 53, 49, 52, 84, 
    29, 27, 57, 48, 84, 0, 0, 2, 43, 88, 81, 69, 70, 70, 58, 
    0, 27, 19, 45, 65, 46, 55, 73, 49, 33, 17, 13, 17, 32, 43, 
    0, 88, 45, 63, 75, 82, 82, 65, 52, 58, 60, 60, 51, 46, 37, 
    48, 39, 40, 39, 38, 40, 39, 23, 32, 12, 24, 12, 8, 13, 21, 
    0, 0, 0, 0, 0, 0, 1, 3, 5, 0, 0, 0, 0, 10, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 23, 15, 20, 
    0, 0, 0, 0, 0, 0, 0, 33, 27, 25, 11, 0, 0, 16, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 21, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 14, 21, 30, 47, 
    
    -- channel=98
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 23, 31, 46, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 20, 0, 0, 0, 0, 0, 0, 0, 1, 40, 40, 38, 23, 0, 
    0, 0, 0, 8, 0, 13, 47, 91, 44, 0, 0, 0, 0, 0, 0, 
    12, 34, 0, 0, 23, 58, 35, 0, 0, 10, 38, 54, 51, 55, 3, 
    74, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 15, 0, 
    0, 0, 0, 0, 0, 0, 87, 83, 70, 69, 70, 29, 0, 0, 20, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 8, 12, 
    0, 3, 0, 1, 2, 2, 0, 0, 0, 14, 47, 9, 0, 6, 1, 
    2, 18, 16, 15, 17, 20, 10, 21, 47, 19, 0, 0, 4, 5, 4, 
    
    -- channel=99
    21, 21, 21, 21, 21, 21, 21, 20, 20, 23, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 20, 23, 39, 32, 22, 20, 21, 21, 
    24, 22, 21, 21, 20, 22, 23, 34, 44, 33, 43, 28, 22, 22, 21, 
    22, 22, 23, 21, 20, 27, 27, 16, 8, 1, 0, 19, 25, 24, 23, 
    68, 63, 35, 23, 23, 13, 17, 16, 19, 31, 55, 64, 65, 44, 27, 
    0, 0, 20, 41, 42, 77, 77, 68, 47, 20, 3, 0, 0, 13, 27, 
    70, 60, 48, 13, 19, 12, 5, 0, 10, 39, 57, 64, 57, 57, 50, 
    5, 3, 21, 30, 14, 0, 0, 34, 43, 24, 9, 0, 0, 0, 21, 
    0, 3, 0, 3, 25, 38, 53, 36, 24, 43, 39, 50, 59, 59, 41, 
    51, 60, 61, 57, 51, 42, 31, 25, 30, 24, 35, 26, 22, 25, 20, 
    36, 31, 40, 51, 60, 64, 62, 57, 51, 42, 34, 23, 8, 6, 13, 
    10, 15, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 12, 4, 4, 
    0, 14, 10, 4, 1, 1, 24, 0, 0, 0, 14, 0, 0, 5, 14, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 17, 24, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 15, 17, 23, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 14, 0, 0, 0, 0, 0, 0, 
    12, 18, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 27, 0, 0, 0, 8, 42, 0, 0, 0, 2, 0, 0, 0, 8, 
    0, 14, 16, 1, 5, 12, 76, 0, 0, 0, 0, 0, 3, 9, 11, 
    0, 12, 14, 10, 12, 13, 30, 23, 0, 9, 17, 18, 3, 6, 8, 
    0, 7, 13, 12, 13, 13, 15, 28, 20, 29, 10, 0, 6, 3, 4, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 32, 42, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 5, 0, 0, 0, 0, 0, 0, 
    85, 90, 18, 0, 0, 0, 0, 0, 0, 0, 20, 60, 59, 56, 0, 
    0, 0, 0, 0, 5, 0, 0, 12, 43, 0, 0, 0, 0, 0, 0, 
    0, 69, 0, 0, 0, 68, 114, 15, 0, 0, 0, 0, 19, 36, 38, 
    84, 31, 68, 58, 7, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 2, 
    0, 0, 16, 23, 3, 0, 50, 93, 50, 50, 65, 75, 22, 0, 11, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 15, 
    6, 1, 0, 0, 0, 0, 0, 0, 0, 0, 28, 45, 0, 1, 0, 
    0, 23, 19, 13, 14, 16, 6, 0, 31, 58, 17, 0, 3, 8, 6, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 2, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    25, 1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 27, 27, 37, 47, 43, 25, 15, 6, 0, 0, 0, 0, 0, 0, 
    0, 22, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 29, 6, 5, 10, 102, 2, 0, 1, 17, 5, 0, 0, 0, 
    0, 7, 10, 4, 7, 7, 45, 18, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 1, 0, 12, 3, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=103
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 26, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 
    0, 0, 0, 0, 0, 0, 23, 18, 12, 0, 0, 0, 0, 9, 0, 
    19, 45, 14, 0, 0, 0, 0, 0, 8, 0, 0, 0, 6, 0, 25, 
    46, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 
    49, 11, 14, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    6, 31, 13, 30, 40, 45, 36, 34, 20, 12, 12, 11, 8, 0, 4, 
    0, 41, 0, 0, 0, 19, 31, 0, 0, 0, 0, 0, 2, 0, 5, 
    0, 21, 29, 4, 4, 10, 130, 22, 17, 15, 23, 25, 2, 2, 4, 
    0, 6, 14, 8, 8, 9, 79, 78, 55, 39, 12, 5, 0, 1, 2, 
    0, 0, 0, 0, 0, 0, 25, 39, 11, 17, 0, 0, 0, 0, 0, 
    
    -- channel=104
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 31, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    69, 40, 0, 0, 0, 0, 0, 0, 0, 0, 19, 48, 58, 0, 0, 
    0, 0, 0, 17, 7, 65, 53, 38, 9, 0, 0, 0, 0, 0, 0, 
    75, 55, 18, 0, 0, 43, 0, 0, 0, 0, 26, 49, 32, 43, 9, 
    0, 0, 6, 0, 0, 0, 0, 0, 45, 37, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 8, 12, 0, 0, 0, 8, 22, 44, 33, 
    0, 54, 48, 47, 39, 30, 28, 9, 6, 10, 13, 17, 0, 0, 0, 
    51, 29, 52, 61, 66, 66, 62, 58, 51, 48, 29, 7, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 23, 27, 3, 0, 0, 11, 0, 7, 47, 34, 0, 0, 0, 
    34, 0, 0, 1, 0, 0, 0, 24, 68, 22, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 8, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 2, 0, 0, 0, 0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 27, 3, 36, 27, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    95, 105, 25, 0, 0, 0, 0, 0, 0, 0, 14, 50, 69, 84, 0, 
    0, 0, 0, 30, 17, 73, 92, 79, 57, 0, 0, 0, 0, 0, 0, 
    99, 128, 63, 0, 0, 0, 7, 0, 0, 0, 34, 58, 61, 50, 78, 
    70, 0, 12, 52, 0, 0, 0, 0, 46, 27, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 20, 0, 0, 5, 2, 9, 46, 63, 44, 
    51, 81, 81, 77, 67, 49, 20, 15, 21, 7, 28, 19, 10, 13, 15, 
    68, 73, 75, 102, 119, 131, 114, 104, 79, 69, 56, 40, 19, 0, 6, 
    8, 49, 0, 0, 2, 26, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 29, 48, 25, 11, 11, 132, 34, 13, 23, 58, 56, 0, 0, 0, 
    0, 5, 13, 9, 7, 7, 57, 33, 64, 38, 0, 0, 0, 5, 6, 
    0, 0, 0, 0, 0, 0, 14, 20, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 20, 38, 46, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 56, 0, 0, 0, 0, 0, 0, 0, 0, 33, 54, 70, 17, 0, 
    0, 0, 0, 0, 15, 35, 3, 31, 12, 0, 0, 0, 0, 0, 0, 
    0, 54, 0, 0, 0, 70, 72, 7, 0, 0, 3, 21, 27, 37, 16, 
    10, 5, 45, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 20, 31, 10, 0, 43, 111, 68, 62, 63, 51, 0, 0, 0, 
    39, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 4, 2, 0, 
    50, 7, 0, 2, 4, 4, 0, 0, 0, 0, 26, 20, 0, 0, 0, 
    25, 31, 24, 20, 20, 21, 5, 0, 33, 24, 6, 0, 0, 0, 0, 
    
    -- channel=108
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 13, 0, 0, 0, 
    8, 1, 0, 0, 0, 0, 11, 0, 17, 18, 38, 58, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 27, 0, 15, 0, 0, 0, 0, 3, 0, 
    44, 62, 21, 0, 0, 0, 0, 0, 0, 0, 12, 36, 18, 83, 6, 
    0, 0, 0, 15, 0, 0, 28, 68, 78, 0, 0, 0, 0, 0, 0, 
    38, 59, 0, 33, 0, 27, 80, 0, 0, 0, 0, 15, 40, 42, 41, 
    174, 14, 38, 45, 16, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 13, 20, 
    0, 32, 0, 0, 0, 11, 95, 52, 46, 48, 63, 48, 10, 0, 36, 
    0, 5, 0, 0, 0, 1, 82, 0, 0, 0, 0, 0, 17, 35, 43, 
    0, 1, 4, 0, 0, 1, 51, 0, 0, 0, 45, 50, 12, 27, 31, 
    0, 9, 12, 9, 11, 15, 32, 22, 45, 65, 18, 3, 19, 27, 33, 
    
    -- channel=109
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 17, 26, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 7, 3, 0, 0, 0, 0, 0, 
    68, 70, 8, 0, 0, 0, 0, 0, 0, 0, 18, 43, 56, 14, 0, 
    0, 0, 0, 0, 15, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 39, 0, 0, 0, 57, 72, 24, 0, 0, 0, 0, 0, 11, 14, 
    0, 13, 57, 39, 9, 0, 0, 0, 26, 10, 6, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    5, 0, 34, 30, 9, 0, 24, 56, 21, 23, 33, 38, 24, 0, 0, 
    25, 0, 0, 0, 0, 2, 0, 14, 36, 20, 0, 0, 0, 3, 0, 
    41, 2, 0, 0, 1, 1, 0, 0, 0, 0, 4, 21, 0, 0, 0, 
    15, 19, 10, 9, 9, 7, 0, 0, 11, 28, 8, 0, 0, 0, 0, 
    
    -- channel=110
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 36, 35, 23, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 90, 64, 13, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=111
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 32, 45, 18, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 3, 0, 0, 0, 0, 0, 0, 
    81, 83, 0, 0, 0, 0, 0, 0, 0, 0, 34, 61, 55, 45, 0, 
    0, 0, 0, 12, 0, 0, 0, 35, 38, 0, 0, 0, 0, 0, 0, 
    0, 67, 0, 0, 0, 82, 101, 0, 0, 0, 0, 10, 25, 46, 21, 
    105, 22, 73, 44, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 19, 12, 0, 0, 84, 77, 46, 50, 67, 61, 0, 0, 17, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 31, 0, 3, 0, 
    0, 19, 15, 11, 13, 14, 8, 0, 44, 47, 6, 0, 5, 9, 7, 
    
    -- channel=112
    5, 6, 6, 6, 5, 5, 5, 7, 7, 4, 3, 5, 6, 6, 6, 
    5, 6, 6, 6, 6, 6, 5, 6, 4, 0, 0, 6, 6, 6, 6, 
    4, 5, 6, 6, 6, 5, 2, 0, 0, 0, 0, 0, 6, 5, 5, 
    0, 0, 4, 6, 6, 7, 4, 5, 0, 1, 2, 2, 0, 1, 3, 
    0, 0, 0, 6, 5, 9, 8, 6, 1, 0, 0, 0, 0, 0, 1, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 4, 8, 4, 0, 
    0, 0, 0, 0, 3, 0, 0, 12, 10, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 12, 7, 9, 8, 0, 0, 0, 1, 6, 6, 8, 0, 
    4, 8, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 
    7, 7, 12, 14, 14, 11, 20, 18, 15, 15, 21, 18, 10, 11, 13, 
    18, 10, 20, 19, 15, 16, 30, 54, 56, 46, 29, 29, 25, 15, 6, 
    14, 18, 19, 18, 17, 17, 37, 105, 84, 55, 43, 26, 14, 8, 2, 
    13, 22, 20, 19, 21, 19, 23, 57, 47, 38, 22, 10, 10, 5, 1, 
    
    -- channel=113
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 31, 37, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 43, 0, 0, 0, 
    1, 28, 34, 0, 0, 0, 15, 0, 2, 0, 0, 0, 0, 53, 4, 
    0, 14, 15, 0, 0, 0, 11, 12, 25, 0, 0, 0, 0, 54, 9, 
    0, 38, 13, 16, 0, 0, 18, 37, 52, 0, 0, 0, 1, 0, 36, 
    66, 19, 0, 56, 1, 0, 20, 0, 0, 0, 0, 0, 10, 6, 18, 
    151, 4, 0, 16, 13, 0, 0, 0, 0, 0, 1, 0, 0, 2, 0, 
    66, 0, 6, 1, 1, 0, 0, 0, 0, 0, 0, 0, 2, 7, 20, 
    0, 17, 0, 4, 13, 20, 8, 7, 0, 0, 0, 8, 22, 5, 23, 
    0, 53, 0, 0, 0, 16, 59, 0, 0, 5, 20, 14, 12, 7, 28, 
    0, 13, 10, 0, 0, 2, 149, 0, 0, 0, 0, 8, 7, 24, 33, 
    0, 0, 6, 0, 0, 2, 74, 14, 0, 6, 16, 24, 7, 23, 32, 
    0, 0, 0, 0, 1, 3, 29, 24, 11, 39, 7, 3, 15, 21, 28, 
    
    -- channel=114
    17, 17, 17, 17, 17, 17, 17, 18, 18, 16, 15, 17, 17, 17, 17, 
    17, 17, 17, 17, 17, 17, 17, 17, 15, 7, 12, 17, 17, 17, 17, 
    18, 18, 17, 17, 17, 16, 16, 9, 4, 1, 4, 16, 17, 17, 17, 
    10, 11, 15, 19, 18, 13, 17, 11, 4, 0, 0, 0, 12, 14, 15, 
    0, 0, 17, 20, 17, 18, 14, 17, 10, 5, 0, 0, 0, 13, 14, 
    5, 5, 3, 17, 13, 11, 12, 14, 14, 5, 3, 4, 0, 1, 11, 
    0, 0, 7, 16, 1, 0, 0, 0, 1, 9, 10, 9, 15, 4, 9, 
    1, 0, 0, 9, 11, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 13, 11, 6, 4, 4, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    13, 11, 14, 7, 7, 6, 0, 0, 0, 0, 0, 0, 9, 11, 15, 
    10, 10, 18, 18, 15, 13, 24, 61, 58, 49, 35, 28, 25, 17, 13, 
    16, 15, 16, 15, 15, 14, 44, 97, 82, 51, 37, 26, 20, 16, 12, 
    20, 18, 15, 15, 16, 14, 22, 42, 39, 35, 27, 21, 20, 15, 11, 
    
    -- channel=115
    106, 106, 106, 106, 106, 106, 106, 106, 106, 105, 105, 106, 106, 106, 106, 
    106, 106, 106, 106, 106, 106, 106, 106, 104, 89, 96, 106, 106, 106, 106, 
    105, 106, 106, 106, 106, 106, 106, 98, 86, 74, 82, 102, 106, 107, 107, 
    103, 103, 107, 107, 107, 97, 103, 93, 85, 79, 76, 98, 107, 106, 107, 
    61, 75, 104, 106, 107, 103, 104, 104, 102, 97, 88, 78, 73, 97, 107, 
    76, 82, 96, 92, 95, 84, 83, 89, 98, 95, 85, 81, 68, 90, 107, 
    45, 60, 81, 87, 84, 22, 32, 51, 88, 99, 90, 80, 84, 77, 90, 
    28, 50, 46, 78, 89, 77, 86, 78, 70, 62, 50, 51, 56, 67, 74, 
    49, 90, 80, 90, 96, 94, 95, 80, 70, 70, 71, 64, 61, 59, 57, 
    55, 53, 54, 55, 55, 59, 51, 45, 49, 35, 37, 30, 31, 37, 46, 
    0, 3, 0, 0, 5, 12, 14, 17, 16, 11, 11, 14, 24, 35, 49, 
    0, 8, 5, 0, 0, 0, 15, 4, 4, 6, 19, 34, 42, 44, 60, 
    0, 0, 0, 0, 0, 0, 34, 51, 49, 45, 37, 37, 45, 55, 72, 
    0, 0, 0, 0, 0, 0, 6, 36, 30, 24, 34, 45, 51, 60, 78, 
    5, 0, 0, 0, 0, 0, 0, 19, 21, 42, 51, 51, 57, 66, 80, 
    
    -- channel=116
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 1, 5, 1, 0, 
    0, 0, 0, 0, 0, 14, 44, 73, 22, 0, 0, 0, 0, 0, 0, 
    9, 15, 10, 11, 13, 8, 0, 0, 0, 17, 33, 33, 27, 19, 0, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    20, 29, 17, 7, 0, 0, 0, 0, 0, 0, 0, 0, 18, 13, 0, 
    0, 0, 0, 0, 2, 3, 50, 63, 60, 57, 55, 17, 0, 2, 4, 
    2, 3, 3, 2, 3, 3, 0, 0, 0, 0, 0, 16, 11, 0, 0, 
    0, 3, 0, 0, 2, 2, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 11, 10, 10, 12, 13, 7, 6, 11, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 19, 38, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 23, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 4, 0, 0, 0, 0, 15, 31, 30, 0, 0, 
    0, 0, 0, 0, 0, 49, 11, 0, 0, 7, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 11, 117, 0, 0, 0, 0, 14, 35, 12, 18, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 19, 27, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 11, 4, 19, 20, 
    0, 27, 10, 15, 8, 8, 21, 0, 0, 22, 0, 26, 0, 0, 0, 
    41, 0, 34, 35, 30, 22, 27, 27, 32, 36, 19, 0, 0, 0, 0, 
    41, 0, 17, 25, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 0, 3, 38, 16, 0, 0, 24, 0, 10, 27, 12, 0, 0, 0, 
    117, 0, 0, 8, 1, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 
    118, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=118
    11, 12, 12, 12, 12, 12, 12, 12, 13, 11, 10, 12, 12, 12, 12, 
    11, 12, 12, 12, 12, 12, 12, 12, 12, 4, 8, 11, 12, 12, 12, 
    12, 12, 12, 12, 12, 12, 11, 7, 2, 0, 0, 10, 11, 12, 11, 
    6, 7, 10, 13, 12, 9, 12, 7, 0, 0, 0, 0, 8, 9, 10, 
    0, 0, 10, 14, 12, 13, 11, 11, 5, 0, 0, 0, 0, 8, 8, 
    0, 0, 4, 10, 11, 4, 5, 6, 7, 2, 0, 0, 0, 0, 7, 
    0, 0, 1, 8, 0, 0, 0, 0, 0, 4, 2, 1, 6, 1, 4, 
    0, 0, 0, 8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 3, 7, 4, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 9, 
    2, 2, 10, 9, 5, 4, 13, 35, 34, 30, 23, 22, 17, 13, 9, 
    2, 6, 8, 6, 6, 6, 24, 76, 71, 48, 30, 20, 15, 11, 9, 
    6, 9, 7, 5, 7, 6, 14, 42, 32, 26, 22, 15, 14, 11, 8, 
    
    -- channel=119
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 2, 13, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 15, 18, 14, 13, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 8, 5, 0, 4, 2, 0, 0, 0, 0, 0, 0, 
    19, 24, 20, 10, 10, 13, 31, 0, 0, 0, 5, 8, 0, 0, 0, 
    3, 13, 13, 9, 12, 11, 35, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 16, 15, 15, 14, 13, 27, 10, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=120
    6, 7, 7, 7, 7, 7, 7, 6, 6, 7, 10, 7, 6, 7, 7, 
    6, 6, 6, 6, 7, 6, 7, 6, 3, 7, 24, 9, 6, 6, 6, 
    9, 8, 7, 6, 6, 4, 11, 5, 21, 20, 29, 31, 6, 7, 7, 
    11, 10, 7, 6, 6, 0, 13, 2, 16, 13, 11, 8, 10, 9, 8, 
    31, 34, 22, 8, 7, 4, 5, 6, 12, 12, 30, 36, 29, 41, 12, 
    19, 19, 11, 10, 13, 27, 48, 46, 47, 19, 7, 6, 3, 11, 15, 
    44, 53, 26, 24, 9, 7, 23, 6, 0, 14, 27, 34, 36, 37, 41, 
    55, 3, 12, 16, 13, 1, 8, 14, 26, 17, 6, 3, 6, 4, 11, 
    24, 18, 13, 14, 25, 23, 23, 30, 33, 44, 49, 44, 53, 48, 33, 
    62, 58, 59, 58, 56, 50, 45, 37, 37, 36, 43, 39, 37, 36, 32, 
    17, 32, 28, 40, 44, 56, 65, 67, 60, 56, 51, 47, 40, 15, 19, 
    6, 19, 9, 1, 3, 11, 39, 0, 10, 12, 10, 2, 22, 15, 7, 
    0, 4, 0, 0, 0, 1, 25, 0, 0, 0, 8, 4, 0, 4, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 12, 
    
    -- channel=121
    24, 24, 24, 24, 25, 24, 24, 25, 24, 25, 25, 24, 24, 24, 25, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 20, 18, 25, 25, 24, 25, 
    23, 24, 24, 24, 25, 25, 23, 22, 11, 6, 22, 22, 24, 24, 25, 
    27, 26, 25, 24, 26, 22, 21, 15, 23, 26, 29, 40, 24, 25, 25, 
    0, 0, 21, 22, 24, 16, 31, 22, 31, 28, 21, 9, 4, 8, 25, 
    31, 40, 37, 13, 17, 4, 3, 6, 12, 18, 20, 28, 26, 46, 27, 
    0, 0, 8, 13, 25, 0, 6, 20, 43, 27, 16, 7, 4, 10, 10, 
    0, 36, 1, 20, 10, 21, 43, 31, 6, 1, 4, 10, 17, 22, 34, 
    39, 28, 27, 37, 35, 24, 22, 6, 23, 22, 21, 19, 13, 5, 2, 
    39, 7, 14, 14, 17, 15, 18, 17, 20, 12, 16, 4, 11, 11, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 2, 10, 13, 11, 
    0, 0, 0, 0, 0, 0, 11, 20, 14, 15, 19, 26, 16, 0, 7, 
    0, 0, 0, 0, 0, 0, 14, 4, 10, 5, 0, 0, 0, 4, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 3, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 5, 16, 
    
    -- channel=122
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 13, 0, 0, 6, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 13, 0, 0, 0, 0, 0, 
    
    -- channel=123
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 17, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 7, 0, 22, 0, 0, 
    0, 0, 0, 0, 16, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 20, 0, 0, 0, 4, 5, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 27, 19, 5, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 14, 7, 0, 0, 19, 6, 1, 0, 4, 0, 0, 0, 
    64, 0, 0, 4, 0, 0, 0, 0, 5, 8, 0, 0, 0, 0, 0, 
    63, 7, 1, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 13, 0, 0, 0, 24, 50, 66, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 5, 38, 49, 38, 26, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 10, 18, 7, 1, 0, 0, 0, 0, 0, 
    31, 30, 24, 10, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 32, 35, 27, 9, 0, 0, 0, 0, 
    0, 4, 10, 1, 0, 0, 0, 0, 0, 0, 0, 12, 1, 0, 0, 
    0, 0, 2, 2, 0, 0, 18, 4, 0, 33, 14, 0, 0, 0, 0, 
    0, 0, 1, 4, 4, 5, 26, 46, 14, 0, 0, 0, 0, 0, 0, 
    
    -- channel=125
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 15, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 3, 0, 0, 22, 0, 0, 
    0, 0, 0, 0, 18, 77, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 8, 0, 0, 1, 0, 18, 0, 3, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 9, 0, 4, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 13, 25, 10, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 12, 5, 0, 0, 0, 1, 9, 11, 0, 0, 0, 0, 
    77, 0, 0, 2, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 
    67, 7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=126
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 0, 18, 13, 29, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 32, 0, 0, 0, 0, 0, 0, 0, 10, 27, 36, 63, 0, 0, 
    0, 0, 0, 0, 24, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 25, 0, 0, 0, 62, 34, 7, 0, 0, 7, 9, 3, 15, 0, 
    0, 0, 35, 1, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    14, 0, 34, 35, 11, 0, 17, 71, 35, 31, 27, 16, 0, 0, 0, 
    37, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    78, 5, 0, 3, 3, 3, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    57, 25, 15, 14, 13, 11, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    
    -- channel=127
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 0, 0, 
    0, 0, 0, 3, 0, 27, 19, 11, 0, 0, 0, 0, 0, 0, 0, 
    33, 26, 0, 0, 0, 14, 0, 0, 0, 0, 4, 20, 11, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 
    0, 20, 12, 14, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 17, 31, 38, 42, 41, 36, 30, 24, 25, 11, 0, 0, 0, 0, 
    16, 0, 0, 0, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 7, 29, 29, 13, 7, 0, 74, 62, 61, 64, 41, 0, 0, 0, 
    17, 5, 8, 10, 6, 5, 25, 116, 122, 53, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=128
    5, 11, 7, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 9, 6, 0, 0, 0, 0, 0, 0, 12, 26, 0, 0, 0, 0, 
    0, 10, 3, 0, 0, 0, 0, 21, 12, 12, 26, 18, 0, 0, 0, 
    6, 3, 5, 4, 0, 0, 0, 0, 51, 59, 57, 89, 60, 15, 18, 
    55, 46, 50, 54, 50, 48, 43, 35, 14, 10, 20, 0, 0, 1, 33, 
    3, 0, 0, 4, 0, 0, 4, 16, 10, 0, 0, 0, 0, 0, 0, 
    14, 15, 21, 20, 21, 4, 0, 0, 0, 0, 0, 3, 0, 4, 9, 
    0, 0, 0, 0, 0, 0, 0, 7, 19, 24, 35, 5, 0, 0, 0, 
    25, 48, 39, 23, 26, 39, 40, 19, 0, 0, 0, 0, 1, 0, 13, 
    13, 0, 6, 30, 23, 0, 0, 17, 31, 8, 2, 4, 26, 35, 33, 
    27, 18, 19, 27, 44, 39, 24, 37, 23, 26, 39, 38, 23, 18, 15, 
    34, 28, 29, 32, 14, 18, 24, 12, 21, 23, 22, 29, 13, 16, 11, 
    32, 41, 42, 32, 44, 47, 20, 11, 26, 32, 12, 14, 15, 9, 4, 
    40, 38, 26, 17, 17, 23, 26, 21, 0, 1, 15, 10, 9, 4, 1, 
    4, 4, 6, 6, 2, 0, 8, 13, 19, 11, 9, 7, 6, 5, 10, 
    
    -- channel=129
    48, 9, 40, 38, 44, 33, 40, 49, 35, 42, 37, 38, 34, 45, 30, 
    43, 6, 34, 33, 43, 31, 41, 49, 33, 56, 9, 35, 33, 46, 27, 
    41, 0, 25, 28, 38, 29, 45, 30, 24, 65, 0, 36, 40, 42, 29, 
    40, 0, 28, 30, 34, 27, 35, 33, 28, 23, 0, 0, 25, 42, 18, 
    20, 3, 12, 9, 18, 18, 19, 40, 18, 14, 7, 0, 0, 26, 0, 
    0, 0, 14, 0, 5, 0, 17, 19, 8, 10, 0, 8, 8, 29, 0, 
    7, 0, 4, 0, 9, 17, 14, 8, 2, 6, 0, 15, 33, 0, 6, 
    7, 7, 9, 13, 25, 29, 33, 31, 34, 35, 9, 8, 13, 5, 0, 
    21, 28, 11, 33, 37, 40, 34, 23, 7, 24, 0, 8, 14, 10, 18, 
    7, 4, 27, 28, 24, 18, 24, 30, 20, 26, 17, 25, 23, 16, 0, 
    29, 23, 25, 31, 28, 31, 37, 4, 0, 23, 26, 19, 6, 0, 0, 
    11, 21, 34, 1, 0, 3, 36, 14, 0, 4, 4, 3, 0, 0, 0, 
    7, 24, 30, 14, 9, 3, 0, 0, 1, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=130
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 19, 6, 12, 9, 12, 0, 0, 0, 
    5, 0, 10, 5, 1, 0, 0, 0, 48, 46, 22, 83, 66, 28, 31, 
    62, 44, 51, 62, 63, 62, 46, 39, 0, 0, 0, 0, 0, 0, 33, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 24, 0, 0, 0, 0, 
    6, 32, 3, 0, 1, 17, 10, 0, 0, 0, 0, 0, 0, 0, 25, 
    0, 0, 0, 1, 0, 0, 0, 16, 23, 0, 0, 1, 34, 43, 31, 
    0, 0, 0, 15, 40, 15, 3, 15, 0, 25, 43, 38, 23, 14, 19, 
    0, 0, 0, 0, 0, 0, 33, 5, 2, 11, 23, 16, 3, 8, 6, 
    22, 42, 50, 29, 35, 34, 6, 2, 25, 21, 3, 7, 11, 0, 0, 
    31, 31, 17, 10, 14, 19, 14, 8, 0, 0, 6, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 7, 6, 0, 0, 0, 0, 15, 
    
    -- channel=131
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 0, 0, 0, 0, 8, 
    
    -- channel=132
    66, 68, 79, 73, 73, 66, 67, 62, 68, 68, 57, 63, 60, 66, 64, 
    58, 59, 70, 60, 64, 56, 62, 63, 63, 48, 57, 67, 57, 63, 62, 
    50, 50, 60, 49, 55, 50, 53, 52, 57, 25, 69, 62, 49, 54, 60, 
    42, 44, 52, 47, 43, 47, 42, 45, 31, 28, 39, 30, 55, 46, 41, 
    34, 31, 35, 41, 36, 39, 41, 42, 41, 44, 43, 42, 43, 29, 30, 
    48, 45, 38, 40, 54, 53, 63, 49, 45, 43, 53, 59, 23, 47, 18, 
    54, 37, 38, 56, 62, 56, 64, 57, 58, 56, 59, 46, 30, 34, 0, 
    61, 59, 72, 80, 77, 73, 71, 63, 59, 36, 38, 44, 42, 11, 38, 
    64, 51, 67, 75, 71, 61, 52, 48, 55, 42, 56, 49, 46, 39, 37, 
    52, 76, 72, 62, 58, 62, 60, 50, 43, 52, 53, 46, 33, 22, 24, 
    67, 66, 64, 53, 56, 55, 42, 25, 45, 50, 35, 27, 23, 20, 22, 
    67, 56, 45, 39, 48, 67, 40, 33, 34, 32, 26, 21, 23, 19, 13, 
    55, 45, 37, 36, 30, 27, 32, 33, 28, 23, 21, 24, 17, 20, 19, 
    20, 19, 21, 26, 25, 22, 24, 20, 31, 23, 20, 20, 18, 21, 20, 
    16, 18, 19, 20, 23, 24, 24, 16, 31, 10, 22, 19, 20, 22, 7, 
    
    -- channel=133
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=134
    38, 0, 14, 13, 17, 10, 11, 24, 4, 9, 4, 7, 13, 16, 6, 
    29, 0, 0, 10, 11, 6, 5, 12, 2, 13, 0, 0, 10, 11, 0, 
    25, 0, 0, 11, 5, 7, 14, 0, 0, 41, 0, 0, 7, 1, 0, 
    14, 0, 0, 0, 0, 0, 10, 17, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 16, 5, 21, 0, 15, 0, 
    12, 4, 28, 6, 30, 14, 16, 19, 12, 23, 12, 44, 52, 8, 15, 
    7, 6, 6, 0, 0, 30, 30, 43, 44, 35, 1, 0, 37, 0, 19, 
    31, 44, 51, 42, 33, 28, 27, 20, 7, 12, 0, 0, 7, 59, 57, 
    5, 0, 0, 7, 9, 1, 0, 11, 5, 52, 19, 9, 7, 13, 0, 
    31, 24, 21, 5, 11, 20, 18, 1, 0, 7, 7, 9, 0, 0, 0, 
    10, 17, 12, 9, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 24, 4, 12, 0, 10, 14, 0, 0, 0, 0, 4, 1, 7, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 4, 0, 10, 4, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 3, 3, 6, 7, 9, 
    6, 3, 3, 2, 5, 8, 2, 4, 0, 20, 4, 6, 5, 5, 10, 
    
    -- channel=135
    47, 40, 36, 36, 30, 24, 18, 18, 15, 16, 13, 11, 16, 14, 11, 
    39, 29, 24, 25, 17, 16, 13, 10, 13, 21, 6, 5, 12, 10, 8, 
    30, 22, 13, 12, 9, 9, 12, 11, 10, 27, 10, 5, 9, 4, 4, 
    15, 11, 1, 0, 0, 0, 6, 12, 19, 26, 21, 21, 0, 0, 0, 
    12, 8, 10, 3, 0, 0, 6, 23, 32, 37, 30, 23, 9, 4, 3, 
    26, 29, 29, 20, 21, 33, 35, 43, 33, 32, 24, 8, 15, 0, 26, 
    35, 30, 34, 25, 34, 37, 45, 42, 40, 38, 18, 6, 4, 17, 13, 
    41, 36, 34, 41, 41, 43, 46, 46, 36, 33, 5, 0, 5, 9, 8, 
    49, 37, 38, 41, 49, 45, 41, 35, 31, 25, 13, 13, 14, 15, 10, 
    49, 43, 42, 44, 42, 43, 39, 36, 22, 22, 20, 21, 19, 19, 13, 
    42, 50, 48, 43, 39, 30, 38, 33, 28, 25, 24, 26, 24, 24, 19, 
    39, 45, 46, 40, 37, 37, 37, 28, 25, 29, 31, 26, 28, 23, 21, 
    38, 40, 41, 35, 32, 31, 30, 32, 30, 26, 29, 27, 25, 23, 22, 
    29, 28, 29, 30, 28, 25, 27, 28, 24, 34, 23, 22, 23, 23, 23, 
    19, 19, 23, 23, 26, 27, 29, 24, 18, 31, 21, 21, 23, 21, 20, 
    
    -- channel=136
    48, 17, 27, 23, 22, 12, 9, 16, 3, 6, 0, 1, 5, 9, 0, 
    37, 6, 9, 12, 9, 4, 6, 7, 0, 26, 0, 0, 2, 4, 0, 
    26, 0, 0, 2, 0, 0, 9, 0, 0, 44, 0, 0, 2, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 13, 17, 23, 14, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 18, 25, 29, 20, 6, 0, 12, 0, 
    19, 7, 28, 8, 25, 20, 30, 35, 24, 28, 0, 6, 27, 0, 8, 
    25, 23, 24, 17, 22, 39, 41, 43, 41, 32, 0, 0, 8, 0, 17, 
    35, 35, 33, 35, 36, 37, 37, 36, 25, 30, 0, 0, 0, 29, 18, 
    36, 28, 19, 32, 38, 36, 34, 29, 13, 29, 2, 3, 6, 6, 0, 
    46, 32, 34, 35, 36, 32, 27, 21, 5, 14, 10, 14, 8, 10, 0, 
    36, 41, 38, 34, 20, 20, 42, 27, 0, 9, 12, 17, 15, 11, 10, 
    19, 33, 52, 32, 30, 12, 26, 22, 15, 16, 17, 18, 18, 15, 12, 
    13, 22, 25, 22, 19, 15, 18, 17, 14, 17, 17, 8, 18, 12, 13, 
    13, 12, 14, 11, 13, 11, 14, 17, 7, 24, 13, 12, 13, 12, 11, 
    9, 8, 11, 11, 13, 14, 14, 12, 0, 25, 10, 12, 11, 9, 12, 
    
    -- channel=137
    10, 0, 0, 0, 2, 3, 6, 20, 1, 9, 11, 7, 12, 13, 3, 
    16, 0, 0, 7, 8, 11, 14, 13, 4, 41, 0, 2, 16, 17, 4, 
    21, 0, 0, 13, 14, 13, 29, 11, 0, 69, 0, 0, 22, 18, 4, 
    27, 0, 12, 13, 26, 15, 29, 23, 26, 34, 0, 3, 0, 18, 5, 
    15, 2, 18, 6, 20, 13, 11, 27, 7, 3, 0, 0, 0, 41, 9, 
    0, 0, 11, 0, 0, 0, 0, 6, 0, 0, 0, 0, 40, 6, 31, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 8, 42, 25, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 3, 16, 39, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 7, 10, 14, 19, 
    3, 0, 0, 0, 0, 0, 0, 6, 0, 0, 4, 19, 17, 27, 9, 
    0, 0, 0, 3, 0, 0, 21, 18, 0, 0, 13, 22, 10, 7, 9, 
    0, 0, 16, 0, 0, 0, 19, 1, 0, 5, 5, 3, 7, 1, 10, 
    0, 0, 10, 0, 0, 3, 2, 0, 0, 3, 2, 0, 12, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 2, 0, 10, 1, 1, 1, 0, 1, 
    2, 0, 0, 0, 0, 0, 0, 5, 0, 20, 0, 2, 0, 0, 19, 
    
    -- channel=138
    0, 16, 18, 12, 10, 11, 13, 0, 17, 12, 16, 12, 0, 4, 12, 
    0, 17, 26, 4, 13, 6, 10, 14, 16, 0, 43, 22, 0, 9, 15, 
    0, 19, 28, 0, 10, 1, 0, 34, 36, 0, 65, 56, 4, 15, 22, 
    0, 14, 29, 29, 13, 12, 0, 0, 4, 0, 10, 35, 85, 36, 51, 
    26, 22, 18, 44, 35, 41, 30, 2, 0, 0, 2, 0, 20, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    2, 0, 0, 10, 4, 0, 0, 0, 0, 0, 8, 15, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 34, 12, 0, 0, 0, 
    2, 24, 25, 16, 11, 20, 12, 0, 0, 0, 0, 0, 0, 0, 20, 
    0, 0, 10, 7, 0, 0, 0, 10, 32, 6, 0, 0, 8, 0, 1, 
    19, 0, 0, 4, 36, 34, 0, 0, 10, 23, 16, 0, 0, 0, 0, 
    36, 4, 0, 0, 0, 22, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 23, 15, 10, 12, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 36, 0, 0, 0, 
    37, 27, 0, 30, 12, 6, 0, 0, 9, 13, 51, 5, 0, 0, 0, 
    17, 12, 5, 26, 0, 4, 10, 25, 29, 17, 7, 0, 0, 0, 0, 
    26, 28, 31, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    27, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 9, 2, 
    18, 0, 0, 16, 29, 2, 0, 2, 8, 0, 0, 11, 18, 26, 32, 
    9, 0, 0, 4, 1, 2, 13, 16, 4, 11, 23, 30, 20, 41, 45, 
    22, 25, 31, 35, 25, 20, 23, 25, 49, 19, 32, 33, 41, 47, 43, 
    42, 47, 46, 45, 44, 42, 34, 28, 37, 19, 38, 41, 46, 48, 24, 
    
    -- channel=140
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    3, 8, 0, 3, 1, 4, 0, 0, 0, 0, 17, 10, 7, 0, 0, 
    0, 1, 0, 2, 0, 0, 0, 0, 9, 3, 13, 0, 0, 0, 0, 
    0, 5, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 1, 2, 
    0, 3, 3, 4, 4, 4, 1, 0, 5, 0, 0, 0, 1, 0, 0, 
    
    -- channel=141
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 2, 1, 1, 3, 
    3, 3, 3, 3, 1, 0, 0, 3, 0, 3, 2, 2, 1, 0, 14, 
    
    -- channel=142
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 13, 13, 20, 20, 1, 0, 0, 
    11, 0, 20, 18, 8, 0, 0, 0, 39, 45, 17, 68, 74, 38, 31, 
    63, 44, 53, 62, 68, 64, 51, 42, 8, 0, 0, 0, 0, 3, 37, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 21, 27, 5, 0, 0, 0, 
    11, 28, 8, 0, 5, 17, 10, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 19, 24, 0, 0, 9, 33, 42, 33, 
    0, 0, 0, 18, 36, 20, 5, 9, 0, 27, 41, 37, 25, 16, 18, 
    0, 0, 0, 0, 0, 0, 34, 11, 3, 12, 21, 15, 4, 8, 8, 
    21, 39, 45, 28, 27, 26, 8, 4, 22, 20, 6, 7, 11, 2, 0, 
    21, 24, 13, 8, 14, 17, 11, 8, 0, 0, 7, 2, 1, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 12, 5, 5, 1, 0, 0, 0, 10, 
    
    -- channel=143
    0, 18, 16, 0, 0, 0, 0, 0, 7, 0, 0, 1, 0, 0, 0, 
    0, 15, 19, 0, 2, 0, 0, 0, 2, 0, 35, 11, 0, 0, 5, 
    0, 10, 21, 0, 0, 0, 0, 2, 15, 0, 70, 18, 0, 0, 11, 
    0, 9, 2, 5, 0, 0, 0, 0, 0, 0, 17, 18, 63, 0, 12, 
    0, 1, 0, 17, 1, 5, 1, 0, 0, 0, 1, 14, 19, 0, 6, 
    23, 9, 0, 18, 5, 0, 0, 0, 0, 0, 41, 17, 0, 26, 0, 
    8, 0, 0, 33, 21, 0, 0, 0, 0, 0, 34, 5, 0, 0, 0, 
    0, 0, 6, 7, 2, 0, 0, 0, 0, 0, 26, 15, 0, 0, 8, 
    0, 0, 36, 14, 0, 0, 0, 0, 6, 0, 16, 0, 0, 0, 0, 
    0, 22, 2, 0, 8, 1, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 1, 22, 0, 0, 41, 2, 0, 0, 0, 0, 0, 
    48, 1, 0, 0, 9, 32, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    3, 7, 3, 9, 0, 0, 3, 0, 23, 0, 0, 0, 0, 1, 0, 
    0, 6, 4, 6, 4, 0, 0, 0, 41, 0, 0, 0, 0, 6, 0, 
    
    -- channel=144
    27, 34, 28, 18, 14, 6, 2, 0, 1, 0, 0, 0, 0, 0, 0, 
    11, 20, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 26, 23, 30, 22, 0, 0, 
    30, 36, 25, 19, 31, 30, 37, 21, 25, 28, 47, 51, 11, 0, 2, 
    35, 17, 6, 29, 16, 28, 37, 44, 51, 43, 35, 0, 0, 0, 0, 
    49, 50, 70, 76, 55, 45, 40, 32, 18, 0, 0, 0, 0, 0, 29, 
    31, 8, 13, 28, 26, 14, 4, 4, 19, 19, 37, 8, 0, 2, 0, 
    26, 64, 52, 20, 18, 35, 33, 13, 1, 5, 6, 0, 0, 0, 0, 
    37, 37, 31, 19, 12, 7, 0, 0, 11, 1, 0, 0, 0, 0, 3, 
    34, 21, 11, 7, 24, 32, 3, 20, 13, 0, 3, 0, 6, 10, 2, 
    29, 13, 3, 17, 1, 0, 4, 21, 11, 0, 10, 17, 5, 15, 19, 
    0, 0, 7, 17, 17, 10, 6, 5, 28, 25, 10, 14, 14, 21, 21, 
    14, 18, 18, 19, 23, 28, 23, 10, 18, 3, 17, 14, 20, 21, 3, 
    
    -- channel=145
    22, 0, 0, 8, 15, 11, 20, 36, 15, 26, 22, 22, 24, 31, 13, 
    28, 0, 2, 18, 24, 20, 30, 29, 17, 66, 0, 16, 28, 35, 12, 
    33, 0, 2, 23, 33, 24, 47, 19, 6, 85, 0, 3, 35, 34, 15, 
    34, 0, 20, 14, 35, 22, 38, 42, 32, 18, 0, 0, 0, 32, 5, 
    6, 0, 8, 0, 13, 9, 5, 32, 0, 1, 0, 0, 0, 44, 3, 
    0, 0, 10, 0, 0, 0, 0, 1, 0, 0, 0, 0, 48, 15, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 40, 18, 23, 
    0, 0, 0, 0, 0, 0, 1, 9, 3, 35, 0, 1, 14, 20, 0, 
    0, 0, 0, 0, 5, 4, 2, 2, 0, 17, 0, 8, 8, 14, 17, 
    0, 0, 0, 0, 0, 0, 4, 18, 0, 4, 4, 25, 20, 20, 0, 
    0, 0, 0, 6, 0, 0, 31, 1, 0, 9, 15, 15, 7, 0, 4, 
    0, 0, 19, 0, 0, 0, 22, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 3, 
    
    -- channel=146
    3, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 1, 8, 7, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 29, 36, 0, 0, 
    0, 0, 0, 0, 0, 2, 1, 16, 21, 11, 0, 0, 13, 0, 0, 
    0, 15, 24, 15, 5, 0, 0, 0, 0, 0, 0, 0, 0, 41, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=147
    54, 38, 60, 65, 71, 68, 72, 74, 68, 76, 69, 73, 74, 77, 72, 
    54, 37, 56, 64, 66, 64, 69, 68, 67, 72, 37, 71, 75, 75, 71, 
    53, 33, 51, 60, 62, 60, 63, 46, 49, 56, 22, 52, 67, 63, 66, 
    45, 31, 50, 50, 55, 53, 51, 53, 27, 0, 0, 0, 7, 44, 37, 
    0, 0, 0, 3, 9, 13, 15, 19, 8, 7, 0, 1, 12, 32, 10, 
    0, 0, 9, 0, 16, 12, 21, 12, 2, 2, 1, 39, 46, 14, 12, 
    1, 0, 0, 0, 15, 26, 27, 23, 25, 24, 29, 40, 37, 17, 0, 
    15, 21, 29, 40, 43, 45, 45, 43, 34, 29, 6, 25, 34, 23, 12, 
    20, 9, 14, 36, 43, 33, 26, 23, 25, 31, 28, 34, 31, 29, 14, 
    11, 20, 30, 29, 23, 30, 34, 30, 13, 28, 34, 34, 16, 1, 0, 
    13, 25, 27, 20, 13, 14, 28, 0, 0, 15, 11, 0, 0, 0, 0, 
    0, 16, 19, 0, 0, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=148
    0, 0, 8, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 45, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 31, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 
    18, 4, 0, 6, 9, 1, 1, 0, 0, 0, 23, 18, 0, 29, 0, 
    11, 0, 0, 18, 13, 0, 0, 0, 0, 4, 27, 0, 0, 0, 0, 
    0, 0, 6, 13, 3, 0, 0, 0, 0, 0, 6, 3, 0, 0, 7, 
    0, 0, 16, 3, 0, 0, 0, 0, 2, 0, 19, 0, 0, 0, 0, 
    0, 19, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 1, 0, 0, 19, 3, 0, 0, 0, 0, 0, 
    39, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 1, 2, 2, 2, 0, 0, 0, 23, 0, 0, 0, 0, 2, 0, 
    
    -- channel=149
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 12, 0, 9, 5, 0, 3, 0, 3, 0, 0, 58, 0, 31, 
    0, 0, 1, 0, 0, 9, 9, 22, 26, 16, 0, 0, 12, 0, 28, 
    3, 13, 1, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 68, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 14, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 18, 5, 2, 0, 0, 0, 0, 0, 0, 2, 10, 5, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 13, 5, 11, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 24, 3, 5, 9, 6, 8, 
    8, 4, 7, 6, 5, 5, 2, 7, 0, 33, 4, 7, 5, 2, 25, 
    
    -- channel=150
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 41, 35, 1, 29, 0, 0, 0, 
    32, 27, 21, 16, 26, 21, 15, 20, 1, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 62, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 0, 15, 0, 
    0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 25, 37, 17, 
    0, 0, 0, 8, 6, 0, 7, 23, 0, 0, 25, 27, 18, 14, 19, 
    0, 0, 7, 0, 0, 0, 26, 12, 0, 0, 14, 14, 5, 11, 17, 
    0, 19, 32, 19, 19, 14, 0, 0, 15, 14, 2, 1, 23, 5, 3, 
    21, 19, 9, 0, 5, 10, 5, 5, 0, 9, 8, 8, 7, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 14, 0, 30, 5, 7, 2, 0, 33, 
    
    -- channel=151
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 27, 14, 0, 0, 
    1, 12, 0, 15, 4, 7, 0, 0, 0, 0, 0, 0, 4, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 3, 
    10, 10, 2, 3, 0, 3, 2, 0, 0, 0, 1, 2, 3, 5, 0, 
    6, 10, 5, 3, 0, 0, 0, 0, 28, 0, 6, 6, 7, 8, 0, 
    
    -- channel=152
    56, 49, 72, 76, 82, 80, 85, 83, 84, 90, 84, 88, 83, 88, 85, 
    59, 50, 75, 75, 82, 77, 84, 84, 83, 81, 63, 88, 85, 90, 86, 
    61, 47, 72, 71, 80, 72, 75, 72, 74, 56, 55, 79, 80, 83, 84, 
    59, 46, 75, 75, 77, 73, 67, 59, 42, 14, 15, 27, 56, 72, 71, 
    25, 19, 22, 33, 38, 43, 40, 34, 12, 10, 5, 3, 26, 40, 29, 
    0, 0, 8, 0, 11, 9, 20, 14, 8, 5, 7, 38, 30, 37, 7, 
    10, 4, 1, 10, 27, 23, 24, 15, 15, 19, 39, 59, 41, 36, 0, 
    12, 13, 19, 33, 43, 47, 47, 47, 47, 40, 33, 44, 43, 1, 0, 
    29, 26, 32, 48, 53, 47, 40, 31, 35, 25, 30, 39, 38, 34, 38, 
    7, 20, 35, 39, 32, 35, 42, 44, 32, 40, 43, 44, 32, 15, 3, 
    24, 30, 34, 30, 37, 36, 32, 3, 8, 36, 29, 13, 0, 0, 0, 
    23, 28, 21, 0, 0, 29, 26, 5, 4, 5, 0, 0, 0, 0, 0, 
    14, 21, 14, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=153
    9, 0, 8, 0, 1, 0, 0, 4, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 22, 8, 0, 0, 
    19, 14, 16, 13, 35, 17, 15, 0, 3, 17, 35, 66, 23, 15, 0, 
    6, 0, 0, 2, 0, 15, 20, 34, 45, 35, 18, 0, 4, 0, 0, 
    27, 43, 61, 55, 33, 23, 17, 1, 0, 0, 0, 0, 0, 18, 64, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 33, 36, 8, 0, 0, 0, 
    6, 33, 20, 0, 0, 14, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 5, 0, 0, 0, 5, 3, 
    1, 5, 4, 4, 8, 11, 3, 0, 0, 0, 0, 0, 2, 5, 0, 
    
    -- channel=154
    53, 42, 57, 50, 49, 40, 38, 38, 37, 36, 23, 33, 34, 39, 35, 
    41, 28, 41, 33, 35, 25, 24, 29, 31, 10, 0, 30, 26, 30, 27, 
    29, 13, 26, 23, 24, 17, 18, 1, 4, 0, 1, 5, 11, 15, 19, 
    2, 0, 0, 0, 0, 3, 8, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 21, 8, 0, 0, 
    20, 17, 13, 13, 38, 29, 28, 20, 14, 19, 38, 57, 18, 10, 0, 
    23, 1, 2, 16, 29, 39, 55, 58, 64, 57, 38, 6, 6, 0, 0, 
    46, 51, 66, 71, 62, 56, 53, 38, 24, 0, 0, 0, 2, 4, 46, 
    22, 1, 20, 38, 35, 20, 19, 26, 32, 35, 38, 17, 10, 2, 0, 
    40, 56, 47, 28, 33, 46, 36, 7, 0, 17, 18, 4, 0, 0, 0, 
    31, 43, 32, 12, 0, 8, 12, 0, 1, 0, 0, 0, 0, 0, 0, 
    26, 23, 20, 10, 25, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=155
    59, 51, 51, 53, 48, 46, 41, 42, 38, 39, 41, 37, 41, 38, 38, 
    54, 43, 43, 44, 39, 38, 34, 35, 37, 40, 31, 32, 39, 35, 34, 
    46, 38, 33, 36, 30, 33, 30, 31, 31, 49, 17, 32, 35, 29, 28, 
    33, 25, 17, 18, 20, 21, 29, 24, 36, 41, 31, 27, 11, 18, 18, 
    23, 20, 21, 13, 14, 14, 23, 35, 37, 35, 34, 24, 17, 17, 9, 
    26, 26, 30, 28, 27, 32, 35, 44, 36, 35, 30, 21, 23, 6, 30, 
    34, 32, 35, 29, 39, 47, 49, 50, 45, 41, 24, 23, 27, 15, 25, 
    44, 39, 36, 42, 47, 51, 54, 51, 45, 41, 22, 15, 22, 33, 11, 
    44, 45, 43, 49, 53, 54, 54, 49, 38, 38, 20, 24, 27, 23, 21, 
    54, 37, 46, 51, 52, 48, 43, 40, 38, 35, 32, 29, 28, 26, 19, 
    47, 53, 49, 46, 40, 43, 46, 42, 26, 28, 33, 33, 25, 24, 15, 
    37, 49, 51, 44, 38, 29, 40, 32, 29, 30, 28, 30, 22, 19, 16, 
    31, 38, 40, 33, 33, 33, 28, 26, 26, 27, 23, 21, 22, 16, 15, 
    22, 23, 23, 21, 21, 22, 24, 24, 20, 26, 19, 16, 17, 15, 13, 
    12, 12, 16, 17, 19, 19, 21, 18, 12, 30, 13, 14, 14, 14, 12, 
    
    -- channel=156
    13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 7, 0, 2, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    10, 7, 0, 2, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 
    2, 4, 0, 0, 0, 0, 0, 7, 11, 9, 10, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 15, 19, 15, 18, 7, 9, 1, 
    14, 18, 22, 18, 13, 18, 9, 18, 20, 23, 16, 8, 38, 0, 32, 
    12, 23, 18, 9, 4, 20, 18, 27, 29, 22, 6, 0, 6, 3, 38, 
    19, 21, 12, 12, 8, 10, 12, 15, 4, 17, 0, 0, 1, 41, 27, 
    8, 7, 0, 0, 5, 6, 13, 17, 11, 22, 8, 6, 5, 11, 0, 
    28, 8, 7, 10, 14, 16, 12, 9, 5, 4, 4, 5, 8, 13, 11, 
    7, 14, 12, 11, 0, 1, 20, 26, 13, 0, 7, 15, 20, 24, 19, 
    0, 14, 24, 24, 21, 0, 10, 21, 20, 18, 22, 26, 26, 26, 28, 
    3, 9, 11, 16, 18, 17, 19, 22, 21, 22, 28, 24, 28, 26, 28, 
    22, 21, 25, 23, 24, 23, 24, 27, 23, 34, 25, 26, 28, 27, 27, 
    27, 28, 30, 29, 29, 30, 29, 27, 13, 38, 23, 26, 27, 25, 30, 
    
    -- channel=157
    6, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 4, 0, 11, 2, 6, 0, 0, 3, 2, 16, 0, 0, 0, 
    9, 0, 0, 2, 0, 2, 11, 10, 20, 17, 5, 0, 0, 0, 0, 
    9, 12, 18, 24, 14, 10, 7, 2, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 16, 15, 0, 0, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 2, 0, 1, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=158
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=159
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=160
    10, 0, 11, 0, 1, 0, 0, 9, 0, 0, 0, 0, 0, 7, 0, 
    5, 0, 0, 0, 10, 0, 4, 15, 0, 8, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 14, 0, 23, 0, 0, 7, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 
    21, 0, 10, 0, 36, 0, 10, 0, 0, 7, 0, 30, 6, 80, 0, 
    10, 0, 0, 0, 7, 3, 16, 3, 19, 22, 0, 0, 4, 0, 0, 
    0, 12, 20, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 0, 
    0, 17, 5, 0, 0, 3, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 13, 0, 0, 4, 0, 0, 0, 0, 2, 
    22, 0, 17, 0, 7, 13, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 
    1, 0, 3, 2, 3, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    
    -- channel=161
    68, 35, 74, 76, 82, 75, 85, 90, 82, 89, 83, 86, 79, 91, 78, 
    70, 35, 75, 73, 87, 72, 83, 90, 79, 89, 43, 83, 79, 94, 74, 
    72, 29, 69, 71, 88, 69, 85, 71, 65, 76, 35, 77, 79, 88, 76, 
    64, 18, 65, 64, 78, 67, 77, 60, 33, 16, 0, 2, 51, 76, 58, 
    19, 2, 18, 23, 29, 31, 28, 44, 12, 17, 7, 0, 18, 45, 5, 
    0, 0, 17, 0, 16, 8, 20, 21, 12, 13, 0, 47, 32, 64, 4, 
    12, 0, 0, 0, 22, 21, 27, 18, 19, 28, 31, 54, 58, 27, 0, 
    13, 14, 21, 30, 44, 48, 52, 48, 52, 49, 27, 37, 37, 2, 1, 
    25, 26, 17, 44, 52, 50, 45, 39, 35, 40, 28, 35, 36, 30, 47, 
    4, 17, 38, 38, 32, 40, 47, 47, 30, 44, 40, 46, 34, 17, 0, 
    25, 32, 35, 35, 36, 36, 43, 2, 0, 42, 32, 19, 3, 0, 0, 
    23, 27, 32, 0, 0, 26, 39, 7, 1, 9, 5, 0, 0, 0, 0, 
    12, 22, 24, 4, 4, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=162
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    21, 5, 0, 20, 33, 15, 0, 0, 0, 6, 31, 29, 0, 15, 0, 
    0, 0, 0, 9, 13, 25, 29, 41, 47, 33, 9, 0, 3, 0, 0, 
    13, 26, 32, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 32, 84, 
    0, 0, 0, 0, 0, 0, 0, 11, 8, 17, 13, 0, 0, 0, 0, 
    30, 22, 0, 0, 11, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 2, 0, 
    0, 3, 6, 9, 9, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    
    -- channel=163
    25, 26, 27, 29, 26, 25, 25, 22, 24, 27, 29, 23, 22, 22, 20, 
    27, 27, 28, 29, 26, 26, 29, 24, 24, 41, 31, 22, 24, 25, 22, 
    26, 27, 27, 22, 26, 23, 27, 37, 37, 33, 42, 39, 31, 27, 26, 
    28, 25, 33, 25, 24, 22, 20, 28, 50, 30, 34, 61, 54, 40, 37, 
    43, 41, 37, 46, 42, 46, 40, 38, 24, 24, 23, 0, 14, 16, 38, 
    5, 12, 15, 2, 0, 9, 20, 24, 21, 15, 0, 0, 5, 2, 13, 
    20, 22, 17, 16, 18, 10, 8, 0, 0, 3, 14, 24, 3, 31, 24, 
    7, 0, 0, 1, 12, 19, 24, 33, 35, 41, 31, 19, 13, 0, 0, 
    38, 38, 30, 29, 39, 45, 41, 25, 20, 0, 1, 12, 16, 20, 25, 
    5, 10, 23, 33, 24, 21, 28, 44, 39, 23, 20, 28, 41, 37, 29, 
    27, 26, 33, 39, 50, 37, 35, 24, 27, 43, 45, 36, 33, 23, 26, 
    32, 32, 31, 21, 11, 33, 39, 27, 26, 28, 37, 25, 19, 20, 11, 
    39, 49, 45, 39, 40, 35, 22, 26, 35, 27, 22, 23, 17, 12, 7, 
    30, 29, 25, 24, 27, 29, 25, 22, 8, 18, 15, 14, 11, 9, 11, 
    10, 9, 11, 11, 11, 14, 20, 20, 22, 16, 12, 9, 11, 9, 14, 
    
    -- channel=164
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 6, 0, 42, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 2, 
    2, 6, 5, 4, 3, 0, 0, 0, 16, 0, 3, 0, 1, 4, 0, 
    
    -- channel=165
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 18, 0, 0, 
    3, 20, 5, 0, 26, 19, 5, 0, 0, 1, 35, 70, 34, 0, 1, 
    3, 0, 0, 0, 0, 0, 15, 28, 49, 40, 33, 0, 0, 0, 0, 
    24, 38, 63, 66, 31, 18, 9, 0, 0, 0, 0, 0, 0, 0, 63, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 44, 2, 0, 0, 0, 
    0, 41, 18, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=166
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 51, 30, 0, 6, 
    10, 7, 13, 28, 18, 18, 1, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 4, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 9, 1, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    
    -- channel=167
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 47, 10, 0, 0, 0, 
    0, 1, 3, 4, 0, 0, 0, 0, 0, 0, 8, 22, 60, 1, 16, 
    13, 14, 11, 30, 20, 22, 11, 0, 0, 0, 0, 0, 10, 0, 11, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 10, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 6, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    3, 0, 0, 0, 5, 7, 0, 0, 16, 1, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    5, 6, 1, 4, 0, 1, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 30, 0, 1, 0, 0, 3, 0, 
    
    -- channel=168
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 9, 0, 74, 0, 0, 4, 0, 0, 
    18, 0, 0, 0, 8, 0, 9, 0, 64, 72, 20, 59, 13, 17, 11, 
    52, 36, 46, 38, 53, 47, 40, 49, 5, 0, 0, 0, 0, 18, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 11, 61, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 6, 0, 0, 17, 0, 
    0, 20, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 3, 6, 0, 0, 5, 33, 51, 26, 
    0, 0, 0, 7, 9, 0, 23, 34, 0, 2, 37, 44, 25, 15, 16, 
    0, 0, 17, 4, 0, 0, 29, 2, 0, 8, 17, 19, 5, 6, 11, 
    0, 16, 33, 10, 22, 25, 4, 0, 12, 18, 2, 0, 17, 0, 0, 
    19, 18, 7, 0, 0, 6, 6, 6, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 25, 0, 0, 0, 0, 23, 
    
    -- channel=169
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=170
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 20, 4, 0, 0, 0, 0, 0, 0, 0, 58, 0, 0, 0, 2, 
    0, 32, 12, 0, 0, 0, 0, 35, 37, 0, 69, 42, 0, 0, 10, 
    0, 33, 21, 25, 6, 8, 0, 0, 35, 42, 44, 105, 111, 27, 62, 
    67, 65, 57, 77, 70, 75, 62, 22, 7, 0, 15, 0, 12, 0, 54, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 8, 17, 9, 0, 0, 0, 0, 0, 0, 10, 0, 27, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 51, 22, 0, 0, 0, 
    11, 36, 39, 10, 6, 21, 18, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 7, 3, 0, 0, 8, 44, 0, 0, 0, 27, 32, 42, 
    12, 0, 0, 12, 43, 37, 0, 19, 40, 28, 38, 30, 19, 17, 11, 
    32, 13, 0, 14, 0, 18, 15, 7, 16, 16, 20, 18, 3, 11, 7, 
    40, 40, 38, 31, 40, 44, 19, 8, 25, 24, 7, 18, 7, 9, 1, 
    40, 45, 27, 24, 19, 24, 23, 13, 9, 0, 12, 9, 7, 3, 0, 
    6, 7, 3, 3, 0, 0, 4, 7, 44, 0, 8, 8, 6, 6, 1, 
    
    -- channel=171
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 
    4, 3, 11, 0, 27, 16, 1, 0, 0, 7, 12, 40, 63, 0, 15, 
    0, 0, 0, 0, 0, 16, 22, 37, 52, 38, 7, 0, 0, 0, 0, 
    18, 36, 41, 38, 15, 9, 4, 0, 0, 0, 0, 0, 0, 46, 78, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 21, 1, 0, 0, 0, 
    18, 16, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 2, 5, 
    0, 1, 3, 4, 5, 6, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    
    -- channel=172
    0, 28, 18, 3, 1, 0, 1, 0, 11, 0, 0, 4, 0, 0, 9, 
    0, 21, 16, 0, 0, 0, 0, 0, 6, 0, 8, 11, 0, 0, 8, 
    0, 15, 15, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 8, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 38, 0, 0, 
    26, 26, 0, 25, 31, 20, 13, 0, 0, 0, 58, 58, 0, 11, 0, 
    14, 0, 0, 35, 15, 6, 17, 21, 36, 29, 51, 1, 0, 0, 0, 
    20, 26, 47, 53, 28, 16, 5, 0, 0, 0, 0, 1, 0, 0, 44, 
    0, 0, 10, 5, 0, 0, 0, 0, 13, 0, 47, 11, 0, 0, 0, 
    0, 43, 21, 0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 3, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 11, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 1, 0, 
    0, 5, 4, 6, 6, 6, 0, 0, 26, 0, 0, 0, 0, 4, 0, 
    
    -- channel=173
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 11, 0, 0, 
    0, 4, 16, 0, 9, 3, 4, 0, 0, 5, 14, 44, 59, 0, 12, 
    0, 0, 0, 0, 0, 5, 3, 19, 28, 20, 14, 0, 0, 0, 10, 
    15, 28, 36, 41, 20, 12, 8, 10, 0, 0, 0, 0, 0, 34, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 24, 5, 0, 4, 0, 
    0, 10, 13, 0, 0, 3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    
    -- channel=174
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=175
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 
    13, 15, 0, 7, 29, 14, 0, 0, 0, 6, 46, 70, 17, 0, 0, 
    0, 0, 0, 0, 0, 7, 15, 33, 49, 37, 28, 0, 0, 0, 0, 
    22, 42, 62, 51, 26, 13, 6, 0, 0, 0, 0, 0, 0, 5, 78, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 38, 0, 0, 0, 0, 
    1, 37, 5, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=176
    0, 0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 4, 0, 4, 2, 
    0, 0, 0, 0, 2, 0, 3, 5, 2, 0, 0, 6, 2, 7, 2, 
    0, 0, 2, 5, 12, 4, 10, 3, 0, 0, 0, 0, 1, 12, 6, 
    0, 0, 7, 9, 18, 13, 14, 3, 0, 0, 0, 0, 1, 7, 8, 
    0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 6, 19, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 17, 13, 37, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 20, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 10, 8, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 5, 3, 3, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 4, 
    5, 4, 2, 1, 0, 0, 0, 0, 0, 0, 4, 3, 1, 2, 10, 
    
    -- channel=177
    0, 26, 17, 3, 2, 2, 2, 0, 12, 0, 0, 3, 0, 0, 7, 
    0, 22, 23, 0, 3, 0, 0, 0, 8, 0, 36, 14, 0, 0, 9, 
    0, 21, 25, 0, 0, 0, 0, 11, 20, 0, 69, 30, 0, 0, 14, 
    0, 16, 9, 10, 0, 2, 0, 0, 0, 0, 12, 14, 55, 3, 25, 
    0, 3, 0, 19, 1, 8, 1, 0, 0, 0, 7, 13, 39, 0, 1, 
    19, 17, 0, 21, 1, 0, 1, 0, 0, 0, 45, 22, 0, 22, 0, 
    14, 0, 0, 31, 18, 0, 0, 0, 0, 0, 38, 12, 0, 1, 0, 
    3, 0, 9, 17, 9, 2, 0, 0, 0, 0, 26, 14, 0, 0, 0, 
    0, 1, 31, 12, 0, 0, 0, 0, 9, 0, 23, 1, 0, 0, 5, 
    0, 20, 14, 0, 1, 1, 0, 0, 11, 3, 1, 0, 0, 0, 0, 
    21, 1, 0, 0, 10, 21, 0, 0, 36, 7, 0, 0, 0, 0, 0, 
    48, 1, 0, 0, 3, 34, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 1, 0, 8, 2, 2, 2, 0, 19, 0, 0, 0, 0, 1, 0, 
    0, 4, 3, 4, 2, 2, 0, 0, 40, 0, 0, 0, 0, 6, 0, 
    
    -- channel=178
    0, 0, 0, 0, 0, 1, 8, 9, 9, 11, 14, 16, 12, 12, 15, 
    0, 0, 0, 3, 8, 10, 12, 14, 13, 4, 15, 18, 16, 16, 16, 
    1, 3, 11, 16, 19, 18, 16, 15, 16, 3, 10, 18, 18, 23, 21, 
    13, 14, 23, 31, 33, 28, 26, 15, 0, 0, 0, 0, 27, 28, 33, 
    7, 6, 6, 12, 19, 18, 11, 3, 0, 0, 0, 7, 11, 14, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 9, 36, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 30, 17, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 23, 20, 13, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 9, 9, 14, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 6, 7, 6, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 
    4, 2, 0, 0, 0, 0, 0, 1, 1, 0, 1, 1, 0, 0, 5, 
    
    -- channel=179
    70, 68, 88, 91, 96, 97, 104, 102, 105, 108, 105, 111, 105, 108, 108, 
    75, 73, 94, 93, 101, 96, 101, 105, 105, 91, 92, 111, 105, 110, 107, 
    79, 72, 95, 95, 104, 96, 95, 93, 98, 66, 82, 104, 100, 106, 107, 
    76, 66, 87, 93, 98, 95, 94, 78, 52, 38, 32, 39, 86, 92, 93, 
    44, 40, 46, 55, 60, 64, 63, 55, 36, 33, 31, 39, 54, 57, 52, 
    26, 35, 33, 34, 46, 42, 43, 36, 34, 35, 45, 75, 48, 80, 35, 
    31, 27, 25, 34, 49, 47, 47, 43, 45, 49, 66, 81, 76, 56, 16, 
    37, 41, 50, 54, 62, 65, 66, 60, 64, 51, 59, 74, 70, 36, 39, 
    39, 39, 47, 62, 62, 59, 57, 57, 62, 58, 63, 66, 64, 58, 65, 
    28, 45, 52, 49, 52, 58, 62, 58, 58, 66, 66, 62, 51, 37, 30, 
    44, 47, 47, 44, 46, 57, 46, 26, 36, 57, 48, 37, 27, 18, 14, 
    42, 45, 35, 24, 29, 48, 44, 29, 29, 32, 26, 17, 12, 6, 1, 
    33, 33, 30, 22, 21, 23, 23, 22, 19, 16, 12, 11, 6, 1, 0, 
    4, 6, 6, 9, 13, 12, 11, 10, 18, 10, 6, 3, 1, 1, 0, 
    0, 1, 2, 4, 7, 8, 8, 5, 17, 4, 2, 0, 0, 2, 0, 
    
    -- channel=180
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 19, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 7, 0, 
    5, 0, 0, 7, 4, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 2, 7, 7, 12, 15, 17, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 45, 
    0, 0, 4, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 16, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 
    0, 0, 0, 0, 0, 9, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 9, 3, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 
    0, 2, 5, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=181
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 133, 0, 0, 4, 0, 0, 
    29, 0, 0, 0, 0, 0, 11, 2, 53, 80, 0, 2, 0, 0, 0, 
    27, 5, 16, 0, 13, 0, 6, 50, 23, 3, 0, 0, 0, 19, 0, 
    0, 0, 7, 0, 0, 0, 0, 16, 0, 0, 0, 0, 35, 0, 53, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 0, 116, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 0, 0, 84, 0, 
    0, 8, 0, 0, 0, 2, 4, 0, 0, 15, 0, 0, 0, 1, 0, 
    3, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 9, 32, 58, 15, 
    0, 0, 0, 15, 0, 0, 43, 52, 0, 0, 30, 53, 35, 27, 17, 
    0, 0, 39, 12, 0, 0, 50, 18, 0, 7, 25, 27, 17, 12, 28, 
    0, 10, 44, 10, 13, 16, 9, 0, 10, 19, 18, 0, 36, 2, 2, 
    12, 14, 9, 0, 0, 3, 2, 14, 0, 21, 9, 3, 9, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 19, 0, 67, 0, 3, 0, 0, 44, 
    
    -- channel=182
    0, 0, 0, 0, 0, 0, 2, 4, 5, 5, 7, 10, 6, 7, 8, 
    0, 0, 0, 0, 3, 4, 8, 10, 8, 1, 9, 13, 9, 12, 11, 
    0, 0, 5, 8, 14, 12, 11, 11, 11, 0, 4, 12, 11, 17, 15, 
    5, 3, 14, 21, 24, 21, 19, 9, 0, 0, 0, 0, 17, 21, 24, 
    2, 0, 5, 10, 15, 15, 10, 0, 0, 0, 0, 0, 6, 13, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 2, 28, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 20, 14, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 14, 2, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 4, 4, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=183
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 25, 47, 0, 0, 0, 
    0, 1, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 5, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    
    -- channel=184
    36, 44, 40, 34, 28, 24, 18, 11, 17, 13, 17, 12, 10, 10, 13, 
    25, 33, 29, 19, 17, 13, 10, 14, 13, 6, 21, 11, 7, 7, 11, 
    17, 26, 19, 7, 3, 6, 0, 15, 17, 3, 26, 30, 6, 4, 10, 
    15, 17, 9, 10, 0, 2, 0, 0, 22, 14, 24, 11, 27, 9, 11, 
    24, 25, 12, 15, 10, 15, 20, 19, 29, 31, 38, 10, 16, 0, 0, 
    24, 20, 19, 23, 14, 13, 32, 33, 32, 24, 25, 8, 0, 0, 0, 
    34, 26, 23, 39, 30, 32, 30, 30, 20, 16, 15, 6, 0, 0, 10, 
    36, 26, 31, 39, 41, 40, 39, 37, 40, 21, 22, 3, 1, 0, 0, 
    41, 54, 44, 48, 47, 52, 43, 27, 18, 10, 7, 5, 10, 3, 9, 
    32, 36, 50, 43, 40, 30, 29, 30, 43, 23, 16, 11, 21, 14, 14, 
    59, 45, 40, 43, 48, 51, 24, 21, 20, 26, 30, 19, 16, 17, 12, 
    49, 44, 34, 31, 29, 28, 33, 35, 28, 17, 20, 27, 9, 17, 8, 
    44, 46, 44, 44, 38, 27, 20, 22, 28, 25, 13, 21, 17, 14, 14, 
    23, 23, 22, 23, 23, 25, 23, 16, 21, 12, 18, 14, 15, 14, 10, 
    11, 12, 12, 12, 13, 16, 18, 13, 27, 12, 15, 13, 14, 16, 4, 
    
    -- channel=185
    29, 28, 38, 34, 35, 30, 30, 26, 30, 31, 22, 27, 25, 30, 27, 
    23, 22, 31, 26, 27, 23, 26, 24, 26, 21, 10, 28, 23, 27, 26, 
    17, 14, 24, 17, 22, 16, 19, 13, 15, 1, 20, 18, 16, 18, 23, 
    9, 10, 18, 10, 10, 13, 6, 15, 2, 0, 5, 0, 0, 8, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 1, 12, 4, 0, 
    6, 4, 5, 0, 15, 12, 20, 8, 6, 4, 12, 26, 13, 1, 0, 
    16, 3, 0, 15, 18, 17, 24, 19, 24, 22, 27, 14, 0, 2, 0, 
    20, 19, 28, 40, 35, 32, 29, 27, 19, 8, 0, 4, 5, 0, 7, 
    22, 9, 19, 29, 29, 21, 14, 9, 16, 6, 22, 14, 9, 6, 0, 
    11, 30, 32, 23, 16, 23, 23, 15, 2, 12, 15, 11, 0, 0, 0, 
    19, 24, 23, 13, 15, 10, 11, 0, 5, 10, 0, 0, 0, 0, 0, 
    23, 15, 12, 0, 7, 25, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=186
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=187
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 68, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 7, 0, 0, 27, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 9, 0, 0, 0, 0, 13, 0, 
    0, 0, 9, 0, 0, 0, 0, 5, 0, 2, 0, 0, 21, 3, 10, 
    0, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 45, 0, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 60, 9, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 30, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 17, 13, 0, 0, 0, 11, 5, 6, 0, 
    0, 0, 19, 0, 0, 0, 16, 6, 0, 0, 0, 9, 2, 0, 11, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 2, 3, 0, 15, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 2, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 3, 0, 29, 0, 0, 0, 0, 17, 
    
    -- channel=188
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 41, 47, 52, 0, 0, 0, 
    0, 4, 18, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 
    2, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 6, 0, 2, 1, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 22, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=189
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 72, 0, 0, 2, 0, 0, 
    12, 0, 0, 0, 0, 0, 3, 5, 24, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 4, 2, 0, 0, 0, 12, 0, 
    0, 0, 10, 0, 0, 0, 0, 8, 0, 0, 0, 0, 48, 0, 40, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 2, 59, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 62, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 1, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 19, 0, 
    0, 0, 0, 3, 0, 0, 23, 22, 0, 0, 4, 14, 9, 6, 5, 
    0, 0, 21, 1, 0, 0, 15, 7, 0, 0, 4, 6, 4, 2, 10, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 1, 0, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 35, 0, 0, 0, 0, 24, 
    
    -- channel=190
    17, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 0, 20, 0, 
    0, 0, 18, 0, 11, 0, 0, 1, 0, 9, 0, 19, 72, 0, 14, 
    0, 0, 0, 0, 0, 13, 9, 26, 30, 20, 0, 0, 22, 0, 35, 
    6, 25, 18, 11, 2, 1, 1, 2, 0, 7, 0, 0, 0, 70, 57, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 3, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 1, 0, 5, 
    2, 0, 0, 0, 0, 1, 0, 1, 0, 23, 0, 0, 0, 0, 11, 
    
    -- channel=191
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    1, 0, 0, 5, 2, 0, 0, 0, 21, 29, 0, 29, 9, 4, 13, 
    27, 21, 21, 20, 32, 28, 20, 11, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 8, 44, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 22, 14, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 8, 12, 5, 1, 3, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 4, 0, 0, 2, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 10, 
    
    -- channel=192
    1, 3, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 15, 1, 0, 0, 19, 15, 10, 12, 13, 13, 6, 1, 1, 0, 
    10, 12, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 
    0, 9, 4, 1, 9, 14, 11, 7, 9, 9, 6, 4, 0, 3, 4, 
    0, 5, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 
    0, 0, 0, 60, 57, 17, 2, 0, 0, 0, 1, 1, 4, 8, 8, 
    0, 0, 0, 0, 0, 59, 38, 6, 2, 2, 0, 0, 0, 1, 3, 
    0, 0, 0, 0, 0, 4, 46, 74, 53, 25, 13, 0, 2, 4, 4, 
    0, 0, 0, 0, 9, 18, 4, 0, 14, 61, 94, 79, 51, 21, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    44, 53, 59, 63, 68, 44, 24, 40, 55, 30, 36, 22, 37, 52, 47, 
    0, 0, 0, 0, 0, 0, 0, 14, 23, 29, 34, 39, 43, 44, 48, 
    21, 31, 28, 20, 15, 14, 12, 9, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    
    -- channel=193
    23, 35, 25, 17, 16, 23, 22, 15, 16, 16, 20, 18, 15, 26, 29, 
    27, 34, 38, 7, 13, 22, 21, 17, 23, 26, 24, 10, 36, 33, 30, 
    25, 35, 45, 0, 17, 6, 1, 2, 10, 16, 13, 7, 29, 34, 33, 
    24, 34, 37, 0, 2, 0, 0, 0, 0, 6, 2, 17, 0, 35, 33, 
    33, 33, 33, 36, 23, 21, 19, 20, 26, 25, 20, 19, 29, 34, 33, 
    39, 37, 35, 43, 26, 26, 26, 30, 29, 29, 27, 29, 34, 32, 30, 
    36, 33, 5, 0, 35, 44, 33, 35, 34, 35, 33, 36, 36, 36, 34, 
    37, 38, 36, 25, 0, 7, 40, 40, 34, 35, 31, 34, 34, 33, 32, 
    38, 38, 36, 38, 19, 0, 0, 11, 40, 46, 35, 34, 33, 34, 33, 
    38, 35, 36, 44, 37, 0, 0, 0, 0, 0, 0, 30, 45, 44, 35, 
    36, 33, 34, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 19, 
    42, 47, 48, 48, 46, 51, 37, 35, 42, 38, 36, 38, 37, 36, 35, 
    1, 5, 4, 4, 2, 3, 3, 5, 16, 12, 15, 13, 16, 20, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    
    -- channel=194
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 31, 29, 22, 26, 24, 25, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 73, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 72, 36, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 46, 101, 81, 28, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 20, 4, 0, 5, 63, 112, 121, 76, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    72, 84, 93, 99, 104, 83, 50, 46, 61, 30, 36, 19, 25, 40, 38, 
    0, 0, 0, 0, 0, 0, 0, 17, 33, 42, 48, 55, 60, 62, 64, 
    25, 33, 29, 20, 17, 14, 11, 9, 5, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 
    
    -- channel=195
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    
    -- channel=196
    72, 77, 56, 55, 62, 63, 58, 59, 58, 59, 60, 59, 65, 69, 65, 
    75, 75, 68, 36, 54, 42, 35, 43, 41, 43, 41, 46, 70, 67, 67, 
    70, 73, 69, 41, 55, 68, 55, 64, 68, 71, 67, 68, 69, 68, 70, 
    70, 74, 58, 55, 60, 59, 55, 66, 59, 53, 58, 62, 70, 67, 69, 
    69, 73, 69, 63, 62, 60, 59, 64, 63, 57, 60, 74, 75, 69, 70, 
    67, 68, 57, 69, 71, 72, 74, 74, 71, 69, 70, 72, 69, 68, 70, 
    69, 52, 34, 45, 60, 67, 72, 72, 70, 67, 69, 68, 68, 68, 70, 
    73, 69, 60, 34, 33, 58, 64, 66, 67, 66, 67, 67, 69, 68, 72, 
    71, 67, 64, 59, 3, 27, 31, 44, 51, 57, 68, 69, 68, 67, 70, 
    69, 66, 66, 59, 0, 18, 24, 24, 21, 21, 39, 42, 51, 60, 69, 
    73, 67, 66, 47, 46, 28, 38, 65, 52, 32, 45, 34, 74, 67, 69, 
    58, 51, 46, 45, 45, 40, 50, 61, 59, 59, 64, 65, 68, 69, 67, 
    39, 44, 43, 38, 34, 34, 39, 44, 36, 35, 34, 35, 35, 32, 28, 
    12, 18, 16, 13, 8, 13, 15, 13, 11, 9, 11, 12, 12, 11, 29, 
    7, 14, 15, 15, 11, 18, 15, 14, 12, 12, 11, 8, 14, 35, 6, 
    
    -- channel=197
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 23, 23, 0, 4, 15, 18, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=198
    0, 21, 34, 14, 5, 19, 19, 13, 18, 14, 16, 15, 13, 18, 15, 
    0, 7, 29, 28, 0, 0, 0, 0, 0, 0, 0, 0, 12, 13, 12, 
    0, 7, 20, 22, 44, 36, 37, 27, 42, 45, 38, 25, 2, 15, 13, 
    6, 10, 38, 37, 20, 21, 31, 23, 17, 27, 15, 30, 0, 10, 7, 
    21, 11, 22, 32, 11, 6, 8, 10, 9, 15, 8, 1, 24, 14, 12, 
    18, 11, 0, 30, 38, 38, 35, 37, 40, 35, 31, 19, 15, 16, 14, 
    11, 47, 33, 0, 0, 8, 17, 20, 22, 22, 15, 17, 14, 11, 7, 
    5, 20, 50, 109, 0, 0, 0, 13, 15, 17, 15, 18, 18, 19, 13, 
    4, 13, 16, 31, 83, 0, 0, 0, 0, 0, 6, 21, 16, 13, 12, 
    3, 10, 13, 16, 61, 0, 0, 5, 0, 0, 0, 0, 0, 0, 13, 
    0, 14, 11, 53, 89, 114, 44, 25, 87, 68, 77, 54, 9, 19, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    3, 18, 22, 19, 15, 15, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    3, 2, 4, 0, 3, 9, 13, 7, 12, 11, 6, 1, 4, 7, 0, 
    
    -- channel=199
    18, 25, 29, 17, 14, 15, 15, 15, 16, 15, 15, 15, 14, 14, 18, 
    26, 34, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 17, 17, 
    25, 35, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 18, 
    27, 34, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 23, 
    28, 33, 33, 26, 19, 19, 22, 19, 20, 20, 16, 17, 18, 26, 26, 
    24, 35, 33, 22, 30, 26, 25, 24, 25, 27, 24, 24, 25, 23, 25, 
    19, 26, 26, 29, 12, 16, 24, 25, 25, 26, 24, 25, 25, 24, 23, 
    17, 26, 24, 12, 28, 15, 5, 16, 21, 20, 21, 23, 24, 25, 27, 
    16, 20, 20, 19, 30, 4, 6, 12, 8, 12, 15, 22, 25, 25, 27, 
    11, 15, 17, 23, 24, 7, 0, 0, 3, 13, 15, 12, 8, 12, 21, 
    12, 16, 19, 14, 12, 17, 9, 3, 7, 22, 5, 15, 7, 14, 20, 
    15, 17, 16, 16, 16, 22, 18, 11, 23, 20, 24, 22, 23, 26, 23, 
    14, 17, 20, 18, 17, 19, 19, 21, 24, 24, 23, 24, 25, 23, 21, 
    10, 8, 9, 7, 6, 6, 7, 6, 7, 6, 6, 6, 6, 4, 17, 
    6, 7, 6, 5, 4, 5, 7, 3, 6, 7, 8, 6, 3, 29, 23, 
    
    -- channel=200
    7, 22, 31, 12, 8, 16, 16, 10, 13, 12, 14, 13, 7, 9, 9, 
    12, 25, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 10, 10, 
    14, 26, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 12, 
    19, 25, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 15, 
    26, 25, 26, 28, 16, 14, 15, 12, 15, 16, 10, 2, 16, 18, 18, 
    20, 23, 14, 24, 26, 24, 21, 22, 24, 24, 19, 18, 20, 18, 17, 
    13, 40, 35, 0, 0, 13, 18, 19, 19, 20, 16, 19, 17, 17, 15, 
    9, 21, 24, 47, 1, 0, 0, 12, 17, 17, 15, 17, 19, 20, 20, 
    7, 11, 13, 14, 51, 0, 0, 0, 0, 2, 9, 19, 19, 18, 19, 
    5, 7, 11, 20, 44, 0, 0, 0, 0, 0, 0, 0, 0, 1, 14, 
    2, 11, 10, 31, 26, 50, 16, 0, 26, 19, 24, 20, 0, 6, 8, 
    0, 0, 0, 0, 0, 4, 0, 0, 11, 17, 11, 17, 17, 18, 16, 
    0, 10, 12, 7, 4, 5, 4, 0, 7, 2, 3, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 4, 
    
    -- channel=201
    0, 0, 19, 12, 4, 9, 14, 8, 11, 10, 11, 12, 3, 5, 7, 
    0, 0, 8, 55, 33, 35, 45, 34, 42, 37, 36, 20, 6, 10, 8, 
    0, 0, 14, 41, 45, 31, 45, 31, 31, 36, 33, 21, 9, 6, 5, 
    0, 0, 27, 43, 30, 31, 32, 32, 32, 46, 34, 33, 8, 6, 3, 
    2, 0, 3, 26, 10, 8, 8, 10, 12, 17, 11, 0, 10, 4, 4, 
    3, 7, 5, 1, 4, 0, 1, 7, 8, 4, 2, 0, 6, 7, 3, 
    0, 23, 31, 13, 0, 0, 6, 9, 9, 11, 7, 8, 7, 7, 5, 
    0, 7, 17, 37, 21, 0, 0, 8, 14, 13, 8, 8, 7, 7, 3, 
    0, 6, 10, 22, 80, 3, 0, 1, 0, 8, 1, 11, 10, 7, 4, 
    0, 9, 10, 31, 92, 8, 3, 7, 8, 22, 0, 4, 0, 0, 5, 
    0, 10, 10, 39, 20, 37, 2, 0, 8, 20, 0, 9, 0, 0, 4, 
    1, 17, 18, 17, 15, 28, 5, 0, 18, 7, 8, 6, 6, 12, 8, 
    4, 10, 12, 9, 7, 8, 4, 3, 15, 11, 12, 10, 12, 17, 14, 
    18, 15, 17, 11, 14, 11, 8, 7, 10, 9, 5, 6, 6, 0, 0, 
    16, 9, 8, 5, 7, 3, 8, 2, 8, 6, 6, 6, 0, 0, 3, 
    
    -- channel=202
    18, 6, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    21, 18, 0, 0, 7, 28, 15, 21, 19, 22, 23, 29, 15, 7, 5, 
    23, 12, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 7, 7, 
    12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 8, 10, 
    0, 8, 0, 0, 0, 0, 0, 0, 2, 0, 0, 18, 0, 5, 7, 
    5, 5, 26, 6, 0, 0, 0, 0, 0, 0, 0, 3, 5, 1, 3, 
    9, 0, 0, 37, 80, 32, 5, 1, 0, 0, 6, 5, 8, 9, 12, 
    18, 1, 0, 0, 0, 79, 75, 16, 1, 0, 2, 1, 2, 0, 4, 
    22, 8, 3, 0, 0, 0, 33, 75, 79, 44, 25, 0, 0, 4, 5, 
    21, 8, 4, 0, 0, 0, 0, 0, 0, 9, 73, 88, 81, 44, 11, 
    22, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    70, 62, 63, 66, 72, 40, 46, 62, 41, 22, 38, 23, 33, 32, 35, 
    0, 0, 0, 0, 0, 0, 0, 16, 9, 20, 21, 28, 31, 27, 30, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    
    -- channel=203
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 13, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 33, 55, 61, 18, 38, 53, 43, 32, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 7, 11, 12, 11, 16, 20, 19, 20, 28, 51, 
    11, 21, 21, 21, 20, 33, 26, 29, 23, 28, 22, 22, 43, 32, 0, 
    
    -- channel=204
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 20, 16, 28, 17, 18, 25, 19, 22, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 2, 2, 5, 32, 
    4, 1, 1, 4, 3, 8, 6, 9, 7, 9, 6, 7, 14, 31, 0, 
    
    -- channel=205
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 8, 0, 0, 1, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 11, 0, 0, 1, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 4, 4, 6, 10, 7, 7, 7, 8, 8, 8, 8, 7, 6, 0, 
    7, 7, 7, 8, 9, 6, 11, 10, 12, 12, 13, 10, 0, 1, 7, 
    
    -- channel=206
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 27, 24, 18, 22, 22, 19, 5, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 51, 66, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 64, 42, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 32, 88, 79, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 22, 17, 12, 0, 1, 45, 92, 111, 77, 23, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    68, 82, 90, 95, 98, 86, 58, 51, 63, 44, 43, 34, 31, 45, 44, 
    0, 0, 0, 0, 0, 0, 2, 16, 29, 36, 40, 44, 49, 50, 48, 
    15, 25, 23, 16, 14, 11, 10, 7, 6, 2, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    
    -- channel=207
    30, 2, 0, 0, 11, 0, 0, 1, 0, 0, 0, 0, 8, 0, 0, 
    30, 9, 0, 0, 16, 7, 0, 11, 0, 2, 0, 12, 14, 0, 0, 
    28, 6, 0, 0, 0, 1, 0, 10, 0, 0, 0, 3, 19, 0, 0, 
    19, 7, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 35, 0, 0, 
    5, 7, 0, 0, 0, 0, 1, 0, 0, 0, 1, 23, 0, 0, 0, 
    6, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 13, 41, 16, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 58, 41, 4, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 14, 35, 38, 24, 5, 13, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 1, 15, 6, 8, 5, 47, 26, 24, 12, 2, 
    26, 0, 0, 0, 0, 0, 11, 65, 0, 0, 0, 0, 65, 13, 10, 
    13, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 5, 4, 0, 3, 
    0, 5, 1, 6, 0, 1, 3, 5, 0, 0, 2, 0, 0, 6, 40, 
    0, 0, 0, 2, 0, 11, 0, 7, 0, 0, 0, 0, 21, 21, 0, 
    
    -- channel=208
    21, 20, 11, 3, 1, 3, 0, 1, 3, 0, 0, 0, 7, 13, 9, 
    25, 20, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 1, 4, 
    21, 20, 12, 0, 0, 8, 0, 1, 10, 14, 14, 16, 4, 7, 7, 
    24, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 
    23, 21, 17, 8, 5, 1, 2, 3, 4, 0, 1, 9, 19, 11, 11, 
    17, 18, 4, 18, 34, 36, 34, 30, 31, 32, 29, 26, 8, 8, 11, 
    12, 5, 0, 0, 0, 5, 10, 11, 12, 12, 11, 10, 9, 5, 4, 
    12, 11, 16, 40, 8, 0, 0, 1, 2, 2, 7, 9, 11, 10, 13, 
    10, 5, 3, 0, 0, 0, 0, 0, 0, 0, 3, 9, 8, 7, 10, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    4, 0, 1, 0, 34, 56, 27, 46, 59, 37, 59, 32, 46, 24, 3, 
    0, 0, 0, 0, 0, 0, 7, 2, 0, 0, 1, 9, 5, 0, 0, 
    13, 14, 20, 20, 21, 21, 25, 16, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    0, 0, 1, 1, 0, 7, 8, 7, 5, 7, 7, 1, 12, 45, 0, 
    
    -- channel=209
    0, 2, 14, 9, 0, 6, 13, 3, 7, 6, 10, 9, 0, 10, 11, 
    0, 0, 10, 26, 11, 12, 21, 13, 20, 18, 20, 0, 5, 9, 11, 
    0, 3, 14, 10, 14, 1, 10, 0, 3, 14, 7, 5, 1, 11, 10, 
    0, 0, 17, 0, 0, 0, 2, 0, 0, 12, 0, 5, 0, 9, 8, 
    7, 2, 4, 24, 4, 3, 0, 3, 7, 9, 5, 0, 8, 9, 7, 
    12, 21, 8, 0, 6, 2, 1, 6, 7, 6, 4, 4, 8, 9, 7, 
    9, 20, 29, 5, 0, 0, 6, 10, 11, 15, 9, 12, 11, 11, 8, 
    7, 15, 21, 40, 10, 0, 0, 9, 16, 14, 10, 11, 10, 10, 6, 
    9, 17, 18, 24, 74, 0, 0, 0, 0, 9, 0, 11, 13, 11, 8, 
    12, 17, 17, 47, 75, 0, 0, 0, 0, 7, 0, 4, 0, 0, 6, 
    8, 13, 15, 36, 0, 23, 0, 0, 5, 0, 0, 0, 0, 0, 3, 
    12, 22, 23, 23, 17, 28, 6, 0, 13, 5, 3, 2, 1, 1, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    
    -- channel=210
    0, 0, 17, 0, 0, 6, 8, 4, 9, 5, 6, 5, 7, 10, 5, 
    0, 0, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 37, 33, 33, 27, 43, 42, 34, 22, 0, 0, 0, 
    0, 0, 24, 38, 12, 12, 31, 19, 11, 18, 6, 18, 0, 0, 0, 
    0, 0, 2, 10, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 5, 21, 21, 19, 21, 22, 16, 15, 2, 0, 0, 0, 
    0, 28, 18, 0, 0, 0, 0, 2, 4, 3, 0, 0, 0, 0, 0, 
    0, 4, 31, 92, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 2, 13, 54, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 31, 88, 104, 38, 30, 78, 63, 70, 50, 10, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=211
    41, 57, 54, 44, 48, 52, 52, 48, 51, 51, 53, 52, 53, 64, 63, 
    41, 52, 56, 47, 45, 48, 48, 48, 51, 52, 51, 43, 65, 62, 64, 
    38, 51, 54, 54, 53, 54, 48, 54, 57, 60, 57, 60, 57, 63, 63, 
    43, 49, 56, 54, 50, 48, 49, 50, 54, 53, 49, 53, 52, 58, 62, 
    51, 51, 53, 57, 42, 41, 40, 47, 48, 43, 41, 45, 63, 60, 61, 
    53, 55, 41, 50, 59, 57, 60, 63, 62, 57, 56, 61, 58, 59, 61, 
    54, 56, 39, 8, 17, 50, 62, 65, 64, 63, 60, 61, 59, 60, 60, 
    55, 65, 58, 57, 15, 2, 32, 60, 64, 61, 59, 60, 60, 60, 60, 
    57, 64, 65, 60, 43, 0, 0, 0, 19, 43, 53, 65, 63, 59, 59, 
    56, 63, 65, 68, 22, 0, 0, 0, 0, 0, 0, 0, 19, 42, 60, 
    54, 64, 64, 59, 43, 42, 2, 9, 45, 19, 22, 14, 21, 49, 54, 
    25, 32, 28, 25, 22, 17, 17, 27, 32, 34, 33, 36, 39, 39, 38, 
    9, 14, 14, 8, 6, 2, 2, 4, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=212
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 11, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 38, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 7, 21, 17, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 6, 0, 0, 0, 19, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 14, 56, 0, 0, 5, 0, 63, 15, 1, 
    9, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 
    0, 0, 0, 0, 0, 5, 0, 2, 0, 0, 0, 0, 9, 28, 0, 
    
    -- channel=213
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 8, 0, 0, 5, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 27, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 85, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 27, 60, 122, 55, 0, 56, 73, 57, 67, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 1, 1, 5, 0, 
    13, 5, 5, 3, 8, 7, 15, 8, 17, 16, 11, 7, 0, 0, 3, 
    
    -- channel=214
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 35, 0, 19, 26, 11, 21, 13, 20, 4, 0, 0, 0, 
    0, 0, 0, 32, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 58, 0, 4, 21, 20, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 103, 16, 0, 0, 2, 33, 33, 41, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 43, 47, 49, 52, 52, 25, 13, 30, 17, 12, 6, 9, 16, 14, 
    0, 0, 0, 0, 0, 0, 0, 5, 24, 25, 31, 30, 34, 42, 44, 
    21, 21, 20, 13, 14, 10, 7, 5, 3, 4, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 
    
    -- channel=215
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 35, 29, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 20, 15, 5, 12, 20, 53, 21, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 6, 5, 2, 12, 
    12, 13, 8, 12, 6, 10, 9, 10, 1, 5, 8, 6, 8, 9, 0, 
    4, 6, 4, 7, 4, 3, 0, 1, 0, 0, 0, 1, 9, 0, 0, 
    
    -- channel=216
    51, 59, 48, 50, 56, 54, 53, 51, 52, 54, 56, 54, 56, 67, 68, 
    53, 63, 62, 58, 80, 86, 81, 82, 85, 86, 83, 75, 79, 72, 73, 
    53, 61, 65, 55, 48, 45, 42, 50, 43, 47, 48, 54, 75, 72, 73, 
    54, 60, 60, 48, 56, 54, 45, 52, 62, 60, 61, 59, 66, 72, 73, 
    57, 60, 57, 53, 46, 46, 46, 51, 54, 46, 47, 56, 64, 69, 70, 
    63, 65, 58, 56, 56, 54, 59, 61, 59, 57, 57, 66, 67, 67, 69, 
    66, 48, 30, 46, 61, 68, 71, 73, 72, 71, 71, 70, 70, 71, 72, 
    70, 71, 55, 22, 16, 48, 67, 74, 73, 69, 68, 68, 68, 67, 68, 
    74, 76, 75, 66, 11, 0, 21, 50, 63, 68, 69, 72, 71, 69, 69, 
    74, 76, 76, 78, 7, 0, 0, 0, 3, 12, 31, 54, 61, 66, 71, 
    72, 74, 75, 55, 15, 0, 0, 5, 19, 0, 0, 0, 26, 52, 66, 
    63, 67, 64, 62, 61, 45, 40, 54, 58, 48, 53, 49, 56, 58, 59, 
    15, 18, 15, 11, 9, 7, 9, 19, 20, 19, 19, 21, 23, 23, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=217
    12, 11, 5, 0, 0, 2, 1, 1, 5, 1, 1, 0, 8, 12, 8, 
    6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 15, 25, 13, 19, 31, 30, 30, 18, 0, 0, 0, 
    6, 1, 0, 2, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 1, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 
    13, 0, 0, 17, 30, 31, 29, 27, 28, 27, 26, 10, 0, 0, 1, 
    11, 14, 0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 
    8, 4, 32, 83, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    7, 1, 0, 10, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 13, 79, 99, 51, 67, 100, 68, 95, 60, 51, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 2, 6, 8, 8, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 45, 
    0, 0, 1, 1, 2, 14, 13, 14, 15, 15, 8, 6, 27, 42, 0, 
    
    -- channel=218
    29, 48, 39, 26, 26, 34, 32, 32, 34, 33, 33, 31, 38, 41, 36, 
    35, 43, 42, 1, 0, 0, 0, 0, 0, 0, 0, 0, 27, 31, 33, 
    32, 41, 33, 0, 14, 15, 5, 11, 23, 26, 20, 15, 22, 35, 34, 
    36, 43, 32, 0, 8, 15, 11, 11, 6, 3, 3, 13, 17, 31, 33, 
    42, 43, 44, 35, 22, 19, 23, 27, 22, 21, 22, 34, 40, 39, 37, 
    40, 34, 10, 41, 57, 54, 55, 54, 53, 52, 50, 44, 38, 38, 41, 
    36, 47, 26, 0, 0, 21, 41, 43, 42, 39, 37, 35, 35, 32, 31, 
    37, 45, 53, 55, 0, 0, 0, 28, 34, 32, 35, 36, 39, 39, 40, 
    37, 37, 35, 40, 0, 0, 0, 0, 0, 0, 24, 41, 38, 35, 36, 
    32, 31, 32, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 32, 
    29, 35, 34, 39, 69, 69, 49, 64, 74, 58, 67, 54, 59, 46, 34, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 
    0, 6, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 
    
    -- channel=219
    27, 42, 44, 31, 29, 34, 33, 32, 33, 33, 32, 33, 31, 31, 35, 
    33, 47, 46, 24, 0, 6, 7, 4, 5, 5, 11, 16, 27, 37, 37, 
    34, 48, 42, 14, 1, 0, 0, 0, 0, 0, 0, 0, 24, 38, 39, 
    35, 46, 41, 0, 6, 10, 7, 0, 6, 8, 4, 6, 10, 39, 42, 
    38, 45, 48, 39, 31, 32, 34, 32, 32, 35, 29, 32, 33, 43, 43, 
    36, 43, 45, 41, 41, 40, 38, 39, 39, 40, 39, 38, 43, 42, 42, 
    34, 51, 38, 24, 24, 38, 42, 42, 42, 42, 41, 42, 42, 42, 41, 
    33, 44, 43, 32, 21, 14, 25, 38, 40, 40, 39, 41, 41, 43, 43, 
    31, 40, 41, 41, 39, 4, 8, 13, 20, 29, 37, 41, 41, 42, 44, 
    27, 36, 38, 35, 44, 5, 1, 2, 7, 16, 13, 16, 23, 32, 39, 
    28, 38, 39, 45, 29, 27, 15, 6, 20, 31, 16, 23, 8, 28, 34, 
    20, 29, 28, 27, 27, 31, 23, 22, 35, 30, 33, 32, 35, 38, 36, 
    15, 21, 20, 18, 15, 16, 17, 18, 22, 21, 22, 21, 22, 22, 22, 
    12, 11, 11, 9, 8, 8, 7, 7, 7, 7, 5, 4, 5, 8, 11, 
    6, 6, 5, 3, 4, 4, 5, 4, 6, 6, 4, 4, 9, 13, 27, 
    
    -- channel=220
    0, 0, 14, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 3, 0, 0, 1, 2, 0, 0, 0, 0, 0, 
    0, 18, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 42, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 56, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 46, 11, 6, 10, 13, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 28, 59, 30, 3, 27, 45, 33, 40, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 5, 8, 9, 12, 12, 8, 1, 4, 2, 2, 0, 0, 0, 3, 
    18, 10, 12, 16, 20, 18, 17, 19, 21, 25, 23, 22, 22, 26, 31, 
    28, 22, 21, 21, 24, 22, 25, 24, 28, 28, 27, 28, 31, 30, 34, 
    
    -- channel=221
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 13, 10, 24, 4, 24, 13, 16, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 3, 
    
    -- channel=222
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 2, 0, 3, 4, 3, 1, 2, 0, 2, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=223
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=224
    16, 10, 0, 0, 0, 4, 6, 0, 0, 0, 5, 0, 0, 2, 0, 
    15, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    9, 0, 0, 0, 0, 4, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    9, 2, 7, 0, 0, 0, 0, 2, 0, 5, 13, 26, 0, 0, 0, 
    19, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 13, 2, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    22, 3, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 3, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 17, 12, 32, 41, 31, 48, 0, 52, 18, 47, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 1, 0, 0, 9, 4, 2, 4, 4, 0, 0, 0, 26, 0, 
    
    -- channel=225
    42, 60, 46, 44, 42, 50, 49, 44, 44, 46, 49, 47, 47, 62, 64, 
    46, 61, 61, 35, 45, 51, 51, 46, 53, 55, 55, 42, 64, 65, 65, 
    47, 57, 67, 30, 39, 26, 22, 25, 31, 39, 37, 32, 63, 67, 65, 
    46, 56, 57, 4, 23, 26, 20, 19, 24, 29, 28, 40, 26, 65, 63, 
    54, 56, 57, 56, 41, 39, 38, 42, 47, 44, 43, 46, 57, 64, 63, 
    66, 65, 55, 59, 56, 51, 54, 58, 56, 58, 56, 57, 63, 62, 62, 
    65, 49, 26, 29, 48, 60, 63, 67, 66, 66, 64, 65, 64, 65, 63, 
    69, 70, 70, 37, 0, 30, 59, 67, 65, 63, 62, 63, 63, 62, 60, 
    74, 73, 73, 74, 18, 0, 0, 33, 55, 61, 57, 63, 65, 64, 61, 
    73, 70, 70, 77, 23, 0, 0, 0, 0, 0, 6, 45, 56, 60, 61, 
    66, 68, 70, 71, 16, 0, 0, 0, 25, 0, 0, 0, 13, 37, 55, 
    56, 61, 58, 56, 53, 52, 39, 38, 46, 36, 43, 39, 40, 39, 44, 
    5, 12, 12, 12, 11, 8, 7, 11, 18, 16, 16, 16, 19, 20, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 17, 
    
    -- channel=226
    4, 0, 6, 2, 6, 11, 14, 17, 16, 17, 15, 14, 18, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 30, 19, 17, 16, 17, 20, 18, 22, 24, 19, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    2, 0, 0, 4, 8, 8, 5, 3, 3, 2, 2, 0, 0, 0, 0, 
    4, 28, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 16, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 95, 79, 93, 98, 68, 75, 90, 85, 68, 20, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 46, 
    1, 1, 3, 1, 4, 20, 15, 18, 19, 20, 6, 0, 30, 20, 0, 
    
    -- channel=227
    18, 13, 10, 11, 9, 8, 8, 6, 5, 6, 8, 8, 5, 10, 15, 
    23, 27, 17, 0, 5, 14, 13, 11, 11, 14, 13, 9, 14, 17, 17, 
    24, 28, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 20, 19, 
    21, 24, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 23, 
    17, 24, 18, 12, 15, 18, 15, 12, 18, 13, 12, 12, 8, 21, 21, 
    19, 33, 42, 10, 5, 4, 3, 3, 3, 8, 7, 16, 20, 17, 18, 
    19, 1, 8, 55, 53, 23, 15, 16, 15, 18, 19, 21, 22, 24, 23, 
    22, 19, 1, 0, 19, 53, 40, 19, 18, 17, 17, 18, 18, 18, 20, 
    23, 21, 20, 8, 3, 11, 39, 66, 59, 37, 18, 14, 18, 22, 22, 
    21, 20, 20, 34, 16, 14, 9, 2, 15, 40, 68, 77, 59, 32, 18, 
    21, 16, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    61, 63, 68, 70, 71, 57, 46, 44, 47, 38, 37, 30, 32, 37, 38, 
    14, 6, 7, 11, 15, 14, 15, 24, 32, 36, 38, 42, 44, 43, 43, 
    23, 22, 22, 18, 18, 15, 15, 15, 13, 12, 11, 10, 9, 4, 0, 
    6, 5, 4, 6, 5, 0, 0, 0, 0, 0, 5, 8, 0, 19, 46, 
    
    -- channel=228
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 11, 12, 9, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 5, 12, 6, 4, 0, 7, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 6, 26, 0, 0, 2, 0, 33, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 2, 3, 4, 4, 2, 6, 6, 6, 6, 19, 
    0, 2, 5, 7, 4, 9, 4, 9, 5, 5, 4, 6, 11, 18, 0, 
    
    -- channel=229
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 5, 12, 17, 11, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 24, 23, 18, 20, 20, 18, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 73, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 69, 118, 64, 83, 109, 81, 107, 78, 73, 31, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 
    0, 0, 0, 0, 0, 3, 11, 10, 10, 13, 8, 1, 11, 49, 0, 
    
    -- channel=230
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 9, 4, 6, 4, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 45, 53, 16, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 6, 0, 13, 41, 67, 43, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 5, 10, 15, 18, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 10, 11, 9, 13, 
    13, 17, 12, 12, 11, 11, 8, 8, 2, 2, 3, 2, 2, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    
    -- channel=231
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 22, 18, 8, 18, 11, 12, 9, 15, 0, 0, 0, 
    4, 0, 0, 0, 0, 4, 0, 12, 0, 0, 0, 1, 8, 0, 0, 
    0, 0, 0, 0, 1, 4, 0, 10, 4, 0, 9, 0, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 47, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 60, 39, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 35, 51, 40, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 18, 7, 7, 13, 60, 52, 40, 9, 0, 
    1, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 15, 0, 0, 
    29, 15, 15, 19, 25, 0, 13, 31, 7, 0, 8, 0, 5, 6, 7, 
    0, 0, 0, 0, 0, 0, 0, 12, 2, 11, 11, 18, 19, 14, 19, 
    0, 11, 5, 8, 0, 4, 6, 6, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    
    -- channel=232
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 30, 0, 15, 26, 8, 17, 12, 16, 2, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 36, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 52, 0, 16, 44, 32, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 111, 12, 0, 0, 6, 56, 55, 61, 29, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 50, 59, 62, 64, 62, 15, 9, 43, 18, 13, 5, 10, 26, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 17, 24, 24, 29, 37, 40, 
    30, 29, 29, 18, 21, 16, 10, 8, 7, 5, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    
    -- channel=233
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=234
    5, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 2, 0, 0, 29, 52, 43, 48, 41, 42, 44, 54, 0, 0, 0, 
    11, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 1, 
    0, 0, 0, 0, 0, 6, 3, 0, 4, 0, 0, 11, 0, 0, 0, 
    0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 89, 107, 18, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 109, 76, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 72, 127, 104, 43, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 22, 6, 22, 69, 147, 136, 98, 37, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    83, 78, 85, 92, 102, 69, 48, 60, 62, 37, 40, 26, 30, 49, 50, 
    7, 0, 0, 0, 0, 1, 7, 30, 36, 51, 54, 65, 70, 67, 77, 
    40, 47, 40, 36, 25, 27, 25, 25, 14, 10, 12, 8, 8, 7, 0, 
    5, 4, 2, 3, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    
    -- channel=235
    0, 0, 15, 0, 0, 0, 3, 0, 7, 2, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 6, 11, 7, 2, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 17, 14, 12, 15, 13, 10, 0, 0, 0, 0, 
    0, 25, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 102, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 90, 150, 80, 53, 102, 97, 105, 95, 36, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 
    4, 0, 0, 0, 0, 12, 18, 13, 19, 20, 11, 4, 10, 31, 0, 
    
    -- channel=236
    35, 13, 0, 0, 15, 5, 2, 10, 10, 10, 7, 5, 20, 17, 9, 
    30, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 3, 
    24, 7, 0, 0, 0, 25, 5, 29, 24, 18, 20, 24, 15, 0, 4, 
    22, 9, 0, 6, 11, 8, 5, 19, 6, 0, 6, 5, 38, 0, 1, 
    12, 10, 0, 0, 0, 0, 0, 2, 0, 0, 3, 23, 11, 1, 2, 
    10, 0, 0, 2, 18, 19, 22, 15, 12, 14, 17, 18, 0, 1, 8, 
    16, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 
    21, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 
    19, 2, 0, 0, 0, 5, 1, 0, 0, 0, 2, 0, 0, 0, 1, 
    18, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 2, 
    23, 0, 0, 0, 28, 32, 63, 107, 59, 38, 75, 56, 102, 46, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 50, 
    0, 0, 0, 2, 0, 15, 8, 16, 9, 10, 3, 0, 31, 38, 0, 
    
    -- channel=237
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 5, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 17, 13, 26, 6, 21, 26, 20, 27, 0, 0, 0, 
    0, 0, 7, 17, 0, 0, 5, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 21, 23, 20, 18, 21, 19, 17, 10, 0, 0, 0, 
    0, 13, 16, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 13, 95, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 53, 110, 28, 13, 80, 58, 72, 47, 9, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 8, 8, 10, 10, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 3, 9, 5, 8, 9, 7, 2, 0, 13, 3, 
    
    -- channel=238
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=239
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 16, 0, 11, 17, 17, 15, 8, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 23, 24, 22, 17, 18, 18, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 79, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 96, 104, 66, 96, 105, 81, 110, 74, 72, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 
    0, 0, 0, 0, 0, 10, 10, 12, 10, 14, 4, 0, 19, 47, 0, 
    
    -- channel=240
    0, 0, 0, 8, 2, 4, 7, 6, 6, 7, 7, 5, 4, 4, 1, 
    0, 0, 0, 32, 43, 28, 30, 30, 30, 27, 25, 21, 1, 0, 0, 
    0, 0, 0, 29, 36, 39, 42, 42, 34, 37, 31, 23, 8, 0, 0, 
    0, 0, 7, 43, 36, 32, 32, 39, 34, 40, 43, 39, 24, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 15, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 6, 3, 17, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 0, 0, 0, 14, 15, 18, 15, 9, 0, 0, 0, 0, 0, 
    4, 1, 1, 12, 25, 27, 34, 34, 27, 22, 29, 28, 26, 11, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 5, 3, 4, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 14, 14, 13, 15, 14, 15, 16, 15, 15, 15, 15, 14, 14, 8, 
    14, 16, 16, 16, 17, 20, 21, 21, 20, 20, 17, 16, 12, 1, 0, 
    
    -- channel=241
    28, 8, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 9, 4, 2, 
    28, 12, 0, 0, 7, 8, 0, 11, 0, 0, 3, 21, 7, 0, 1, 
    26, 8, 0, 0, 0, 4, 0, 15, 1, 0, 0, 6, 24, 0, 2, 
    17, 9, 0, 0, 0, 3, 0, 3, 0, 0, 3, 0, 29, 0, 2, 
    1, 8, 0, 0, 0, 0, 0, 2, 0, 0, 3, 26, 0, 0, 0, 
    4, 0, 0, 5, 0, 0, 2, 0, 0, 0, 0, 6, 0, 0, 2, 
    10, 0, 0, 20, 42, 16, 2, 0, 0, 0, 0, 0, 0, 0, 1, 
    19, 0, 0, 0, 0, 61, 45, 5, 0, 0, 0, 0, 0, 0, 0, 
    21, 2, 0, 0, 0, 12, 35, 38, 30, 10, 16, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 5, 13, 6, 7, 0, 43, 27, 30, 18, 4, 
    23, 0, 0, 0, 0, 0, 0, 55, 0, 0, 0, 0, 57, 17, 10, 
    24, 0, 0, 0, 5, 0, 5, 28, 0, 0, 7, 0, 6, 0, 1, 
    1, 0, 0, 0, 0, 0, 4, 16, 0, 4, 3, 9, 8, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 1, 0, 0, 6, 27, 
    0, 0, 0, 1, 0, 6, 0, 5, 0, 0, 0, 0, 20, 13, 0, 
    
    -- channel=242
    1, 0, 0, 6, 3, 3, 4, 5, 4, 3, 5, 5, 8, 9, 7, 
    0, 0, 0, 26, 35, 34, 34, 35, 35, 33, 31, 29, 5, 5, 5, 
    0, 0, 0, 39, 35, 37, 45, 40, 36, 36, 30, 28, 13, 4, 3, 
    0, 0, 8, 37, 31, 23, 28, 31, 25, 31, 35, 28, 17, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 11, 13, 0, 7, 14, 3, 0, 2, 1, 0, 0, 0, 0, 
    5, 5, 5, 11, 8, 14, 6, 13, 20, 11, 3, 0, 0, 0, 0, 
    8, 8, 6, 5, 11, 15, 20, 22, 11, 0, 2, 15, 18, 10, 0, 
    8, 5, 5, 7, 19, 1, 1, 17, 14, 5, 10, 1, 10, 1, 0, 
    13, 8, 10, 11, 9, 14, 11, 3, 0, 3, 0, 1, 0, 0, 0, 
    11, 7, 7, 10, 13, 11, 9, 3, 3, 4, 3, 2, 2, 3, 1, 
    12, 10, 11, 13, 16, 14, 14, 15, 17, 17, 18, 19, 17, 17, 8, 
    22, 17, 16, 18, 19, 17, 16, 20, 18, 18, 19, 21, 16, 5, 3, 
    
    -- channel=243
    75, 81, 67, 68, 75, 77, 76, 76, 75, 76, 78, 77, 83, 89, 91, 
    70, 80, 77, 59, 68, 73, 71, 73, 73, 76, 75, 80, 88, 90, 91, 
    71, 75, 73, 73, 72, 70, 63, 74, 74, 73, 74, 72, 88, 89, 91, 
    68, 74, 72, 64, 69, 69, 68, 66, 70, 68, 73, 75, 78, 87, 88, 
    71, 74, 78, 69, 66, 66, 67, 70, 71, 68, 70, 82, 81, 84, 85, 
    82, 75, 72, 79, 77, 76, 79, 81, 78, 78, 80, 80, 84, 84, 85, 
    86, 66, 46, 53, 75, 81, 84, 86, 86, 84, 84, 84, 84, 85, 86, 
    89, 88, 89, 55, 29, 59, 85, 88, 86, 84, 84, 84, 84, 83, 83, 
    92, 93, 93, 92, 27, 27, 35, 60, 76, 79, 83, 84, 84, 83, 83, 
    93, 92, 93, 84, 25, 18, 23, 27, 28, 25, 40, 64, 76, 82, 83, 
    91, 90, 92, 81, 62, 25, 25, 56, 58, 35, 40, 31, 64, 71, 81, 
    74, 72, 69, 68, 67, 62, 56, 61, 63, 60, 61, 62, 59, 60, 64, 
    40, 40, 38, 37, 37, 34, 32, 34, 33, 33, 31, 32, 34, 32, 32, 
    19, 21, 20, 21, 20, 16, 16, 18, 20, 15, 16, 17, 16, 19, 32, 
    16, 17, 17, 16, 16, 17, 18, 21, 20, 19, 17, 17, 24, 36, 26, 
    
    -- channel=244
    0, 0, 0, 0, 0, 0, 2, 3, 4, 6, 3, 1, 0, 0, 0, 
    0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 6, 7, 6, 3, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 29, 29, 59, 39, 7, 32, 31, 48, 23, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 11, 11, 10, 6, 7, 6, 6, 2, 1, 1, 0, 0, 4, 14, 
    0, 1, 0, 0, 1, 13, 9, 10, 12, 12, 1, 0, 8, 0, 0, 
    
    -- channel=245
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 42, 0, 0, 14, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 172, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 227, 0, 0, 0, 0, 18, 0, 4, 0, 0, 0, 
    0, 0, 0, 43, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 32, 32, 29, 69, 1, 0, 18, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 9, 16, 10, 15, 29, 21, 
    24, 12, 20, 9, 18, 7, 2, 0, 6, 7, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 
    
    -- channel=246
    3, 0, 0, 0, 2, 0, 1, 2, 1, 1, 1, 2, 4, 4, 4, 
    0, 0, 0, 11, 19, 19, 19, 22, 21, 20, 21, 21, 2, 0, 1, 
    0, 0, 0, 25, 29, 35, 37, 40, 34, 31, 28, 21, 13, 0, 0, 
    0, 0, 0, 23, 22, 17, 21, 21, 15, 19, 25, 20, 16, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 2, 1, 0, 3, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 1, 0, 5, 0, 7, 5, 8, 9, 3, 0, 0, 0, 0, 0, 
    9, 4, 2, 0, 0, 8, 12, 13, 8, 1, 0, 5, 8, 3, 0, 
    10, 0, 0, 2, 7, 0, 1, 13, 7, 2, 3, 1, 8, 1, 0, 
    10, 0, 2, 2, 2, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 4, 5, 7, 10, 9, 7, 8, 10, 9, 10, 10, 10, 10, 7, 
    14, 9, 9, 10, 11, 11, 9, 12, 11, 10, 10, 12, 11, 2, 0, 
    
    -- channel=247
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 31, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 21, 40, 26, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 19, 14, 16, 19, 16, 12, 13, 8, 11, 9, 7, 8, 7, 0, 
    7, 7, 5, 8, 8, 5, 7, 9, 11, 10, 9, 7, 0, 0, 23, 
    
    -- channel=248
    28, 32, 18, 9, 19, 15, 9, 10, 8, 9, 8, 9, 11, 13, 17, 
    33, 38, 26, 0, 0, 10, 3, 3, 3, 8, 8, 12, 27, 21, 20, 
    33, 36, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 22, 23, 
    29, 36, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 26, 
    25, 33, 31, 20, 22, 23, 22, 18, 23, 19, 16, 24, 22, 26, 28, 
    23, 25, 42, 36, 22, 24, 24, 23, 23, 24, 22, 27, 26, 23, 23, 
    22, 16, 0, 7, 52, 44, 26, 25, 24, 23, 25, 26, 27, 27, 28, 
    22, 23, 11, 0, 0, 32, 51, 29, 20, 21, 21, 23, 25, 25, 28, 
    19, 19, 19, 11, 0, 3, 11, 23, 44, 42, 36, 23, 23, 25, 28, 
    16, 15, 18, 6, 0, 2, 2, 1, 2, 4, 26, 37, 50, 44, 30, 
    19, 18, 18, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 15, 
    39, 42, 42, 42, 45, 38, 44, 52, 41, 42, 43, 42, 46, 43, 42, 
    13, 17, 16, 18, 16, 17, 23, 29, 29, 32, 34, 34, 37, 37, 34, 
    0, 4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 14, 
    
    -- channel=249
    25, 31, 22, 21, 22, 24, 21, 20, 22, 22, 23, 21, 24, 30, 27, 
    30, 31, 28, 13, 23, 13, 9, 16, 15, 15, 14, 13, 30, 26, 27, 
    28, 31, 31, 3, 14, 21, 15, 18, 20, 25, 22, 25, 28, 29, 29, 
    30, 31, 23, 13, 17, 19, 12, 22, 20, 15, 16, 20, 26, 28, 28, 
    31, 32, 25, 24, 20, 19, 18, 22, 22, 15, 19, 24, 33, 30, 30, 
    28, 30, 17, 23, 32, 31, 34, 33, 32, 30, 30, 36, 28, 28, 31, 
    28, 21, 14, 7, 6, 24, 31, 32, 31, 30, 29, 28, 29, 28, 28, 
    31, 31, 17, 14, 11, 9, 14, 26, 29, 26, 27, 28, 29, 29, 31, 
    31, 29, 27, 19, 0, 0, 0, 0, 0, 14, 24, 31, 30, 28, 29, 
    29, 27, 27, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 28, 
    29, 28, 28, 13, 9, 17, 10, 19, 25, 4, 19, 10, 31, 33, 29, 
    9, 7, 2, 0, 0, 0, 4, 17, 10, 11, 17, 15, 25, 21, 19, 
    3, 5, 6, 1, 0, 0, 2, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=250
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 30, 19, 36, 31, 19, 36, 21, 21, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=251
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 67, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 88, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 47, 37, 50, 0, 0, 16, 16, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    
    -- channel=252
    0, 0, 0, 0, 0, 0, 1, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 26, 9, 9, 12, 19, 20, 28, 21, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 37, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 8, 36, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 17, 60, 21, 0, 17, 13, 44, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 13, 9, 7, 7, 9, 5, 1, 0, 0, 0, 0, 0, 7, 2, 
    0, 0, 0, 0, 0, 3, 0, 0, 1, 0, 0, 0, 3, 0, 0, 
    
    -- channel=253
    0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 8, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 6, 0, 0, 4, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 59, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 120, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 127, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 31, 17, 65, 0, 0, 6, 29, 0, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    
    -- channel=254
    0, 0, 21, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 6, 0, 1, 7, 0, 0, 0, 0, 0, 
    0, 0, 22, 26, 0, 0, 14, 0, 0, 13, 0, 3, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 10, 4, 7, 11, 7, 4, 0, 0, 0, 0, 
    0, 36, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 79, 134, 44, 0, 78, 72, 72, 60, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    7, 0, 0, 0, 2, 7, 12, 5, 13, 12, 6, 4, 0, 2, 0, 
    
    -- channel=255
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 44, 30, 45, 47, 41, 46, 39, 39, 30, 0, 0, 0, 
    0, 0, 0, 46, 16, 3, 24, 11, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 30, 15, 10, 14, 16, 18, 31, 22, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 20, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 27, 0, 11, 31, 25, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 62, 14, 5, 2, 4, 31, 39, 41, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 27, 32, 34, 36, 35, 9, 3, 20, 11, 2, 1, 0, 11, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 16, 17, 20, 25, 28, 
    25, 23, 21, 15, 15, 14, 11, 8, 5, 4, 1, 0, 1, 0, 0, 
    11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=256
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 12, 0, 5, 0, 0, 0, 0, 12, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 9, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 14, 3, 3, 4, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 32, 0, 0, 0, 0, 0, 5, 19, 0, 0, 0, 0, 8, 1, 
    0, 48, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 27, 22, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    
    -- channel=257
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 24, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 24, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 36, 
    0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 4, 36, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 9, 25, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 9, 0, 0, 8, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 7, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 7, 3, 0, 1, 0, 0, 0, 0, 
    0, 10, 16, 0, 0, 0, 1, 8, 0, 3, 0, 0, 0, 0, 0, 
    4, 0, 7, 11, 0, 0, 0, 0, 0, 2, 2, 0, 3, 0, 0, 
    6, 0, 0, 2, 16, 0, 0, 0, 0, 3, 8, 0, 0, 0, 0, 
    
    -- channel=258
    0, 0, 0, 0, 5, 0, 0, 0, 9, 15, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 4, 10, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 16, 0, 9, 1, 0, 0, 0, 7, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 29, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 18, 
    8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 19, 12, 25, 0, 0, 0, 0, 0, 0, 0, 27, 26, 0, 
    0, 24, 7, 5, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    54, 53, 0, 0, 0, 0, 7, 48, 32, 0, 0, 0, 0, 13, 11, 
    0, 77, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 
    9, 0, 46, 42, 0, 0, 0, 0, 16, 25, 47, 0, 0, 0, 0, 
    
    -- channel=259
    0, 16, 1, 11, 29, 1, 14, 12, 15, 14, 20, 0, 25, 0, 5, 
    0, 18, 13, 7, 35, 7, 8, 6, 8, 13, 16, 0, 4, 0, 6, 
    19, 15, 6, 12, 33, 0, 8, 26, 5, 28, 0, 0, 0, 4, 3, 
    15, 0, 10, 9, 13, 2, 38, 33, 0, 13, 0, 6, 0, 0, 6, 
    26, 0, 5, 18, 0, 9, 22, 0, 5, 7, 18, 19, 0, 0, 23, 
    28, 0, 0, 16, 0, 0, 0, 0, 9, 7, 1, 3, 10, 0, 27, 
    20, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 
    0, 0, 8, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 
    4, 11, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 18, 0, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    10, 0, 3, 24, 18, 0, 0, 0, 0, 0, 0, 0, 0, 8, 28, 
    14, 24, 0, 0, 20, 23, 11, 0, 0, 0, 0, 0, 10, 12, 0, 
    25, 17, 10, 0, 0, 11, 22, 13, 14, 0, 0, 0, 5, 0, 0, 
    
    -- channel=260
    12, 0, 11, 4, 0, 9, 1, 1, 0, 0, 0, 14, 0, 5, 3, 
    8, 0, 1, 8, 0, 5, 0, 5, 0, 5, 0, 24, 0, 22, 6, 
    2, 0, 4, 3, 0, 5, 4, 0, 2, 0, 5, 24, 6, 6, 12, 
    0, 23, 8, 0, 0, 7, 0, 0, 17, 0, 14, 9, 9, 13, 3, 
    0, 35, 0, 2, 8, 1, 0, 8, 1, 3, 0, 0, 5, 18, 0, 
    0, 34, 15, 0, 13, 5, 5, 20, 0, 0, 0, 8, 0, 17, 0, 
    0, 25, 18, 10, 0, 5, 7, 11, 8, 15, 17, 12, 0, 13, 0, 
    0, 18, 16, 17, 22, 4, 20, 21, 13, 17, 19, 33, 12, 10, 0, 
    10, 16, 6, 6, 29, 16, 28, 23, 22, 21, 15, 23, 16, 3, 0, 
    18, 0, 0, 12, 6, 37, 23, 34, 29, 25, 19, 17, 4, 9, 15, 
    0, 11, 0, 16, 11, 2, 47, 30, 29, 25, 18, 16, 6, 9, 19, 
    15, 25, 0, 5, 2, 20, 30, 27, 28, 18, 29, 19, 0, 9, 0, 
    9, 15, 0, 0, 0, 22, 22, 10, 26, 24, 32, 11, 5, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 28, 30, 23, 12, 0, 12, 0, 
    0, 0, 8, 7, 3, 0, 0, 0, 0, 21, 18, 0, 0, 2, 27, 
    
    -- channel=261
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 2, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 0, 0, 12, 1, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 4, 18, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 20, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 0, 1, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 16, 0, 0, 
    
    -- channel=262
    15, 12, 0, 0, 21, 0, 1, 0, 0, 0, 6, 0, 45, 0, 0, 
    3, 1, 0, 0, 19, 0, 0, 0, 5, 0, 11, 0, 64, 0, 12, 
    0, 0, 0, 0, 14, 0, 2, 0, 0, 0, 0, 0, 35, 0, 10, 
    10, 0, 2, 15, 0, 0, 0, 0, 0, 33, 0, 0, 6, 0, 24, 
    7, 0, 48, 0, 0, 0, 23, 0, 2, 0, 0, 0, 0, 0, 47, 
    5, 0, 0, 61, 0, 0, 12, 9, 0, 0, 0, 0, 0, 0, 61, 
    26, 0, 0, 6, 0, 0, 17, 0, 0, 0, 11, 0, 0, 0, 50, 
    0, 0, 0, 0, 42, 0, 0, 1, 26, 23, 0, 0, 36, 0, 13, 
    1, 0, 0, 0, 0, 65, 0, 9, 6, 0, 0, 0, 0, 0, 37, 
    0, 0, 0, 0, 0, 0, 21, 15, 1, 17, 2, 5, 28, 2, 0, 
    7, 0, 8, 0, 0, 17, 0, 11, 17, 0, 3, 7, 13, 0, 0, 
    24, 38, 34, 0, 1, 0, 0, 0, 0, 19, 16, 4, 2, 0, 0, 
    0, 0, 16, 3, 0, 0, 0, 0, 0, 18, 0, 18, 14, 0, 0, 
    11, 0, 0, 0, 11, 0, 0, 25, 0, 0, 7, 1, 8, 0, 0, 
    14, 21, 0, 0, 0, 15, 0, 0, 0, 0, 0, 3, 34, 10, 0, 
    
    -- channel=263
    10, 15, 15, 24, 28, 6, 15, 11, 14, 6, 18, 0, 20, 0, 11, 
    16, 17, 21, 22, 26, 6, 8, 9, 10, 14, 17, 0, 12, 10, 18, 
    17, 1, 18, 24, 18, 4, 17, 26, 9, 22, 1, 1, 11, 17, 21, 
    19, 2, 24, 11, 11, 10, 23, 10, 13, 6, 5, 8, 9, 14, 25, 
    24, 5, 17, 22, 0, 10, 16, 6, 12, 10, 14, 1, 12, 17, 32, 
    21, 6, 18, 19, 14, 0, 3, 0, 8, 1, 4, 0, 16, 15, 28, 
    16, 11, 15, 15, 0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 26, 
    16, 10, 14, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 24, 
    12, 19, 22, 15, 4, 0, 0, 0, 0, 0, 0, 0, 1, 7, 12, 
    22, 14, 17, 9, 0, 1, 0, 0, 0, 0, 0, 0, 0, 7, 15, 
    20, 0, 23, 10, 28, 0, 0, 0, 0, 0, 0, 0, 0, 13, 19, 
    6, 0, 15, 24, 15, 15, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    10, 0, 0, 14, 17, 10, 0, 0, 0, 0, 0, 0, 0, 5, 27, 
    12, 9, 0, 0, 13, 11, 7, 2, 4, 0, 0, 0, 0, 9, 5, 
    22, 3, 6, 0, 0, 7, 13, 7, 6, 0, 0, 0, 8, 11, 0, 
    
    -- channel=264
    3, 0, 0, 3, 19, 0, 0, 0, 0, 0, 9, 0, 27, 0, 0, 
    0, 0, 0, 4, 13, 0, 0, 0, 0, 0, 6, 0, 24, 0, 7, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 3, 0, 0, 15, 0, 5, 
    10, 0, 0, 8, 0, 0, 0, 0, 0, 5, 0, 0, 2, 0, 29, 
    6, 0, 28, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 40, 
    4, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 15, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    12, 0, 2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 2, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=265
    2, 1, 0, 0, 25, 0, 0, 0, 0, 0, 16, 0, 66, 0, 0, 
    0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 17, 0, 57, 0, 2, 
    5, 0, 0, 0, 16, 0, 0, 0, 0, 15, 0, 0, 34, 0, 4, 
    11, 0, 9, 10, 0, 0, 1, 12, 0, 6, 0, 0, 18, 0, 48, 
    4, 0, 21, 13, 0, 0, 39, 0, 0, 0, 0, 0, 6, 0, 73, 
    20, 0, 0, 19, 0, 0, 22, 0, 0, 0, 11, 0, 18, 0, 73, 
    10, 0, 0, 0, 21, 14, 18, 17, 23, 12, 11, 6, 11, 0, 51, 
    5, 0, 0, 0, 9, 30, 7, 21, 22, 20, 26, 0, 39, 0, 44, 
    0, 0, 0, 0, 0, 28, 9, 21, 23, 23, 27, 14, 49, 14, 18, 
    0, 1, 2, 0, 0, 0, 17, 13, 25, 33, 21, 30, 44, 3, 0, 
    28, 0, 11, 0, 0, 0, 0, 28, 26, 38, 24, 30, 33, 0, 0, 
    0, 0, 17, 0, 0, 0, 0, 25, 26, 36, 22, 31, 35, 0, 0, 
    0, 0, 4, 0, 2, 0, 7, 48, 0, 24, 25, 43, 40, 0, 0, 
    21, 0, 0, 0, 11, 0, 0, 13, 0, 19, 17, 45, 57, 0, 0, 
    30, 3, 0, 0, 0, 0, 0, 0, 9, 18, 20, 21, 17, 0, 0, 
    
    -- channel=266
    0, 0, 0, 0, 0, 6, 0, 0, 0, 6, 0, 31, 0, 11, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 42, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 40, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 43, 0, 0, 2, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 
    0, 57, 0, 0, 0, 0, 0, 2, 0, 0, 0, 9, 0, 6, 0, 
    0, 15, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 4, 8, 30, 0, 1, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 5, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 9, 0, 0, 0, 0, 0, 0, 3, 0, 
    36, 79, 0, 0, 0, 15, 15, 0, 46, 0, 0, 0, 0, 16, 0, 
    0, 46, 86, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 62, 80, 0, 0, 0, 0, 0, 14, 28, 0, 0, 0, 30, 
    
    -- channel=267
    15, 39, 32, 29, 13, 67, 14, 33, 0, 0, 0, 48, 0, 28, 27, 
    13, 27, 3, 20, 18, 36, 17, 45, 3, 16, 0, 49, 0, 46, 0, 
    0, 3, 13, 8, 27, 73, 43, 0, 15, 0, 19, 39, 0, 1, 0, 
    9, 52, 0, 17, 61, 23, 0, 6, 41, 30, 19, 8, 0, 0, 0, 
    11, 19, 0, 0, 46, 0, 0, 70, 3, 18, 0, 0, 0, 0, 0, 
    0, 8, 0, 21, 8, 0, 0, 2, 0, 0, 0, 20, 0, 0, 0, 
    15, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 28, 
    0, 14, 0, 15, 4, 6, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    36, 0, 0, 5, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 20, 26, 
    0, 33, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 29, 2, 
    
    -- channel=268
    10, 15, 24, 20, 0, 31, 16, 21, 16, 18, 10, 36, 0, 13, 26, 
    11, 29, 12, 18, 1, 15, 4, 36, 15, 27, 4, 39, 0, 32, 15, 
    10, 18, 18, 7, 7, 33, 36, 19, 12, 2, 18, 34, 4, 25, 18, 
    2, 33, 14, 13, 26, 37, 24, 0, 38, 13, 20, 49, 0, 17, 0, 
    15, 24, 9, 5, 44, 22, 0, 50, 17, 39, 27, 25, 9, 14, 0, 
    5, 18, 12, 25, 31, 12, 8, 20, 25, 15, 4, 51, 14, 8, 0, 
    19, 18, 14, 13, 5, 4, 14, 6, 5, 4, 9, 22, 4, 25, 0, 
    17, 19, 32, 9, 7, 1, 10, 8, 3, 13, 13, 0, 16, 13, 0, 
    22, 27, 5, 6, 1, 26, 0, 0, 8, 2, 0, 11, 0, 2, 17, 
    21, 5, 17, 24, 5, 0, 16, 8, 0, 0, 7, 0, 0, 17, 30, 
    0, 27, 17, 10, 32, 27, 4, 0, 0, 0, 0, 0, 2, 15, 23, 
    32, 32, 28, 33, 4, 16, 9, 0, 0, 0, 4, 0, 4, 22, 21, 
    8, 3, 25, 38, 28, 15, 0, 0, 0, 0, 0, 0, 0, 23, 28, 
    4, 15, 17, 27, 34, 35, 22, 17, 29, 0, 3, 0, 0, 49, 26, 
    0, 25, 23, 23, 21, 41, 36, 28, 9, 0, 0, 0, 29, 16, 43, 
    
    -- channel=269
    11, 20, 15, 11, 25, 11, 15, 11, 18, 12, 18, 2, 30, 14, 13, 
    10, 19, 14, 11, 25, 16, 14, 13, 12, 12, 18, 0, 24, 10, 11, 
    10, 7, 9, 13, 22, 14, 19, 19, 6, 27, 10, 0, 14, 10, 9, 
    23, 8, 18, 12, 20, 20, 26, 24, 12, 13, 21, 11, 7, 4, 15, 
    18, 0, 12, 23, 0, 16, 32, 15, 18, 14, 16, 12, 10, 0, 23, 
    17, 0, 0, 16, 28, 16, 9, 0, 18, 21, 26, 11, 11, 0, 29, 
    16, 5, 3, 4, 14, 7, 10, 15, 13, 3, 0, 7, 17, 5, 19, 
    14, 4, 2, 1, 0, 21, 3, 6, 1, 10, 10, 0, 6, 6, 26, 
    7, 8, 7, 5, 0, 0, 4, 0, 4, 5, 8, 0, 1, 0, 13, 
    3, 7, 14, 4, 4, 4, 0, 0, 0, 0, 3, 5, 10, 14, 5, 
    15, 10, 17, 5, 10, 1, 0, 0, 0, 2, 0, 8, 13, 3, 6, 
    4, 11, 31, 16, 12, 3, 0, 0, 0, 2, 0, 6, 13, 2, 12, 
    5, 0, 11, 26, 18, 5, 0, 4, 0, 0, 0, 4, 17, 10, 16, 
    23, 20, 0, 9, 29, 24, 22, 12, 6, 0, 0, 9, 17, 8, 6, 
    22, 17, 23, 0, 4, 20, 31, 24, 21, 0, 0, 0, 19, 22, 19, 
    
    -- channel=270
    0, 0, 0, 0, 3, 0, 0, 0, 8, 15, 4, 0, 0, 7, 0, 
    0, 0, 0, 0, 2, 7, 11, 0, 0, 0, 2, 0, 0, 0, 0, 
    34, 23, 0, 2, 0, 0, 0, 0, 6, 14, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 17, 0, 0, 0, 0, 3, 0, 18, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 17, 
    3, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 10, 11, 29, 0, 0, 0, 0, 0, 0, 0, 33, 21, 0, 
    0, 18, 8, 16, 4, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    50, 56, 0, 0, 0, 0, 16, 46, 39, 0, 0, 0, 0, 0, 13, 
    4, 62, 64, 0, 0, 0, 0, 0, 0, 4, 0, 4, 24, 5, 0, 
    12, 0, 36, 47, 0, 0, 0, 0, 14, 37, 50, 7, 0, 0, 0, 
    
    -- channel=271
    0, 0, 16, 4, 0, 58, 0, 19, 0, 10, 0, 71, 0, 39, 7, 
    0, 0, 0, 2, 0, 33, 2, 36, 0, 9, 0, 89, 0, 35, 0, 
    0, 5, 0, 0, 0, 51, 18, 0, 21, 0, 36, 77, 0, 0, 0, 
    0, 63, 0, 0, 8, 39, 0, 0, 63, 0, 44, 48, 0, 0, 0, 
    0, 82, 0, 0, 50, 0, 0, 53, 0, 19, 0, 26, 0, 0, 0, 
    0, 83, 2, 0, 33, 3, 0, 23, 0, 0, 0, 51, 0, 6, 0, 
    0, 47, 31, 0, 0, 0, 0, 3, 0, 2, 1, 10, 0, 13, 0, 
    0, 36, 17, 0, 0, 0, 25, 0, 0, 0, 0, 21, 0, 5, 0, 
    8, 10, 0, 0, 21, 0, 9, 0, 0, 3, 0, 3, 0, 0, 0, 
    0, 0, 0, 24, 0, 28, 2, 4, 0, 0, 0, 0, 0, 0, 40, 
    0, 38, 0, 28, 8, 0, 63, 0, 0, 0, 0, 0, 0, 8, 4, 
    19, 10, 0, 19, 0, 27, 22, 2, 0, 0, 8, 0, 0, 18, 0, 
    9, 53, 0, 0, 0, 22, 0, 0, 39, 0, 0, 0, 0, 26, 0, 
    0, 33, 80, 1, 0, 0, 0, 0, 31, 6, 1, 0, 0, 48, 29, 
    0, 0, 70, 71, 0, 0, 0, 0, 0, 8, 0, 0, 0, 12, 77, 
    
    -- channel=272
    12, 9, 28, 16, 0, 24, 11, 9, 0, 0, 0, 15, 0, 0, 4, 
    7, 13, 8, 15, 0, 9, 0, 10, 4, 14, 0, 21, 0, 40, 14, 
    0, 0, 2, 1, 0, 22, 32, 13, 0, 0, 0, 22, 0, 9, 6, 
    0, 27, 8, 0, 7, 29, 0, 0, 13, 2, 18, 13, 0, 4, 0, 
    6, 23, 3, 0, 23, 7, 0, 28, 15, 17, 0, 0, 0, 0, 0, 
    0, 12, 0, 14, 23, 0, 0, 32, 2, 0, 0, 17, 0, 0, 0, 
    8, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 6, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 17, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 3, 0, 10, 7, 1, 0, 0, 0, 0, 0, 0, 0, 3, 25, 
    16, 41, 2, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 13, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 8, 19, 
    
    -- channel=273
    7, 0, 0, 0, 29, 0, 11, 0, 16, 0, 37, 0, 94, 0, 0, 
    0, 0, 12, 0, 20, 0, 0, 0, 13, 0, 35, 0, 78, 0, 21, 
    22, 0, 1, 1, 5, 0, 0, 22, 0, 27, 0, 0, 69, 6, 32, 
    17, 0, 21, 9, 0, 0, 46, 8, 0, 0, 0, 0, 57, 14, 79, 
    13, 0, 46, 14, 0, 14, 52, 0, 11, 0, 36, 0, 40, 19, 89, 
    19, 0, 14, 24, 1, 7, 12, 0, 23, 21, 29, 0, 52, 7, 90, 
    11, 0, 0, 25, 27, 8, 6, 14, 16, 8, 0, 5, 32, 5, 63, 
    12, 0, 0, 21, 16, 5, 0, 17, 11, 8, 14, 0, 45, 17, 47, 
    0, 2, 9, 6, 0, 25, 0, 9, 17, 16, 20, 11, 40, 15, 25, 
    14, 12, 18, 4, 7, 0, 5, 9, 14, 33, 10, 29, 42, 6, 0, 
    42, 0, 25, 0, 3, 6, 0, 26, 26, 30, 13, 23, 31, 0, 14, 
    0, 17, 49, 1, 26, 0, 6, 27, 18, 27, 17, 27, 31, 0, 15, 
    17, 0, 45, 47, 33, 1, 14, 49, 0, 15, 19, 27, 44, 0, 29, 
    41, 0, 0, 30, 57, 29, 23, 23, 0, 18, 13, 38, 48, 0, 0, 
    51, 7, 0, 0, 35, 45, 46, 32, 28, 17, 19, 7, 12, 0, 0, 
    
    -- channel=274
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    1, 0, 0, 0, 0, 0, 7, 0, 0, 0, 2, 0, 0, 0, 12, 
    0, 0, 0, 0, 29, 0, 0, 0, 15, 22, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 0, 51, 0, 0, 4, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 12, 12, 0, 8, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 2, 11, 0, 0, 0, 0, 0, 0, 
    17, 30, 18, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 7, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    
    -- channel=275
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 1, 4, 0, 5, 7, 11, 0, 0, 0, 
    0, 0, 0, 0, 16, 0, 2, 14, 14, 16, 17, 14, 29, 0, 0, 
    0, 0, 0, 0, 0, 31, 11, 18, 26, 21, 15, 20, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 22, 32, 25, 34, 18, 19, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 35, 38, 22, 18, 15, 8, 0, 0, 
    0, 20, 0, 0, 0, 0, 14, 29, 29, 24, 25, 21, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 4, 13, 0, 25, 25, 20, 9, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 19, 24, 19, 0, 0, 0, 
    0, 0, 0, 0, 6, 8, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    
    -- channel=276
    5, 0, 23, 7, 0, 40, 3, 8, 14, 3, 0, 43, 0, 31, 0, 
    0, 0, 0, 6, 0, 30, 1, 22, 0, 12, 0, 64, 0, 40, 0, 
    0, 0, 0, 0, 0, 33, 24, 2, 10, 0, 26, 62, 0, 5, 5, 
    0, 59, 0, 0, 0, 44, 0, 0, 56, 0, 52, 41, 0, 2, 0, 
    0, 75, 0, 0, 23, 11, 0, 31, 19, 25, 8, 16, 0, 2, 0, 
    0, 75, 3, 0, 45, 10, 0, 23, 0, 1, 0, 31, 0, 6, 0, 
    0, 52, 23, 0, 0, 0, 0, 9, 0, 0, 0, 2, 0, 17, 0, 
    0, 33, 10, 6, 0, 0, 13, 0, 0, 0, 0, 9, 0, 0, 0, 
    3, 19, 0, 0, 33, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 18, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 30, 
    0, 21, 0, 32, 18, 0, 59, 0, 0, 0, 0, 0, 0, 0, 13, 
    8, 28, 0, 27, 0, 35, 23, 0, 0, 0, 8, 0, 0, 0, 0, 
    11, 31, 0, 0, 0, 26, 13, 0, 12, 0, 4, 0, 0, 0, 1, 
    0, 29, 48, 0, 0, 0, 10, 0, 39, 6, 0, 0, 0, 25, 11, 
    0, 0, 70, 54, 0, 0, 0, 10, 0, 10, 0, 0, 0, 23, 80, 
    
    -- channel=277
    18, 33, 4, 5, 55, 0, 11, 0, 0, 0, 29, 0, 81, 0, 8, 
    12, 24, 15, 3, 56, 0, 0, 0, 11, 0, 31, 0, 83, 0, 23, 
    0, 0, 4, 4, 46, 0, 13, 10, 0, 29, 0, 0, 40, 7, 12, 
    38, 0, 28, 26, 14, 0, 15, 30, 0, 39, 0, 0, 3, 0, 46, 
    33, 0, 61, 22, 0, 0, 68, 0, 11, 0, 0, 0, 0, 0, 86, 
    35, 0, 0, 85, 0, 0, 1, 0, 8, 0, 7, 0, 14, 0, 99, 
    48, 0, 0, 6, 2, 0, 9, 0, 0, 0, 0, 0, 1, 0, 77, 
    21, 0, 0, 0, 10, 17, 0, 0, 3, 15, 4, 0, 34, 0, 68, 
    0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 53, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 17, 0, 
    37, 0, 29, 0, 0, 21, 0, 0, 0, 0, 0, 0, 13, 0, 0, 
    10, 19, 67, 0, 11, 0, 0, 0, 0, 10, 0, 0, 6, 0, 0, 
    0, 0, 10, 34, 29, 0, 0, 0, 0, 0, 0, 14, 19, 0, 0, 
    34, 0, 0, 0, 41, 21, 0, 31, 0, 0, 0, 5, 34, 0, 0, 
    37, 35, 0, 0, 0, 33, 32, 15, 0, 0, 0, 0, 56, 28, 0, 
    
    -- channel=278
    0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 
    0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 33, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 2, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 54, 
    30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 62, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 11, 5, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 0, 7, 0, 0, 
    3, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 64, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 8, 0, 0, 0, 
    
    -- channel=279
    0, 0, 0, 0, 0, 32, 0, 14, 0, 1, 0, 35, 0, 29, 0, 
    0, 0, 0, 0, 0, 33, 4, 15, 0, 0, 0, 42, 0, 0, 0, 
    0, 1, 0, 0, 0, 15, 0, 0, 6, 0, 0, 36, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 1, 13, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 14, 0, 0, 6, 0, 0, 0, 15, 0, 0, 0, 
    0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 34, 0, 
    0, 51, 24, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 3, 0, 
    0, 0, 59, 16, 0, 0, 0, 0, 0, 1, 10, 0, 0, 0, 0, 
    
    -- channel=280
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 5, 5, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 9, 0, 
    0, 7, 6, 0, 0, 0, 2, 9, 5, 5, 2, 0, 8, 5, 0, 
    0, 0, 8, 11, 15, 14, 4, 18, 17, 18, 14, 25, 13, 7, 0, 
    0, 0, 2, 15, 12, 2, 16, 25, 17, 15, 22, 30, 25, 16, 0, 
    0, 0, 2, 0, 21, 15, 26, 27, 32, 33, 26, 31, 30, 8, 0, 
    4, 0, 0, 0, 0, 20, 25, 36, 37, 40, 25, 27, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 29, 45, 42, 35, 30, 25, 11, 0, 5, 
    0, 18, 0, 0, 0, 3, 32, 47, 42, 28, 33, 31, 10, 7, 0, 
    19, 28, 18, 1, 0, 5, 21, 31, 23, 33, 39, 24, 14, 0, 0, 
    0, 0, 17, 15, 5, 0, 0, 0, 0, 36, 34, 26, 0, 0, 0, 
    0, 0, 0, 19, 22, 10, 0, 0, 5, 22, 28, 0, 0, 0, 13, 
    
    -- channel=281
    31, 20, 36, 19, 3, 22, 22, 9, 3, 0, 6, 13, 15, 0, 17, 
    23, 21, 20, 17, 0, 0, 0, 11, 26, 18, 12, 16, 44, 49, 30, 
    0, 0, 9, 0, 0, 42, 50, 11, 5, 0, 20, 20, 33, 24, 26, 
    9, 51, 11, 11, 15, 45, 4, 0, 8, 30, 42, 14, 13, 21, 0, 
    11, 30, 40, 0, 37, 28, 7, 41, 46, 39, 22, 0, 13, 12, 0, 
    0, 5, 22, 56, 33, 0, 13, 54, 24, 6, 1, 23, 9, 9, 9, 
    24, 21, 0, 14, 0, 4, 24, 1, 0, 0, 19, 12, 0, 15, 19, 
    0, 14, 10, 0, 47, 0, 4, 6, 31, 33, 1, 6, 21, 3, 0, 
    29, 25, 0, 0, 0, 46, 2, 9, 8, 0, 0, 0, 0, 0, 23, 
    8, 0, 0, 0, 3, 0, 22, 19, 0, 10, 0, 0, 6, 8, 24, 
    0, 15, 16, 30, 9, 23, 3, 8, 5, 0, 0, 0, 7, 21, 31, 
    54, 89, 52, 18, 10, 5, 9, 0, 0, 0, 19, 0, 0, 7, 8, 
    0, 0, 38, 38, 21, 10, 0, 0, 0, 10, 0, 1, 0, 0, 0, 
    1, 0, 0, 32, 42, 27, 2, 40, 17, 0, 2, 0, 0, 5, 37, 
    6, 36, 0, 0, 30, 54, 38, 19, 0, 0, 0, 0, 42, 48, 26, 
    
    -- channel=282
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    22, 46, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 15, 5, 
    
    -- channel=283
    9, 16, 5, 21, 25, 0, 11, 11, 11, 14, 18, 6, 20, 2, 9, 
    23, 16, 20, 20, 24, 0, 11, 6, 15, 12, 20, 0, 25, 3, 17, 
    11, 9, 17, 21, 21, 2, 11, 14, 19, 20, 5, 7, 23, 21, 18, 
    23, 2, 18, 13, 13, 3, 17, 26, 0, 20, 4, 8, 23, 23, 24, 
    24, 7, 30, 15, 0, 18, 28, 0, 18, 10, 12, 20, 21, 25, 34, 
    24, 4, 31, 34, 6, 8, 3, 2, 16, 14, 16, 2, 23, 26, 32, 
    20, 10, 24, 24, 9, 0, 0, 0, 0, 0, 0, 0, 18, 22, 35, 
    22, 13, 18, 23, 0, 4, 0, 0, 0, 0, 0, 0, 4, 16, 35, 
    19, 21, 29, 27, 8, 0, 0, 0, 0, 0, 0, 0, 8, 13, 22, 
    18, 27, 19, 8, 16, 5, 0, 0, 1, 0, 0, 0, 5, 7, 18, 
    30, 3, 23, 18, 20, 14, 0, 6, 2, 2, 0, 0, 2, 19, 18, 
    22, 8, 24, 20, 25, 17, 0, 0, 4, 7, 0, 0, 0, 5, 37, 
    13, 11, 19, 23, 25, 12, 9, 0, 0, 2, 0, 0, 0, 11, 26, 
    15, 0, 2, 15, 26, 21, 17, 16, 2, 0, 0, 0, 9, 0, 32, 
    19, 2, 0, 4, 16, 27, 24, 20, 10, 0, 0, 7, 13, 21, 0, 
    
    -- channel=284
    32, 49, 40, 47, 53, 31, 41, 37, 36, 35, 46, 24, 56, 23, 40, 
    38, 55, 45, 41, 58, 27, 32, 39, 41, 40, 45, 18, 53, 33, 44, 
    33, 35, 39, 39, 56, 40, 52, 48, 32, 47, 25, 21, 38, 44, 36, 
    49, 26, 42, 44, 50, 43, 56, 54, 27, 49, 29, 39, 27, 34, 36, 
    54, 9, 54, 38, 34, 40, 57, 40, 45, 47, 45, 35, 33, 31, 52, 
    53, 3, 32, 74, 35, 23, 23, 22, 44, 32, 32, 34, 42, 27, 61, 
    56, 21, 23, 34, 25, 9, 18, 16, 12, 3, 10, 20, 28, 36, 57, 
    49, 26, 36, 24, 9, 24, 0, 0, 9, 15, 14, 0, 28, 28, 60, 
    37, 38, 34, 30, 1, 22, 0, 0, 6, 0, 3, 7, 3, 24, 61, 
    34, 38, 46, 26, 25, 0, 9, 0, 0, 2, 6, 6, 22, 33, 32, 
    46, 24, 54, 27, 44, 42, 0, 1, 1, 0, 3, 3, 20, 35, 37, 
    38, 35, 69, 48, 39, 22, 0, 0, 0, 10, 0, 2, 20, 26, 53, 
    19, 0, 43, 63, 61, 18, 8, 2, 0, 1, 0, 13, 15, 35, 51, 
    42, 20, 0, 31, 65, 62, 42, 42, 21, 0, 0, 10, 32, 30, 50, 
    47, 51, 16, 4, 28, 62, 64, 50, 29, 0, 0, 18, 53, 47, 19, 
    
    -- channel=285
    6, 0, 16, 7, 0, 2, 5, 0, 4, 0, 0, 0, 2, 0, 0, 
    1, 0, 6, 8, 0, 2, 0, 0, 2, 3, 0, 0, 1, 15, 11, 
    0, 0, 0, 0, 0, 5, 16, 8, 0, 0, 2, 0, 6, 6, 8, 
    0, 20, 3, 0, 0, 27, 9, 0, 6, 0, 24, 3, 0, 2, 5, 
    0, 20, 5, 0, 0, 11, 0, 0, 18, 8, 9, 0, 0, 0, 0, 
    0, 13, 0, 0, 28, 0, 0, 16, 4, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 32, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 3, 0, 0, 0, 11, 11, 7, 0, 0, 0, 0, 0, 18, 24, 
    
    -- channel=286
    0, 6, 0, 0, 0, 1, 0, 4, 0, 4, 0, 3, 0, 5, 1, 
    0, 2, 0, 0, 2, 1, 1, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 13, 4, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 17, 0, 0, 26, 0, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 2, 1, 0, 0, 0, 13, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 11, 0, 1, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 14, 3, 0, 2, 1, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 
    0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 4, 0, 22, 0, 
    0, 12, 5, 0, 0, 2, 0, 2, 0, 0, 0, 0, 15, 0, 10, 
    0, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 16, 6, 0, 0, 
    
    -- channel=287
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=288
    34, 0, 35, 2, 2, 3, 12, 0, 5, 0, 16, 0, 49, 6, 0, 
    0, 0, 0, 8, 0, 4, 5, 0, 16, 0, 24, 0, 59, 15, 20, 
    0, 0, 0, 0, 0, 19, 15, 0, 0, 0, 60, 0, 57, 0, 37, 
    7, 57, 0, 0, 0, 40, 13, 0, 27, 0, 59, 0, 42, 2, 56, 
    0, 52, 30, 0, 0, 1, 4, 0, 26, 4, 17, 0, 18, 5, 36, 
    0, 40, 11, 0, 41, 0, 0, 22, 0, 0, 0, 0, 2, 5, 28, 
    0, 28, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 7, 39, 0, 14, 0, 0, 4, 0, 0, 11, 5, 0, 
    0, 0, 0, 0, 0, 20, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 11, 0, 0, 10, 0, 12, 0, 0, 18, 10, 0, 
    0, 22, 0, 21, 0, 0, 24, 0, 5, 0, 0, 4, 2, 0, 27, 
    0, 61, 8, 0, 2, 0, 16, 13, 0, 0, 31, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    29, 0, 10, 9, 2, 0, 0, 13, 0, 10, 0, 0, 0, 13, 0, 
    14, 33, 0, 1, 2, 0, 5, 18, 0, 2, 0, 0, 0, 33, 38, 
    
    -- channel=289
    1, 0, 0, 0, 0, 0, 0, 0, 12, 1, 8, 0, 35, 0, 0, 
    2, 0, 1, 0, 0, 0, 0, 0, 8, 0, 12, 0, 38, 0, 14, 
    4, 0, 0, 0, 0, 0, 0, 4, 0, 0, 8, 0, 58, 13, 29, 
    0, 0, 4, 0, 0, 18, 21, 0, 0, 0, 27, 7, 63, 26, 46, 
    0, 25, 28, 0, 0, 23, 6, 0, 25, 9, 35, 7, 46, 30, 32, 
    0, 24, 40, 0, 22, 7, 3, 29, 28, 22, 28, 0, 40, 35, 24, 
    0, 12, 24, 39, 23, 12, 4, 16, 14, 13, 8, 15, 35, 29, 15, 
    0, 9, 9, 38, 29, 0, 12, 23, 21, 12, 9, 29, 28, 32, 0, 
    4, 16, 19, 25, 23, 11, 20, 26, 24, 25, 28, 16, 38, 16, 0, 
    19, 13, 0, 14, 17, 31, 13, 30, 33, 40, 17, 28, 21, 0, 0, 
    20, 8, 4, 17, 4, 0, 34, 45, 39, 36, 22, 27, 22, 1, 38, 
    4, 51, 32, 8, 29, 13, 34, 47, 35, 28, 31, 29, 23, 10, 31, 
    28, 51, 61, 39, 17, 30, 36, 34, 12, 31, 44, 21, 21, 0, 28, 
    17, 0, 41, 56, 51, 24, 27, 9, 0, 34, 29, 24, 6, 0, 7, 
    20, 0, 0, 43, 64, 49, 44, 32, 14, 24, 29, 7, 0, 8, 37, 
    
    -- channel=290
    14, 18, 13, 6, 0, 14, 0, 0, 0, 0, 0, 16, 0, 3, 26, 
    14, 16, 0, 4, 0, 0, 1, 17, 5, 0, 0, 17, 27, 29, 0, 
    0, 0, 11, 0, 0, 43, 31, 0, 0, 0, 22, 17, 8, 10, 4, 
    9, 49, 1, 6, 35, 11, 0, 0, 19, 28, 27, 7, 0, 5, 0, 
    0, 10, 20, 0, 15, 3, 7, 52, 7, 19, 0, 0, 0, 0, 0, 
    0, 0, 5, 44, 19, 7, 3, 0, 0, 1, 6, 15, 0, 0, 0, 
    16, 6, 0, 0, 0, 0, 22, 7, 2, 0, 8, 10, 1, 0, 1, 
    1, 12, 8, 0, 25, 0, 10, 4, 8, 35, 10, 1, 5, 0, 0, 
    24, 4, 0, 0, 0, 24, 0, 1, 5, 9, 4, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 0, 0, 10, 1, 0, 5, 0, 1, 19, 31, 
    0, 18, 3, 15, 0, 11, 13, 0, 1, 0, 0, 6, 2, 19, 0, 
    66, 45, 30, 12, 0, 6, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 13, 13, 9, 0, 0, 0, 0, 7, 0, 2, 0, 0, 0, 
    0, 0, 0, 19, 14, 10, 1, 37, 13, 0, 2, 0, 0, 0, 40, 
    0, 15, 0, 0, 7, 25, 19, 15, 0, 0, 0, 3, 49, 52, 18, 
    
    -- channel=291
    10, 5, 18, 30, 23, 18, 25, 25, 43, 41, 35, 26, 26, 24, 14, 
    13, 17, 28, 30, 20, 29, 25, 23, 25, 32, 29, 26, 1, 9, 26, 
    52, 39, 28, 32, 16, 0, 17, 44, 33, 41, 22, 25, 20, 30, 31, 
    22, 7, 25, 16, 2, 33, 60, 28, 30, 2, 15, 49, 36, 30, 40, 
    27, 32, 17, 25, 19, 32, 18, 6, 23, 29, 47, 50, 38, 35, 29, 
    28, 44, 34, 0, 29, 18, 3, 14, 30, 30, 23, 35, 43, 40, 19, 
    12, 28, 44, 35, 18, 3, 0, 5, 11, 7, 0, 7, 28, 43, 15, 
    29, 30, 35, 41, 0, 3, 0, 0, 0, 0, 0, 3, 2, 39, 32, 
    16, 30, 46, 41, 34, 0, 0, 0, 0, 2, 1, 10, 19, 37, 17, 
    41, 42, 43, 46, 32, 32, 0, 0, 0, 0, 0, 5, 0, 17, 16, 
    38, 28, 28, 19, 35, 20, 8, 3, 2, 8, 3, 0, 4, 11, 42, 
    0, 0, 16, 40, 36, 25, 15, 7, 5, 1, 0, 2, 12, 35, 52, 
    70, 60, 29, 38, 38, 43, 24, 34, 24, 0, 1, 0, 9, 35, 68, 
    32, 72, 67, 34, 33, 43, 45, 5, 11, 10, 3, 11, 19, 47, 19, 
    35, 12, 57, 69, 37, 28, 42, 41, 44, 25, 35, 6, 0, 0, 41, 
    
    -- channel=292
    17, 0, 30, 11, 0, 39, 12, 12, 21, 14, 0, 29, 0, 37, 6, 
    2, 0, 7, 12, 0, 37, 16, 18, 12, 14, 3, 42, 0, 29, 7, 
    0, 7, 4, 0, 0, 35, 21, 7, 18, 0, 44, 32, 1, 7, 11, 
    0, 54, 0, 0, 0, 50, 12, 0, 43, 0, 56, 24, 10, 4, 0, 
    0, 64, 0, 0, 25, 18, 0, 26, 27, 19, 18, 13, 9, 2, 0, 
    0, 64, 7, 0, 46, 9, 0, 31, 6, 13, 10, 22, 0, 10, 0, 
    0, 42, 17, 0, 0, 9, 2, 12, 4, 8, 1, 7, 1, 12, 0, 
    0, 29, 5, 4, 12, 0, 25, 8, 2, 5, 0, 15, 0, 13, 0, 
    5, 11, 0, 3, 10, 0, 10, 1, 4, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 11, 24, 0, 5, 0, 0, 0, 0, 0, 5, 20, 
    0, 33, 0, 32, 2, 0, 45, 0, 0, 0, 0, 3, 0, 0, 21, 
    1, 31, 0, 11, 0, 16, 22, 10, 0, 0, 15, 0, 0, 10, 0, 
    10, 34, 1, 0, 0, 22, 7, 0, 14, 0, 9, 0, 0, 2, 8, 
    3, 25, 59, 17, 0, 4, 12, 0, 13, 13, 2, 0, 0, 34, 17, 
    0, 14, 55, 53, 13, 0, 6, 17, 0, 14, 6, 0, 0, 26, 67, 
    
    -- channel=293
    16, 17, 40, 9, 0, 21, 12, 3, 0, 0, 0, 9, 0, 0, 6, 
    12, 30, 8, 9, 0, 0, 0, 14, 7, 17, 0, 19, 4, 65, 21, 
    0, 0, 0, 0, 0, 36, 57, 15, 0, 0, 0, 30, 8, 16, 12, 
    0, 41, 21, 0, 13, 54, 0, 0, 18, 0, 51, 27, 0, 10, 0, 
    5, 19, 13, 2, 26, 17, 0, 47, 38, 41, 9, 0, 0, 0, 0, 
    0, 0, 0, 37, 51, 0, 8, 48, 21, 0, 0, 37, 0, 0, 0, 
    16, 21, 0, 0, 0, 0, 11, 7, 0, 0, 4, 17, 0, 11, 0, 
    0, 2, 9, 0, 14, 0, 0, 0, 11, 32, 11, 0, 16, 0, 0, 
    18, 31, 0, 0, 0, 8, 12, 0, 4, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 1, 10, 
    0, 1, 7, 10, 19, 0, 0, 0, 0, 0, 0, 0, 0, 7, 38, 
    34, 104, 52, 29, 0, 0, 0, 0, 0, 0, 3, 0, 0, 3, 0, 
    0, 0, 1, 39, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 36, 21, 0, 1, 36, 0, 0, 0, 0, 1, 0, 
    0, 11, 0, 0, 0, 42, 32, 4, 0, 0, 0, 0, 30, 39, 57, 
    
    -- channel=294
    0, 0, 1, 1, 0, 21, 1, 11, 22, 20, 0, 23, 0, 33, 0, 
    0, 0, 0, 1, 0, 34, 15, 13, 0, 8, 0, 32, 0, 0, 0, 
    19, 9, 0, 7, 0, 2, 0, 10, 14, 13, 9, 27, 0, 0, 0, 
    0, 4, 0, 0, 0, 13, 19, 10, 32, 0, 15, 22, 0, 0, 0, 
    0, 25, 0, 5, 0, 5, 0, 0, 0, 0, 8, 33, 0, 0, 0, 
    0, 42, 0, 0, 19, 16, 0, 0, 0, 17, 8, 14, 0, 0, 0, 
    0, 22, 18, 0, 1, 5, 0, 10, 6, 2, 0, 3, 0, 3, 0, 
    0, 12, 0, 0, 0, 3, 7, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 1, 10, 6, 31, 0, 5, 0, 0, 0, 0, 1, 0, 6, 0, 
    0, 8, 1, 17, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 4, 11, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 15, 7, 0, 0, 0, 0, 0, 0, 3, 0, 
    45, 38, 0, 0, 0, 6, 10, 14, 23, 0, 0, 0, 0, 21, 15, 
    0, 82, 58, 0, 0, 1, 10, 0, 11, 4, 0, 0, 0, 22, 0, 
    0, 0, 84, 54, 0, 0, 0, 13, 15, 15, 20, 0, 0, 0, 37, 
    
    -- channel=295
    0, 0, 0, 0, 0, 32, 0, 4, 0, 0, 0, 36, 0, 24, 0, 
    0, 0, 0, 0, 0, 25, 0, 9, 0, 0, 0, 49, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 3, 0, 7, 36, 0, 0, 0, 
    0, 16, 0, 0, 0, 0, 0, 0, 25, 0, 2, 4, 0, 0, 0, 
    0, 38, 0, 0, 20, 0, 0, 8, 0, 0, 0, 2, 0, 0, 0, 
    0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 15, 3, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 16, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 39, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 7, 0, 
    0, 35, 56, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 19, 0, 
    0, 0, 54, 45, 0, 0, 0, 0, 0, 17, 17, 0, 0, 0, 25, 
    
    -- channel=296
    0, 0, 0, 0, 32, 0, 0, 0, 0, 2, 19, 0, 58, 0, 0, 
    0, 0, 0, 0, 32, 0, 9, 0, 0, 0, 20, 0, 33, 0, 0, 
    22, 14, 0, 4, 27, 0, 0, 0, 0, 36, 0, 0, 10, 0, 0, 
    20, 0, 0, 3, 0, 0, 13, 53, 0, 0, 0, 0, 19, 0, 52, 
    3, 0, 6, 6, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 83, 
    31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 17, 0, 71, 
    0, 0, 0, 0, 4, 0, 0, 0, 2, 0, 0, 0, 15, 0, 46, 
    10, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 76, 
    0, 0, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 33, 26, 15, 
    0, 26, 18, 0, 8, 2, 0, 0, 0, 0, 0, 1, 31, 0, 0, 
    47, 0, 1, 0, 0, 0, 0, 0, 0, 13, 0, 1, 3, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 4, 0, 0, 19, 0, 0, 
    19, 10, 0, 0, 0, 0, 0, 57, 8, 0, 0, 9, 20, 0, 0, 
    24, 23, 4, 0, 0, 0, 0, 0, 0, 0, 0, 19, 78, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 15, 10, 34, 27, 0, 0, 0, 
    
    -- channel=297
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 6, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 1, 0, 0, 0, 3, 0, 0, 5, 0, 9, 3, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 2, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 21, 9, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 7, 0, 
    0, 2, 33, 17, 0, 1, 2, 2, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 8, 26, 13, 2, 6, 6, 0, 0, 0, 11, 0, 1, 0, 
    
    -- channel=298
    0, 0, 0, 0, 0, 21, 0, 21, 0, 27, 0, 42, 0, 33, 0, 
    0, 0, 0, 0, 0, 29, 16, 12, 0, 0, 0, 42, 0, 0, 0, 
    15, 28, 0, 9, 0, 0, 0, 0, 27, 0, 0, 39, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 20, 13, 0, 0, 13, 0, 0, 0, 
    0, 16, 0, 0, 4, 0, 0, 0, 0, 0, 0, 51, 0, 0, 0, 
    0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 4, 0, 
    0, 6, 37, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 10, 3, 0, 0, 0, 0, 18, 0, 2, 0, 
    0, 0, 26, 20, 40, 0, 7, 0, 0, 0, 1, 0, 14, 29, 0, 
    0, 23, 1, 12, 5, 77, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 7, 0, 0, 0, 0, 28, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 3, 0, 0, 0, 0, 20, 0, 
    52, 88, 0, 0, 0, 18, 6, 26, 76, 0, 0, 0, 0, 61, 0, 
    0, 93, 92, 0, 0, 0, 0, 0, 0, 7, 0, 0, 4, 15, 0, 
    0, 0, 80, 74, 0, 0, 0, 0, 15, 29, 47, 15, 0, 0, 3, 
    
    -- channel=299
    20, 27, 26, 8, 18, 0, 13, 0, 0, 0, 10, 0, 41, 0, 15, 
    14, 30, 10, 7, 19, 0, 0, 3, 9, 6, 9, 0, 54, 31, 26, 
    0, 0, 4, 0, 13, 23, 41, 10, 0, 0, 0, 0, 32, 17, 16, 
    11, 19, 24, 18, 19, 20, 3, 0, 0, 26, 19, 0, 0, 7, 10, 
    19, 0, 46, 4, 4, 9, 31, 29, 21, 24, 6, 0, 1, 0, 22, 
    8, 0, 0, 78, 26, 0, 10, 15, 21, 0, 0, 5, 5, 0, 43, 
    37, 0, 0, 3, 0, 0, 18, 9, 0, 0, 2, 14, 0, 0, 34, 
    7, 0, 6, 0, 21, 4, 0, 0, 13, 36, 19, 0, 41, 0, 5, 
    13, 17, 0, 0, 0, 43, 0, 0, 11, 0, 0, 0, 0, 0, 34, 
    2, 0, 0, 0, 0, 0, 6, 10, 0, 4, 0, 0, 12, 15, 0, 
    0, 0, 24, 0, 13, 22, 0, 0, 1, 0, 0, 0, 12, 7, 15, 
    37, 73, 71, 16, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 
    0, 0, 14, 45, 29, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 
    10, 0, 0, 0, 49, 26, 0, 29, 14, 0, 0, 0, 0, 0, 2, 
    8, 31, 0, 0, 0, 52, 39, 16, 0, 0, 0, 0, 58, 40, 0, 
    
    -- channel=300
    6, 0, 32, 9, 0, 48, 0, 18, 0, 0, 0, 63, 0, 24, 10, 
    12, 9, 0, 7, 0, 23, 0, 34, 0, 19, 0, 83, 0, 66, 0, 
    0, 0, 0, 0, 0, 54, 46, 0, 8, 0, 5, 90, 0, 14, 0, 
    0, 72, 0, 0, 20, 52, 0, 0, 49, 0, 58, 58, 0, 6, 0, 
    0, 69, 0, 0, 47, 12, 0, 61, 25, 39, 0, 19, 0, 0, 0, 
    0, 54, 0, 0, 53, 7, 0, 43, 0, 1, 0, 62, 0, 1, 0, 
    0, 50, 24, 0, 0, 3, 10, 15, 0, 1, 12, 22, 0, 18, 0, 
    0, 34, 23, 0, 14, 0, 17, 2, 10, 31, 14, 23, 0, 0, 0, 
    21, 29, 0, 0, 10, 0, 28, 4, 12, 0, 0, 15, 0, 0, 0, 
    3, 0, 0, 0, 0, 9, 5, 21, 2, 0, 0, 0, 0, 0, 35, 
    0, 25, 0, 32, 17, 0, 53, 1, 0, 0, 0, 0, 0, 17, 23, 
    39, 68, 0, 39, 0, 24, 24, 0, 0, 0, 14, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 5, 0, 0, 12, 0, 
    0, 0, 3, 1, 0, 8, 0, 0, 59, 1, 0, 0, 0, 20, 20, 
    0, 0, 42, 18, 0, 5, 0, 7, 0, 0, 0, 0, 2, 39, 88, 
    
    -- channel=301
    9, 15, 12, 0, 12, 0, 12, 0, 0, 0, 3, 0, 27, 0, 0, 
    6, 19, 3, 1, 15, 0, 0, 0, 4, 6, 3, 0, 26, 19, 19, 
    0, 0, 0, 0, 14, 1, 20, 10, 0, 0, 0, 0, 14, 9, 9, 
    0, 0, 12, 16, 3, 8, 4, 0, 0, 24, 0, 0, 0, 8, 4, 
    17, 0, 35, 0, 12, 12, 15, 5, 13, 13, 6, 0, 0, 0, 10, 
    11, 0, 0, 58, 5, 5, 6, 34, 23, 7, 0, 10, 0, 0, 28, 
    29, 0, 0, 11, 13, 5, 19, 4, 0, 0, 15, 16, 0, 0, 23, 
    3, 0, 3, 0, 35, 0, 0, 0, 25, 25, 8, 0, 40, 0, 3, 
    5, 12, 0, 0, 0, 58, 0, 2, 13, 0, 0, 13, 0, 0, 29, 
    5, 0, 0, 0, 0, 0, 25, 18, 0, 12, 1, 1, 7, 0, 0, 
    1, 0, 13, 0, 0, 34, 0, 8, 9, 0, 0, 0, 2, 0, 12, 
    18, 58, 43, 0, 0, 0, 7, 0, 0, 8, 12, 1, 0, 0, 0, 
    0, 0, 18, 31, 17, 0, 0, 0, 0, 5, 0, 8, 6, 0, 0, 
    5, 0, 0, 0, 30, 15, 0, 8, 11, 0, 1, 0, 0, 0, 0, 
    4, 25, 0, 0, 0, 40, 20, 4, 0, 0, 0, 0, 28, 6, 0, 
    
    -- channel=302
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=303
    18, 18, 31, 10, 0, 28, 9, 6, 0, 0, 0, 22, 0, 0, 17, 
    15, 25, 1, 9, 0, 0, 0, 19, 12, 12, 0, 27, 19, 56, 13, 
    0, 0, 1, 0, 0, 49, 52, 0, 0, 0, 15, 27, 13, 17, 18, 
    0, 55, 5, 0, 25, 45, 0, 0, 19, 20, 41, 22, 0, 12, 0, 
    1, 27, 22, 0, 40, 18, 0, 64, 31, 43, 4, 0, 0, 0, 0, 
    0, 0, 8, 50, 38, 0, 13, 44, 23, 0, 0, 42, 0, 0, 0, 
    18, 14, 0, 7, 0, 0, 19, 0, 0, 0, 13, 13, 0, 11, 0, 
    0, 7, 11, 0, 36, 0, 0, 6, 20, 34, 3, 0, 14, 0, 0, 
    27, 23, 0, 0, 0, 42, 0, 0, 2, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 13, 15, 0, 0, 0, 0, 0, 3, 30, 
    0, 16, 7, 17, 11, 15, 3, 0, 0, 0, 0, 0, 0, 14, 21, 
    67, 95, 47, 14, 0, 5, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 23, 35, 9, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 38, 17, 0, 22, 25, 0, 0, 0, 0, 9, 26, 
    0, 25, 0, 0, 9, 51, 33, 8, 0, 0, 0, 0, 41, 42, 42, 
    
    -- channel=304
    15, 11, 11, 0, 4, 8, 5, 2, 3, 0, 3, 0, 19, 10, 7, 
    8, 4, 1, 0, 1, 8, 6, 3, 6, 0, 8, 3, 27, 15, 6, 
    0, 0, 0, 0, 0, 17, 12, 0, 0, 0, 14, 3, 19, 0, 5, 
    7, 17, 10, 7, 8, 12, 0, 0, 11, 8, 26, 1, 9, 2, 7, 
    0, 6, 5, 10, 3, 4, 12, 12, 14, 9, 3, 0, 10, 0, 9, 
    0, 3, 0, 5, 19, 20, 23, 13, 6, 11, 20, 2, 4, 0, 13, 
    5, 8, 0, 0, 20, 33, 39, 36, 30, 29, 28, 25, 15, 0, 6, 
    0, 4, 0, 2, 34, 27, 35, 38, 40, 46, 36, 29, 26, 3, 0, 
    5, 2, 0, 0, 11, 21, 36, 35, 37, 38, 37, 26, 24, 1, 1, 
    0, 0, 0, 0, 5, 24, 22, 32, 35, 33, 30, 33, 31, 11, 4, 
    0, 11, 3, 8, 0, 0, 34, 31, 30, 33, 31, 39, 33, 8, 0, 
    14, 32, 21, 0, 0, 8, 24, 38, 28, 29, 38, 38, 31, 6, 0, 
    0, 1, 11, 10, 4, 4, 16, 23, 18, 32, 39, 35, 34, 0, 0, 
    9, 0, 2, 9, 13, 6, 12, 17, 18, 33, 31, 31, 19, 0, 0, 
    6, 13, 4, 2, 7, 6, 5, 10, 14, 20, 17, 20, 20, 22, 21, 
    
    -- channel=305
    0, 0, 11, 4, 0, 52, 0, 26, 4, 14, 0, 72, 0, 38, 0, 
    4, 0, 0, 2, 0, 35, 3, 32, 0, 13, 0, 89, 0, 38, 0, 
    0, 0, 0, 0, 0, 42, 18, 0, 24, 0, 19, 88, 0, 1, 0, 
    0, 51, 0, 0, 10, 35, 0, 0, 49, 0, 43, 48, 0, 0, 0, 
    0, 77, 0, 0, 42, 5, 0, 40, 11, 21, 0, 44, 0, 0, 0, 
    0, 79, 3, 0, 30, 9, 0, 28, 0, 0, 0, 48, 0, 10, 0, 
    0, 49, 40, 0, 0, 8, 0, 6, 0, 6, 3, 9, 0, 15, 0, 
    0, 35, 14, 0, 0, 0, 20, 0, 0, 0, 0, 24, 0, 0, 0, 
    9, 16, 3, 9, 39, 0, 26, 2, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 14, 0, 54, 0, 3, 2, 0, 0, 0, 0, 0, 37, 
    0, 25, 0, 34, 14, 0, 66, 0, 0, 0, 0, 0, 0, 10, 6, 
    15, 13, 0, 23, 0, 34, 28, 1, 0, 0, 5, 0, 0, 16, 0, 
    17, 56, 0, 0, 0, 29, 18, 0, 41, 0, 8, 0, 0, 29, 0, 
    0, 41, 71, 0, 0, 0, 3, 0, 41, 10, 0, 0, 0, 23, 27, 
    0, 0, 82, 72, 0, 0, 0, 0, 0, 11, 4, 0, 0, 14, 77, 
    
    -- channel=306
    20, 19, 14, 7, 11, 17, 19, 19, 21, 25, 20, 24, 26, 21, 20, 
    17, 19, 14, 9, 13, 16, 19, 18, 25, 17, 22, 22, 34, 20, 14, 
    15, 25, 15, 8, 16, 20, 19, 13, 18, 12, 27, 24, 28, 15, 21, 
    15, 20, 14, 16, 21, 20, 21, 22, 15, 27, 22, 26, 29, 21, 13, 
    13, 18, 19, 18, 29, 27, 22, 24, 26, 27, 26, 36, 28, 16, 12, 
    16, 16, 19, 16, 17, 38, 41, 31, 26, 35, 34, 32, 28, 17, 20, 
    20, 14, 17, 24, 42, 49, 50, 37, 41, 46, 45, 35, 36, 16, 23, 
    17, 17, 13, 25, 49, 33, 47, 52, 53, 45, 36, 48, 32, 22, 14, 
    21, 15, 15, 20, 29, 45, 42, 49, 42, 46, 52, 38, 38, 25, 23, 
    13, 17, 16, 19, 28, 36, 42, 41, 45, 42, 44, 44, 35, 18, 19, 
    15, 29, 20, 18, 10, 24, 40, 39, 41, 40, 43, 47, 38, 21, 13, 
    29, 33, 32, 15, 22, 20, 38, 49, 39, 40, 42, 49, 46, 30, 13, 
    18, 44, 49, 35, 26, 30, 36, 41, 44, 45, 45, 43, 46, 22, 15, 
    19, 17, 44, 50, 36, 30, 34, 34, 24, 43, 47, 43, 33, 18, 22, 
    22, 26, 20, 46, 51, 35, 33, 29, 39, 41, 42, 40, 26, 16, 29, 
    
    -- channel=307
    28, 11, 25, 23, 1, 16, 23, 26, 38, 40, 28, 43, 31, 23, 25, 
    37, 29, 29, 27, 0, 13, 17, 26, 38, 34, 29, 49, 44, 37, 36, 
    29, 30, 28, 23, 0, 18, 33, 29, 33, 17, 37, 57, 65, 47, 47, 
    19, 41, 30, 16, 13, 49, 39, 7, 31, 21, 53, 63, 73, 56, 37, 
    20, 61, 44, 23, 38, 53, 22, 29, 49, 53, 56, 61, 69, 58, 19, 
    17, 57, 65, 29, 51, 47, 46, 58, 56, 53, 53, 61, 64, 60, 19, 
    24, 46, 63, 63, 54, 55, 52, 53, 54, 57, 56, 59, 65, 62, 26, 
    30, 48, 52, 64, 65, 42, 59, 66, 63, 60, 54, 77, 54, 62, 15, 
    46, 50, 51, 55, 65, 52, 65, 68, 66, 69, 71, 61, 63, 44, 24, 
    49, 44, 31, 45, 49, 69, 60, 71, 74, 72, 63, 64, 46, 31, 46, 
    32, 48, 35, 48, 43, 38, 79, 77, 74, 67, 62, 63, 52, 47, 58, 
    56, 77, 56, 51, 52, 53, 70, 80, 74, 63, 66, 65, 56, 55, 58, 
    54, 90, 89, 68, 50, 67, 67, 58, 62, 70, 76, 59, 49, 42, 51, 
    30, 31, 81, 92, 74, 59, 63, 50, 50, 68, 71, 57, 30, 33, 48, 
    30, 12, 41, 85, 98, 80, 72, 61, 53, 59, 59, 51, 30, 40, 79, 
    
    -- channel=308
    0, 5, 0, 0, 0, 5, 0, 0, 0, 0, 0, 3, 0, 4, 9, 
    3, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 5, 1, 0, 0, 
    0, 0, 1, 0, 0, 23, 6, 0, 0, 0, 8, 1, 0, 0, 0, 
    1, 19, 0, 5, 20, 0, 0, 5, 17, 9, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 8, 10, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 12, 6, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 16, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    25, 2, 7, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 2, 0, 0, 0, 0, 0, 27, 
    0, 2, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 17, 32, 2, 
    
    -- channel=309
    0, 21, 0, 0, 89, 0, 0, 0, 0, 0, 55, 0, 142, 0, 0, 
    0, 0, 12, 0, 95, 0, 8, 0, 6, 0, 57, 0, 120, 0, 7, 
    25, 18, 0, 13, 82, 0, 0, 7, 0, 61, 0, 0, 55, 0, 3, 
    57, 0, 10, 33, 0, 0, 36, 90, 0, 52, 0, 0, 38, 0, 98, 
    41, 0, 69, 25, 0, 0, 107, 0, 0, 0, 0, 0, 9, 0, 176, 
    80, 0, 0, 70, 0, 0, 18, 0, 0, 0, 31, 0, 39, 0, 179, 
    49, 0, 0, 12, 21, 0, 0, 0, 1, 0, 0, 0, 31, 0, 142, 
    40, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 26, 0, 148, 
    0, 0, 8, 2, 0, 21, 0, 0, 0, 0, 1, 0, 46, 30, 83, 
    0, 33, 39, 0, 1, 0, 0, 0, 0, 0, 0, 2, 59, 0, 0, 
    91, 0, 41, 0, 0, 5, 0, 0, 0, 10, 0, 2, 21, 0, 0, 
    0, 0, 46, 0, 33, 0, 0, 0, 0, 24, 0, 0, 39, 0, 16, 
    0, 0, 29, 18, 24, 0, 0, 50, 0, 0, 0, 27, 36, 0, 8, 
    57, 0, 0, 0, 35, 0, 0, 25, 0, 0, 0, 31, 119, 0, 0, 
    83, 20, 0, 0, 0, 11, 14, 0, 17, 0, 5, 36, 26, 0, 0, 
    
    -- channel=310
    12, 8, 9, 2, 0, 10, 12, 11, 16, 18, 12, 15, 18, 16, 12, 
    11, 9, 10, 3, 1, 11, 11, 10, 15, 11, 13, 17, 24, 13, 8, 
    6, 13, 9, 2, 3, 13, 12, 8, 12, 4, 19, 18, 22, 11, 13, 
    7, 16, 7, 6, 9, 16, 16, 12, 11, 11, 19, 19, 24, 14, 7, 
    4, 16, 8, 10, 18, 20, 15, 15, 19, 20, 23, 26, 25, 11, 4, 
    5, 15, 14, 5, 16, 25, 29, 22, 20, 26, 27, 24, 24, 10, 7, 
    7, 13, 13, 11, 28, 39, 37, 30, 31, 34, 33, 30, 28, 12, 11, 
    8, 13, 7, 16, 34, 28, 38, 41, 41, 37, 31, 37, 22, 18, 3, 
    13, 11, 11, 14, 24, 27, 34, 38, 35, 38, 41, 31, 31, 19, 8, 
    7, 11, 6, 12, 18, 30, 32, 31, 36, 36, 33, 35, 28, 12, 16, 
    5, 16, 12, 15, 9, 12, 33, 32, 31, 31, 33, 37, 29, 18, 6, 
    18, 26, 21, 13, 11, 16, 29, 39, 33, 29, 36, 37, 36, 24, 9, 
    14, 36, 35, 27, 17, 21, 26, 34, 34, 34, 36, 34, 34, 21, 7, 
    11, 17, 37, 38, 30, 22, 26, 28, 19, 35, 35, 33, 26, 11, 18, 
    14, 15, 22, 39, 40, 29, 27, 24, 25, 32, 32, 33, 17, 15, 23, 
    
    -- channel=311
    0, 15, 5, 9, 15, 11, 8, 14, 22, 20, 9, 16, 9, 27, 8, 
    13, 14, 12, 7, 17, 23, 16, 19, 0, 13, 9, 19, 0, 2, 4, 
    14, 8, 8, 16, 18, 12, 10, 15, 14, 34, 0, 23, 0, 12, 0, 
    15, 5, 14, 9, 20, 14, 26, 39, 20, 1, 19, 26, 0, 1, 2, 
    14, 0, 0, 21, 0, 16, 34, 5, 13, 10, 12, 36, 8, 0, 4, 
    17, 5, 0, 3, 29, 29, 0, 0, 16, 32, 27, 18, 11, 0, 1, 
    3, 13, 14, 0, 16, 14, 3, 31, 17, 2, 0, 21, 10, 8, 0, 
    14, 9, 10, 0, 0, 40, 9, 0, 0, 12, 22, 0, 0, 4, 30, 
    0, 13, 17, 12, 18, 0, 12, 0, 12, 14, 0, 10, 0, 3, 0, 
    1, 19, 16, 3, 5, 13, 0, 0, 0, 0, 5, 4, 0, 8, 5, 
    19, 0, 11, 4, 22, 4, 0, 0, 0, 3, 5, 5, 5, 3, 0, 
    0, 0, 16, 28, 1, 17, 4, 0, 0, 0, 0, 3, 10, 0, 14, 
    26, 3, 0, 20, 24, 0, 6, 10, 0, 0, 0, 6, 4, 27, 15, 
    14, 58, 17, 0, 22, 29, 27, 0, 24, 1, 0, 9, 15, 0, 21, 
    6, 8, 55, 17, 0, 16, 26, 36, 27, 0, 0, 0, 6, 29, 25, 
    
    -- channel=312
    0, 0, 0, 1, 0, 1, 0, 1, 0, 0, 0, 6, 0, 1, 0, 
    0, 0, 0, 1, 0, 2, 0, 0, 0, 0, 0, 6, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 14, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 2, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=313
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 1, 1, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    
    -- channel=314
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 3, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 40, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 8, 16, 
    
    -- channel=315
    9, 12, 0, 0, 44, 0, 0, 0, 0, 0, 25, 0, 79, 0, 0, 
    0, 0, 3, 0, 41, 0, 4, 0, 10, 0, 33, 0, 94, 0, 7, 
    0, 4, 0, 0, 35, 0, 0, 0, 0, 6, 3, 0, 47, 0, 6, 
    33, 0, 0, 21, 0, 0, 0, 39, 0, 46, 0, 0, 31, 0, 49, 
    13, 0, 57, 0, 0, 0, 60, 0, 0, 0, 0, 0, 2, 0, 93, 
    25, 0, 5, 58, 0, 0, 8, 0, 0, 0, 16, 0, 11, 0, 101, 
    27, 0, 0, 5, 5, 0, 7, 0, 0, 0, 0, 0, 13, 0, 84, 
    14, 0, 0, 0, 27, 0, 0, 0, 14, 0, 0, 0, 21, 0, 59, 
    0, 0, 0, 0, 0, 47, 0, 0, 0, 0, 0, 0, 11, 0, 56, 
    0, 2, 0, 0, 8, 0, 1, 0, 0, 5, 0, 1, 43, 0, 0, 
    37, 0, 16, 0, 0, 11, 0, 0, 4, 0, 0, 6, 14, 0, 0, 
    1, 0, 35, 0, 19, 0, 0, 0, 0, 14, 0, 0, 15, 0, 0, 
    0, 0, 34, 6, 7, 0, 0, 1, 0, 8, 0, 17, 20, 0, 0, 
    30, 0, 0, 11, 22, 0, 0, 33, 0, 0, 0, 3, 52, 0, 16, 
    40, 26, 0, 0, 11, 16, 8, 0, 0, 0, 0, 29, 26, 3, 0, 
    
    -- channel=316
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 5, 0, 0, 2, 0, 0, 7, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 11, 16, 0, 
    
    -- channel=317
    0, 16, 0, 0, 47, 0, 0, 0, 0, 0, 22, 0, 81, 0, 0, 
    0, 8, 3, 0, 54, 0, 0, 0, 0, 0, 25, 0, 70, 0, 7, 
    4, 0, 0, 3, 45, 0, 0, 1, 0, 32, 0, 0, 30, 0, 0, 
    26, 0, 10, 18, 0, 0, 10, 38, 0, 27, 0, 0, 5, 0, 51, 
    25, 0, 44, 15, 0, 0, 63, 0, 0, 0, 0, 0, 0, 0, 94, 
    45, 0, 0, 59, 0, 0, 7, 0, 2, 0, 9, 0, 18, 0, 101, 
    34, 0, 0, 3, 13, 0, 0, 0, 0, 0, 0, 0, 7, 0, 78, 
    19, 0, 0, 0, 0, 23, 0, 0, 2, 0, 0, 0, 28, 0, 81, 
    0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 13, 6, 47, 
    0, 10, 14, 0, 0, 0, 0, 0, 0, 4, 0, 3, 35, 0, 0, 
    46, 0, 23, 0, 0, 8, 0, 0, 0, 5, 0, 0, 14, 0, 0, 
    0, 0, 41, 0, 9, 0, 0, 0, 0, 18, 0, 1, 18, 0, 0, 
    0, 0, 10, 15, 16, 0, 0, 22, 0, 0, 0, 21, 23, 0, 0, 
    27, 0, 0, 0, 27, 3, 0, 11, 0, 0, 0, 20, 61, 0, 0, 
    39, 12, 0, 0, 0, 15, 12, 0, 3, 0, 0, 10, 24, 0, 0, 
    
    -- channel=318
    17, 23, 5, 1, 41, 0, 13, 0, 0, 0, 27, 0, 81, 0, 7, 
    7, 17, 6, 0, 42, 0, 0, 0, 14, 0, 29, 0, 90, 0, 25, 
    0, 0, 3, 0, 34, 0, 14, 3, 0, 7, 0, 0, 50, 7, 21, 
    24, 0, 18, 31, 5, 0, 13, 11, 0, 45, 0, 0, 10, 5, 43, 
    25, 0, 69, 1, 0, 2, 55, 0, 9, 5, 4, 0, 3, 0, 76, 
    26, 0, 0, 93, 0, 0, 9, 0, 16, 0, 4, 0, 16, 0, 94, 
    44, 0, 0, 15, 9, 0, 19, 0, 0, 0, 3, 1, 0, 0, 75, 
    19, 0, 0, 0, 36, 0, 0, 0, 21, 25, 6, 0, 54, 0, 45, 
    2, 0, 0, 0, 0, 75, 0, 0, 8, 0, 0, 0, 0, 0, 64, 
    0, 0, 8, 0, 0, 0, 21, 7, 0, 13, 0, 6, 34, 9, 0, 
    28, 0, 29, 0, 0, 39, 0, 4, 10, 0, 0, 4, 17, 0, 0, 
    24, 42, 69, 0, 8, 0, 0, 0, 0, 17, 9, 1, 10, 0, 0, 
    0, 0, 32, 41, 33, 0, 0, 0, 0, 8, 0, 21, 20, 0, 0, 
    29, 0, 0, 2, 49, 22, 0, 36, 0, 0, 0, 5, 21, 0, 6, 
    33, 44, 0, 0, 0, 49, 32, 14, 0, 0, 0, 2, 54, 17, 0, 
    
    -- channel=319
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 18, 
    9, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 4, 8, 1, 0, 10, 7, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 20, 0, 3, 1, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 10, 13, 0, 27, 3, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 4, 4, 8, 8, 17, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 4, 16, 12, 11, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 7, 12, 0, 12, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 38, 19, 5, 3, 18, 17, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 5, 5, 23, 44, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 26, 17, 0, 0, 0, 
    
    -- channel=320
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 25, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 44, 17, 10, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=321
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 3, 0, 13, 0, 0, 0, 0, 
    0, 0, 4, 11, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 8, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=322
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 34, 3, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 43, 35, 66, 73, 11, 0, 0, 0, 
    0, 0, 0, 2, 66, 1, 9, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 5, 8, 0, 66, 37, 42, 43, 4, 24, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 16, 1, 23, 1, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=323
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 4, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=324
    0, 6, 0, 7, 0, 0, 0, 0, 0, 5, 11, 6, 9, 18, 5, 
    4, 0, 0, 1, 1, 0, 0, 0, 0, 0, 14, 13, 15, 8, 9, 
    0, 8, 0, 0, 2, 0, 0, 0, 0, 0, 13, 5, 14, 11, 12, 
    0, 7, 1, 3, 1, 0, 0, 0, 6, 1, 0, 0, 7, 15, 14, 
    3, 10, 3, 0, 0, 3, 12, 18, 3, 13, 6, 0, 13, 11, 13, 
    21, 2, 14, 7, 0, 22, 17, 22, 0, 21, 11, 0, 15, 7, 14, 
    36, 17, 13, 8, 10, 23, 0, 9, 32, 26, 2, 1, 11, 9, 13, 
    4, 37, 12, 11, 26, 15, 9, 29, 22, 20, 6, 1, 10, 21, 4, 
    14, 34, 22, 2, 27, 13, 11, 10, 12, 8, 0, 0, 18, 30, 0, 
    9, 38, 29, 0, 39, 24, 0, 34, 1, 0, 9, 10, 17, 40, 0, 
    16, 27, 19, 0, 10, 9, 8, 25, 0, 0, 8, 12, 15, 42, 1, 
    11, 24, 16, 6, 0, 11, 14, 0, 0, 4, 4, 11, 16, 19, 15, 
    17, 19, 13, 15, 5, 10, 23, 7, 1, 3, 2, 5, 16, 3, 27, 
    18, 26, 11, 8, 3, 15, 26, 7, 13, 11, 5, 14, 4, 12, 8, 
    17, 26, 14, 20, 12, 19, 12, 13, 10, 11, 15, 16, 12, 6, 16, 
    
    -- channel=325
    50, 36, 32, 32, 35, 31, 34, 26, 14, 11, 13, 13, 14, 9, 18, 
    23, 26, 39, 32, 33, 42, 45, 40, 33, 10, 6, 12, 19, 16, 17, 
    7, 17, 33, 32, 32, 36, 40, 37, 47, 49, 32, 31, 13, 17, 20, 
    24, 13, 26, 31, 28, 40, 33, 37, 27, 36, 35, 23, 16, 15, 14, 
    10, 17, 29, 29, 33, 31, 26, 29, 19, 21, 27, 14, 14, 12, 14, 
    15, 19, 18, 24, 23, 26, 4, 0, 21, 16, 5, 4, 2, 14, 11, 
    0, 17, 9, 14, 29, 0, 13, 30, 16, 11, 8, 7, 4, 13, 7, 
    15, 0, 9, 8, 12, 19, 31, 2, 0, 4, 10, 6, 12, 23, 10, 
    28, 13, 10, 6, 0, 2, 0, 0, 0, 0, 0, 0, 4, 4, 11, 
    22, 0, 0, 0, 0, 0, 15, 32, 11, 2, 17, 12, 8, 5, 5, 
    20, 3, 0, 10, 0, 0, 0, 0, 3, 5, 0, 9, 14, 0, 0, 
    25, 11, 1, 45, 35, 44, 35, 5, 0, 0, 0, 0, 3, 0, 0, 
    30, 20, 3, 1, 39, 26, 28, 34, 31, 21, 11, 11, 0, 13, 0, 
    7, 12, 16, 12, 4, 20, 13, 27, 28, 28, 38, 35, 39, 26, 11, 
    24, 20, 29, 29, 36, 21, 18, 22, 20, 26, 29, 27, 28, 24, 28, 
    
    -- channel=326
    38, 15, 5, 11, 14, 4, 10, 0, 15, 0, 9, 14, 8, 0, 22, 
    2, 11, 4, 8, 8, 13, 16, 12, 26, 0, 0, 0, 12, 16, 7, 
    9, 2, 3, 0, 5, 4, 17, 0, 18, 51, 19, 21, 5, 5, 13, 
    8, 0, 0, 0, 1, 2, 6, 5, 0, 11, 8, 17, 9, 1, 5, 
    0, 0, 6, 0, 2, 1, 15, 26, 9, 0, 0, 27, 0, 2, 7, 
    0, 10, 1, 2, 0, 0, 30, 0, 19, 1, 4, 11, 0, 2, 0, 
    0, 0, 7, 13, 1, 0, 4, 59, 31, 18, 26, 18, 0, 4, 0, 
    17, 0, 12, 0, 0, 22, 15, 5, 7, 20, 47, 17, 0, 21, 16, 
    24, 0, 15, 0, 0, 0, 11, 0, 0, 0, 0, 3, 0, 0, 52, 
    26, 0, 12, 46, 0, 0, 27, 34, 28, 0, 21, 27, 0, 0, 84, 
    25, 0, 0, 52, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 62, 
    12, 8, 0, 58, 32, 42, 27, 21, 0, 0, 3, 0, 0, 0, 7, 
    11, 13, 0, 0, 28, 23, 22, 42, 41, 31, 25, 17, 0, 0, 0, 
    11, 0, 18, 0, 13, 16, 0, 33, 24, 32, 36, 33, 38, 16, 18, 
    20, 15, 25, 17, 30, 21, 4, 9, 10, 12, 14, 13, 20, 24, 10, 
    
    -- channel=327
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=328
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=329
    58, 18, 47, 43, 53, 49, 51, 35, 54, 23, 28, 32, 27, 20, 42, 
    35, 50, 42, 48, 48, 51, 58, 47, 64, 33, 19, 31, 30, 42, 33, 
    53, 33, 41, 44, 46, 53, 60, 46, 52, 50, 24, 44, 40, 38, 33, 
    48, 33, 43, 39, 50, 53, 61, 52, 41, 51, 49, 59, 39, 30, 36, 
    24, 31, 43, 45, 48, 52, 46, 42, 55, 37, 41, 70, 23, 34, 33, 
    0, 45, 36, 44, 48, 13, 45, 41, 50, 24, 49, 61, 15, 29, 29, 
    0, 13, 47, 46, 22, 30, 45, 43, 16, 26, 58, 41, 12, 26, 32, 
    51, 0, 48, 34, 11, 43, 43, 31, 34, 35, 66, 41, 2, 14, 49, 
    57, 0, 41, 46, 24, 23, 70, 48, 39, 45, 71, 34, 0, 5, 74, 
    65, 0, 33, 99, 0, 18, 76, 20, 78, 38, 25, 32, 0, 0, 92, 
    64, 17, 41, 96, 8, 22, 34, 37, 65, 31, 20, 19, 10, 0, 82, 
    57, 42, 27, 49, 50, 27, 31, 58, 29, 14, 13, 3, 2, 10, 33, 
    41, 52, 42, 21, 50, 50, 40, 57, 37, 21, 21, 5, 3, 21, 25, 
    58, 29, 64, 30, 48, 38, 35, 66, 39, 38, 34, 24, 34, 25, 41, 
    50, 39, 57, 42, 43, 52, 52, 53, 49, 49, 41, 41, 49, 53, 27, 
    
    -- channel=330
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 
    28, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20, 0, 0, 13, 4, 0, 15, 11, 16, 0, 0, 3, 6, 0, 
    0, 23, 0, 0, 95, 17, 0, 0, 0, 0, 0, 0, 6, 28, 0, 
    0, 16, 0, 0, 0, 13, 0, 24, 0, 0, 0, 0, 0, 59, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 0, 
    0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=331
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 4, 5, 15, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    22, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 25, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 48, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 19, 35, 0, 0, 
    0, 0, 0, 0, 35, 0, 0, 0, 0, 8, 11, 18, 27, 0, 0, 
    0, 0, 0, 0, 0, 28, 15, 0, 18, 33, 36, 37, 30, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 23, 44, 49, 60, 28, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 19, 17, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=332
    3, 20, 0, 4, 0, 0, 0, 5, 0, 0, 0, 3, 4, 2, 0, 
    12, 1, 7, 0, 0, 4, 2, 1, 0, 4, 0, 0, 0, 0, 0, 
    0, 5, 8, 2, 4, 0, 2, 3, 4, 11, 5, 0, 0, 0, 0, 
    6, 0, 2, 5, 2, 2, 0, 4, 0, 0, 2, 0, 0, 2, 0, 
    0, 6, 5, 6, 4, 3, 1, 10, 0, 0, 7, 0, 2, 0, 0, 
    23, 0, 10, 4, 0, 20, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    18, 8, 0, 0, 18, 4, 0, 5, 13, 12, 0, 0, 3, 3, 0, 
    0, 8, 0, 0, 15, 0, 8, 0, 0, 0, 0, 0, 3, 5, 0, 
    0, 9, 0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 15, 6, 0, 
    0, 9, 0, 0, 0, 3, 0, 0, 0, 0, 5, 0, 4, 10, 0, 
    0, 2, 0, 0, 17, 0, 0, 0, 0, 3, 0, 0, 9, 1, 0, 
    0, 1, 0, 15, 0, 7, 3, 0, 3, 2, 0, 3, 4, 1, 0, 
    1, 0, 6, 0, 13, 0, 0, 0, 5, 7, 6, 9, 3, 4, 1, 
    0, 0, 0, 8, 0, 1, 0, 0, 0, 0, 3, 7, 6, 9, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=333
    22, 25, 20, 16, 21, 25, 25, 20, 23, 13, 11, 17, 17, 12, 11, 
    13, 18, 20, 22, 23, 23, 24, 22, 30, 22, 11, 12, 7, 13, 13, 
    21, 16, 20, 21, 19, 26, 26, 24, 20, 22, 21, 15, 11, 10, 10, 
    9, 18, 19, 18, 19, 21, 20, 19, 17, 17, 21, 24, 15, 14, 11, 
    12, 15, 17, 19, 23, 15, 9, 10, 22, 12, 10, 18, 9, 10, 10, 
    0, 19, 20, 16, 21, 2, 9, 6, 1, 5, 13, 17, 12, 13, 10, 
    12, 0, 9, 11, 11, 10, 11, 7, 13, 6, 15, 15, 15, 16, 12, 
    16, 0, 7, 8, 0, 8, 11, 0, 0, 1, 15, 10, 6, 10, 20, 
    11, 0, 3, 12, 0, 3, 15, 2, 0, 3, 11, 14, 10, 1, 17, 
    13, 2, 0, 22, 0, 0, 10, 2, 22, 15, 13, 16, 9, 0, 17, 
    10, 0, 0, 26, 20, 20, 9, 6, 9, 9, 11, 8, 10, 0, 10, 
    6, 6, 5, 16, 23, 15, 15, 18, 23, 19, 15, 13, 7, 9, 0, 
    7, 6, 12, 7, 8, 3, 6, 18, 17, 19, 24, 21, 19, 13, 12, 
    10, 0, 10, 7, 17, 13, 8, 14, 12, 14, 16, 15, 18, 16, 14, 
    11, 10, 9, 8, 7, 14, 11, 8, 11, 11, 11, 10, 12, 16, 10, 
    
    -- channel=334
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 3, 4, 2, 0, 
    16, 0, 0, 0, 0, 0, 0, 40, 23, 0, 0, 12, 9, 0, 0, 
    0, 11, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 1, 24, 7, 13, 47, 44, 63, 67, 15, 0, 0, 0, 
    0, 0, 0, 8, 70, 17, 21, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 13, 4, 0, 59, 49, 46, 50, 9, 28, 11, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 6, 21, 13, 23, 13, 
    0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    0, 8, 1, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=335
    0, 10, 0, 2, 0, 0, 0, 9, 0, 0, 4, 0, 9, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 3, 9, 0, 1, 
    0, 12, 0, 0, 0, 0, 0, 5, 0, 0, 15, 0, 3, 3, 0, 
    0, 2, 0, 6, 0, 0, 0, 0, 3, 0, 0, 0, 0, 15, 5, 
    0, 9, 0, 1, 0, 0, 0, 0, 0, 18, 1, 0, 14, 0, 3, 
    96, 0, 14, 0, 0, 35, 0, 0, 0, 18, 0, 0, 17, 2, 11, 
    75, 37, 0, 0, 14, 2, 0, 0, 17, 4, 0, 0, 13, 8, 2, 
    0, 80, 0, 0, 27, 0, 0, 14, 0, 0, 0, 0, 24, 22, 0, 
    0, 62, 0, 0, 24, 24, 0, 4, 0, 0, 0, 0, 53, 50, 0, 
    0, 72, 0, 0, 76, 12, 0, 30, 0, 0, 0, 0, 41, 81, 0, 
    0, 44, 0, 0, 30, 17, 1, 37, 0, 0, 0, 10, 21, 85, 0, 
    0, 11, 9, 0, 0, 3, 4, 0, 0, 0, 0, 18, 41, 28, 14, 
    4, 2, 0, 15, 0, 0, 15, 0, 0, 0, 0, 15, 23, 9, 35, 
    0, 30, 0, 8, 0, 11, 21, 0, 0, 0, 0, 10, 0, 8, 0, 
    8, 12, 0, 5, 0, 0, 0, 0, 0, 0, 7, 8, 0, 0, 12, 
    
    -- channel=336
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 12, 11, 12, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=337
    23, 4, 18, 14, 23, 19, 20, 3, 29, 0, 0, 0, 0, 0, 7, 
    21, 35, 10, 18, 21, 20, 24, 13, 34, 0, 0, 0, 0, 9, 0, 
    43, 18, 17, 18, 20, 24, 32, 8, 21, 21, 0, 6, 1, 0, 0, 
    17, 17, 21, 15, 27, 25, 29, 20, 12, 18, 10, 29, 1, 0, 0, 
    2, 13, 21, 19, 24, 28, 15, 15, 24, 3, 9, 54, 0, 0, 0, 
    0, 18, 17, 26, 24, 0, 41, 31, 24, 0, 23, 26, 0, 0, 0, 
    0, 0, 34, 33, 0, 32, 25, 25, 1, 8, 34, 8, 0, 0, 0, 
    15, 0, 35, 12, 2, 31, 23, 20, 25, 26, 57, 16, 0, 0, 18, 
    18, 0, 25, 28, 33, 0, 60, 27, 26, 32, 46, 0, 0, 0, 54, 
    22, 0, 24, 95, 0, 4, 44, 0, 50, 0, 0, 3, 0, 0, 87, 
    28, 0, 32, 69, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 79, 
    8, 10, 2, 24, 14, 0, 0, 25, 0, 0, 0, 0, 0, 0, 13, 
    1, 9, 13, 0, 28, 15, 0, 18, 3, 0, 0, 0, 0, 0, 0, 
    24, 0, 30, 0, 25, 3, 0, 27, 0, 5, 0, 0, 0, 0, 12, 
    4, 5, 12, 2, 3, 16, 16, 11, 10, 1, 0, 2, 11, 18, 0, 
    
    -- channel=338
    32, 17, 6, 10, 11, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 8, 9, 10, 11, 18, 17, 12, 13, 0, 0, 0, 0, 0, 0, 
    4, 0, 11, 6, 12, 11, 22, 2, 13, 41, 11, 11, 0, 0, 1, 
    3, 0, 4, 5, 6, 11, 9, 8, 0, 9, 12, 11, 0, 0, 0, 
    0, 2, 9, 5, 11, 9, 20, 30, 11, 0, 0, 8, 0, 0, 0, 
    0, 14, 12, 8, 0, 4, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 13, 12, 0, 0, 51, 30, 17, 10, 0, 0, 0, 0, 
    2, 0, 8, 0, 5, 24, 21, 0, 0, 11, 30, 0, 0, 9, 1, 
    15, 0, 16, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 28, 
    18, 0, 8, 19, 0, 0, 8, 23, 14, 0, 2, 0, 0, 0, 51, 
    18, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    5, 3, 0, 51, 13, 25, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 5, 0, 0, 27, 9, 16, 24, 16, 4, 0, 0, 0, 0, 0, 
    5, 0, 4, 0, 0, 9, 0, 20, 13, 14, 17, 17, 23, 4, 0, 
    11, 17, 20, 14, 26, 15, 0, 0, 0, 6, 7, 8, 14, 13, 5, 
    
    -- channel=339
    1, 6, 4, 9, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 11, 4, 9, 10, 10, 7, 5, 0, 0, 0, 0, 0, 0, 0, 
    17, 4, 10, 10, 14, 11, 13, 2, 5, 6, 0, 0, 0, 0, 0, 
    4, 5, 10, 13, 16, 15, 15, 9, 5, 9, 6, 2, 0, 0, 0, 
    0, 10, 14, 12, 15, 18, 13, 19, 11, 3, 10, 5, 0, 0, 0, 
    0, 15, 17, 18, 8, 10, 33, 9, 0, 2, 9, 0, 0, 0, 0, 
    0, 4, 27, 23, 10, 28, 12, 23, 15, 18, 9, 0, 0, 0, 0, 
    2, 0, 28, 12, 25, 31, 29, 31, 29, 28, 25, 0, 0, 0, 0, 
    13, 12, 30, 16, 20, 11, 36, 6, 9, 4, 0, 0, 0, 0, 11, 
    16, 8, 35, 27, 0, 15, 12, 17, 20, 0, 0, 0, 0, 0, 27, 
    25, 9, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    11, 23, 7, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 16, 17, 0, 16, 5, 5, 6, 0, 0, 0, 0, 0, 0, 0, 
    20, 5, 19, 7, 3, 2, 11, 17, 1, 1, 0, 0, 0, 0, 0, 
    9, 25, 18, 17, 16, 19, 15, 6, 7, 3, 6, 9, 12, 7, 0, 
    
    -- channel=340
    0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 1, 0, 0, 
    0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 6, 0, 0, 
    44, 0, 12, 0, 0, 19, 0, 0, 0, 14, 0, 0, 15, 0, 5, 
    75, 7, 0, 0, 0, 9, 0, 0, 25, 10, 0, 0, 7, 4, 1, 
    0, 56, 0, 0, 15, 0, 0, 8, 0, 0, 0, 0, 8, 18, 0, 
    0, 39, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 34, 39, 0, 
    0, 47, 0, 0, 67, 5, 0, 23, 0, 0, 0, 0, 27, 61, 0, 
    0, 19, 0, 0, 21, 7, 0, 29, 0, 0, 0, 1, 13, 62, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 18, 23, 17, 0, 
    0, 0, 0, 2, 0, 0, 1, 0, 0, 0, 0, 10, 26, 0, 36, 
    0, 8, 0, 0, 0, 4, 17, 0, 0, 0, 0, 7, 0, 6, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=341
    40, 4, 0, 0, 2, 0, 1, 0, 19, 0, 0, 13, 5, 0, 14, 
    0, 2, 0, 0, 0, 1, 8, 0, 29, 17, 0, 0, 0, 6, 0, 
    16, 0, 0, 0, 0, 0, 11, 0, 0, 45, 0, 14, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 29, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 9, 18, 0, 0, 37, 0, 0, 0, 
    0, 13, 0, 0, 0, 0, 28, 0, 2, 0, 4, 29, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 41, 12, 6, 35, 29, 0, 0, 0, 
    13, 0, 0, 0, 0, 2, 1, 0, 0, 0, 50, 23, 0, 0, 31, 
    3, 0, 0, 4, 0, 0, 12, 0, 0, 0, 6, 12, 0, 0, 69, 
    16, 0, 0, 77, 0, 0, 20, 0, 41, 9, 21, 20, 0, 0, 97, 
    8, 0, 0, 74, 2, 0, 0, 0, 3, 10, 0, 0, 0, 0, 53, 
    0, 0, 0, 44, 30, 13, 4, 26, 27, 9, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 21, 4, 0, 32, 35, 34, 36, 17, 0, 2, 0, 
    0, 0, 1, 0, 5, 0, 0, 16, 5, 15, 16, 7, 23, 1, 2, 
    0, 0, 1, 0, 7, 0, 0, 0, 0, 0, 0, 0, 3, 13, 0, 
    
    -- channel=342
    1, 0, 5, 0, 0, 0, 7, 0, 19, 12, 5, 3, 0, 0, 16, 
    0, 1, 0, 0, 0, 0, 3, 0, 11, 12, 0, 9, 0, 10, 3, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 10, 0, 
    10, 0, 0, 0, 0, 3, 8, 8, 0, 0, 2, 15, 14, 0, 2, 
    14, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 37, 0, 11, 5, 
    0, 0, 0, 0, 10, 0, 0, 21, 33, 0, 15, 45, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 29, 27, 0, 0, 8, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 31, 0, 0, 22, 
    2, 0, 0, 22, 0, 0, 25, 24, 22, 52, 90, 33, 0, 0, 40, 
    18, 0, 0, 71, 0, 0, 50, 0, 32, 36, 1, 2, 0, 0, 34, 
    13, 0, 5, 76, 0, 36, 42, 17, 71, 32, 26, 11, 0, 0, 30, 
    26, 0, 0, 0, 11, 0, 0, 36, 26, 14, 20, 11, 0, 8, 0, 
    0, 2, 0, 4, 6, 24, 0, 3, 0, 0, 0, 0, 0, 13, 0, 
    15, 0, 24, 6, 28, 0, 0, 21, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 9, 0, 0, 0, 10, 20, 14, 11, 0, 0, 2, 11, 0, 
    
    -- channel=343
    0, 4, 18, 20, 14, 23, 19, 31, 0, 31, 27, 18, 23, 28, 8, 
    1, 0, 23, 16, 16, 14, 19, 26, 0, 24, 37, 31, 26, 15, 26, 
    0, 5, 15, 19, 15, 17, 9, 37, 16, 0, 12, 17, 32, 31, 22, 
    2, 11, 13, 19, 14, 21, 18, 24, 32, 19, 23, 2, 28, 34, 27, 
    23, 7, 9, 18, 11, 14, 11, 0, 10, 41, 26, 0, 34, 29, 26, 
    84, 5, 1, 6, 17, 8, 0, 7, 3, 28, 12, 6, 36, 30, 32, 
    56, 35, 0, 0, 12, 0, 0, 0, 0, 0, 0, 6, 31, 25, 28, 
    11, 55, 0, 12, 1, 0, 0, 0, 0, 0, 0, 1, 44, 9, 3, 
    8, 43, 0, 1, 0, 28, 0, 28, 15, 23, 6, 23, 57, 26, 0, 
    12, 48, 0, 0, 70, 23, 0, 1, 0, 28, 17, 9, 54, 37, 0, 
    4, 48, 0, 0, 40, 53, 42, 62, 19, 34, 36, 34, 40, 67, 0, 
    27, 19, 12, 0, 4, 7, 14, 9, 25, 29, 24, 47, 57, 61, 3, 
    27, 23, 16, 26, 0, 18, 26, 0, 0, 7, 7, 16, 35, 43, 37, 
    13, 51, 3, 37, 0, 15, 31, 3, 14, 4, 7, 6, 1, 16, 11, 
    20, 16, 14, 20, 10, 11, 23, 27, 25, 28, 27, 25, 15, 8, 28, 
    
    -- channel=344
    0, 10, 12, 15, 13, 12, 8, 6, 0, 0, 0, 0, 0, 1, 0, 
    24, 20, 10, 18, 19, 16, 11, 12, 0, 0, 0, 0, 5, 3, 0, 
    21, 17, 18, 22, 22, 21, 16, 13, 10, 0, 2, 0, 5, 2, 1, 
    9, 22, 21, 25, 28, 27, 25, 18, 18, 21, 11, 0, 0, 0, 4, 
    12, 23, 24, 23, 25, 24, 13, 16, 11, 20, 20, 1, 0, 0, 2, 
    0, 20, 27, 27, 21, 19, 25, 30, 6, 10, 14, 0, 0, 0, 0, 
    14, 26, 37, 28, 16, 43, 27, 8, 12, 18, 3, 0, 0, 0, 0, 
    8, 29, 37, 27, 36, 38, 34, 46, 42, 36, 14, 0, 0, 0, 0, 
    17, 32, 36, 22, 45, 31, 39, 37, 37, 34, 0, 0, 0, 16, 0, 
    16, 34, 42, 12, 17, 36, 18, 27, 17, 0, 0, 0, 0, 24, 2, 
    26, 33, 42, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 28, 19, 
    19, 31, 24, 2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 9, 19, 
    23, 27, 28, 27, 7, 6, 7, 0, 0, 0, 0, 0, 0, 0, 9, 
    25, 22, 27, 18, 12, 8, 26, 18, 3, 2, 0, 0, 0, 0, 1, 
    16, 31, 22, 23, 15, 26, 25, 15, 15, 9, 14, 18, 17, 9, 3, 
    
    -- channel=345
    27, 35, 1, 9, 8, 0, 1, 0, 0, 0, 2, 5, 4, 0, 3, 
    1, 3, 4, 6, 7, 10, 9, 8, 10, 0, 0, 0, 7, 2, 0, 
    0, 6, 4, 0, 6, 0, 7, 0, 19, 41, 28, 10, 0, 0, 6, 
    0, 1, 0, 2, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 
    0, 1, 5, 0, 0, 5, 8, 27, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 7, 4, 0, 32, 17, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 14, 0, 0, 48, 50, 28, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 19, 13, 13, 13, 2, 13, 12, 0, 1, 35, 0, 
    7, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 5, 
    0, 0, 5, 0, 0, 0, 0, 49, 0, 0, 11, 20, 0, 23, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 12, 
    0, 1, 0, 41, 22, 40, 29, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 8, 13, 23, 29, 29, 21, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 1, 16, 22, 30, 40, 35, 20, 6, 
    2, 9, 0, 11, 19, 6, 0, 0, 0, 0, 6, 8, 7, 6, 12, 
    
    -- channel=346
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=347
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=348
    18, 10, 0, 0, 0, 0, 0, 0, 14, 7, 0, 9, 6, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 18, 0, 0, 0, 0, 1, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 23, 1, 6, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 14, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 9, 0, 2, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 16, 3, 5, 15, 20, 8, 3, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 21, 7, 0, 16, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 3, 17, 2, 0, 32, 
    0, 0, 0, 32, 0, 0, 0, 0, 10, 11, 15, 13, 0, 0, 37, 
    0, 0, 0, 25, 17, 0, 0, 0, 0, 18, 8, 0, 3, 0, 16, 
    0, 0, 0, 18, 14, 7, 2, 10, 24, 19, 22, 13, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 7, 25, 29, 33, 26, 6, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 5, 15, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=349
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=350
    34, 10, 27, 24, 30, 31, 33, 30, 19, 19, 17, 19, 17, 9, 16, 
    19, 22, 36, 27, 27, 30, 36, 34, 33, 23, 15, 14, 12, 16, 19, 
    13, 16, 29, 30, 29, 35, 34, 37, 35, 24, 7, 20, 16, 21, 16, 
    30, 13, 27, 28, 27, 38, 31, 36, 29, 31, 37, 26, 23, 19, 17, 
    22, 14, 24, 34, 27, 29, 22, 15, 23, 27, 30, 18, 18, 17, 17, 
    34, 24, 13, 22, 33, 17, 0, 0, 23, 14, 15, 26, 9, 20, 16, 
    0, 24, 7, 14, 24, 0, 20, 5, 0, 0, 12, 17, 11, 16, 14, 
    17, 5, 7, 15, 4, 0, 16, 0, 0, 0, 0, 11, 17, 3, 12, 
    15, 7, 0, 19, 0, 27, 3, 19, 12, 12, 24, 24, 15, 2, 8, 
    25, 8, 0, 7, 0, 8, 20, 0, 13, 28, 13, 3, 11, 0, 0, 
    14, 17, 0, 20, 17, 19, 25, 16, 30, 26, 13, 13, 14, 4, 0, 
    27, 11, 10, 8, 16, 9, 6, 17, 25, 14, 7, 12, 20, 18, 5, 
    22, 20, 17, 10, 16, 21, 19, 16, 12, 12, 9, 7, 4, 31, 4, 
    12, 22, 14, 29, 13, 14, 10, 21, 17, 8, 14, 5, 13, 10, 8, 
    20, 7, 21, 14, 19, 9, 19, 22, 23, 24, 20, 18, 19, 18, 19, 
    
    -- channel=351
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=352
    0, 6, 0, 3, 3, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 1, 8, 0, 2, 0, 4, 0, 0, 
    0, 24, 0, 0, 0, 0, 2, 0, 0, 2, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 0, 4, 0, 0, 0, 6, 0, 0, 5, 0, 0, 
    8, 0, 0, 4, 0, 10, 0, 28, 47, 9, 0, 0, 0, 7, 0, 
    0, 5, 0, 0, 0, 0, 0, 15, 0, 6, 8, 0, 0, 36, 0, 
    1, 1, 0, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 
    0, 0, 4, 1, 7, 0, 0, 62, 0, 0, 0, 23, 0, 30, 43, 
    0, 0, 4, 0, 7, 0, 0, 10, 0, 0, 0, 9, 0, 0, 48, 
    0, 7, 0, 10, 0, 4, 0, 6, 0, 0, 2, 0, 0, 0, 36, 
    0, 0, 0, 0, 0, 0, 13, 0, 0, 2, 8, 17, 6, 0, 21, 
    6, 0, 0, 0, 0, 18, 7, 0, 0, 0, 0, 21, 1, 0, 11, 
    10, 13, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    
    -- channel=353
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 18, 0, 7, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 17, 2, 7, 8, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 22, 9, 10, 14, 6, 7, 0, 0, 5, 0, 0, 0, 0, 0, 
    3, 12, 13, 7, 14, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 17, 14, 10, 8, 28, 26, 2, 0, 0, 0, 0, 0, 0, 
    0, 5, 33, 22, 0, 36, 23, 6, 13, 8, 0, 0, 0, 0, 0, 
    0, 4, 30, 17, 24, 39, 15, 36, 39, 37, 15, 0, 0, 0, 0, 
    0, 6, 28, 2, 47, 6, 28, 22, 23, 18, 2, 0, 0, 3, 0, 
    0, 4, 36, 14, 22, 14, 14, 23, 3, 0, 0, 0, 0, 10, 25, 
    5, 0, 36, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 47, 
    0, 2, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 6, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 2, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=354
    29, 16, 0, 0, 4, 0, 2, 3, 0, 0, 3, 12, 21, 0, 0, 
    0, 0, 6, 5, 6, 9, 1, 6, 17, 4, 0, 0, 0, 0, 7, 
    0, 7, 3, 1, 5, 1, 9, 0, 8, 32, 21, 0, 0, 0, 2, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 12, 5, 3, 10, 0, 
    0, 6, 0, 3, 4, 0, 9, 27, 0, 0, 0, 0, 0, 0, 0, 
    24, 15, 26, 0, 0, 31, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 0, 0, 48, 48, 17, 0, 4, 5, 5, 0, 
    0, 3, 0, 0, 9, 5, 0, 0, 0, 2, 0, 0, 1, 27, 0, 
    4, 5, 6, 0, 0, 7, 0, 0, 0, 0, 0, 0, 9, 11, 0, 
    7, 10, 0, 0, 0, 0, 0, 22, 0, 0, 24, 3, 0, 18, 5, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 2, 41, 5, 31, 8, 0, 8, 5, 0, 0, 5, 0, 1, 
    0, 4, 0, 0, 0, 0, 22, 16, 22, 27, 26, 32, 0, 12, 0, 
    0, 0, 0, 0, 0, 19, 0, 3, 20, 9, 23, 24, 24, 7, 0, 
    21, 6, 7, 6, 14, 2, 0, 0, 0, 5, 3, 6, 4, 3, 14, 
    
    -- channel=355
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 13, 0, 0, 12, 14, 29, 18, 0, 0, 0, 0, 
    0, 0, 0, 6, 18, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 25, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=356
    0, 24, 10, 21, 16, 19, 14, 16, 0, 7, 14, 9, 13, 18, 0, 
    5, 9, 7, 18, 23, 17, 11, 21, 5, 0, 23, 13, 18, 7, 7, 
    0, 30, 12, 17, 18, 15, 14, 17, 16, 0, 25, 0, 15, 13, 10, 
    0, 23, 14, 19, 14, 13, 11, 8, 21, 15, 2, 0, 12, 18, 13, 
    4, 20, 15, 14, 17, 11, 6, 17, 0, 26, 7, 0, 20, 13, 15, 
    42, 4, 27, 12, 6, 27, 0, 6, 0, 24, 2, 0, 27, 13, 19, 
    55, 20, 6, 6, 6, 20, 0, 0, 28, 9, 0, 0, 17, 19, 16, 
    0, 54, 0, 3, 20, 0, 0, 18, 0, 2, 0, 0, 14, 33, 0, 
    4, 39, 2, 0, 44, 1, 0, 15, 12, 0, 0, 0, 29, 40, 0, 
    1, 44, 2, 0, 68, 11, 0, 48, 0, 0, 1, 14, 29, 56, 0, 
    0, 24, 4, 0, 22, 17, 10, 36, 0, 0, 10, 22, 18, 55, 0, 
    0, 15, 14, 0, 0, 10, 13, 2, 0, 11, 10, 21, 29, 18, 29, 
    8, 12, 2, 19, 0, 0, 18, 0, 0, 3, 5, 20, 29, 2, 36, 
    7, 17, 0, 1, 2, 19, 26, 0, 8, 3, 7, 22, 6, 15, 15, 
    15, 19, 1, 10, 0, 17, 9, 8, 7, 2, 17, 18, 4, 5, 11, 
    
    -- channel=357
    5, 61, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 4, 4, 2, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 37, 44, 16, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 8, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 0, 0, 0, 3, 3, 0, 25, 60, 33, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 16, 0, 0, 0, 6, 0, 0, 25, 7, 
    2, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 2, 0, 0, 0, 0, 0, 30, 9, 0, 1, 23, 3, 12, 5, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 3, 0, 31, 33, 48, 49, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 23, 33, 33, 27, 25, 13, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 28, 31, 52, 42, 37, 0, 
    0, 21, 0, 12, 13, 7, 0, 0, 0, 0, 2, 1, 4, 0, 12, 
    
    -- channel=358
    0, 2, 7, 4, 4, 14, 6, 15, 0, 9, 3, 0, 3, 10, 0, 
    0, 0, 4, 7, 7, 2, 3, 8, 0, 6, 16, 9, 3, 0, 0, 
    0, 9, 7, 8, 5, 8, 1, 17, 0, 0, 0, 0, 10, 4, 0, 
    0, 16, 8, 8, 11, 8, 7, 3, 16, 4, 1, 0, 3, 9, 5, 
    8, 6, 5, 11, 7, 0, 0, 0, 1, 19, 2, 0, 11, 8, 5, 
    33, 0, 4, 2, 9, 0, 0, 19, 0, 4, 0, 0, 19, 8, 11, 
    52, 11, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 11, 9, 11, 
    0, 34, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 13, 0, 0, 23, 12, 0, 35, 22, 31, 8, 4, 27, 14, 0, 
    0, 25, 0, 0, 60, 14, 0, 0, 0, 1, 0, 0, 24, 17, 0, 
    0, 22, 4, 0, 30, 54, 22, 52, 0, 2, 19, 5, 10, 45, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 5, 11, 5, 30, 23, 43, 0, 
    0, 0, 8, 13, 0, 0, 0, 0, 0, 0, 0, 0, 26, 6, 42, 
    0, 15, 0, 13, 0, 2, 13, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 1, 5, 1, 3, 0, 0, 0, 0, 0, 0, 
    
    -- channel=359
    0, 2, 6, 16, 5, 11, 4, 14, 0, 14, 16, 3, 10, 22, 0, 
    1, 0, 6, 8, 10, 5, 2, 15, 0, 0, 30, 21, 23, 4, 11, 
    0, 13, 6, 11, 9, 5, 0, 20, 3, 0, 10, 0, 23, 20, 12, 
    0, 11, 6, 15, 7, 11, 8, 8, 24, 11, 0, 0, 14, 24, 18, 
    10, 12, 6, 8, 8, 5, 4, 1, 0, 39, 15, 0, 27, 19, 19, 
    86, 0, 10, 2, 3, 14, 0, 12, 0, 28, 1, 0, 31, 17, 25, 
    67, 41, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 19, 16, 19, 
    0, 71, 0, 5, 15, 0, 0, 8, 0, 0, 0, 0, 30, 16, 0, 
    2, 54, 0, 0, 28, 22, 0, 30, 25, 19, 0, 1, 48, 41, 0, 
    0, 59, 0, 0, 94, 31, 0, 28, 0, 0, 0, 0, 46, 59, 0, 
    0, 47, 0, 0, 22, 37, 33, 63, 0, 5, 21, 28, 28, 79, 0, 
    11, 20, 13, 0, 0, 0, 6, 0, 0, 8, 6, 31, 49, 47, 20, 
    22, 17, 6, 30, 0, 7, 24, 0, 0, 0, 0, 2, 26, 17, 39, 
    9, 47, 0, 20, 0, 13, 34, 0, 4, 0, 0, 4, 0, 9, 2, 
    15, 21, 6, 15, 0, 11, 16, 19, 13, 15, 22, 21, 4, 0, 17, 
    
    -- channel=360
    5, 0, 0, 0, 0, 0, 5, 0, 19, 0, 0, 0, 0, 0, 5, 
    0, 10, 0, 0, 0, 0, 0, 0, 15, 3, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 0, 2, 3, 0, 0, 0, 0, 0, 0, 1, 0, 
    16, 0, 0, 0, 0, 4, 9, 5, 0, 0, 0, 15, 7, 0, 0, 
    12, 0, 0, 0, 0, 4, 1, 0, 9, 0, 0, 43, 0, 1, 0, 
    0, 1, 0, 0, 18, 0, 0, 24, 34, 0, 16, 52, 0, 0, 0, 
    0, 0, 3, 5, 0, 0, 25, 0, 0, 0, 28, 20, 0, 0, 0, 
    4, 0, 9, 3, 0, 0, 0, 0, 0, 0, 17, 20, 0, 0, 9, 
    0, 0, 0, 20, 1, 4, 33, 39, 34, 62, 108, 31, 0, 0, 39, 
    15, 0, 0, 82, 0, 0, 57, 0, 25, 31, 0, 0, 0, 0, 45, 
    6, 0, 19, 92, 0, 48, 44, 23, 78, 21, 19, 2, 0, 0, 52, 
    17, 0, 2, 0, 0, 0, 0, 28, 23, 7, 7, 0, 0, 0, 15, 
    0, 0, 0, 8, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 20, 0, 33, 0, 0, 13, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 2, 12, 5, 0, 0, 0, 0, 3, 0, 
    
    -- channel=361
    15, 0, 16, 15, 18, 16, 16, 10, 0, 1, 2, 0, 0, 0, 0, 
    9, 16, 19, 17, 21, 20, 17, 19, 11, 0, 3, 1, 1, 0, 1, 
    6, 20, 17, 23, 22, 23, 23, 24, 21, 0, 0, 0, 0, 6, 0, 
    8, 14, 19, 21, 17, 24, 21, 19, 23, 20, 15, 2, 7, 4, 2, 
    12, 12, 17, 20, 23, 20, 18, 12, 4, 21, 14, 1, 5, 3, 4, 
    30, 12, 17, 17, 24, 23, 0, 0, 10, 13, 2, 4, 6, 3, 4, 
    0, 21, 6, 10, 15, 0, 6, 0, 0, 0, 0, 0, 0, 3, 1, 
    0, 15, 3, 11, 6, 5, 1, 0, 0, 0, 0, 0, 3, 6, 0, 
    0, 6, 1, 0, 4, 17, 0, 6, 4, 0, 5, 0, 1, 6, 0, 
    6, 8, 0, 0, 29, 0, 5, 13, 0, 4, 0, 0, 2, 11, 0, 
    0, 5, 0, 0, 0, 6, 13, 6, 12, 0, 0, 7, 0, 11, 0, 
    10, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 15, 
    4, 8, 0, 20, 0, 1, 8, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 11, 0, 0, 9, 5, 3, 1, 0, 0, 0, 0, 0, 0, 3, 
    9, 0, 5, 0, 0, 0, 3, 9, 3, 3, 5, 8, 2, 4, 2, 
    
    -- channel=362
    0, 0, 0, 0, 0, 0, 0, 5, 0, 15, 4, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 16, 1, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 6, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 5, 6, 6, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 23, 9, 0, 12, 12, 6, 
    79, 0, 0, 0, 7, 0, 0, 33, 0, 3, 0, 4, 19, 9, 11, 
    28, 38, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 10, 0, 8, 
    0, 45, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 
    0, 18, 0, 4, 2, 44, 0, 48, 43, 63, 45, 18, 35, 10, 0, 
    0, 40, 0, 0, 111, 23, 0, 0, 0, 25, 0, 0, 31, 24, 0, 
    0, 42, 9, 0, 4, 85, 53, 65, 42, 17, 34, 20, 6, 70, 0, 
    16, 0, 19, 0, 0, 0, 0, 0, 10, 17, 9, 32, 41, 58, 18, 
    0, 4, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 12, 20, 26, 
    0, 39, 0, 18, 5, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 13, 3, 5, 0, 0, 0, 0, 0, 
    
    -- channel=363
    32, 39, 0, 1, 4, 1, 1, 1, 9, 0, 0, 13, 9, 0, 8, 
    0, 0, 1, 3, 1, 8, 12, 6, 26, 11, 0, 0, 0, 5, 0, 
    2, 0, 3, 0, 0, 0, 11, 0, 8, 60, 28, 20, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 23, 9, 0, 0, 11, 0, 0, 0, 
    0, 11, 4, 0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 53, 48, 31, 15, 10, 0, 0, 0, 
    13, 0, 0, 0, 0, 4, 15, 0, 0, 2, 38, 6, 0, 16, 20, 
    9, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 
    9, 0, 0, 31, 0, 0, 0, 6, 31, 0, 16, 25, 0, 0, 65, 
    6, 0, 0, 10, 17, 0, 0, 0, 0, 0, 0, 0, 4, 0, 20, 
    0, 3, 0, 56, 33, 42, 34, 12, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 22, 0, 2, 37, 45, 43, 40, 28, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 10, 17, 28, 33, 39, 43, 26, 0, 
    0, 12, 1, 8, 21, 6, 0, 0, 0, 0, 1, 0, 9, 11, 8, 
    
    -- channel=364
    0, 46, 2, 9, 0, 3, 0, 14, 0, 2, 4, 4, 11, 21, 0, 
    0, 0, 7, 6, 8, 6, 0, 11, 0, 0, 10, 0, 10, 0, 3, 
    0, 3, 8, 5, 9, 0, 0, 11, 4, 3, 39, 5, 3, 0, 8, 
    0, 7, 0, 11, 0, 0, 0, 0, 6, 0, 7, 0, 0, 16, 5, 
    0, 9, 2, 8, 1, 4, 1, 19, 0, 9, 1, 0, 7, 0, 3, 
    53, 7, 19, 5, 0, 45, 0, 0, 0, 25, 0, 0, 11, 0, 8, 
    79, 14, 0, 0, 26, 13, 0, 6, 54, 31, 0, 0, 12, 8, 2, 
    0, 66, 0, 0, 36, 0, 8, 16, 0, 0, 0, 0, 18, 37, 0, 
    0, 64, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 44, 44, 0, 
    0, 64, 0, 0, 19, 7, 0, 43, 0, 0, 2, 2, 38, 73, 0, 
    0, 32, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 30, 67, 0, 
    0, 16, 2, 0, 4, 29, 32, 0, 0, 0, 0, 6, 19, 16, 0, 
    12, 4, 3, 0, 0, 0, 17, 0, 3, 16, 10, 25, 31, 5, 14, 
    0, 16, 0, 9, 0, 14, 24, 0, 11, 8, 14, 37, 19, 29, 0, 
    5, 29, 0, 18, 12, 9, 0, 0, 0, 0, 13, 16, 4, 0, 24, 
    
    -- channel=365
    26, 45, 9, 15, 12, 11, 10, 10, 6, 1, 3, 13, 3, 6, 13, 
    14, 12, 13, 10, 9, 16, 23, 20, 16, 4, 0, 0, 11, 13, 2, 
    8, 0, 15, 5, 8, 9, 17, 1, 18, 54, 28, 28, 3, 0, 14, 
    2, 1, 5, 5, 9, 11, 5, 12, 2, 9, 12, 15, 0, 0, 1, 
    0, 3, 11, 6, 4, 6, 8, 19, 14, 0, 3, 17, 0, 0, 2, 
    0, 10, 0, 9, 0, 0, 34, 0, 8, 0, 2, 0, 0, 2, 0, 
    0, 0, 4, 10, 6, 7, 0, 41, 26, 25, 16, 7, 0, 3, 0, 
    15, 0, 6, 0, 10, 15, 32, 1, 4, 11, 34, 14, 0, 17, 17, 
    15, 2, 7, 10, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 36, 
    10, 0, 1, 34, 0, 5, 0, 24, 29, 0, 11, 25, 0, 0, 48, 
    17, 0, 0, 1, 6, 0, 0, 0, 0, 2, 0, 0, 13, 0, 13, 
    0, 13, 0, 48, 37, 46, 41, 9, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 7, 0, 38, 25, 8, 33, 40, 31, 24, 15, 0, 0, 0, 
    2, 0, 5, 11, 0, 10, 0, 19, 17, 36, 36, 41, 43, 32, 1, 
    0, 23, 11, 18, 30, 16, 3, 0, 9, 4, 13, 10, 18, 17, 16, 
    
    -- channel=366
    23, 28, 41, 40, 45, 50, 48, 40, 18, 11, 13, 13, 13, 14, 6, 
    23, 29, 43, 44, 48, 49, 54, 57, 41, 11, 14, 18, 21, 19, 16, 
    15, 24, 40, 46, 43, 53, 53, 54, 48, 23, 26, 25, 26, 23, 19, 
    11, 25, 39, 42, 46, 58, 52, 47, 45, 48, 43, 27, 25, 23, 21, 
    18, 24, 36, 43, 47, 39, 22, 18, 30, 44, 32, 10, 16, 19, 20, 
    20, 28, 27, 31, 37, 5, 0, 0, 11, 17, 17, 4, 9, 17, 20, 
    12, 19, 12, 16, 14, 7, 15, 0, 0, 0, 0, 0, 1, 15, 17, 
    22, 18, 11, 12, 2, 4, 23, 2, 0, 0, 0, 0, 1, 6, 5, 
    28, 16, 1, 6, 1, 16, 13, 24, 17, 12, 5, 0, 5, 6, 0, 
    33, 17, 0, 0, 1, 6, 16, 17, 21, 6, 0, 1, 11, 3, 0, 
    29, 24, 0, 1, 7, 7, 18, 33, 13, 1, 0, 4, 11, 12, 0, 
    35, 26, 7, 4, 25, 19, 22, 14, 0, 0, 0, 0, 9, 20, 5, 
    38, 33, 21, 15, 5, 23, 28, 19, 5, 0, 0, 0, 2, 11, 8, 
    25, 31, 25, 27, 16, 25, 33, 33, 19, 16, 19, 18, 16, 19, 15, 
    34, 32, 32, 30, 24, 35, 37, 34, 35, 33, 35, 34, 30, 27, 23, 
    
    -- channel=367
    19, 48, 0, 5, 1, 0, 0, 0, 0, 0, 0, 1, 6, 1, 0, 
    0, 0, 1, 2, 2, 10, 4, 4, 0, 0, 0, 0, 1, 0, 0, 
    0, 1, 2, 0, 0, 0, 2, 0, 10, 41, 37, 7, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 1, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 0, 27, 3, 0, 0, 1, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 18, 0, 0, 40, 60, 30, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 17, 8, 11, 1, 0, 1, 1, 0, 0, 34, 0, 
    3, 18, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 11, 0, 
    0, 2, 0, 0, 0, 0, 0, 45, 0, 0, 11, 14, 3, 24, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 49, 14, 51, 39, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 10, 19, 29, 30, 21, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 16, 21, 35, 48, 41, 27, 0, 
    0, 13, 0, 11, 19, 3, 0, 0, 0, 0, 5, 4, 3, 0, 14, 
    
    -- channel=368
    63, 65, 68, 71, 74, 75, 72, 62, 51, 39, 48, 47, 50, 49, 43, 
    53, 61, 68, 74, 79, 79, 79, 80, 73, 41, 46, 50, 54, 54, 50, 
    54, 63, 67, 73, 74, 79, 80, 77, 77, 62, 65, 56, 58, 55, 53, 
    41, 60, 67, 71, 72, 78, 78, 70, 70, 76, 69, 60, 57, 57, 55, 
    45, 60, 67, 69, 77, 70, 61, 67, 62, 69, 60, 48, 47, 51, 54, 
    40, 64, 71, 66, 63, 56, 42, 36, 40, 56, 53, 38, 44, 48, 52, 
    44, 48, 55, 56, 53, 50, 46, 52, 58, 47, 42, 34, 37, 49, 50, 
    55, 54, 53, 49, 47, 55, 59, 53, 41, 45, 42, 27, 32, 56, 45, 
    68, 55, 53, 36, 44, 45, 53, 47, 41, 32, 29, 29, 33, 50, 35, 
    70, 58, 40, 35, 39, 36, 51, 72, 60, 34, 37, 44, 38, 52, 40, 
    68, 53, 40, 47, 34, 29, 41, 56, 41, 28, 26, 41, 43, 45, 43, 
    65, 62, 50, 58, 62, 59, 60, 50, 27, 24, 21, 21, 38, 38, 50, 
    68, 71, 52, 51, 45, 54, 68, 64, 46, 39, 35, 35, 38, 37, 45, 
    63, 60, 62, 46, 52, 63, 69, 68, 60, 55, 58, 61, 57, 55, 55, 
    74, 70, 69, 68, 62, 75, 68, 65, 64, 64, 68, 70, 66, 64, 57, 
    
    -- channel=369
    0, 14, 0, 0, 0, 0, 0, 8, 0, 4, 4, 0, 4, 17, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 19, 7, 11, 0, 1, 
    0, 8, 0, 2, 0, 0, 0, 9, 0, 0, 17, 0, 6, 3, 0, 
    0, 13, 0, 8, 0, 0, 0, 0, 8, 0, 0, 0, 0, 11, 4, 
    4, 7, 0, 2, 0, 0, 0, 0, 0, 19, 0, 0, 14, 4, 4, 
    87, 0, 8, 0, 0, 26, 0, 0, 0, 21, 0, 0, 22, 3, 12, 
    80, 35, 0, 0, 12, 6, 0, 0, 14, 6, 0, 0, 14, 7, 5, 
    0, 79, 0, 7, 26, 0, 0, 12, 0, 0, 0, 0, 29, 20, 0, 
    0, 63, 0, 0, 13, 24, 0, 5, 0, 0, 0, 0, 52, 47, 0, 
    0, 67, 0, 0, 91, 22, 0, 25, 0, 0, 0, 0, 46, 78, 0, 
    0, 44, 0, 0, 20, 15, 0, 36, 0, 0, 1, 11, 23, 91, 0, 
    0, 6, 9, 0, 0, 0, 10, 0, 0, 0, 0, 20, 40, 37, 5, 
    3, 4, 0, 25, 0, 0, 9, 0, 0, 0, 0, 9, 28, 7, 29, 
    0, 32, 0, 7, 0, 6, 25, 0, 0, 0, 0, 9, 0, 9, 0, 
    1, 10, 0, 6, 0, 1, 0, 0, 0, 0, 8, 10, 0, 0, 10, 
    
    -- channel=370
    73, 67, 79, 81, 82, 81, 81, 68, 54, 47, 49, 46, 46, 49, 47, 
    74, 79, 82, 81, 87, 89, 88, 87, 72, 43, 47, 54, 57, 54, 53, 
    65, 76, 80, 87, 86, 91, 90, 88, 89, 63, 60, 58, 56, 60, 56, 
    61, 70, 82, 86, 87, 95, 91, 86, 84, 86, 74, 64, 57, 56, 57, 
    63, 72, 81, 82, 92, 85, 74, 72, 67, 82, 76, 61, 55, 56, 57, 
    63, 66, 76, 81, 80, 74, 49, 52, 64, 64, 58, 46, 47, 53, 55, 
    41, 73, 68, 69, 69, 58, 65, 54, 47, 45, 47, 37, 38, 51, 51, 
    51, 62, 67, 65, 63, 71, 73, 61, 52, 54, 47, 35, 40, 55, 43, 
    69, 60, 63, 53, 57, 63, 66, 62, 62, 53, 47, 34, 37, 53, 39, 
    66, 59, 53, 42, 57, 57, 67, 77, 52, 41, 38, 37, 43, 55, 35, 
    69, 60, 50, 50, 20, 32, 53, 54, 61, 36, 31, 46, 43, 54, 45, 
    73, 60, 58, 61, 57, 56, 54, 42, 27, 24, 21, 21, 43, 46, 61, 
    74, 70, 54, 69, 67, 63, 66, 58, 41, 29, 21, 25, 32, 42, 37, 
    64, 68, 68, 56, 64, 60, 66, 69, 59, 54, 55, 54, 53, 53, 54, 
    71, 66, 72, 69, 65, 69, 71, 72, 67, 66, 70, 71, 68, 65, 62, 
    
    -- channel=371
    48, 52, 55, 55, 54, 51, 46, 41, 31, 22, 25, 21, 23, 32, 23, 
    65, 64, 54, 60, 63, 60, 52, 50, 39, 15, 24, 30, 35, 32, 29, 
    60, 64, 61, 66, 67, 66, 58, 57, 56, 32, 41, 31, 33, 35, 34, 
    52, 66, 64, 69, 67, 68, 63, 56, 59, 59, 50, 35, 29, 32, 36, 
    54, 64, 66, 67, 72, 70, 59, 59, 47, 58, 57, 36, 29, 34, 35, 
    46, 61, 73, 70, 67, 78, 61, 60, 44, 52, 46, 20, 26, 27, 33, 
    44, 70, 75, 68, 67, 74, 66, 50, 59, 55, 37, 14, 18, 27, 29, 
    33, 68, 72, 69, 80, 81, 70, 77, 75, 73, 43, 14, 20, 43, 23, 
    45, 67, 74, 53, 72, 73, 64, 59, 61, 53, 26, 3, 19, 55, 20, 
    44, 70, 76, 30, 65, 64, 49, 67, 36, 17, 9, 9, 23, 69, 30, 
    50, 61, 66, 26, 6, 24, 26, 43, 30, 4, 7, 17, 20, 65, 50, 
    51, 52, 63, 44, 32, 26, 30, 21, 0, 0, 0, 0, 19, 34, 59, 
    51, 57, 48, 72, 46, 38, 42, 31, 13, 4, 0, 2, 16, 14, 34, 
    48, 53, 52, 41, 46, 40, 53, 43, 37, 30, 27, 33, 29, 30, 36, 
    49, 54, 51, 51, 47, 53, 51, 48, 42, 39, 45, 51, 47, 41, 38, 
    
    -- channel=372
    7, 4, 0, 0, 0, 0, 0, 6, 2, 0, 0, 10, 18, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 2, 12, 3, 1, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 2, 7, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 13, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 16, 16, 3, 0, 0, 4, 3, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 5, 10, 4, 0, 
    5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 3, 0, 
    0, 0, 0, 0, 30, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 2, 14, 4, 0, 10, 5, 0, 0, 5, 0, 0, 
    0, 2, 4, 0, 0, 0, 8, 5, 12, 19, 24, 26, 2, 14, 3, 
    0, 0, 0, 0, 0, 14, 0, 0, 8, 1, 15, 12, 13, 4, 0, 
    15, 2, 0, 0, 4, 2, 0, 0, 0, 4, 0, 0, 0, 0, 1, 
    
    -- channel=373
    50, 0, 0, 0, 0, 0, 6, 0, 42, 0, 0, 0, 0, 0, 24, 
    0, 13, 0, 0, 0, 0, 0, 0, 36, 7, 0, 0, 0, 0, 0, 
    29, 0, 0, 0, 0, 0, 3, 0, 0, 23, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 80, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 14, 3, 48, 0, 6, 83, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 41, 12, 0, 0, 58, 45, 0, 0, 0, 
    8, 0, 8, 0, 0, 0, 0, 0, 0, 0, 67, 48, 0, 0, 28, 
    0, 0, 0, 26, 0, 0, 45, 6, 6, 34, 136, 45, 0, 0, 107, 
    17, 0, 0, 154, 0, 0, 95, 0, 49, 41, 0, 0, 0, 0, 137, 
    8, 0, 5, 178, 0, 1, 22, 0, 97, 25, 6, 0, 0, 0, 121, 
    14, 0, 0, 16, 20, 0, 0, 37, 35, 7, 9, 0, 0, 0, 1, 
    0, 0, 0, 0, 24, 7, 0, 20, 13, 0, 3, 0, 0, 0, 0, 
    0, 0, 28, 0, 43, 0, 0, 26, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    
    -- channel=374
    57, 52, 66, 65, 69, 67, 65, 56, 43, 36, 38, 35, 35, 37, 34, 
    58, 65, 67, 68, 72, 73, 72, 70, 61, 34, 36, 41, 44, 42, 41, 
    55, 62, 66, 72, 73, 76, 76, 75, 73, 48, 46, 45, 46, 48, 44, 
    50, 58, 67, 71, 72, 79, 76, 73, 70, 71, 62, 52, 46, 45, 45, 
    48, 58, 67, 71, 75, 76, 63, 61, 55, 68, 65, 49, 43, 45, 45, 
    46, 57, 65, 69, 69, 67, 38, 44, 50, 54, 49, 38, 36, 42, 44, 
    35, 60, 58, 58, 58, 49, 49, 43, 39, 39, 36, 27, 26, 40, 41, 
    44, 52, 54, 55, 53, 55, 59, 54, 42, 43, 34, 24, 27, 43, 34, 
    55, 51, 52, 44, 48, 54, 52, 54, 51, 43, 36, 25, 26, 45, 27, 
    56, 53, 44, 31, 48, 47, 52, 61, 46, 34, 25, 26, 30, 50, 25, 
    56, 52, 42, 36, 19, 28, 39, 50, 46, 26, 22, 32, 33, 46, 34, 
    59, 51, 48, 41, 43, 38, 42, 39, 20, 16, 14, 15, 33, 36, 49, 
    58, 60, 45, 57, 51, 52, 54, 44, 28, 19, 12, 16, 24, 32, 36, 
    54, 55, 54, 46, 47, 48, 54, 55, 46, 38, 38, 40, 39, 39, 43, 
    57, 53, 57, 55, 50, 56, 59, 58, 54, 52, 55, 58, 55, 52, 48, 
    
    -- channel=375
    13, 24, 24, 13, 21, 29, 21, 29, 17, 17, 11, 18, 20, 14, 3, 
    11, 16, 25, 26, 23, 22, 25, 24, 22, 27, 16, 10, 5, 12, 12, 
    19, 15, 26, 24, 21, 30, 26, 31, 12, 10, 15, 15, 15, 9, 9, 
    17, 26, 24, 21, 25, 26, 21, 21, 20, 18, 32, 20, 17, 17, 13, 
    20, 15, 20, 31, 23, 16, 8, 3, 28, 17, 12, 6, 10, 11, 11, 
    15, 34, 20, 18, 31, 0, 3, 2, 0, 7, 14, 16, 14, 14, 14, 
    33, 4, 11, 10, 14, 18, 13, 0, 0, 8, 11, 10, 18, 17, 15, 
    24, 13, 5, 14, 2, 0, 13, 0, 0, 0, 0, 2, 14, 1, 19, 
    1, 7, 0, 18, 1, 25, 7, 18, 5, 15, 12, 15, 23, 6, 0, 
    15, 15, 0, 8, 0, 3, 3, 0, 27, 19, 6, 4, 17, 0, 0, 
    4, 15, 5, 6, 47, 44, 17, 31, 0, 12, 15, 0, 16, 14, 0, 
    9, 10, 6, 0, 21, 0, 12, 20, 26, 17, 10, 26, 15, 32, 0, 
    8, 9, 25, 6, 0, 5, 2, 3, 6, 14, 19, 18, 26, 25, 29, 
    9, 10, 4, 26, 5, 15, 14, 6, 5, 5, 7, 6, 10, 15, 6, 
    7, 11, 4, 5, 6, 14, 14, 5, 16, 12, 10, 10, 11, 12, 7, 
    
    -- channel=376
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=377
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=378
    3, 31, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 5, 6, 10, 6, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 1, 4, 3, 6, 5, 4, 15, 18, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 3, 0, 0, 8, 26, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 4, 15, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 18, 12, 6, 0, 
    0, 5, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=379
    45, 0, 0, 0, 11, 0, 12, 0, 23, 0, 0, 4, 0, 0, 18, 
    0, 15, 0, 0, 2, 3, 8, 3, 33, 0, 0, 0, 0, 7, 0, 
    13, 0, 0, 0, 0, 3, 15, 0, 14, 35, 0, 2, 0, 0, 0, 
    18, 0, 0, 0, 0, 1, 4, 2, 0, 8, 2, 15, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 4, 0, 0, 0, 44, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 12, 0, 37, 0, 0, 37, 0, 0, 0, 
    0, 0, 2, 11, 0, 0, 23, 45, 0, 0, 30, 23, 0, 0, 0, 
    8, 0, 10, 0, 0, 13, 0, 0, 0, 13, 43, 19, 0, 0, 6, 
    9, 0, 0, 0, 0, 0, 12, 0, 0, 0, 56, 23, 0, 0, 59, 
    22, 0, 0, 71, 0, 0, 53, 2, 21, 15, 10, 9, 0, 0, 95, 
    12, 0, 0, 105, 0, 0, 6, 0, 42, 3, 0, 9, 0, 0, 90, 
    13, 0, 0, 36, 18, 8, 0, 26, 9, 0, 6, 0, 0, 0, 26, 
    0, 3, 0, 0, 11, 14, 2, 26, 23, 12, 10, 0, 0, 0, 0, 
    0, 0, 18, 0, 31, 0, 0, 28, 5, 9, 15, 0, 11, 0, 22, 
    10, 0, 14, 0, 7, 0, 0, 7, 1, 1, 0, 0, 3, 16, 0, 
    
    -- channel=380
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 0, 
    0, 0, 0, 0, 0, 0, 3, 2, 2, 0, 0, 0, 0, 0, 0, 
    12, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 5, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 31, 20, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 24, 11, 1, 13, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 3, 2, 0, 16, 9, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=381
    37, 0, 4, 0, 5, 1, 6, 0, 25, 0, 0, 4, 0, 0, 17, 
    0, 12, 1, 0, 0, 0, 11, 0, 27, 11, 0, 0, 0, 8, 0, 
    24, 0, 0, 0, 0, 4, 12, 0, 2, 29, 0, 14, 0, 0, 0, 
    22, 0, 0, 0, 0, 3, 6, 7, 0, 0, 10, 27, 2, 0, 0, 
    0, 0, 0, 0, 0, 1, 3, 0, 20, 0, 0, 49, 0, 0, 0, 
    0, 12, 0, 0, 10, 0, 27, 0, 26, 0, 11, 42, 0, 0, 0, 
    0, 0, 5, 8, 0, 0, 17, 21, 0, 0, 43, 29, 0, 0, 0, 
    17, 0, 9, 0, 0, 7, 8, 0, 0, 3, 51, 30, 0, 0, 31, 
    7, 0, 0, 24, 0, 0, 31, 0, 0, 5, 53, 16, 0, 0, 72, 
    21, 0, 0, 98, 0, 0, 50, 0, 50, 19, 5, 7, 0, 0, 93, 
    15, 0, 0, 96, 0, 0, 0, 0, 37, 15, 0, 0, 0, 0, 65, 
    11, 0, 0, 24, 29, 0, 0, 33, 18, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 28, 17, 0, 25, 22, 12, 11, 0, 0, 0, 0, 
    6, 0, 19, 0, 18, 0, 0, 24, 0, 8, 6, 0, 9, 0, 8, 
    0, 0, 8, 0, 6, 0, 0, 2, 4, 2, 0, 0, 5, 15, 0, 
    
    -- channel=382
    46, 20, 3, 6, 15, 6, 10, 0, 21, 0, 1, 15, 6, 0, 20, 
    5, 16, 7, 7, 5, 14, 20, 12, 35, 5, 0, 0, 0, 13, 0, 
    14, 0, 7, 0, 3, 6, 22, 0, 16, 64, 11, 20, 0, 0, 6, 
    15, 0, 1, 0, 1, 4, 3, 6, 0, 6, 11, 28, 2, 0, 0, 
    0, 0, 6, 1, 2, 1, 11, 23, 16, 0, 0, 40, 0, 0, 0, 
    0, 13, 0, 2, 0, 0, 33, 0, 20, 0, 3, 17, 0, 0, 0, 
    0, 0, 2, 15, 0, 0, 3, 61, 21, 17, 33, 22, 0, 1, 0, 
    17, 0, 8, 0, 0, 15, 17, 0, 0, 12, 59, 22, 0, 8, 21, 
    16, 0, 8, 3, 0, 0, 17, 0, 0, 0, 0, 6, 0, 0, 73, 
    21, 0, 0, 79, 0, 0, 25, 2, 38, 0, 19, 25, 0, 0, 106, 
    19, 0, 0, 64, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 66, 
    0, 0, 0, 67, 30, 33, 19, 21, 7, 0, 1, 0, 0, 0, 0, 
    3, 0, 0, 0, 37, 18, 7, 40, 45, 35, 31, 16, 0, 0, 0, 
    3, 0, 9, 0, 5, 11, 0, 29, 15, 27, 32, 26, 38, 14, 2, 
    3, 4, 13, 4, 24, 9, 0, 0, 3, 4, 3, 0, 12, 21, 1, 
    
    -- channel=383
    35, 0, 43, 35, 42, 43, 48, 34, 40, 30, 28, 26, 22, 20, 35, 
    28, 36, 41, 35, 39, 40, 48, 44, 47, 32, 25, 35, 29, 35, 32, 
    34, 21, 34, 41, 37, 46, 48, 47, 42, 22, 7, 36, 38, 41, 31, 
    39, 21, 38, 35, 41, 55, 56, 52, 45, 47, 42, 46, 40, 30, 34, 
    35, 23, 32, 37, 40, 44, 37, 20, 43, 48, 43, 51, 28, 35, 34, 
    14, 30, 18, 33, 45, 1, 9, 36, 49, 23, 41, 55, 20, 32, 31, 
    0, 29, 26, 29, 15, 7, 43, 8, 0, 0, 38, 36, 13, 23, 33, 
    36, 1, 31, 29, 0, 19, 27, 9, 11, 10, 28, 34, 14, 0, 33, 
    45, 0, 19, 40, 9, 36, 51, 52, 51, 63, 83, 40, 2, 0, 41, 
    54, 5, 11, 61, 18, 23, 69, 4, 45, 47, 20, 14, 9, 0, 26, 
    50, 27, 27, 70, 4, 49, 62, 52, 83, 38, 31, 28, 13, 2, 32, 
    62, 31, 26, 12, 29, 12, 15, 40, 32, 20, 15, 13, 22, 33, 29, 
    46, 45, 32, 36, 36, 43, 35, 34, 17, 4, 1, 0, 4, 33, 16, 
    50, 45, 54, 40, 51, 27, 33, 55, 29, 23, 19, 3, 13, 13, 33, 
    43, 28, 51, 34, 31, 35, 50, 54, 48, 50, 38, 36, 40, 41, 27, 
    
    -- channel=384
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 0, 23, 54, 67, 40, 11, 0, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 17, 17, 28, 2, 0, 2, 13, 11, 4, 0, 0, 0, 
    0, 0, 0, 11, 9, 7, 12, 16, 9, 41, 48, 0, 0, 0, 10, 
    0, 63, 7, 5, 4, 0, 0, 9, 30, 66, 67, 82, 25, 31, 59, 
    0, 0, 1, 0, 0, 1, 5, 0, 5, 0, 0, 42, 21, 22, 0, 
    0, 1, 13, 0, 0, 0, 0, 10, 0, 0, 0, 3, 48, 23, 2, 
    0, 0, 37, 39, 77, 112, 119, 121, 65, 19, 23, 4, 41, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 17, 5, 0, 0, 0, 
    
    -- channel=385
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 26, 50, 46, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 26, 55, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 70, 5, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 26, 43, 48, 62, 0, 0, 0, 6, 
    0, 0, 6, 0, 0, 0, 0, 39, 33, 44, 57, 32, 0, 16, 23, 
    0, 27, 54, 0, 0, 0, 0, 34, 66, 8, 0, 19, 46, 35, 23, 
    0, 0, 33, 0, 0, 0, 0, 31, 67, 0, 0, 0, 32, 28, 0, 
    0, 0, 21, 0, 0, 0, 0, 25, 45, 0, 0, 0, 16, 4, 0, 
    0, 0, 12, 0, 1, 25, 32, 35, 44, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    
    -- channel=386
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 6, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 47, 65, 0, 0, 26, 0, 0, 
    0, 0, 0, 0, 0, 41, 61, 78, 43, 0, 0, 0, 0, 33, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 0, 0, 0, 
    0, 0, 0, 16, 29, 20, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 16, 10, 0, 0, 0, 77, 73, 0, 0, 0, 20, 
    0, 102, 2, 1, 4, 0, 0, 0, 45, 72, 65, 78, 20, 45, 90, 
    0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 36, 0, 36, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 40, 6, 
    0, 5, 58, 61, 102, 152, 161, 166, 100, 1, 16, 6, 50, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 30, 8, 0, 0, 0, 
    
    -- channel=387
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 13, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 8, 0, 0, 0, 0, 16, 
    0, 0, 0, 11, 0, 0, 0, 0, 5, 0, 0, 0, 0, 9, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 6, 0, 26, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 10, 0, 0, 12, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 15, 6, 5, 0, 
    
    -- channel=388
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 6, 0, 10, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 32, 11, 5, 8, 0, 
    2, 3, 2, 1, 2, 2, 5, 1, 2, 5, 5, 8, 0, 0, 0, 
    6, 4, 4, 3, 6, 10, 13, 12, 20, 31, 21, 18, 12, 4, 1, 
    4, 5, 4, 3, 10, 33, 65, 60, 55, 39, 58, 0, 22, 13, 5, 
    5, 6, 3, 9, 38, 29, 19, 0, 8, 46, 97, 2, 8, 24, 13, 
    6, 4, 21, 34, 25, 27, 17, 28, 64, 95, 72, 22, 0, 10, 44, 
    7, 14, 25, 34, 12, 15, 43, 97, 70, 65, 49, 0, 38, 60, 64, 
    11, 83, 11, 31, 0, 23, 62, 77, 66, 53, 55, 46, 75, 58, 39, 
    39, 54, 13, 17, 0, 32, 77, 67, 43, 0, 24, 75, 46, 37, 0, 
    24, 23, 48, 2, 19, 56, 76, 66, 0, 20, 14, 46, 52, 3, 1, 
    24, 33, 52, 6, 55, 61, 82, 60, 0, 38, 21, 17, 52, 0, 9, 
    19, 30, 31, 10, 30, 26, 25, 22, 0, 36, 16, 1, 13, 0, 9, 
    21, 17, 21, 22, 19, 20, 17, 13, 7, 31, 16, 0, 5, 5, 10, 
    
    -- channel=389
    114, 105, 99, 97, 90, 82, 78, 76, 60, 28, 47, 46, 0, 10, 43, 
    91, 86, 81, 76, 70, 65, 63, 61, 58, 56, 52, 17, 8, 27, 49, 
    50, 49, 59, 60, 59, 59, 59, 60, 60, 62, 2, 13, 29, 40, 47, 
    49, 57, 58, 59, 62, 63, 65, 64, 62, 49, 0, 0, 37, 42, 49, 
    55, 60, 59, 59, 61, 56, 45, 50, 56, 26, 7, 17, 37, 46, 46, 
    60, 60, 59, 57, 53, 44, 22, 12, 0, 0, 12, 4, 0, 33, 39, 
    60, 59, 54, 54, 18, 0, 0, 0, 0, 0, 0, 16, 0, 0, 24, 
    58, 58, 53, 25, 0, 2, 0, 31, 36, 0, 0, 0, 18, 2, 18, 
    56, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 21, 0, 
    64, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 
    32, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    9, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=390
    17, 6, 0, 0, 0, 0, 0, 3, 0, 0, 3, 4, 3, 0, 17, 
    0, 8, 5, 3, 5, 7, 6, 8, 8, 14, 12, 10, 20, 8, 21, 
    0, 0, 6, 12, 9, 16, 15, 15, 15, 13, 1, 27, 26, 17, 22, 
    11, 15, 17, 19, 17, 19, 27, 26, 21, 9, 8, 0, 12, 6, 14, 
    19, 18, 17, 19, 16, 18, 14, 20, 37, 59, 54, 13, 23, 17, 13, 
    19, 20, 19, 18, 11, 24, 34, 27, 0, 0, 91, 61, 0, 42, 14, 
    18, 20, 21, 14, 4, 0, 0, 0, 0, 0, 0, 157, 2, 0, 13, 
    17, 20, 17, 26, 18, 3, 27, 74, 75, 31, 18, 49, 65, 0, 49, 
    19, 16, 0, 0, 11, 0, 0, 10, 0, 7, 35, 56, 33, 41, 23, 
    12, 38, 80, 0, 16, 0, 0, 0, 6, 0, 0, 112, 47, 23, 4, 
    0, 0, 64, 14, 9, 13, 0, 7, 15, 0, 0, 0, 14, 0, 2, 
    0, 0, 31, 33, 10, 0, 0, 15, 85, 11, 16, 0, 5, 39, 12, 
    0, 0, 10, 46, 18, 53, 0, 7, 92, 2, 51, 0, 0, 33, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 5, 0, 11, 13, 0, 3, 0, 
    15, 17, 21, 39, 18, 22, 18, 16, 12, 0, 4, 17, 6, 5, 2, 
    
    -- channel=391
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 35, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 16, 0, 0, 20, 22, 21, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 10, 18, 31, 46, 4, 2, 0, 
    0, 0, 0, 4, 18, 6, 9, 7, 18, 18, 18, 18, 0, 5, 10, 
    0, 0, 34, 16, 20, 13, 0, 25, 29, 41, 10, 8, 19, 24, 25, 
    0, 9, 26, 21, 12, 5, 20, 28, 41, 23, 21, 4, 31, 35, 19, 
    0, 13, 23, 28, 9, 19, 15, 32, 46, 7, 20, 15, 17, 37, 0, 
    0, 11, 22, 26, 14, 26, 26, 31, 46, 9, 24, 17, 13, 27, 0, 
    0, 5, 28, 26, 26, 25, 23, 23, 20, 5, 17, 19, 14, 11, 4, 
    0, 0, 18, 23, 20, 19, 19, 16, 14, 17, 10, 11, 9, 9, 7, 
    
    -- channel=392
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 34, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 91, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 20, 5, 1, 17, 47, 29, 0, 0, 
    0, 0, 0, 0, 15, 0, 0, 0, 5, 11, 40, 29, 0, 0, 0, 
    0, 0, 46, 0, 13, 0, 0, 12, 18, 12, 0, 41, 15, 17, 16, 
    0, 0, 58, 18, 5, 0, 0, 19, 50, 22, 0, 0, 31, 25, 16, 
    0, 5, 30, 24, 0, 0, 0, 20, 71, 8, 10, 0, 18, 43, 0, 
    0, 1, 19, 30, 3, 28, 4, 22, 74, 0, 29, 0, 0, 30, 0, 
    0, 0, 4, 7, 0, 0, 0, 0, 25, 0, 16, 13, 0, 4, 0, 
    0, 1, 15, 25, 12, 13, 10, 9, 5, 0, 9, 8, 0, 0, 0, 
    
    -- channel=393
    99, 110, 109, 112, 114, 105, 97, 100, 83, 86, 74, 60, 47, 18, 57, 
    107, 104, 108, 106, 100, 92, 87, 86, 77, 73, 55, 58, 38, 10, 66, 
    84, 93, 88, 89, 81, 79, 79, 76, 73, 65, 37, 33, 29, 36, 69, 
    71, 74, 75, 77, 74, 77, 76, 74, 69, 60, 61, 0, 43, 66, 72, 
    70, 76, 77, 79, 73, 70, 58, 60, 45, 65, 37, 0, 56, 65, 64, 
    75, 78, 78, 78, 60, 36, 10, 15, 16, 23, 0, 77, 0, 56, 59, 
    77, 79, 83, 61, 38, 26, 40, 37, 22, 0, 0, 100, 11, 14, 40, 
    77, 80, 48, 44, 46, 1, 21, 0, 0, 0, 3, 94, 46, 0, 0, 
    79, 55, 39, 7, 32, 0, 0, 0, 1, 9, 44, 96, 12, 0, 0, 
    54, 0, 77, 0, 31, 0, 0, 0, 0, 30, 0, 28, 0, 9, 33, 
    20, 13, 54, 16, 14, 0, 0, 0, 58, 52, 0, 0, 24, 33, 66, 
    39, 0, 9, 39, 0, 0, 0, 0, 112, 0, 17, 0, 0, 71, 10, 
    32, 0, 0, 22, 0, 0, 0, 2, 98, 0, 30, 0, 0, 59, 4, 
    31, 6, 7, 8, 0, 5, 8, 15, 55, 0, 25, 25, 3, 13, 2, 
    30, 21, 1, 5, 0, 0, 0, 4, 8, 0, 13, 22, 2, 0, 0, 
    
    -- channel=394
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 51, 54, 0, 0, 17, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 38, 49, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 30, 44, 31, 20, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 4, 73, 34, 8, 31, 90, 0, 0, 0, 0, 
    5, 90, 0, 0, 0, 0, 42, 14, 0, 0, 24, 132, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 56, 4, 0, 0, 0, 71, 14, 0, 0, 
    0, 0, 7, 0, 0, 0, 19, 0, 0, 0, 0, 0, 63, 0, 0, 
    0, 0, 26, 4, 69, 86, 89, 83, 0, 19, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 
    
    -- channel=395
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 58, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 33, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 24, 53, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 17, 0, 27, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 89, 0, 0, 40, 10, 15, 
    0, 0, 0, 0, 0, 27, 10, 105, 105, 33, 0, 0, 20, 59, 73, 
    0, 0, 0, 0, 0, 27, 69, 0, 0, 0, 0, 0, 54, 75, 0, 
    0, 22, 0, 38, 21, 50, 74, 0, 0, 0, 0, 1, 2, 0, 0, 
    0, 0, 0, 24, 47, 91, 77, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 35, 5, 18, 73, 41, 44, 0, 0, 47, 36, 41, 0, 0, 53, 
    3, 23, 10, 44, 89, 53, 6, 0, 0, 56, 32, 42, 0, 0, 48, 
    18, 11, 0, 4, 0, 0, 0, 0, 0, 40, 1, 27, 22, 46, 57, 
    15, 26, 61, 62, 68, 69, 62, 59, 57, 37, 9, 43, 61, 62, 63, 
    
    -- channel=396
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 20, 12, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 15, 2, 0, 0, 14, 3, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 30, 0, 0, 8, 0, 0, 
    0, 0, 0, 7, 0, 8, 0, 32, 47, 48, 0, 0, 0, 2, 20, 
    0, 0, 2, 0, 0, 0, 22, 11, 0, 0, 0, 0, 0, 44, 0, 
    0, 41, 0, 1, 0, 9, 34, 0, 0, 0, 0, 10, 11, 0, 0, 
    17, 0, 0, 0, 2, 24, 40, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 0, 0, 15, 8, 26, 0, 0, 6, 0, 8, 0, 0, 6, 
    0, 0, 0, 4, 29, 17, 11, 0, 0, 3, 3, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 3, 
    0, 0, 7, 15, 9, 10, 8, 4, 3, 0, 0, 0, 5, 6, 9, 
    
    -- channel=397
    50, 47, 49, 49, 47, 41, 40, 38, 32, 28, 31, 22, 9, 12, 28, 
    39, 38, 39, 34, 30, 29, 30, 29, 28, 29, 18, 23, 17, 20, 25, 
    23, 25, 26, 25, 27, 26, 28, 29, 29, 26, 0, 0, 20, 26, 26, 
    25, 25, 24, 26, 26, 25, 20, 27, 28, 20, 10, 14, 29, 27, 27, 
    24, 24, 23, 23, 21, 17, 11, 11, 10, 15, 7, 13, 14, 24, 23, 
    23, 22, 23, 23, 15, 1, 0, 0, 0, 0, 0, 29, 3, 9, 22, 
    23, 22, 22, 16, 0, 0, 0, 12, 9, 0, 0, 1, 25, 7, 11, 
    21, 21, 4, 0, 0, 0, 0, 0, 6, 0, 0, 1, 0, 8, 0, 
    20, 9, 7, 0, 7, 5, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    12, 0, 1, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 12, 0, 0, 0, 0, 0, 6, 0, 0, 0, 7, 
    4, 0, 0, 15, 3, 0, 0, 0, 9, 3, 12, 0, 0, 12, 13, 
    4, 0, 0, 6, 0, 0, 0, 0, 10, 0, 5, 7, 0, 10, 13, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 21, 11, 14, 12, 
    5, 1, 6, 11, 6, 6, 10, 11, 15, 2, 0, 11, 15, 15, 12, 
    
    -- channel=398
    0, 0, 8, 13, 15, 13, 15, 9, 8, 27, 1, 0, 12, 29, 0, 
    6, 0, 13, 14, 14, 10, 9, 4, 1, 0, 0, 0, 0, 0, 0, 
    29, 30, 18, 7, 1, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 15, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 62, 70, 0, 0, 39, 2, 0, 
    0, 0, 0, 0, 0, 35, 52, 65, 40, 0, 0, 0, 0, 43, 19, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 
    0, 0, 0, 24, 22, 18, 0, 0, 1, 2, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 13, 10, 0, 0, 0, 68, 80, 0, 0, 0, 25, 
    0, 76, 23, 2, 6, 0, 0, 0, 45, 62, 48, 76, 23, 49, 72, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 20, 15, 25, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 38, 12, 
    0, 1, 47, 55, 82, 128, 140, 143, 95, 7, 11, 2, 34, 20, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 34, 12, 0, 0, 0, 
    
    -- channel=399
    9, 0, 1, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 29, 0, 
    0, 0, 0, 0, 2, 1, 1, 3, 2, 6, 15, 0, 0, 16, 0, 
    3, 5, 3, 0, 5, 4, 8, 4, 2, 3, 0, 29, 5, 0, 0, 
    5, 4, 3, 1, 8, 7, 6, 8, 24, 0, 0, 0, 0, 0, 0, 
    5, 2, 0, 1, 18, 44, 18, 0, 0, 0, 9, 0, 31, 0, 0, 
    4, 0, 0, 11, 25, 4, 0, 0, 7, 123, 66, 0, 0, 8, 0, 
    3, 0, 24, 0, 0, 15, 0, 37, 61, 60, 0, 0, 0, 21, 40, 
    0, 23, 0, 15, 0, 22, 84, 71, 0, 0, 0, 0, 37, 47, 17, 
    26, 90, 0, 19, 0, 36, 120, 26, 0, 0, 17, 0, 0, 0, 0, 
    73, 9, 0, 0, 0, 58, 118, 8, 0, 0, 33, 121, 0, 0, 0, 
    33, 10, 7, 0, 24, 56, 108, 0, 0, 10, 0, 90, 26, 0, 0, 
    26, 19, 24, 0, 68, 23, 61, 0, 0, 41, 0, 1, 64, 0, 13, 
    14, 21, 1, 0, 30, 15, 10, 0, 0, 54, 0, 0, 21, 0, 10, 
    4, 0, 4, 0, 0, 1, 0, 0, 0, 43, 0, 0, 2, 4, 15, 
    
    -- channel=400
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 33, 39, 7, 0, 57, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 32, 0, 19, 0, 0, 
    0, 0, 0, 0, 0, 6, 4, 40, 83, 113, 20, 0, 2, 13, 34, 
    0, 0, 0, 0, 0, 0, 20, 68, 11, 0, 0, 0, 5, 72, 38, 
    0, 43, 14, 15, 0, 17, 51, 10, 6, 0, 0, 44, 68, 21, 0, 
    0, 0, 0, 11, 0, 40, 67, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 18, 1, 27, 45, 45, 22, 0, 14, 8, 18, 1, 0, 0, 
    0, 13, 20, 12, 61, 61, 49, 3, 0, 29, 23, 17, 0, 0, 0, 
    0, 11, 2, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 10, 
    0, 3, 14, 36, 32, 32, 26, 19, 12, 8, 2, 0, 14, 15, 18, 
    
    -- channel=401
    28, 35, 36, 38, 42, 31, 25, 29, 15, 18, 16, 5, 13, 0, 0, 
    25, 30, 28, 22, 17, 12, 11, 13, 6, 6, 0, 17, 1, 0, 1, 
    16, 16, 6, 6, 2, 2, 3, 5, 5, 0, 9, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 5, 5, 6, 33, 0, 0, 5, 7, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 26, 8, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 21, 15, 3, 56, 0, 8, 0, 
    0, 0, 7, 0, 0, 0, 25, 7, 0, 0, 0, 101, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 14, 111, 20, 0, 0, 
    0, 0, 1, 0, 21, 0, 0, 0, 20, 17, 64, 49, 0, 0, 0, 
    0, 0, 58, 0, 3, 0, 0, 8, 8, 55, 0, 16, 0, 8, 40, 
    0, 5, 50, 3, 0, 0, 0, 7, 93, 13, 0, 0, 32, 41, 41, 
    0, 0, 12, 14, 0, 0, 0, 10, 116, 0, 0, 0, 0, 64, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 98, 0, 10, 0, 0, 30, 0, 
    0, 0, 7, 0, 0, 2, 7, 12, 38, 0, 4, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    
    -- channel=402
    43, 37, 30, 28, 28, 24, 19, 23, 6, 0, 0, 0, 0, 0, 3, 
    35, 40, 32, 28, 23, 21, 17, 17, 13, 11, 19, 0, 0, 0, 12, 
    7, 7, 18, 19, 15, 20, 19, 17, 17, 17, 0, 0, 2, 9, 12, 
    11, 16, 19, 21, 20, 23, 32, 32, 27, 13, 0, 0, 0, 0, 7, 
    18, 19, 19, 19, 21, 20, 15, 27, 60, 69, 30, 4, 18, 8, 7, 
    20, 22, 22, 17, 18, 33, 40, 14, 0, 0, 63, 42, 0, 28, 4, 
    21, 22, 18, 17, 0, 0, 0, 0, 0, 0, 0, 121, 0, 0, 0, 
    20, 22, 22, 23, 0, 0, 0, 67, 90, 44, 4, 0, 21, 0, 42, 
    20, 21, 0, 0, 0, 0, 0, 0, 0, 0, 9, 29, 16, 38, 4, 
    22, 50, 46, 0, 0, 0, 0, 0, 0, 0, 0, 96, 36, 2, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 3, 37, 0, 0, 42, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=403
    21, 17, 14, 13, 13, 8, 5, 3, 0, 0, 0, 0, 0, 0, 0, 
    15, 17, 11, 11, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 0, 1, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 5, 7, 2, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 1, 7, 2, 7, 14, 34, 0, 0, 0, 0, 0, 
    0, 2, 1, 0, 0, 7, 31, 33, 28, 8, 38, 17, 0, 0, 0, 
    1, 3, 3, 0, 11, 0, 0, 0, 0, 0, 45, 58, 0, 0, 0, 
    2, 4, 0, 12, 0, 0, 0, 0, 13, 61, 66, 47, 0, 0, 0, 
    4, 1, 0, 0, 0, 0, 0, 52, 66, 63, 74, 9, 0, 12, 28, 
    0, 39, 25, 0, 0, 0, 0, 46, 53, 50, 16, 56, 45, 37, 32, 
    3, 2, 10, 0, 0, 0, 0, 45, 56, 0, 0, 0, 42, 23, 0, 
    0, 0, 0, 0, 0, 0, 7, 53, 31, 0, 0, 0, 12, 3, 0, 
    0, 0, 0, 0, 0, 18, 36, 48, 31, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=404
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 26, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 9, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 36, 0, 0, 0, 5, 0, 23, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 63, 84, 0, 0, 19, 0, 
    0, 0, 4, 0, 0, 4, 0, 15, 66, 76, 4, 0, 0, 2, 44, 
    0, 0, 0, 0, 0, 7, 43, 82, 0, 0, 0, 0, 28, 33, 38, 
    0, 73, 0, 9, 0, 21, 69, 31, 0, 0, 0, 0, 15, 0, 0, 
    26, 15, 0, 0, 0, 37, 92, 7, 0, 0, 18, 76, 0, 0, 0, 
    1, 0, 21, 0, 11, 57, 70, 0, 0, 0, 0, 66, 5, 0, 0, 
    0, 6, 34, 0, 55, 28, 63, 0, 0, 30, 0, 0, 57, 0, 9, 
    1, 6, 6, 0, 18, 0, 0, 0, 0, 35, 0, 0, 21, 0, 7, 
    0, 0, 0, 0, 1, 3, 0, 0, 0, 45, 0, 0, 1, 2, 11, 
    
    -- channel=405
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 24, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 25, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 5, 3, 0, 28, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 66, 62, 16, 15, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 125, 0, 29, 5, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 161, 45, 0, 8, 
    0, 0, 0, 11, 19, 0, 22, 57, 51, 0, 0, 56, 51, 0, 17, 
    0, 0, 12, 0, 23, 0, 0, 0, 0, 0, 23, 103, 5, 7, 0, 
    0, 0, 114, 0, 40, 0, 0, 0, 0, 0, 0, 53, 13, 0, 0, 
    0, 0, 50, 24, 24, 0, 0, 0, 20, 24, 0, 0, 0, 0, 30, 
    0, 0, 0, 58, 5, 0, 0, 0, 115, 8, 25, 0, 0, 71, 13, 
    0, 0, 0, 66, 0, 28, 0, 0, 122, 0, 57, 4, 0, 60, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 19, 38, 0, 15, 4, 
    0, 18, 31, 51, 26, 27, 28, 25, 25, 0, 0, 29, 15, 14, 5, 
    
    -- channel=406
    16, 35, 35, 43, 47, 44, 39, 45, 35, 49, 33, 25, 37, 20, 30, 
    36, 31, 52, 52, 48, 45, 41, 39, 34, 32, 9, 19, 27, 0, 28, 
    50, 62, 49, 47, 37, 34, 35, 26, 26, 21, 0, 36, 1, 0, 31, 
    35, 33, 32, 33, 28, 29, 17, 11, 9, 12, 45, 5, 23, 35, 36, 
    31, 34, 35, 35, 29, 15, 11, 9, 0, 0, 0, 0, 22, 30, 28, 
    33, 35, 35, 34, 20, 0, 0, 0, 22, 48, 0, 65, 7, 24, 29, 
    32, 36, 40, 26, 0, 37, 48, 73, 34, 0, 0, 42, 17, 25, 33, 
    35, 38, 0, 0, 8, 0, 5, 0, 0, 0, 0, 90, 47, 0, 0, 
    39, 13, 8, 2, 47, 8, 0, 0, 0, 0, 5, 93, 0, 0, 0, 
    21, 0, 48, 0, 54, 0, 0, 0, 0, 43, 17, 0, 0, 0, 16, 
    0, 42, 44, 18, 33, 0, 0, 0, 40, 100, 19, 0, 21, 30, 119, 
    13, 0, 0, 47, 0, 0, 0, 0, 99, 0, 5, 0, 0, 83, 17, 
    9, 0, 0, 19, 0, 0, 0, 0, 77, 0, 0, 8, 0, 96, 13, 
    6, 0, 24, 54, 39, 75, 83, 92, 108, 0, 33, 37, 24, 34, 8, 
    7, 6, 0, 0, 0, 0, 0, 0, 5, 0, 37, 41, 5, 3, 0, 
    
    -- channel=407
    73, 83, 92, 97, 89, 90, 90, 80, 86, 73, 63, 51, 32, 57, 49, 
    98, 79, 88, 94, 91, 85, 84, 76, 74, 67, 63, 31, 17, 49, 54, 
    84, 85, 84, 83, 80, 74, 73, 68, 64, 68, 27, 14, 26, 40, 46, 
    73, 75, 74, 71, 73, 71, 67, 57, 55, 51, 8, 51, 41, 57, 60, 
    71, 76, 77, 73, 76, 59, 54, 56, 37, 0, 0, 26, 42, 61, 62, 
    74, 75, 72, 72, 77, 46, 0, 0, 4, 0, 0, 0, 58, 21, 60, 
    76, 73, 66, 74, 42, 51, 4, 22, 22, 78, 0, 0, 12, 31, 52, 
    76, 70, 65, 26, 8, 22, 0, 0, 0, 0, 0, 0, 0, 40, 0, 
    73, 73, 32, 20, 0, 35, 60, 0, 0, 0, 0, 0, 17, 0, 0, 
    88, 2, 0, 20, 0, 44, 75, 0, 0, 0, 0, 0, 0, 0, 0, 
    98, 40, 0, 0, 16, 26, 47, 0, 0, 0, 46, 53, 0, 0, 0, 
    73, 15, 0, 0, 22, 14, 19, 0, 0, 7, 0, 89, 0, 0, 18, 
    65, 14, 0, 0, 4, 0, 0, 0, 0, 20, 0, 26, 24, 0, 40, 
    46, 24, 4, 13, 48, 42, 39, 35, 0, 30, 0, 0, 44, 16, 34, 
    34, 18, 0, 0, 6, 2, 4, 8, 12, 50, 4, 12, 24, 25, 28, 
    
    -- channel=408
    39, 32, 33, 30, 27, 20, 18, 10, 10, 14, 0, 0, 0, 0, 0, 
    24, 21, 18, 16, 12, 7, 7, 2, 0, 0, 0, 0, 0, 0, 0, 
    11, 8, 4, 3, 0, 1, 3, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 0, 2, 2, 3, 7, 7, 8, 3, 3, 0, 0, 3, 4, 0, 
    0, 4, 6, 6, 7, 12, 8, 9, 2, 5, 0, 0, 0, 0, 0, 
    5, 5, 4, 3, 3, 3, 19, 24, 43, 30, 23, 0, 0, 0, 0, 
    5, 7, 7, 0, 12, 11, 16, 0, 0, 0, 73, 2, 0, 0, 0, 
    7, 7, 0, 0, 0, 0, 0, 0, 0, 49, 73, 44, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 70, 82, 79, 77, 0, 0, 0, 35, 
    0, 26, 0, 0, 0, 0, 3, 68, 64, 75, 56, 19, 27, 37, 41, 
    17, 47, 0, 0, 0, 0, 12, 59, 65, 0, 2, 46, 52, 39, 0, 
    5, 0, 6, 0, 0, 0, 31, 62, 13, 0, 0, 0, 29, 0, 0, 
    0, 0, 8, 0, 0, 4, 49, 56, 2, 0, 0, 0, 19, 0, 0, 
    0, 0, 7, 0, 8, 26, 32, 32, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=409
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 14, 7, 17, 9, 0, 
    0, 0, 0, 0, 0, 0, 6, 9, 10, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 6, 10, 43, 54, 42, 14, 4, 0, 0, 
    0, 0, 0, 0, 0, 40, 69, 49, 0, 0, 108, 0, 0, 15, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 3, 22, 62, 0, 0, 0, 
    0, 0, 21, 28, 4, 7, 18, 95, 139, 106, 14, 0, 13, 11, 70, 
    0, 11, 0, 0, 0, 0, 5, 66, 0, 0, 0, 0, 39, 80, 42, 
    7, 98, 26, 0, 0, 0, 11, 0, 0, 0, 0, 90, 71, 15, 0, 
    0, 0, 0, 0, 0, 49, 24, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 0, 27, 18, 18, 9, 0, 8, 3, 0, 0, 0, 0, 
    0, 2, 15, 17, 67, 76, 26, 0, 0, 24, 31, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    9, 12, 21, 39, 26, 29, 20, 12, 7, 0, 0, 0, 9, 10, 14, 
    
    -- channel=410
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 60, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 30, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 55, 119, 104, 54, 0, 0, 0, 30, 
    0, 0, 0, 0, 0, 0, 0, 67, 26, 27, 20, 0, 18, 51, 46, 
    0, 35, 2, 0, 0, 0, 0, 39, 32, 0, 0, 50, 67, 34, 0, 
    0, 0, 0, 0, 0, 7, 41, 38, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 19, 0, 0, 13, 31, 43, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 18, 1, 45, 77, 63, 33, 1, 5, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=411
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 21, 32, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 18, 1, 7, 24, 45, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 16, 12, 8, 47, 48, 10, 1, 0, 
    0, 0, 0, 4, 17, 6, 13, 10, 38, 46, 42, 41, 0, 0, 18, 
    0, 0, 33, 10, 17, 0, 5, 36, 45, 39, 35, 33, 20, 32, 24, 
    0, 11, 37, 13, 8, 3, 12, 43, 38, 42, 9, 13, 45, 34, 33, 
    0, 7, 20, 25, 3, 7, 20, 46, 59, 5, 10, 4, 26, 40, 0, 
    0, 4, 22, 33, 13, 31, 27, 46, 54, 9, 18, 4, 6, 32, 0, 
    0, 0, 15, 19, 14, 23, 24, 26, 32, 1, 22, 10, 4, 5, 0, 
    0, 0, 17, 12, 12, 11, 10, 8, 4, 0, 6, 9, 0, 0, 0, 
    
    -- channel=412
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 33, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 76, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 9, 1, 0, 66, 41, 0, 0, 
    0, 0, 0, 0, 8, 7, 22, 41, 30, 7, 0, 18, 38, 24, 6, 
    0, 0, 2, 0, 22, 15, 4, 0, 0, 0, 7, 49, 0, 15, 0, 
    0, 0, 55, 14, 39, 14, 0, 0, 0, 0, 0, 29, 8, 8, 8, 
    0, 0, 33, 29, 37, 23, 0, 0, 11, 37, 9, 0, 9, 9, 27, 
    0, 24, 3, 44, 28, 2, 0, 4, 48, 23, 29, 0, 0, 38, 26, 
    0, 9, 0, 53, 18, 24, 0, 7, 58, 9, 38, 29, 0, 47, 15, 
    0, 0, 3, 22, 0, 0, 0, 0, 15, 4, 18, 36, 12, 32, 23, 
    0, 21, 33, 41, 36, 35, 35, 33, 33, 4, 15, 39, 31, 31, 27, 
    
    -- channel=413
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 43, 53, 2, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 11, 14, 
    0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 22, 1, 0, 
    0, 0, 0, 0, 0, 7, 13, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 0, 0, 19, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 21, 30, 26, 0, 0, 1, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 3, 5, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=414
    83, 95, 95, 102, 97, 90, 85, 83, 74, 55, 60, 43, 17, 26, 41, 
    95, 83, 84, 83, 77, 71, 67, 66, 60, 57, 48, 30, 19, 14, 43, 
    66, 69, 66, 65, 63, 57, 57, 57, 54, 54, 3, 15, 22, 20, 41, 
    53, 54, 54, 55, 55, 53, 51, 50, 50, 45, 13, 18, 29, 46, 50, 
    47, 54, 54, 54, 53, 42, 37, 43, 39, 6, 0, 0, 28, 46, 46, 
    52, 54, 53, 54, 51, 27, 0, 0, 0, 0, 0, 0, 10, 18, 41, 
    55, 53, 50, 50, 9, 13, 0, 15, 9, 12, 0, 0, 1, 0, 26, 
    54, 53, 38, 10, 4, 0, 0, 0, 0, 0, 0, 0, 6, 12, 0, 
    51, 50, 15, 0, 0, 6, 4, 0, 0, 0, 0, 16, 0, 0, 0, 
    58, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 0, 0, 0, 14, 0, 0, 0, 0, 26, 0, 0, 0, 0, 10, 
    34, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 9, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 6, 
    11, 8, 0, 0, 0, 0, 0, 0, 1, 0, 0, 15, 5, 5, 4, 
    
    -- channel=415
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=416
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 15, 2, 
    0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 5, 0, 18, 61, 11, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 19, 36, 0, 0, 0, 96, 0, 0, 20, 0, 
    0, 0, 0, 0, 18, 0, 9, 0, 16, 0, 78, 36, 0, 20, 0, 
    0, 0, 0, 1, 9, 0, 2, 56, 77, 55, 2, 0, 0, 0, 75, 
    0, 0, 0, 0, 0, 0, 0, 87, 0, 0, 33, 0, 41, 13, 30, 
    0, 99, 0, 0, 0, 0, 0, 39, 0, 0, 0, 1, 22, 3, 0, 
    0, 0, 25, 7, 0, 27, 0, 14, 43, 0, 0, 8, 0, 0, 0, 
    0, 0, 98, 0, 2, 41, 0, 0, 13, 15, 3, 0, 32, 0, 0, 
    0, 6, 73, 0, 35, 53, 35, 0, 0, 10, 19, 0, 55, 0, 0, 
    3, 4, 9, 0, 0, 0, 0, 0, 0, 27, 0, 0, 10, 0, 0, 
    5, 0, 11, 30, 2, 13, 10, 7, 5, 0, 0, 0, 3, 1, 1, 
    
    -- channel=417
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 25, 40, 50, 46, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 84, 35, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 74, 89, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 77, 80, 79, 86, 0, 0, 0, 41, 
    0, 0, 0, 0, 0, 0, 0, 76, 60, 78, 65, 26, 27, 41, 40, 
    0, 48, 20, 0, 0, 0, 0, 65, 81, 0, 0, 37, 56, 44, 4, 
    0, 0, 34, 0, 0, 0, 5, 65, 64, 0, 0, 0, 31, 24, 0, 
    0, 0, 27, 0, 0, 10, 40, 53, 36, 0, 0, 0, 23, 0, 0, 
    0, 0, 16, 0, 0, 19, 23, 22, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=418
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 4, 8, 4, 
    0, 0, 0, 0, 0, 1, 0, 3, 3, 9, 0, 0, 16, 5, 0, 
    1, 1, 0, 2, 2, 3, 17, 18, 13, 1, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 22, 84, 80, 51, 4, 1, 0, 0, 
    1, 0, 0, 0, 13, 61, 25, 0, 0, 0, 49, 0, 0, 0, 0, 
    1, 0, 0, 10, 0, 0, 0, 0, 0, 66, 11, 41, 0, 0, 0, 
    0, 0, 28, 7, 0, 4, 11, 135, 168, 58, 0, 0, 0, 21, 74, 
    0, 27, 0, 0, 0, 0, 41, 1, 0, 0, 0, 22, 75, 76, 3, 
    28, 80, 0, 0, 0, 0, 9, 0, 0, 0, 0, 36, 18, 0, 0, 
    0, 0, 0, 0, 3, 60, 38, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 10, 0, 32, 3, 24, 0, 0, 17, 11, 0, 0, 0, 13, 
    0, 2, 5, 34, 78, 76, 25, 8, 0, 23, 22, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    2, 15, 50, 40, 22, 27, 20, 16, 13, 0, 0, 0, 7, 7, 11, 
    
    -- channel=419
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 39, 31, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 11, 34, 38, 19, 0, 16, 0, 3, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 45, 0, 0, 0, 
    0, 0, 0, 8, 20, 18, 0, 11, 37, 28, 29, 0, 0, 0, 0, 
    0, 0, 0, 10, 11, 16, 16, 29, 29, 78, 48, 0, 0, 11, 39, 
    0, 52, 19, 14, 3, 0, 8, 26, 65, 30, 54, 57, 40, 51, 36, 
    0, 7, 8, 4, 0, 15, 16, 25, 20, 0, 0, 35, 23, 26, 0, 
    0, 3, 12, 0, 0, 0, 13, 25, 12, 0, 0, 15, 44, 18, 0, 
    0, 7, 46, 46, 72, 89, 96, 95, 44, 16, 9, 8, 26, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 24, 4, 0, 0, 0, 
    
    -- channel=420
    40, 33, 48, 41, 38, 34, 40, 27, 32, 23, 24, 19, 3, 18, 18, 
    37, 30, 28, 28, 29, 25, 31, 25, 25, 22, 28, 8, 0, 28, 20, 
    25, 19, 22, 22, 26, 23, 25, 27, 25, 24, 28, 0, 7, 32, 18, 
    24, 23, 22, 20, 25, 23, 27, 26, 25, 18, 0, 12, 19, 20, 20, 
    23, 21, 20, 20, 24, 27, 28, 22, 22, 6, 0, 2, 17, 20, 22, 
    21, 20, 19, 21, 25, 30, 26, 0, 0, 0, 12, 0, 20, 9, 18, 
    21, 18, 18, 23, 29, 7, 0, 0, 10, 25, 48, 0, 0, 27, 11, 
    19, 16, 22, 5, 0, 6, 0, 12, 32, 31, 0, 0, 0, 7, 37, 
    17, 21, 0, 8, 0, 12, 10, 52, 0, 0, 0, 0, 23, 11, 16, 
    18, 59, 0, 6, 0, 16, 27, 11, 0, 0, 0, 0, 0, 0, 0, 
    28, 15, 0, 0, 0, 29, 32, 0, 0, 0, 9, 55, 0, 0, 0, 
    29, 0, 29, 0, 12, 39, 27, 0, 0, 8, 0, 28, 4, 0, 0, 
    21, 9, 31, 0, 31, 8, 25, 0, 0, 22, 0, 0, 51, 0, 19, 
    17, 15, 11, 0, 13, 0, 0, 0, 0, 31, 0, 0, 27, 0, 14, 
    14, 0, 1, 0, 3, 6, 4, 3, 6, 30, 0, 0, 12, 13, 17, 
    
    -- channel=421
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 13, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 7, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 28, 61, 35, 34, 0, 0, 0, 
    0, 0, 0, 0, 0, 24, 77, 45, 0, 0, 59, 41, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 27, 16, 32, 0, 0, 
    0, 0, 6, 32, 0, 2, 0, 71, 169, 180, 7, 0, 0, 11, 58, 
    0, 0, 0, 0, 0, 0, 0, 78, 0, 0, 0, 0, 28, 112, 50, 
    0, 96, 24, 0, 0, 0, 15, 0, 0, 0, 0, 48, 92, 11, 0, 
    7, 0, 0, 0, 0, 34, 66, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 31, 13, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 71, 83, 56, 0, 0, 14, 29, 4, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 8, 46, 27, 27, 22, 11, 5, 0, 0, 0, 5, 6, 9, 
    
    -- channel=422
    33, 35, 46, 47, 41, 37, 39, 28, 34, 35, 24, 7, 0, 19, 13, 
    31, 21, 30, 28, 24, 21, 26, 19, 19, 15, 8, 0, 0, 24, 11, 
    29, 27, 20, 17, 19, 16, 17, 17, 15, 11, 0, 0, 0, 17, 8, 
    20, 17, 15, 12, 16, 13, 6, 4, 7, 4, 0, 30, 22, 23, 15, 
    16, 15, 15, 12, 14, 5, 7, 0, 0, 0, 0, 0, 0, 9, 15, 
    15, 12, 11, 12, 7, 0, 0, 0, 1, 0, 0, 0, 21, 0, 11, 
    13, 12, 9, 5, 0, 27, 21, 29, 22, 10, 0, 0, 0, 18, 6, 
    13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 20, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 19, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 43, 0, 0, 0, 0, 13, 0, 0, 0, 61, 50, 0, 0, 1, 
    18, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 62, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 42, 0, 18, 
    8, 6, 24, 8, 61, 68, 65, 63, 0, 20, 0, 0, 46, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 4, 4, 4, 
    
    -- channel=423
    50, 48, 62, 58, 51, 52, 57, 41, 52, 41, 33, 29, 6, 41, 26, 
    60, 44, 49, 56, 56, 50, 53, 43, 43, 38, 41, 1, 0, 41, 31, 
    53, 51, 54, 50, 49, 45, 45, 40, 38, 40, 29, 0, 1, 35, 22, 
    46, 47, 45, 42, 46, 45, 46, 34, 32, 29, 0, 34, 30, 33, 34, 
    46, 48, 48, 45, 52, 45, 42, 39, 22, 0, 0, 10, 28, 34, 37, 
    48, 47, 45, 45, 53, 39, 12, 4, 24, 11, 0, 0, 47, 13, 33, 
    47, 46, 41, 49, 42, 34, 4, 0, 19, 74, 27, 0, 0, 33, 33, 
    48, 43, 47, 14, 0, 20, 0, 0, 0, 0, 0, 0, 0, 14, 13, 
    47, 48, 4, 20, 0, 23, 50, 32, 0, 0, 0, 0, 19, 2, 0, 
    56, 48, 0, 17, 0, 35, 86, 3, 0, 0, 33, 0, 0, 0, 0, 
    84, 46, 0, 0, 0, 24, 63, 0, 0, 0, 37, 106, 0, 0, 0, 
    54, 2, 0, 0, 10, 34, 59, 0, 0, 5, 0, 79, 11, 0, 3, 
    42, 15, 10, 0, 17, 0, 13, 0, 0, 25, 0, 5, 60, 0, 27, 
    29, 24, 16, 3, 51, 50, 49, 42, 0, 44, 0, 0, 31, 0, 16, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 44, 3, 0, 5, 6, 12, 
    
    -- channel=424
    0, 16, 24, 36, 43, 36, 30, 36, 25, 47, 26, 11, 31, 6, 4, 
    29, 22, 36, 35, 32, 27, 21, 23, 15, 11, 0, 16, 16, 0, 2, 
    37, 49, 29, 24, 15, 8, 7, 4, 1, 0, 0, 23, 0, 0, 8, 
    12, 3, 3, 4, 0, 0, 0, 0, 0, 0, 56, 0, 0, 12, 16, 
    0, 2, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 4, 12, 6, 
    0, 2, 4, 7, 0, 0, 0, 0, 8, 52, 0, 37, 0, 2, 7, 
    1, 3, 12, 0, 0, 35, 73, 87, 48, 0, 0, 47, 0, 17, 11, 
    3, 8, 0, 0, 14, 0, 4, 0, 0, 0, 0, 105, 24, 0, 0, 
    6, 0, 9, 9, 45, 7, 0, 0, 0, 0, 34, 99, 0, 0, 0, 
    0, 0, 40, 0, 40, 0, 0, 0, 0, 52, 29, 0, 0, 0, 23, 
    0, 56, 60, 7, 18, 0, 0, 0, 66, 112, 28, 0, 30, 43, 126, 
    1, 0, 0, 32, 0, 0, 0, 0, 120, 0, 0, 0, 0, 88, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 89, 0, 0, 0, 0, 88, 0, 
    0, 0, 23, 40, 37, 92, 105, 115, 123, 0, 36, 26, 24, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 27, 0, 0, 0, 
    
    -- channel=425
    48, 61, 73, 79, 76, 67, 65, 58, 47, 36, 30, 25, 0, 12, 13, 
    75, 62, 60, 59, 53, 46, 44, 41, 34, 28, 35, 5, 0, 0, 16, 
    44, 44, 42, 37, 34, 29, 30, 30, 28, 29, 1, 0, 0, 6, 15, 
    28, 25, 25, 25, 27, 25, 27, 27, 26, 20, 0, 0, 3, 19, 23, 
    20, 23, 23, 23, 26, 23, 23, 29, 30, 0, 0, 0, 15, 21, 22, 
    22, 23, 23, 23, 28, 22, 0, 0, 0, 0, 0, 0, 11, 2, 16, 
    24, 21, 20, 28, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 
    23, 22, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=426
    0, 6, 14, 20, 16, 19, 21, 13, 25, 43, 16, 13, 10, 34, 1, 
    18, 2, 12, 21, 21, 18, 17, 13, 13, 8, 1, 0, 0, 4, 0, 
    31, 35, 26, 19, 18, 9, 9, 5, 3, 6, 3, 0, 0, 0, 0, 
    16, 13, 10, 7, 6, 5, 0, 0, 0, 1, 6, 44, 6, 14, 9, 
    7, 11, 12, 10, 12, 1, 1, 0, 0, 0, 0, 0, 0, 4, 8, 
    10, 10, 8, 10, 17, 0, 0, 0, 37, 62, 0, 0, 64, 0, 7, 
    11, 9, 7, 15, 4, 59, 54, 73, 51, 80, 0, 0, 0, 39, 10, 
    13, 9, 9, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 21, 0, 
    12, 15, 8, 42, 4, 47, 69, 0, 0, 6, 0, 0, 0, 0, 0, 
    28, 0, 0, 24, 4, 46, 83, 4, 0, 43, 97, 0, 0, 0, 0, 
    62, 113, 0, 0, 13, 0, 38, 0, 0, 60, 86, 158, 5, 13, 44, 
    45, 19, 0, 0, 0, 10, 42, 0, 0, 0, 0, 107, 19, 0, 12, 
    33, 17, 0, 0, 0, 0, 0, 0, 0, 10, 0, 17, 72, 2, 23, 
    9, 33, 48, 60, 111, 149, 157, 157, 62, 33, 13, 0, 56, 25, 13, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 54, 22, 8, 2, 3, 6, 
    
    -- channel=427
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 16, 6, 1, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 22, 7, 3, 
    0, 0, 0, 0, 0, 0, 6, 16, 12, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 45, 91, 63, 16, 2, 0, 0, 
    0, 0, 0, 0, 0, 23, 34, 0, 0, 0, 58, 92, 0, 13, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 117, 36, 0, 0, 
    0, 0, 1, 29, 3, 0, 13, 98, 144, 100, 2, 0, 29, 7, 53, 
    0, 1, 9, 0, 0, 0, 0, 3, 0, 0, 1, 22, 29, 82, 13, 
    0, 58, 77, 0, 0, 0, 0, 0, 0, 0, 0, 75, 61, 8, 0, 
    0, 0, 4, 8, 0, 28, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 21, 18, 0, 0, 0, 26, 8, 13, 0, 0, 1, 0, 
    0, 0, 0, 45, 46, 74, 15, 0, 52, 0, 54, 5, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    2, 17, 28, 57, 28, 30, 27, 21, 16, 0, 0, 0, 9, 9, 7, 
    
    -- channel=428
    21, 2, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 28, 1, 
    0, 0, 0, 0, 1, 3, 3, 5, 7, 17, 24, 0, 10, 26, 0, 
    0, 5, 7, 4, 10, 9, 17, 17, 17, 20, 0, 4, 0, 0, 0, 
    9, 7, 6, 3, 12, 13, 13, 22, 62, 36, 0, 29, 1, 0, 2, 
    9, 7, 4, 2, 27, 63, 68, 21, 0, 0, 38, 0, 8, 0, 0, 
    9, 5, 0, 18, 35, 0, 0, 0, 0, 104, 75, 0, 7, 0, 0, 
    6, 2, 39, 31, 0, 19, 0, 82, 156, 162, 17, 0, 0, 32, 70, 
    2, 35, 10, 0, 0, 3, 77, 98, 3, 0, 0, 0, 56, 103, 53, 
    41, 127, 0, 13, 0, 21, 116, 19, 0, 0, 0, 0, 70, 8, 0, 
    68, 0, 0, 0, 0, 71, 142, 9, 0, 0, 0, 29, 0, 0, 0, 
    28, 4, 0, 0, 34, 64, 94, 6, 0, 10, 0, 70, 0, 0, 0, 
    22, 14, 14, 0, 104, 76, 92, 0, 0, 47, 0, 7, 10, 0, 3, 
    18, 9, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 9, 
    12, 6, 16, 14, 20, 21, 13, 5, 0, 25, 0, 0, 5, 7, 18, 
    
    -- channel=429
    41, 22, 9, 5, 3, 2, 0, 4, 0, 0, 1, 0, 0, 0, 15, 
    0, 11, 8, 0, 0, 0, 1, 3, 5, 10, 4, 4, 6, 20, 16, 
    0, 0, 0, 0, 2, 10, 9, 11, 14, 13, 0, 9, 24, 24, 18, 
    3, 9, 12, 13, 16, 15, 18, 20, 19, 13, 0, 0, 21, 3, 5, 
    15, 14, 12, 12, 11, 11, 11, 7, 18, 35, 27, 30, 12, 9, 8, 
    14, 14, 13, 10, 4, 0, 24, 42, 3, 0, 63, 76, 0, 34, 7, 
    13, 14, 11, 5, 0, 0, 0, 0, 0, 0, 0, 97, 24, 0, 3, 
    13, 12, 0, 23, 0, 2, 5, 46, 62, 84, 5, 0, 53, 0, 33, 
    12, 0, 0, 0, 0, 0, 0, 21, 3, 0, 8, 1, 0, 54, 18, 
    0, 26, 66, 0, 3, 0, 0, 0, 0, 0, 0, 81, 55, 12, 0, 
    0, 0, 7, 9, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 6, 0, 0, 3, 16, 4, 0, 0, 0, 2, 0, 
    0, 0, 0, 26, 16, 40, 1, 0, 34, 0, 35, 8, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 4, 0, 30, 15, 16, 14, 9, 4, 0, 0, 1, 4, 4, 2, 
    
    -- channel=430
    176, 172, 177, 177, 166, 151, 145, 133, 118, 92, 93, 63, 0, 17, 64, 
    157, 141, 144, 141, 128, 115, 114, 105, 97, 92, 68, 28, 2, 33, 73, 
    104, 108, 107, 106, 102, 97, 100, 96, 93, 89, 1, 0, 15, 55, 71, 
    90, 94, 94, 94, 99, 100, 95, 91, 85, 65, 0, 4, 67, 80, 81, 
    90, 98, 98, 96, 97, 79, 63, 66, 44, 1, 0, 0, 40, 71, 73, 
    97, 96, 95, 93, 82, 28, 0, 0, 0, 0, 0, 0, 0, 25, 63, 
    97, 96, 91, 78, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    96, 93, 48, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    94, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=431
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 17, 20, 0, 
    0, 0, 0, 0, 0, 0, 5, 12, 10, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 1, 49, 57, 36, 27, 0, 0, 0, 
    0, 0, 0, 0, 0, 42, 73, 25, 0, 0, 96, 0, 0, 4, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 21, 14, 41, 0, 0, 0, 
    0, 0, 15, 18, 0, 4, 0, 114, 182, 135, 2, 0, 0, 10, 85, 
    0, 4, 0, 0, 0, 0, 19, 65, 0, 0, 0, 0, 44, 109, 36, 
    5, 109, 0, 0, 0, 0, 22, 0, 0, 0, 0, 80, 67, 1, 0, 
    0, 0, 0, 0, 0, 52, 51, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 27, 14, 30, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 80, 86, 32, 0, 0, 21, 26, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 42, 24, 27, 18, 8, 3, 0, 0, 0, 3, 5, 10, 
    
    -- channel=432
    160, 154, 158, 154, 149, 139, 136, 127, 117, 100, 98, 83, 39, 42, 81, 
    148, 140, 138, 135, 128, 119, 117, 112, 106, 101, 89, 65, 33, 55, 90, 
    106, 109, 113, 114, 111, 108, 110, 108, 104, 101, 54, 22, 53, 79, 90, 
    100, 105, 106, 106, 109, 111, 112, 110, 106, 87, 32, 26, 76, 90, 94, 
    102, 108, 108, 107, 108, 102, 88, 94, 94, 78, 28, 31, 75, 90, 90, 
    107, 108, 107, 106, 98, 82, 49, 18, 0, 0, 11, 10, 22, 61, 84, 
    109, 108, 104, 96, 67, 24, 11, 3, 19, 7, 15, 10, 14, 28, 55, 
    106, 106, 86, 58, 29, 24, 20, 32, 50, 18, 0, 2, 6, 21, 40, 
    105, 92, 38, 12, 8, 5, 2, 10, 0, 0, 3, 19, 52, 27, 21, 
    100, 63, 5, 6, 5, 5, 0, 0, 0, 0, 0, 1, 12, 1, 0, 
    66, 3, 0, 6, 7, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    67, 0, 12, 7, 12, 5, 0, 0, 4, 11, 14, 0, 0, 3, 19, 
    53, 10, 8, 1, 13, 14, 5, 0, 0, 12, 14, 4, 4, 0, 24, 
    52, 21, 0, 0, 0, 0, 0, 0, 0, 4, 11, 12, 12, 9, 18, 
    48, 24, 13, 13, 7, 9, 12, 14, 17, 12, 1, 7, 17, 16, 17, 
    
    -- channel=433
    12, 0, 5, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 9, 0, 0, 37, 0, 
    0, 0, 0, 0, 1, 0, 1, 0, 0, 8, 0, 0, 0, 22, 0, 
    2, 4, 3, 0, 5, 4, 5, 0, 1, 2, 0, 29, 7, 0, 0, 
    7, 4, 3, 0, 10, 4, 8, 9, 14, 0, 0, 16, 0, 0, 0, 
    5, 2, 0, 0, 17, 31, 21, 5, 12, 0, 0, 0, 39, 0, 0, 
    3, 0, 0, 11, 16, 15, 0, 0, 0, 109, 72, 0, 0, 16, 2, 
    3, 0, 20, 0, 0, 17, 0, 14, 46, 62, 7, 0, 0, 24, 27, 
    0, 18, 0, 10, 0, 20, 87, 75, 8, 0, 0, 0, 32, 34, 36, 
    28, 58, 0, 20, 0, 36, 123, 30, 0, 0, 35, 0, 10, 0, 0, 
    63, 38, 0, 0, 0, 45, 120, 11, 0, 0, 26, 112, 0, 0, 0, 
    22, 0, 0, 0, 18, 55, 100, 1, 0, 1, 0, 103, 10, 0, 0, 
    17, 12, 21, 0, 59, 18, 63, 0, 0, 43, 0, 3, 58, 0, 16, 
    9, 15, 8, 0, 39, 22, 13, 3, 0, 45, 0, 0, 24, 0, 11, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 0, 1, 3, 14, 
    
    -- channel=434
    163, 166, 173, 175, 168, 155, 150, 141, 125, 101, 101, 88, 39, 52, 77, 
    163, 154, 148, 145, 135, 124, 121, 116, 109, 101, 90, 59, 33, 51, 84, 
    120, 117, 118, 113, 109, 105, 105, 105, 102, 101, 55, 36, 46, 72, 88, 
    98, 100, 101, 101, 105, 106, 106, 104, 102, 88, 27, 29, 75, 88, 91, 
    95, 102, 103, 102, 104, 100, 93, 92, 82, 52, 19, 35, 73, 89, 88, 
    101, 101, 102, 100, 94, 72, 56, 45, 36, 30, 18, 0, 37, 59, 81, 
    103, 102, 98, 93, 66, 30, 8, 4, 15, 10, 0, 10, 4, 31, 58, 
    102, 100, 84, 52, 23, 30, 16, 9, 11, 1, 0, 7, 19, 15, 28, 
    99, 86, 28, 18, 7, 8, 14, 12, 4, 5, 0, 19, 27, 14, 13, 
    94, 51, 1, 1, 9, 11, 5, 0, 0, 0, 23, 17, 1, 0, 4, 
    69, 12, 3, 0, 12, 5, 0, 0, 0, 0, 0, 12, 0, 0, 9, 
    56, 5, 0, 1, 10, 0, 0, 0, 0, 7, 8, 0, 1, 0, 25, 
    45, 7, 0, 0, 0, 0, 0, 0, 0, 8, 2, 2, 3, 8, 23, 
    43, 18, 0, 3, 0, 0, 0, 0, 14, 3, 6, 8, 2, 15, 16, 
    43, 14, 0, 0, 1, 1, 2, 4, 8, 6, 11, 14, 13, 13, 14, 
    
    -- channel=435
    69, 68, 73, 70, 65, 56, 56, 48, 42, 38, 29, 33, 12, 7, 16, 
    67, 59, 53, 47, 44, 38, 39, 35, 31, 28, 33, 17, 0, 10, 22, 
    42, 37, 36, 31, 31, 29, 30, 30, 31, 33, 40, 12, 8, 26, 24, 
    23, 26, 27, 27, 29, 32, 36, 39, 38, 38, 7, 2, 23, 28, 24, 
    24, 26, 27, 28, 32, 40, 42, 46, 53, 42, 12, 14, 25, 21, 22, 
    27, 27, 27, 28, 34, 49, 70, 66, 67, 66, 65, 0, 20, 15, 17, 
    28, 28, 27, 30, 40, 33, 27, 3, 7, 35, 99, 29, 0, 18, 9, 
    28, 29, 39, 32, 18, 24, 21, 20, 51, 80, 91, 56, 0, 3, 28, 
    27, 35, 19, 25, 11, 10, 35, 98, 97, 98, 79, 14, 27, 35, 65, 
    36, 70, 8, 10, 0, 3, 43, 86, 83, 74, 88, 61, 60, 61, 49, 
    40, 60, 21, 0, 0, 5, 46, 80, 54, 4, 9, 77, 62, 45, 8, 
    24, 8, 35, 0, 0, 25, 64, 82, 29, 4, 0, 21, 52, 13, 0, 
    12, 16, 37, 2, 26, 43, 72, 77, 22, 20, 6, 0, 39, 0, 0, 
    7, 17, 22, 5, 17, 30, 34, 33, 13, 15, 14, 0, 0, 0, 0, 
    14, 5, 2, 0, 0, 0, 0, 0, 0, 6, 4, 0, 0, 0, 0, 
    
    -- channel=436
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 9, 19, 6, 
    0, 0, 0, 0, 0, 0, 3, 4, 3, 4, 0, 0, 10, 10, 0, 
    3, 4, 3, 3, 4, 4, 8, 9, 4, 0, 0, 22, 19, 7, 3, 
    5, 3, 2, 1, 1, 0, 0, 3, 37, 29, 9, 0, 0, 0, 0, 
    5, 2, 1, 0, 3, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 2, 0, 0, 0, 0, 1, 16, 20, 48, 0, 0, 1, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 78, 78, 0, 0, 0, 0, 15, 26, 
    0, 7, 0, 0, 0, 2, 16, 0, 0, 0, 0, 35, 42, 18, 0, 
    10, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 29, 17, 0, 0, 15, 12, 0, 0, 0, 0, 
    0, 9, 0, 0, 12, 0, 6, 0, 0, 11, 6, 0, 0, 0, 12, 
    0, 0, 0, 15, 31, 32, 11, 2, 0, 5, 8, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 2, 3, 8, 1, 
    0, 6, 29, 12, 4, 8, 10, 12, 11, 0, 0, 0, 4, 4, 4, 
    
    -- channel=437
    0, 0, 0, 0, 4, 0, 0, 9, 0, 20, 8, 0, 20, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 46, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 0, 137, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 56, 93, 34, 0, 0, 219, 8, 0, 0, 
    0, 0, 0, 0, 19, 0, 21, 0, 0, 0, 0, 203, 103, 0, 0, 
    0, 0, 0, 0, 69, 0, 0, 0, 0, 0, 55, 219, 0, 0, 0, 
    0, 0, 144, 0, 87, 0, 0, 0, 0, 47, 0, 25, 0, 0, 32, 
    0, 0, 146, 23, 47, 0, 0, 0, 94, 170, 0, 0, 47, 59, 181, 
    0, 0, 0, 89, 0, 0, 0, 0, 255, 0, 21, 0, 0, 166, 22, 
    0, 0, 0, 66, 0, 0, 0, 0, 231, 0, 30, 0, 0, 177, 0, 
    0, 0, 2, 54, 0, 37, 52, 71, 182, 0, 57, 61, 0, 51, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 32, 66, 0, 0, 0, 
    
    -- channel=438
    136, 144, 151, 155, 149, 136, 131, 124, 108, 92, 84, 74, 38, 33, 60, 
    146, 136, 130, 128, 119, 108, 105, 101, 92, 85, 79, 53, 21, 31, 67, 
    106, 101, 100, 98, 94, 89, 89, 88, 86, 85, 57, 22, 31, 54, 72, 
    81, 83, 84, 84, 86, 88, 87, 89, 87, 79, 26, 9, 52, 72, 76, 
    77, 84, 84, 85, 87, 86, 79, 79, 74, 51, 13, 18, 58, 73, 73, 
    83, 84, 84, 84, 82, 69, 51, 38, 31, 23, 8, 0, 28, 44, 65, 
    86, 84, 83, 81, 61, 29, 7, 0, 7, 7, 5, 0, 0, 23, 41, 
    84, 84, 76, 49, 23, 17, 11, 5, 12, 0, 0, 0, 2, 10, 19, 
    83, 79, 32, 13, 1, 6, 9, 10, 1, 1, 0, 0, 24, 7, 10, 
    86, 53, 0, 0, 0, 4, 0, 0, 0, 0, 12, 6, 0, 0, 0, 
    68, 16, 0, 0, 1, 3, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    55, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    42, 4, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 3, 0, 12, 
    34, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 8, 
    34, 13, 0, 0, 0, 0, 0, 0, 0, 5, 0, 1, 5, 5, 7, 
    
    -- channel=439
    58, 59, 61, 63, 57, 51, 49, 44, 43, 45, 35, 18, 2, 16, 27, 
    48, 41, 49, 41, 34, 33, 35, 32, 31, 28, 23, 14, 9, 31, 26, 
    31, 35, 30, 27, 31, 28, 31, 31, 30, 29, 0, 0, 18, 27, 23, 
    30, 28, 29, 27, 30, 27, 21, 26, 25, 19, 5, 30, 34, 36, 26, 
    27, 27, 27, 25, 25, 10, 13, 16, 17, 0, 0, 16, 14, 22, 25, 
    27, 25, 26, 25, 21, 0, 0, 0, 0, 0, 0, 34, 6, 5, 23, 
    26, 25, 22, 19, 0, 14, 15, 38, 18, 8, 0, 0, 33, 2, 11, 
    25, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    23, 10, 15, 0, 2, 19, 0, 0, 0, 0, 0, 19, 0, 0, 0, 
    17, 0, 0, 1, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 8, 0, 0, 0, 0, 17, 47, 0, 0, 0, 19, 
    7, 0, 0, 7, 0, 0, 0, 0, 0, 0, 1, 29, 0, 3, 4, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 17, 
    9, 0, 0, 0, 13, 12, 8, 8, 0, 0, 1, 11, 31, 6, 12, 
    0, 1, 3, 0, 0, 0, 5, 8, 11, 16, 0, 5, 11, 11, 9, 
    
    -- channel=440
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 19, 42, 18, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 5, 3, 2, 28, 18, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 21, 0, 0, 8, 0, 
    0, 0, 0, 6, 8, 13, 20, 22, 29, 27, 10, 0, 0, 0, 11, 
    0, 0, 0, 14, 0, 12, 54, 28, 26, 22, 61, 11, 6, 14, 2, 
    0, 41, 17, 4, 1, 13, 27, 29, 5, 21, 12, 62, 33, 14, 16, 
    0, 8, 18, 0, 7, 21, 42, 26, 0, 8, 0, 33, 33, 1, 0, 
    0, 14, 27, 2, 13, 6, 19, 21, 0, 19, 0, 3, 34, 5, 0, 
    0, 9, 28, 31, 46, 50, 53, 51, 29, 27, 11, 0, 11, 2, 0, 
    0, 0, 0, 0, 6, 4, 1, 0, 0, 8, 18, 3, 0, 0, 0, 
    
    -- channel=441
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 11, 7, 0, 18, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 69, 35, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 53, 33, 22, 27, 0, 0, 23, 26, 
    0, 27, 0, 0, 0, 0, 13, 33, 24, 19, 0, 7, 38, 21, 11, 
    0, 2, 0, 0, 0, 0, 34, 26, 22, 0, 0, 4, 11, 3, 0, 
    0, 0, 5, 0, 0, 16, 27, 28, 0, 0, 0, 6, 5, 0, 0, 
    0, 0, 8, 0, 10, 26, 47, 22, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=442
    60, 40, 33, 26, 19, 14, 13, 9, 1, 0, 0, 0, 0, 0, 0, 
    24, 23, 12, 7, 2, 1, 2, 1, 0, 0, 9, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 3, 4, 7, 7, 10, 0, 0, 0, 13, 0, 
    0, 2, 4, 5, 8, 10, 17, 20, 17, 3, 0, 0, 0, 0, 0, 
    4, 5, 4, 3, 7, 7, 3, 9, 39, 28, 0, 0, 0, 0, 0, 
    6, 4, 4, 1, 6, 23, 22, 0, 0, 0, 8, 0, 0, 0, 0, 
    6, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 1, 9, 0, 0, 0, 0, 39, 94, 57, 0, 0, 0, 0, 26, 
    0, 4, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 10, 33, 0, 
    10, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 15, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=443
    0, 4, 2, 3, 12, 6, 2, 13, 0, 10, 11, 3, 2, 0, 11, 
    3, 6, 8, 6, 6, 6, 3, 8, 3, 9, 0, 1, 30, 0, 8, 
    0, 11, 6, 7, 3, 5, 5, 6, 5, 0, 0, 36, 9, 0, 14, 
    4, 1, 2, 5, 1, 3, 4, 5, 1, 0, 32, 0, 2, 4, 13, 
    0, 1, 0, 4, 0, 0, 0, 3, 0, 10, 31, 0, 5, 8, 3, 
    1, 2, 3, 4, 0, 0, 0, 0, 0, 25, 42, 44, 0, 25, 3, 
    0, 2, 8, 0, 0, 0, 7, 8, 8, 0, 0, 168, 0, 0, 5, 
    0, 5, 0, 0, 14, 0, 25, 24, 0, 0, 0, 86, 73, 0, 0, 
    2, 0, 0, 0, 28, 0, 0, 0, 0, 0, 30, 103, 0, 0, 0, 
    0, 0, 72, 0, 32, 0, 0, 0, 0, 0, 0, 68, 0, 0, 0, 
    0, 0, 97, 6, 19, 0, 0, 0, 22, 65, 0, 0, 14, 6, 71, 
    0, 0, 19, 42, 0, 0, 0, 0, 138, 0, 11, 0, 0, 73, 14, 
    0, 0, 0, 41, 0, 0, 0, 0, 126, 0, 28, 0, 0, 80, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 86, 0, 29, 21, 0, 22, 0, 
    0, 6, 7, 8, 0, 0, 0, 2, 5, 0, 11, 34, 0, 0, 0, 
    
    -- channel=444
    0, 0, 0, 0, 0, 1, 1, 0, 1, 6, 0, 0, 0, 18, 0, 
    12, 3, 4, 8, 7, 6, 5, 3, 2, 0, 11, 0, 0, 1, 0, 
    0, 12, 13, 7, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 3, 2, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 55, 52, 14, 4, 19, 7, 0, 
    0, 0, 0, 0, 7, 21, 0, 0, 0, 0, 0, 7, 4, 10, 4, 
    0, 0, 0, 5, 0, 0, 21, 41, 29, 30, 0, 0, 13, 8, 17, 
    0, 0, 0, 0, 11, 0, 0, 58, 44, 0, 0, 0, 0, 0, 25, 
    0, 8, 20, 4, 0, 12, 3, 0, 0, 0, 0, 43, 30, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 16, 1, 0, 0, 23, 29, 0, 0, 0, 0, 
    0, 1, 0, 0, 3, 0, 0, 0, 0, 8, 2, 0, 0, 0, 3, 
    0, 0, 0, 19, 17, 13, 0, 0, 0, 0, 3, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 5, 8, 7, 0, 
    0, 6, 34, 15, 5, 9, 8, 8, 8, 0, 0, 0, 0, 0, 0, 
    
    -- channel=445
    1, 12, 2, 7, 13, 9, 2, 15, 0, 6, 6, 2, 17, 0, 10, 
    3, 8, 18, 10, 7, 8, 3, 8, 4, 6, 0, 17, 18, 0, 10, 
    3, 14, 7, 9, 2, 4, 4, 3, 2, 0, 0, 29, 10, 0, 13, 
    1, 1, 3, 5, 1, 1, 0, 1, 0, 0, 34, 0, 0, 7, 9, 
    0, 2, 3, 4, 0, 0, 0, 0, 0, 15, 27, 0, 12, 6, 3, 
    1, 4, 5, 4, 0, 0, 0, 0, 0, 1, 0, 125, 0, 22, 6, 
    1, 4, 9, 0, 0, 0, 9, 28, 0, 0, 0, 151, 28, 0, 7, 
    2, 6, 0, 0, 13, 0, 15, 0, 0, 0, 0, 107, 60, 0, 0, 
    5, 0, 3, 0, 35, 0, 0, 0, 0, 0, 37, 124, 0, 0, 0, 
    0, 0, 110, 0, 48, 0, 0, 0, 0, 16, 0, 43, 0, 0, 18, 
    0, 0, 66, 18, 22, 0, 0, 0, 49, 70, 0, 0, 21, 21, 84, 
    0, 0, 0, 59, 0, 0, 0, 0, 146, 0, 11, 0, 0, 95, 6, 
    0, 0, 0, 52, 0, 0, 0, 0, 138, 0, 33, 0, 0, 90, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 59, 0, 22, 34, 0, 15, 0, 
    0, 6, 0, 10, 0, 0, 0, 3, 6, 0, 9, 32, 0, 0, 0, 
    
    -- channel=446
    17, 7, 0, 0, 0, 0, 0, 4, 0, 0, 3, 0, 0, 0, 13, 
    0, 6, 1, 0, 0, 0, 0, 1, 1, 7, 1, 11, 19, 0, 14, 
    0, 0, 0, 0, 0, 4, 3, 6, 7, 2, 0, 19, 25, 6, 14, 
    0, 0, 3, 6, 5, 6, 14, 17, 12, 1, 6, 0, 9, 1, 7, 
    4, 3, 2, 4, 0, 1, 0, 6, 29, 68, 57, 7, 17, 8, 3, 
    3, 4, 5, 4, 0, 0, 0, 0, 0, 0, 68, 106, 0, 42, 5, 
    3, 4, 8, 0, 0, 0, 0, 0, 0, 0, 0, 188, 15, 0, 4, 
    1, 6, 0, 14, 13, 0, 17, 73, 58, 9, 0, 43, 78, 0, 33, 
    3, 0, 0, 0, 7, 0, 0, 0, 0, 0, 34, 83, 7, 24, 0, 
    0, 0, 103, 0, 24, 0, 0, 0, 0, 0, 0, 100, 23, 5, 1, 
    0, 0, 70, 17, 14, 0, 0, 0, 22, 9, 0, 0, 0, 0, 8, 
    0, 0, 6, 40, 2, 0, 0, 0, 103, 7, 15, 0, 0, 50, 12, 
    0, 0, 0, 55, 0, 37, 0, 0, 117, 0, 57, 0, 0, 47, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 0, 6, 0, 
    1, 12, 17, 45, 15, 20, 19, 17, 14, 0, 0, 23, 5, 5, 0, 
    
    -- channel=447
    110, 128, 132, 141, 141, 132, 123, 122, 110, 100, 89, 76, 42, 40, 66, 
    133, 123, 131, 134, 125, 115, 107, 104, 95, 85, 67, 50, 33, 23, 73, 
    112, 122, 116, 109, 100, 95, 93, 86, 83, 80, 24, 32, 21, 36, 74, 
    91, 92, 91, 91, 90, 92, 82, 76, 71, 65, 42, 19, 61, 81, 84, 
    85, 94, 96, 95, 92, 76, 64, 66, 33, 8, 0, 3, 55, 75, 77, 
    93, 95, 94, 92, 81, 24, 0, 0, 13, 28, 0, 24, 22, 44, 72, 
    94, 96, 95, 83, 32, 38, 42, 58, 38, 0, 0, 14, 3, 25, 52, 
    96, 97, 57, 26, 17, 4, 1, 0, 0, 0, 0, 38, 32, 1, 0, 
    97, 72, 29, 13, 17, 6, 0, 0, 0, 0, 0, 80, 0, 0, 0, 
    84, 0, 15, 0, 31, 0, 0, 0, 0, 15, 15, 0, 0, 0, 5, 
    50, 25, 23, 1, 23, 0, 0, 0, 8, 70, 16, 0, 1, 11, 71, 
    56, 6, 0, 15, 0, 0, 0, 0, 39, 0, 2, 0, 0, 35, 21, 
    42, 0, 0, 2, 0, 0, 0, 0, 32, 0, 0, 2, 0, 56, 15, 
    35, 8, 3, 28, 16, 48, 56, 64, 72, 0, 19, 20, 11, 27, 4, 
    30, 12, 0, 0, 0, 0, 0, 0, 0, 0, 20, 25, 0, 0, 0, 
    
    -- channel=448
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 34, 12, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 14, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=449
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 6, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 21, 31, 65, 3, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 51, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    56, 39, 9, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=450
    0, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 7, 6, 0, 8, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 26, 5, 0, 0, 0, 0, 0, 0, 3, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 14, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 40, 53, 41, 50, 19, 20, 0, 2, 3, 0, 0, 0, 0, 
    90, 78, 1, 0, 0, 10, 0, 0, 9, 0, 0, 0, 0, 0, 0, 
    26, 19, 2, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 33, 16, 0, 0, 1, 4, 25, 35, 3, 5, 0, 0, 
    20, 30, 9, 0, 0, 0, 0, 0, 0, 0, 5, 18, 6, 0, 0, 
    
    -- channel=451
    0, 0, 0, 0, 2, 4, 4, 0, 0, 1, 2, 4, 4, 0, 0, 
    0, 0, 0, 5, 13, 22, 22, 16, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 11, 25, 34, 37, 33, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 34, 32, 33, 35, 29, 8, 5, 3, 0, 0, 0, 
    0, 0, 0, 32, 36, 17, 22, 42, 39, 39, 29, 17, 0, 0, 0, 
    0, 0, 0, 28, 17, 7, 30, 41, 31, 41, 42, 28, 1, 0, 0, 
    0, 0, 0, 9, 8, 20, 37, 33, 19, 34, 41, 37, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 26, 21, 34, 42, 43, 21, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 30, 25, 32, 39, 45, 28, 21, 3, 
    0, 0, 0, 0, 0, 0, 0, 34, 28, 30, 34, 48, 38, 19, 0, 
    0, 0, 13, 0, 24, 28, 30, 29, 28, 32, 30, 39, 33, 0, 0, 
    0, 0, 0, 0, 28, 38, 10, 22, 20, 26, 19, 28, 26, 0, 0, 
    0, 0, 0, 0, 0, 19, 11, 19, 24, 21, 15, 32, 26, 0, 0, 
    0, 0, 2, 5, 0, 0, 6, 16, 25, 25, 18, 33, 29, 7, 0, 
    3, 2, 0, 0, 0, 0, 5, 5, 1, 4, 10, 12, 10, 0, 0, 
    
    -- channel=452
    17, 14, 20, 17, 1, 0, 3, 8, 10, 9, 7, 5, 4, 8, 6, 
    16, 13, 17, 1, 0, 0, 0, 0, 1, 6, 6, 8, 12, 16, 13, 
    13, 13, 8, 0, 0, 0, 0, 0, 0, 12, 12, 12, 13, 14, 7, 
    11, 13, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 9, 4, 
    28, 35, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 6, 6, 
    36, 33, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 
    31, 29, 25, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 11, 9, 
    27, 31, 28, 16, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    32, 39, 43, 21, 19, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    65, 68, 50, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    62, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    28, 17, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    14, 14, 14, 15, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    11, 13, 3, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=453
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 3, 0, 0, 0, 6, 10, 8, 5, 
    0, 0, 0, 0, 0, 9, 7, 15, 18, 6, 3, 0, 0, 0, 0, 
    0, 0, 1, 0, 6, 10, 17, 19, 11, 0, 0, 0, 0, 0, 6, 
    4, 7, 0, 19, 4, 9, 16, 21, 21, 18, 9, 11, 6, 13, 16, 
    0, 0, 0, 9, 14, 1, 0, 13, 15, 21, 18, 8, 6, 9, 4, 
    0, 0, 0, 15, 0, 0, 5, 13, 7, 14, 17, 14, 6, 0, 0, 
    0, 0, 0, 8, 29, 8, 10, 14, 5, 9, 17, 14, 3, 0, 5, 
    0, 0, 2, 3, 4, 0, 6, 16, 0, 3, 15, 15, 7, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 0, 2, 10, 15, 6, 7, 14, 
    0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 4, 11, 11, 21, 19, 
    0, 0, 0, 0, 0, 0, 4, 1, 0, 1, 6, 11, 15, 10, 24, 
    0, 0, 0, 0, 6, 14, 0, 8, 6, 8, 0, 4, 27, 13, 14, 
    0, 0, 0, 0, 0, 6, 9, 0, 5, 0, 0, 1, 5, 19, 7, 
    0, 0, 2, 13, 15, 4, 9, 17, 17, 11, 1, 0, 10, 18, 14, 
    
    -- channel=454
    0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 0, 2, 3, 4, 12, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 6, 10, 17, 21, 22, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 12, 10, 3, 5, 3, 
    0, 2, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 10, 
    25, 32, 52, 6, 0, 0, 0, 0, 0, 0, 0, 0, 3, 15, 14, 
    7, 0, 46, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 
    0, 0, 16, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 7, 18, 74, 0, 1, 0, 0, 0, 0, 0, 0, 0, 9, 
    5, 14, 50, 26, 41, 39, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 28, 0, 47, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    8, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 12, 
    0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 22, 11, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=455
    13, 13, 8, 10, 3, 0, 9, 10, 10, 10, 11, 12, 10, 7, 8, 
    13, 13, 8, 9, 0, 0, 0, 0, 7, 3, 3, 3, 3, 2, 3, 
    13, 11, 13, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    10, 8, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 6, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 5, 7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 4, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 4, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 12, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 11, 5, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 6, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=456
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=457
    1, 3, 0, 5, 3, 2, 10, 8, 6, 5, 7, 8, 6, 2, 7, 
    1, 5, 0, 2, 4, 0, 5, 7, 9, 5, 6, 5, 3, 4, 10, 
    1, 3, 15, 0, 4, 0, 0, 0, 0, 3, 5, 12, 13, 17, 21, 
    0, 0, 23, 0, 0, 0, 0, 0, 3, 1, 3, 21, 16, 18, 17, 
    0, 0, 35, 15, 0, 0, 0, 4, 1, 0, 0, 5, 12, 23, 21, 
    0, 6, 50, 14, 0, 0, 2, 2, 0, 0, 2, 0, 6, 27, 30, 
    7, 11, 18, 45, 1, 0, 3, 0, 0, 3, 6, 0, 9, 18, 30, 
    1, 3, 16, 14, 41, 0, 13, 0, 0, 3, 3, 0, 0, 8, 18, 
    0, 0, 6, 21, 17, 39, 8, 11, 0, 0, 0, 0, 0, 6, 35, 
    0, 0, 19, 53, 9, 48, 2, 18, 0, 0, 0, 3, 0, 26, 31, 
    13, 33, 64, 28, 0, 18, 0, 0, 0, 0, 3, 4, 1, 18, 36, 
    31, 36, 23, 15, 23, 0, 0, 18, 0, 0, 0, 6, 17, 11, 43, 
    13, 7, 12, 9, 22, 9, 0, 13, 0, 0, 0, 3, 20, 22, 24, 
    8, 6, 16, 27, 22, 20, 10, 11, 3, 0, 0, 0, 14, 28, 23, 
    19, 27, 26, 28, 16, 20, 22, 31, 27, 20, 9, 14, 26, 27, 33, 
    
    -- channel=458
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 0, 22, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 1, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=459
    6, 7, 9, 0, 0, 0, 0, 8, 13, 15, 19, 24, 33, 41, 44, 
    7, 8, 5, 16, 0, 0, 0, 0, 9, 23, 29, 36, 38, 35, 28, 
    7, 8, 0, 17, 0, 0, 0, 0, 9, 14, 7, 1, 0, 0, 1, 
    13, 17, 27, 26, 9, 8, 5, 0, 0, 0, 0, 0, 1, 6, 12, 
    32, 22, 0, 14, 6, 7, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 13, 20, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 
    0, 0, 0, 0, 0, 0, 4, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 7, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=460
    5, 6, 6, 0, 9, 15, 8, 3, 5, 5, 3, 2, 3, 6, 7, 
    5, 5, 4, 9, 13, 19, 18, 16, 5, 6, 11, 14, 14, 11, 8, 
    5, 3, 0, 14, 19, 30, 28, 32, 24, 16, 11, 8, 5, 0, 0, 
    7, 8, 8, 19, 31, 37, 39, 33, 31, 12, 13, 5, 3, 1, 4, 
    22, 22, 3, 21, 33, 31, 35, 35, 36, 35, 28, 19, 6, 6, 8, 
    6, 2, 0, 19, 30, 35, 27, 34, 36, 37, 39, 30, 12, 3, 2, 
    0, 0, 0, 19, 15, 20, 25, 32, 31, 34, 33, 40, 20, 1, 0, 
    5, 7, 2, 0, 9, 33, 26, 34, 33, 30, 34, 40, 22, 10, 6, 
    9, 12, 16, 33, 12, 15, 14, 31, 33, 30, 37, 37, 30, 16, 0, 
    21, 10, 0, 0, 0, 0, 11, 30, 35, 32, 34, 36, 33, 8, 0, 
    0, 0, 0, 0, 15, 4, 25, 20, 32, 29, 26, 35, 29, 9, 0, 
    0, 0, 3, 0, 20, 31, 27, 21, 27, 33, 33, 29, 17, 6, 6, 
    0, 0, 0, 6, 3, 22, 13, 19, 31, 38, 28, 25, 21, 10, 0, 
    5, 7, 0, 0, 0, 4, 18, 12, 23, 23, 11, 27, 16, 5, 5, 
    0, 0, 0, 3, 7, 3, 12, 3, 8, 11, 14, 8, 5, 4, 1, 
    
    -- channel=461
    3, 4, 0, 3, 12, 15, 14, 7, 8, 10, 10, 12, 12, 12, 14, 
    3, 5, 5, 11, 23, 25, 23, 24, 14, 12, 16, 15, 13, 9, 10, 
    5, 5, 12, 13, 33, 39, 44, 42, 19, 7, 8, 9, 6, 5, 9, 
    8, 7, 15, 35, 40, 44, 46, 46, 37, 23, 16, 16, 7, 12, 15, 
    4, 0, 8, 27, 37, 25, 31, 46, 47, 45, 39, 25, 11, 15, 15, 
    0, 0, 5, 28, 30, 32, 36, 41, 41, 49, 49, 37, 20, 10, 10, 
    0, 0, 0, 19, 29, 18, 34, 41, 34, 40, 48, 40, 23, 7, 8, 
    0, 0, 0, 0, 16, 29, 36, 39, 29, 36, 47, 45, 32, 19, 16, 
    0, 0, 0, 10, 0, 14, 16, 39, 31, 35, 43, 48, 35, 23, 17, 
    0, 0, 0, 0, 5, 13, 20, 37, 35, 35, 40, 48, 38, 28, 19, 
    0, 0, 6, 22, 24, 28, 28, 30, 33, 33, 36, 46, 39, 20, 23, 
    0, 0, 0, 8, 33, 42, 24, 30, 38, 35, 30, 37, 37, 17, 19, 
    2, 0, 3, 7, 12, 20, 23, 26, 33, 26, 24, 34, 31, 25, 17, 
    8, 9, 12, 16, 17, 18, 25, 34, 34, 29, 25, 35, 36, 25, 20, 
    12, 16, 22, 24, 18, 17, 22, 26, 28, 29, 30, 31, 30, 25, 20, 
    
    -- channel=462
    0, 0, 0, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 3, 15, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 15, 11, 7, 0, 4, 0, 0, 0, 0, 0, 0, 1, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    5, 2, 0, 0, 11, 30, 9, 0, 0, 0, 0, 0, 5, 10, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 21, 
    0, 0, 15, 16, 20, 7, 1, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 5, 27, 47, 39, 42, 22, 25, 1, 5, 5, 0, 0, 0, 0, 
    80, 71, 19, 0, 0, 11, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    27, 18, 5, 0, 0, 0, 8, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 13, 29, 15, 0, 0, 3, 4, 21, 32, 8, 12, 5, 3, 
    20, 27, 12, 0, 0, 0, 0, 4, 0, 0, 4, 18, 11, 3, 2, 
    
    -- channel=463
    0, 0, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 3, 0, 0, 10, 0, 0, 0, 0, 0, 2, 1, 1, 0, 
    0, 0, 0, 7, 0, 2, 4, 9, 13, 1, 0, 0, 0, 0, 0, 
    0, 3, 0, 2, 5, 5, 5, 4, 7, 15, 4, 0, 0, 0, 0, 
    17, 12, 0, 0, 2, 26, 0, 0, 0, 3, 12, 0, 3, 0, 0, 
    4, 0, 0, 0, 3, 38, 0, 0, 0, 0, 0, 13, 10, 0, 0, 
    0, 0, 0, 0, 8, 21, 0, 0, 7, 0, 0, 16, 0, 4, 0, 
    5, 6, 0, 0, 0, 25, 0, 8, 9, 0, 0, 0, 2, 4, 0, 
    9, 20, 3, 0, 0, 0, 4, 0, 10, 0, 0, 0, 11, 0, 0, 
    13, 1, 0, 0, 0, 0, 15, 0, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 22, 0, 20, 13, 2, 0, 0, 19, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 9, 27, 0, 0, 0, 3, 6, 
    2, 2, 0, 0, 2, 2, 0, 0, 0, 12, 9, 0, 0, 0, 11, 
    0, 0, 0, 0, 15, 11, 0, 0, 0, 1, 10, 0, 0, 0, 0, 
    
    -- channel=464
    4, 3, 3, 0, 0, 0, 0, 0, 3, 2, 1, 2, 4, 8, 8, 
    4, 3, 1, 0, 0, 0, 0, 0, 0, 0, 3, 11, 19, 21, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 7, 1, 0, 0, 0, 
    1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 37, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 2, 14, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=465
    0, 0, 0, 0, 3, 8, 12, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 15, 10, 20, 14, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 12, 13, 18, 17, 0, 2, 1, 6, 2, 3, 3, 
    0, 0, 7, 0, 5, 13, 12, 17, 20, 12, 10, 19, 2, 1, 0, 
    0, 0, 54, 4, 7, 0, 19, 26, 27, 24, 20, 21, 3, 4, 4, 
    5, 14, 60, 0, 3, 0, 28, 29, 24, 24, 33, 13, 5, 10, 12, 
    11, 12, 17, 36, 6, 0, 33, 22, 20, 25, 33, 10, 21, 9, 14, 
    4, 4, 26, 7, 35, 0, 26, 14, 21, 34, 30, 25, 22, 3, 2, 
    2, 0, 8, 26, 38, 54, 16, 26, 20, 29, 29, 32, 13, 13, 19, 
    3, 20, 40, 85, 23, 72, 5, 36, 21, 24, 30, 37, 18, 21, 0, 
    31, 58, 60, 42, 26, 36, 24, 13, 22, 26, 29, 32, 18, 9, 5, 
    53, 37, 26, 23, 32, 7, 4, 18, 5, 8, 17, 29, 20, 0, 20, 
    15, 7, 3, 4, 20, 13, 5, 22, 4, 0, 29, 28, 28, 6, 4, 
    0, 3, 16, 17, 0, 6, 0, 19, 12, 10, 17, 24, 28, 8, 0, 
    12, 8, 3, 1, 0, 3, 12, 10, 3, 6, 1, 11, 15, 0, 2, 
    
    -- channel=466
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 20, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 13, 53, 34, 24, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    47, 30, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=467
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 23, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 16, 12, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 16, 23, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 29, 44, 39, 25, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    63, 77, 67, 52, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    78, 77, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 15, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=468
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 11, 0, 0, 0, 0, 0, 0, 3, 3, 0, 
    0, 0, 0, 0, 0, 5, 8, 11, 12, 6, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 3, 12, 12, 14, 9, 13, 0, 0, 0, 0, 0, 
    15, 17, 0, 0, 10, 28, 9, 0, 8, 6, 14, 5, 6, 0, 0, 
    5, 0, 0, 0, 0, 41, 0, 0, 11, 2, 4, 20, 17, 0, 0, 
    0, 0, 0, 0, 15, 13, 0, 6, 17, 0, 0, 22, 8, 5, 0, 
    0, 2, 0, 0, 0, 25, 0, 11, 17, 0, 0, 8, 14, 7, 0, 
    7, 11, 2, 0, 0, 0, 2, 0, 16, 0, 0, 0, 22, 4, 0, 
    21, 11, 0, 0, 7, 0, 15, 0, 13, 6, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 7, 6, 0, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 5, 29, 0, 14, 16, 10, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 10, 28, 5, 0, 0, 4, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 4, 0, 0, 0, 5, 
    0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    
    -- channel=469
    0, 3, 0, 0, 0, 1, 9, 0, 8, 6, 5, 10, 11, 8, 20, 
    0, 7, 0, 0, 1, 0, 1, 9, 4, 9, 18, 20, 19, 16, 17, 
    0, 1, 3, 0, 6, 3, 0, 0, 0, 6, 8, 6, 1, 2, 5, 
    1, 5, 46, 10, 6, 13, 11, 0, 0, 0, 0, 8, 0, 10, 10, 
    13, 10, 46, 33, 1, 0, 11, 24, 5, 2, 0, 0, 0, 9, 8, 
    0, 0, 45, 35, 20, 0, 7, 16, 7, 12, 9, 0, 0, 0, 3, 
    0, 0, 1, 86, 0, 0, 6, 3, 0, 19, 15, 0, 0, 0, 3, 
    0, 0, 0, 0, 81, 8, 24, 0, 0, 19, 18, 7, 0, 0, 9, 
    0, 0, 23, 42, 14, 44, 0, 18, 0, 12, 18, 19, 0, 0, 1, 
    0, 0, 0, 24, 0, 25, 0, 23, 0, 2, 10, 22, 1, 22, 7, 
    0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 4, 19, 9, 12, 21, 
    0, 0, 4, 9, 38, 0, 0, 35, 0, 0, 2, 22, 16, 0, 32, 
    0, 0, 0, 0, 11, 16, 0, 17, 0, 0, 9, 11, 27, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 6, 13, 1, 0, 
    0, 0, 0, 6, 0, 0, 4, 8, 3, 2, 0, 0, 5, 0, 0, 
    
    -- channel=470
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 7, 4, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 0, 21, 0, 6, 0, 0, 0, 0, 0, 0, 0, 10, 12, 
    0, 0, 78, 10, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    53, 48, 10, 0, 6, 0, 0, 5, 0, 0, 0, 0, 0, 0, 11, 
    7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 30, 18, 0, 0, 0, 0, 0, 0, 0, 0, 9, 1, 
    17, 31, 15, 10, 0, 0, 0, 14, 6, 0, 0, 4, 12, 9, 12, 
    
    -- channel=471
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 7, 13, 6, 
    0, 0, 0, 12, 0, 7, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 4, 8, 3, 1, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 15, 5, 0, 2, 7, 11, 7, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 5, 2, 0, 0, 0, 3, 6, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 8, 12, 4, 1, 
    0, 0, 0, 0, 8, 20, 0, 0, 0, 0, 0, 13, 0, 13, 4, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 15, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 1, 2, 25, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 9, 0, 0, 12, 2, 0, 0, 4, 28, 0, 
    0, 0, 0, 0, 0, 0, 14, 0, 2, 4, 0, 0, 0, 26, 15, 
    0, 0, 0, 11, 25, 2, 15, 0, 9, 16, 2, 0, 0, 26, 34, 
    5, 21, 22, 21, 41, 19, 6, 18, 28, 19, 28, 20, 14, 33, 34, 
    
    -- channel=472
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 35, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 3, 
    29, 28, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 25, 31, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 35, 36, 26, 24, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 79, 85, 51, 26, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    91, 90, 30, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    70, 44, 14, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 8, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=473
    5, 2, 2, 0, 0, 9, 1, 2, 5, 3, 0, 0, 2, 7, 13, 
    5, 5, 1, 0, 3, 0, 9, 9, 1, 9, 17, 27, 34, 33, 26, 
    0, 2, 0, 0, 0, 8, 1, 7, 27, 35, 24, 18, 6, 0, 0, 
    5, 11, 25, 0, 8, 19, 20, 14, 3, 0, 4, 0, 4, 4, 9, 
    51, 61, 44, 6, 10, 29, 39, 18, 16, 9, 0, 12, 14, 14, 18, 
    19, 3, 15, 0, 32, 26, 3, 12, 24, 17, 15, 8, 1, 6, 3, 
    0, 0, 8, 29, 0, 0, 7, 15, 24, 19, 17, 10, 4, 0, 0, 
    6, 13, 4, 17, 64, 29, 23, 17, 25, 20, 17, 13, 11, 2, 8, 
    20, 32, 65, 32, 48, 30, 25, 15, 13, 15, 22, 21, 17, 1, 0, 
    68, 47, 0, 4, 0, 9, 0, 11, 17, 15, 21, 19, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 5, 13, 10, 22, 6, 
    0, 0, 0, 13, 0, 0, 26, 5, 0, 7, 24, 23, 1, 1, 13, 
    0, 0, 0, 0, 21, 28, 0, 13, 17, 25, 30, 9, 19, 0, 6, 
    0, 1, 0, 0, 0, 6, 9, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    
    -- channel=474
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 34, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 25, 56, 26, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    68, 54, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=475
    15, 14, 10, 12, 7, 4, 8, 9, 9, 7, 8, 7, 5, 3, 4, 
    15, 14, 8, 12, 1, 0, 0, 1, 5, 6, 3, 1, 1, 0, 0, 
    13, 12, 8, 0, 0, 0, 0, 0, 0, 1, 2, 0, 0, 1, 0, 
    10, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    11, 12, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 18, 27, 9, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 19, 22, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 16, 14, 14, 12, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    16, 18, 22, 19, 7, 2, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    20, 22, 30, 27, 15, 11, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    36, 34, 42, 17, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 36, 18, 12, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 15, 13, 5, 3, 0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 
    7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=476
    26, 27, 19, 20, 29, 32, 32, 28, 29, 27, 28, 30, 30, 28, 32, 
    26, 28, 20, 32, 35, 32, 40, 41, 32, 28, 31, 31, 30, 26, 26, 
    26, 25, 24, 30, 44, 48, 47, 44, 32, 30, 25, 22, 19, 16, 18, 
    27, 27, 39, 41, 53, 52, 49, 40, 40, 24, 29, 28, 16, 20, 21, 
    27, 24, 31, 56, 48, 34, 46, 55, 47, 47, 41, 33, 16, 17, 16, 
    11, 10, 26, 51, 46, 36, 50, 56, 45, 49, 50, 38, 14, 6, 8, 
    8, 9, 14, 60, 22, 22, 47, 49, 42, 51, 50, 44, 28, 4, 11, 
    15, 13, 13, 14, 53, 34, 42, 40, 41, 53, 56, 52, 35, 24, 19, 
    12, 9, 17, 43, 19, 34, 18, 50, 43, 52, 57, 57, 42, 26, 11, 
    5, 0, 0, 23, 12, 19, 22, 54, 47, 50, 52, 61, 47, 29, 8, 
    0, 0, 46, 19, 28, 36, 39, 31, 42, 44, 46, 55, 41, 17, 15, 
    0, 3, 21, 25, 55, 46, 28, 52, 36, 42, 42, 47, 33, 3, 22, 
    15, 16, 17, 18, 26, 38, 24, 41, 47, 41, 43, 47, 38, 12, 4, 
    20, 18, 17, 14, 12, 14, 31, 26, 36, 30, 28, 48, 32, 12, 4, 
    15, 12, 12, 14, 5, 6, 21, 16, 16, 20, 21, 18, 19, 7, 5, 
    
    -- channel=477
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=478
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 1, 2, 3, 
    0, 0, 0, 9, 3, 14, 16, 15, 5, 0, 3, 0, 0, 0, 0, 
    0, 0, 0, 11, 19, 27, 32, 34, 16, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 12, 30, 28, 31, 30, 36, 16, 7, 9, 1, 0, 6, 
    0, 0, 0, 26, 21, 12, 11, 29, 35, 38, 31, 19, 7, 6, 7, 
    0, 0, 0, 17, 16, 9, 17, 27, 26, 34, 36, 31, 16, 10, 6, 
    0, 0, 0, 5, 0, 14, 20, 27, 17, 23, 31, 33, 20, 8, 6, 
    0, 0, 0, 0, 0, 5, 11, 23, 14, 15, 30, 34, 19, 17, 6, 
    0, 0, 0, 0, 0, 0, 0, 25, 18, 16, 24, 29, 23, 14, 17, 
    0, 0, 0, 0, 0, 0, 7, 30, 18, 16, 18, 28, 28, 23, 20, 
    0, 0, 15, 3, 11, 24, 25, 26, 19, 18, 24, 31, 26, 14, 18, 
    0, 0, 0, 0, 14, 30, 9, 19, 22, 24, 12, 18, 27, 17, 21, 
    0, 0, 0, 0, 0, 2, 12, 17, 17, 16, 0, 14, 27, 25, 16, 
    0, 0, 0, 15, 25, 8, 21, 13, 26, 20, 14, 22, 21, 31, 24, 
    2, 18, 24, 22, 24, 13, 17, 27, 29, 23, 24, 22, 26, 28, 27, 
    
    -- channel=479
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=480
    0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 
    0, 0, 8, 0, 1, 0, 0, 0, 0, 1, 3, 8, 7, 8, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 6, 0, 0, 0, 
    0, 4, 19, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 20, 55, 0, 0, 17, 11, 0, 0, 0, 0, 2, 2, 0, 0, 
    0, 0, 38, 0, 14, 14, 0, 0, 8, 0, 1, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 12, 0, 1, 0, 0, 2, 0, 
    0, 0, 4, 0, 13, 0, 6, 0, 8, 0, 0, 0, 18, 0, 0, 
    0, 7, 33, 0, 47, 30, 31, 0, 0, 0, 0, 0, 1, 0, 0, 
    21, 10, 0, 15, 0, 46, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 
    0, 0, 0, 0, 0, 0, 24, 0, 4, 0, 3, 6, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 18, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    
    -- channel=481
    0, 0, 0, 3, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 1, 0, 0, 0, 
    0, 14, 40, 0, 0, 1, 7, 0, 0, 0, 4, 3, 0, 0, 0, 
    34, 40, 52, 0, 0, 3, 11, 4, 0, 0, 0, 0, 0, 0, 0, 
    32, 31, 35, 0, 0, 4, 15, 5, 7, 1, 3, 0, 0, 0, 0, 
    26, 29, 39, 27, 7, 0, 7, 3, 14, 14, 3, 0, 0, 0, 0, 
    32, 34, 46, 20, 51, 26, 24, 6, 10, 15, 5, 1, 0, 0, 0, 
    59, 78, 88, 88, 52, 61, 19, 9, 10, 14, 14, 6, 0, 0, 0, 
    91, 98, 31, 41, 18, 26, 2, 0, 12, 11, 11, 1, 0, 0, 0, 
    78, 51, 18, 24, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 0, 
    17, 13, 8, 8, 12, 0, 3, 0, 0, 0, 22, 14, 0, 0, 0, 
    0, 3, 9, 0, 0, 0, 0, 0, 0, 0, 17, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=482
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 8, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 10, 22, 29, 26, 19, 12, 
    0, 0, 0, 0, 0, 0, 0, 5, 17, 12, 5, 2, 0, 0, 0, 
    1, 10, 35, 4, 4, 19, 20, 3, 0, 0, 0, 0, 6, 2, 5, 
    50, 42, 0, 0, 0, 7, 13, 2, 3, 0, 0, 0, 8, 13, 10, 
    0, 0, 0, 2, 24, 21, 0, 1, 12, 5, 1, 4, 1, 1, 0, 
    0, 0, 7, 27, 0, 0, 0, 4, 12, 7, 1, 0, 0, 0, 0, 
    6, 12, 0, 0, 32, 44, 12, 5, 3, 0, 2, 1, 3, 6, 14, 
    12, 39, 74, 22, 13, 4, 14, 0, 1, 3, 9, 5, 5, 0, 0, 
    47, 4, 0, 0, 0, 0, 0, 0, 5, 4, 5, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 7, 18, 2, 
    0, 0, 0, 0, 0, 1, 21, 0, 7, 13, 13, 8, 1, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 6, 1, 11, 5, 0, 4, 0, 4, 
    4, 0, 0, 0, 0, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 
    
    -- channel=483
    18, 19, 15, 20, 25, 20, 20, 16, 13, 15, 14, 12, 9, 2, 0, 
    18, 16, 18, 17, 28, 38, 29, 22, 14, 4, 0, 0, 0, 0, 0, 
    21, 18, 24, 25, 30, 31, 36, 29, 11, 2, 3, 3, 5, 7, 6, 
    16, 10, 0, 16, 32, 25, 22, 25, 29, 31, 24, 15, 1, 0, 0, 
    0, 0, 5, 13, 33, 25, 20, 26, 28, 32, 37, 23, 0, 0, 0, 
    12, 20, 9, 11, 10, 22, 39, 35, 25, 25, 31, 31, 10, 0, 0, 
    25, 22, 9, 0, 26, 41, 40, 32, 27, 26, 28, 35, 22, 7, 7, 
    16, 9, 19, 2, 0, 0, 12, 25, 34, 33, 31, 35, 28, 9, 0, 
    8, 0, 0, 2, 3, 6, 5, 22, 40, 37, 32, 34, 31, 22, 7, 
    0, 5, 45, 35, 39, 20, 23, 27, 40, 39, 34, 37, 36, 8, 0, 
    24, 36, 43, 49, 59, 52, 46, 33, 38, 41, 35, 32, 24, 0, 0, 
    76, 56, 26, 17, 24, 36, 18, 16, 34, 33, 25, 22, 12, 0, 0, 
    36, 30, 17, 13, 6, 10, 26, 19, 29, 30, 31, 35, 9, 0, 0, 
    12, 14, 24, 22, 6, 0, 3, 18, 25, 42, 47, 37, 24, 0, 0, 
    20, 14, 0, 0, 0, 0, 4, 0, 0, 0, 12, 17, 3, 0, 0, 
    
    -- channel=484
    1, 0, 6, 0, 8, 12, 0, 2, 1, 6, 2, 1, 4, 9, 5, 
    1, 0, 10, 0, 16, 24, 15, 11, 1, 8, 7, 9, 9, 9, 4, 
    2, 4, 1, 10, 18, 28, 34, 32, 18, 10, 6, 8, 2, 1, 1, 
    6, 8, 0, 13, 29, 34, 34, 38, 29, 24, 13, 2, 4, 1, 6, 
    11, 9, 0, 0, 28, 44, 29, 17, 36, 32, 32, 21, 12, 6, 9, 
    1, 0, 0, 0, 25, 47, 17, 18, 35, 32, 35, 37, 20, 10, 4, 
    0, 0, 0, 0, 26, 33, 19, 30, 34, 20, 31, 35, 18, 16, 0, 
    0, 0, 0, 0, 0, 22, 19, 33, 34, 16, 24, 32, 33, 16, 6, 
    4, 4, 0, 0, 8, 0, 27, 11, 32, 19, 23, 28, 36, 13, 3, 
    0, 0, 0, 0, 10, 2, 21, 2, 32, 24, 25, 21, 28, 3, 11, 
    0, 0, 0, 9, 11, 12, 20, 18, 32, 24, 22, 24, 24, 19, 4, 
    0, 0, 0, 1, 0, 31, 38, 0, 39, 32, 27, 22, 11, 28, 0, 
    0, 0, 0, 2, 0, 7, 32, 10, 28, 34, 22, 15, 9, 19, 23, 
    4, 7, 6, 2, 8, 19, 12, 26, 23, 28, 30, 18, 20, 15, 23, 
    4, 5, 13, 11, 19, 26, 12, 9, 17, 23, 27, 25, 16, 18, 18, 
    
    -- channel=485
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 25, 36, 37, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 33, 20, 13, 1, 0, 0, 
    0, 0, 8, 13, 0, 3, 10, 7, 0, 0, 0, 0, 0, 0, 1, 
    52, 69, 46, 0, 8, 7, 27, 12, 1, 0, 0, 0, 2, 11, 17, 
    15, 0, 0, 7, 16, 29, 0, 0, 5, 5, 2, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 0, 0, 8, 7, 0, 2, 0, 0, 0, 
    0, 3, 1, 0, 50, 50, 19, 10, 9, 4, 1, 3, 0, 0, 0, 
    10, 19, 53, 66, 20, 28, 2, 15, 0, 0, 7, 7, 2, 0, 0, 
    80, 56, 0, 0, 0, 0, 0, 0, 3, 0, 6, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 8, 
    0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 9, 7, 0, 0, 0, 
    0, 0, 0, 0, 5, 29, 0, 0, 13, 13, 16, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=486
    0, 0, 0, 0, 9, 3, 2, 0, 0, 1, 2, 1, 1, 2, 0, 
    0, 0, 3, 5, 12, 34, 12, 13, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 12, 22, 31, 42, 36, 7, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 19, 29, 30, 30, 38, 40, 30, 10, 7, 0, 0, 0, 
    0, 0, 0, 0, 30, 25, 9, 20, 35, 39, 41, 16, 4, 0, 0, 
    0, 0, 0, 0, 5, 31, 26, 19, 27, 32, 37, 39, 23, 0, 0, 
    0, 0, 0, 0, 31, 39, 19, 30, 24, 17, 29, 43, 23, 12, 0, 
    0, 0, 0, 0, 0, 7, 8, 29, 23, 12, 25, 37, 27, 18, 0, 
    0, 0, 0, 0, 0, 0, 0, 14, 31, 17, 19, 27, 34, 23, 18, 
    0, 0, 0, 0, 18, 0, 24, 5, 29, 23, 21, 24, 36, 17, 6, 
    0, 0, 0, 30, 34, 35, 33, 28, 30, 30, 27, 24, 30, 1, 2, 
    8, 9, 0, 0, 8, 37, 20, 8, 40, 31, 15, 15, 22, 24, 0, 
    3, 6, 0, 0, 0, 1, 34, 2, 23, 26, 6, 18, 5, 23, 7, 
    1, 3, 15, 24, 22, 3, 11, 27, 31, 50, 39, 23, 27, 20, 26, 
    16, 24, 20, 12, 19, 15, 12, 16, 18, 21, 36, 38, 23, 22, 16, 
    
    -- channel=487
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 5, 1, 0, 
    0, 0, 0, 0, 3, 18, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 21, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 9, 10, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 4, 1, 0, 0, 6, 20, 
    0, 6, 7, 4, 23, 14, 0, 0, 5, 3, 9, 5, 0, 14, 16, 
    
    -- channel=488
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 10, 0, 7, 0, 0, 0, 0, 0, 0, 1, 9, 
    0, 0, 0, 0, 2, 0, 0, 0, 1, 3, 0, 9, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 36, 5, 0, 0, 5, 9, 0, 0, 3, 0, 0, 0, 0, 
    0, 1, 0, 7, 0, 1, 16, 0, 0, 0, 7, 0, 1, 6, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 6, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 3, 0, 0, 31, 
    0, 0, 5, 50, 13, 42, 0, 16, 0, 0, 0, 8, 0, 20, 4, 
    0, 11, 100, 61, 30, 52, 18, 20, 0, 1, 14, 10, 0, 0, 0, 
    84, 88, 25, 9, 23, 10, 0, 9, 5, 0, 0, 0, 8, 0, 7, 
    25, 17, 7, 0, 0, 0, 0, 7, 0, 0, 0, 4, 6, 0, 0, 
    0, 0, 9, 35, 21, 0, 0, 3, 3, 6, 23, 12, 14, 10, 0, 
    16, 33, 18, 4, 0, 0, 0, 13, 4, 0, 1, 15, 19, 2, 7, 
    
    -- channel=489
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 23, 29, 29, 9, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 25, 30, 33, 36, 25, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 27, 20, 26, 37, 31, 26, 17, 0, 0, 0, 
    0, 0, 0, 0, 17, 18, 16, 27, 35, 38, 38, 34, 11, 2, 0, 
    0, 0, 0, 0, 1, 22, 22, 30, 27, 25, 34, 34, 16, 4, 0, 
    0, 0, 0, 0, 0, 1, 13, 29, 24, 19, 31, 32, 26, 8, 0, 
    0, 0, 0, 0, 0, 0, 11, 17, 25, 22, 28, 32, 28, 6, 0, 
    0, 0, 0, 0, 0, 0, 8, 19, 25, 22, 25, 29, 27, 10, 5, 
    0, 0, 0, 5, 9, 20, 18, 31, 26, 22, 26, 32, 24, 12, 0, 
    0, 0, 0, 0, 4, 32, 22, 0, 28, 30, 21, 22, 18, 14, 0, 
    0, 0, 0, 0, 0, 0, 15, 11, 15, 24, 9, 17, 17, 10, 14, 
    0, 0, 0, 0, 6, 5, 6, 12, 18, 16, 22, 23, 22, 17, 10, 
    0, 1, 8, 7, 8, 6, 3, 11, 13, 11, 13, 16, 18, 14, 10, 
    
    -- channel=490
    0, 0, 7, 10, 10, 0, 0, 3, 0, 0, 4, 4, 2, 1, 0, 
    0, 0, 2, 23, 0, 24, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    5, 1, 7, 23, 7, 2, 10, 4, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 8, 5, 0, 0, 0, 7, 30, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 0, 0, 
    9, 6, 0, 0, 14, 38, 0, 0, 0, 0, 0, 11, 0, 16, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 2, 3, 15, 
    0, 0, 13, 0, 25, 0, 18, 0, 0, 0, 0, 0, 1, 0, 3, 
    0, 0, 10, 40, 38, 40, 18, 25, 0, 0, 0, 0, 0, 0, 0, 
    67, 67, 1, 0, 0, 14, 0, 0, 21, 8, 0, 0, 0, 17, 0, 
    30, 25, 14, 0, 0, 0, 17, 0, 0, 4, 0, 0, 0, 7, 6, 
    7, 1, 12, 29, 33, 0, 0, 0, 8, 30, 37, 0, 0, 8, 20, 
    16, 32, 20, 5, 19, 7, 0, 2, 5, 1, 18, 21, 6, 11, 11, 
    
    -- channel=491
    0, 0, 0, 0, 0, 0, 5, 0, 3, 0, 0, 0, 2, 6, 17, 
    0, 2, 0, 0, 0, 0, 0, 6, 0, 6, 20, 30, 33, 32, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 27, 16, 13, 2, 0, 0, 
    0, 5, 40, 8, 0, 10, 12, 0, 0, 0, 0, 0, 1, 6, 9, 
    45, 50, 52, 17, 1, 0, 22, 17, 2, 0, 0, 0, 4, 16, 17, 
    5, 0, 14, 20, 23, 8, 0, 4, 7, 7, 6, 0, 0, 0, 1, 
    0, 0, 0, 75, 0, 0, 0, 0, 6, 13, 7, 0, 0, 0, 0, 
    0, 3, 2, 0, 81, 37, 26, 2, 1, 12, 9, 5, 0, 0, 9, 
    5, 18, 59, 70, 28, 50, 3, 17, 0, 3, 14, 13, 0, 0, 0, 
    53, 27, 0, 0, 0, 0, 0, 12, 0, 1, 9, 13, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 14, 15, 
    0, 0, 0, 0, 19, 0, 0, 26, 0, 0, 8, 16, 5, 0, 24, 
    0, 0, 0, 0, 8, 26, 0, 5, 3, 0, 16, 0, 17, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 
    
    -- channel=492
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 11, 18, 24, 25, 13, 
    0, 0, 0, 0, 0, 0, 0, 1, 26, 22, 11, 6, 0, 0, 0, 
    0, 7, 0, 8, 0, 8, 12, 9, 5, 1, 0, 0, 0, 0, 0, 
    49, 54, 0, 0, 4, 22, 16, 0, 1, 2, 2, 0, 13, 5, 9, 
    20, 2, 0, 0, 11, 46, 0, 0, 6, 0, 0, 12, 15, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 17, 0, 0, 0, 
    7, 14, 0, 0, 0, 52, 0, 12, 15, 0, 0, 3, 1, 9, 0, 
    24, 42, 45, 17, 0, 0, 0, 0, 9, 0, 0, 0, 15, 0, 0, 
    68, 46, 0, 0, 0, 0, 8, 0, 10, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 0, 
    0, 0, 0, 0, 0, 0, 25, 0, 0, 8, 10, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 12, 33, 5, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 14, 4, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    
    -- channel=493
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 1, 3, 8, 
    0, 2, 0, 0, 0, 0, 0, 4, 0, 1, 9, 17, 24, 27, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 24, 19, 14, 8, 2, 0, 
    0, 1, 20, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 5, 10, 
    25, 37, 47, 20, 0, 0, 17, 14, 0, 0, 0, 0, 9, 15, 19, 
    11, 0, 6, 16, 14, 0, 0, 3, 2, 4, 2, 0, 0, 5, 5, 
    0, 0, 0, 62, 0, 0, 1, 0, 0, 7, 1, 0, 0, 0, 0, 
    0, 2, 6, 0, 70, 12, 17, 0, 0, 10, 4, 1, 0, 0, 5, 
    7, 10, 30, 50, 33, 45, 3, 12, 0, 0, 7, 5, 0, 7, 0, 
    43, 38, 0, 18, 0, 0, 0, 10, 0, 0, 4, 7, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 16, 16, 
    0, 0, 0, 8, 7, 0, 0, 20, 0, 0, 1, 13, 8, 0, 25, 
    0, 0, 0, 0, 14, 37, 0, 1, 0, 0, 10, 0, 24, 2, 0, 
    0, 1, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 9, 5, 3, 2, 0, 0, 0, 0, 0, 
    
    -- channel=494
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 10, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 15, 19, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 15, 19, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 12, 16, 7, 8, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 8, 9, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 7, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 16, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 23, 12, 
    0, 0, 0, 2, 11, 0, 0, 2, 3, 0, 0, 0, 3, 26, 22, 
    0, 6, 15, 17, 20, 9, 6, 22, 25, 17, 15, 16, 20, 29, 25, 
    
    -- channel=495
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 14, 28, 35, 33, 23, 
    0, 0, 0, 0, 0, 0, 0, 2, 19, 29, 18, 11, 0, 0, 0, 
    0, 3, 20, 2, 2, 14, 20, 10, 0, 0, 0, 0, 0, 0, 4, 
    59, 69, 32, 1, 7, 23, 33, 14, 8, 1, 0, 0, 3, 14, 17, 
    12, 0, 0, 0, 30, 29, 0, 4, 16, 14, 6, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 8, 15, 13, 6, 6, 0, 0, 0, 
    0, 8, 0, 6, 49, 46, 22, 15, 14, 10, 9, 5, 0, 0, 4, 
    15, 31, 72, 49, 36, 20, 20, 11, 1, 5, 16, 11, 6, 0, 0, 
    79, 45, 0, 0, 0, 0, 0, 1, 7, 7, 14, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 6, 5, 16, 0, 
    0, 0, 0, 0, 0, 0, 20, 0, 0, 1, 18, 15, 0, 0, 5, 
    0, 0, 0, 0, 10, 26, 0, 1, 13, 22, 19, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=496
    6, 6, 10, 10, 13, 18, 17, 12, 10, 12, 11, 12, 13, 16, 18, 
    6, 8, 12, 9, 19, 18, 21, 24, 16, 18, 23, 26, 26, 25, 24, 
    6, 8, 10, 9, 21, 24, 28, 33, 28, 21, 22, 25, 21, 20, 23, 
    10, 13, 23, 23, 19, 25, 30, 37, 35, 28, 21, 25, 25, 26, 31, 
    22, 22, 24, 12, 17, 21, 24, 28, 35, 35, 31, 30, 34, 40, 41, 
    13, 10, 19, 11, 24, 27, 18, 19, 28, 33, 33, 30, 37, 42, 37, 
    6, 8, 16, 17, 21, 11, 18, 25, 26, 25, 32, 26, 29, 32, 25, 
    12, 16, 16, 21, 32, 31, 30, 30, 22, 19, 26, 27, 29, 30, 33, 
    16, 22, 31, 18, 27, 28, 34, 28, 18, 17, 23, 26, 25, 24, 34, 
    22, 15, 1, 5, 16, 31, 28, 24, 19, 16, 21, 23, 21, 31, 46, 
    5, 5, 0, 16, 9, 18, 13, 18, 21, 18, 22, 25, 28, 43, 48, 
    0, 0, 1, 12, 12, 17, 25, 16, 22, 21, 20, 26, 36, 45, 45, 
    4, 6, 15, 19, 21, 17, 24, 24, 20, 16, 16, 20, 36, 46, 48, 
    18, 20, 21, 25, 32, 40, 30, 31, 22, 14, 13, 14, 31, 46, 46, 
    21, 28, 38, 44, 45, 43, 35, 43, 47, 42, 33, 32, 39, 50, 50, 
    
    -- channel=497
    0, 0, 10, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 4, 4, 0, 15, 0, 0, 0, 0, 0, 0, 1, 2, 0, 
    0, 0, 0, 7, 0, 3, 7, 7, 13, 2, 0, 0, 0, 0, 0, 
    0, 2, 0, 7, 3, 2, 4, 10, 7, 15, 6, 0, 0, 0, 0, 
    14, 14, 0, 0, 5, 27, 1, 0, 0, 4, 13, 0, 6, 0, 0, 
    10, 1, 0, 0, 0, 39, 0, 0, 0, 0, 0, 15, 16, 0, 0, 
    1, 0, 0, 0, 9, 28, 0, 2, 8, 0, 0, 20, 0, 6, 0, 
    6, 6, 0, 0, 0, 24, 0, 11, 10, 0, 0, 0, 2, 7, 0, 
    12, 19, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 15, 0, 0, 
    17, 12, 0, 0, 14, 0, 25, 0, 7, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 20, 0, 14, 13, 2, 0, 0, 23, 0, 
    0, 0, 0, 0, 0, 0, 19, 0, 12, 31, 0, 0, 0, 6, 4, 
    0, 3, 0, 0, 0, 0, 2, 0, 0, 14, 9, 0, 0, 0, 11, 
    0, 0, 0, 0, 17, 9, 0, 0, 0, 0, 10, 1, 0, 2, 0, 
    
    -- channel=498
    14, 15, 17, 18, 26, 35, 25, 20, 17, 18, 17, 16, 16, 16, 16, 
    14, 15, 18, 20, 35, 44, 47, 39, 25, 22, 24, 24, 25, 24, 24, 
    15, 16, 18, 29, 41, 51, 55, 60, 50, 29, 31, 32, 29, 27, 28, 
    18, 18, 19, 26, 44, 50, 57, 68, 60, 49, 40, 38, 31, 28, 35, 
    21, 22, 22, 32, 44, 51, 52, 59, 68, 65, 61, 56, 43, 44, 46, 
    22, 21, 24, 27, 42, 42, 44, 55, 60, 66, 67, 61, 56, 52, 46, 
    20, 20, 25, 21, 32, 46, 53, 58, 54, 55, 63, 62, 56, 46, 35, 
    22, 24, 25, 42, 31, 32, 47, 59, 53, 51, 59, 61, 55, 41, 37, 
    25, 26, 27, 22, 44, 35, 51, 53, 50, 49, 56, 59, 54, 48, 46, 
    25, 24, 24, 37, 37, 48, 44, 56, 50, 48, 54, 58, 54, 49, 50, 
    19, 19, 13, 27, 43, 47, 48, 56, 54, 53, 54, 57, 57, 55, 48, 
    16, 14, 29, 30, 27, 47, 51, 29, 43, 51, 48, 53, 59, 57, 52, 
    21, 20, 22, 29, 38, 38, 43, 45, 42, 48, 41, 50, 63, 57, 58, 
    26, 29, 34, 40, 43, 47, 41, 47, 48, 43, 42, 47, 57, 61, 54, 
    33, 39, 48, 51, 53, 49, 49, 57, 56, 52, 48, 52, 58, 60, 56, 
    
    -- channel=499
    31, 28, 31, 33, 37, 40, 31, 28, 22, 19, 14, 10, 6, 5, 3, 
    30, 27, 30, 25, 38, 42, 41, 32, 24, 21, 18, 19, 20, 20, 19, 
    28, 27, 21, 23, 33, 35, 39, 41, 38, 38, 36, 36, 31, 27, 21, 
    26, 27, 16, 19, 32, 33, 38, 46, 42, 47, 47, 38, 30, 26, 24, 
    44, 54, 46, 18, 31, 45, 50, 44, 47, 44, 50, 47, 37, 37, 36, 
    66, 69, 55, 19, 30, 50, 50, 46, 47, 47, 45, 47, 46, 46, 41, 
    63, 62, 60, 20, 33, 46, 48, 48, 52, 46, 45, 47, 43, 42, 30, 
    60, 64, 64, 63, 33, 37, 43, 51, 57, 50, 46, 42, 43, 33, 29, 
    69, 78, 85, 64, 74, 50, 58, 50, 55, 52, 48, 44, 45, 35, 24, 
    100, 108, 106, 85, 79, 67, 59, 51, 53, 54, 53, 46, 40, 21, 17, 
    115, 107, 52, 58, 53, 53, 46, 45, 52, 53, 50, 45, 36, 31, 19, 
    84, 68, 53, 48, 27, 33, 42, 23, 40, 46, 50, 46, 33, 39, 24, 
    46, 42, 41, 43, 42, 29, 40, 34, 40, 52, 54, 51, 37, 31, 39, 
    35, 38, 38, 31, 27, 35, 30, 36, 32, 36, 49, 44, 37, 27, 31, 
    29, 24, 24, 21, 24, 35, 31, 26, 24, 25, 27, 31, 26, 23, 22, 
    
    -- channel=500
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 11, 
    0, 0, 0, 1, 0, 0, 0, 2, 2, 6, 14, 15, 9, 4, 1, 
    0, 0, 0, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 
    0, 4, 23, 7, 2, 8, 6, 0, 0, 0, 0, 0, 2, 2, 3, 
    18, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 
    0, 0, 0, 0, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 6, 24, 0, 0, 0, 0, 0, 0, 0, 3, 9, 
    0, 15, 26, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 6, 2, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 7, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 3, 0, 0, 0, 0, 3, 4, 1, 0, 1, 0, 0, 
    
    -- channel=501
    0, 0, 0, 0, 0, 0, 8, 6, 5, 2, 9, 15, 9, 0, 1, 
    0, 4, 0, 6, 8, 0, 22, 9, 8, 0, 0, 0, 0, 0, 0, 
    0, 2, 21, 0, 22, 4, 5, 0, 0, 0, 0, 0, 0, 3, 16, 
    0, 0, 26, 0, 9, 0, 0, 0, 0, 0, 0, 20, 0, 6, 1, 
    0, 0, 23, 55, 0, 0, 0, 19, 2, 1, 0, 4, 0, 0, 0, 
    0, 0, 90, 42, 0, 0, 13, 32, 0, 6, 6, 0, 0, 0, 0, 
    0, 0, 11, 85, 0, 0, 37, 7, 0, 12, 21, 0, 0, 0, 25, 
    0, 0, 0, 14, 60, 0, 7, 0, 0, 25, 26, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 27, 0, 16, 0, 21, 16, 20, 0, 0, 33, 
    0, 0, 0, 114, 0, 80, 0, 50, 0, 3, 9, 33, 0, 36, 4, 
    0, 14, 163, 58, 21, 62, 12, 16, 0, 4, 21, 30, 3, 0, 6, 
    72, 86, 60, 28, 57, 6, 0, 32, 0, 0, 0, 16, 20, 0, 34, 
    28, 12, 7, 0, 28, 3, 0, 31, 0, 0, 0, 20, 31, 0, 0, 
    0, 0, 10, 36, 16, 0, 0, 7, 6, 0, 12, 27, 24, 7, 0, 
    17, 32, 18, 7, 0, 0, 5, 21, 3, 0, 0, 7, 26, 0, 0, 
    
    -- channel=502
    7, 7, 10, 8, 16, 24, 16, 12, 9, 9, 9, 7, 7, 8, 8, 
    7, 7, 10, 11, 24, 33, 33, 28, 17, 13, 15, 15, 15, 14, 14, 
    7, 9, 10, 16, 29, 39, 44, 48, 38, 21, 20, 22, 21, 18, 18, 
    10, 10, 10, 17, 34, 41, 47, 54, 50, 39, 28, 28, 22, 18, 23, 
    14, 15, 14, 19, 35, 41, 42, 46, 57, 52, 50, 44, 32, 31, 34, 
    16, 15, 16, 15, 30, 36, 36, 43, 52, 55, 58, 51, 44, 41, 37, 
    13, 14, 16, 8, 26, 36, 40, 46, 46, 44, 52, 52, 45, 39, 27, 
    14, 16, 17, 27, 20, 26, 38, 49, 46, 39, 48, 50, 46, 33, 26, 
    19, 21, 22, 15, 31, 26, 38, 43, 43, 38, 45, 48, 46, 36, 35, 
    19, 18, 16, 20, 31, 36, 36, 44, 43, 39, 44, 46, 44, 37, 39, 
    14, 13, 6, 25, 29, 39, 41, 44, 44, 43, 44, 47, 45, 42, 36, 
    9, 10, 13, 21, 23, 38, 40, 23, 36, 42, 40, 42, 46, 47, 39, 
    11, 11, 14, 18, 25, 26, 36, 33, 33, 39, 33, 38, 46, 46, 47, 
    16, 19, 23, 28, 33, 35, 32, 37, 39, 36, 35, 37, 45, 49, 46, 
    22, 28, 36, 38, 41, 41, 36, 43, 44, 40, 38, 40, 44, 47, 46, 
    
    -- channel=503
    0, 3, 2, 1, 15, 14, 14, 4, 5, 6, 8, 9, 10, 11, 11, 
    1, 1, 4, 19, 19, 31, 20, 28, 15, 11, 15, 9, 4, 1, 1, 
    5, 3, 10, 14, 36, 43, 54, 49, 16, 0, 1, 3, 4, 2, 9, 
    6, 7, 9, 39, 46, 50, 50, 50, 52, 27, 16, 21, 5, 9, 12, 
    0, 0, 0, 26, 41, 22, 26, 49, 50, 54, 47, 25, 14, 11, 10, 
    0, 0, 0, 29, 27, 39, 44, 41, 42, 53, 54, 48, 28, 9, 7, 
    0, 0, 0, 10, 29, 25, 31, 47, 35, 41, 47, 52, 30, 9, 7, 
    0, 0, 0, 0, 1, 35, 34, 42, 29, 34, 48, 53, 34, 29, 11, 
    0, 0, 0, 9, 0, 1, 1, 43, 38, 36, 42, 49, 41, 28, 23, 
    0, 0, 0, 0, 17, 0, 29, 36, 40, 39, 39, 48, 48, 36, 16, 
    0, 0, 31, 34, 32, 36, 38, 33, 36, 38, 42, 49, 46, 15, 21, 
    0, 6, 0, 0, 40, 51, 22, 41, 46, 43, 27, 38, 43, 21, 14, 
    2, 7, 9, 3, 0, 15, 32, 19, 35, 33, 18, 36, 28, 32, 10, 
    10, 7, 15, 26, 29, 11, 31, 34, 40, 47, 31, 40, 40, 29, 28, 
    15, 27, 29, 25, 23, 16, 23, 30, 31, 30, 42, 40, 35, 30, 22, 
    
    -- channel=504
    0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=505
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 7, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 36, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=506
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 
    9, 15, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=507
    0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 1, 4, 3, 0, 6, 
    0, 1, 0, 0, 1, 0, 12, 0, 0, 4, 1, 1, 0, 0, 1, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 4, 6, 
    0, 0, 29, 22, 0, 0, 0, 3, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 68, 4, 11, 0, 0, 12, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 15, 55, 0, 0, 17, 1, 0, 3, 8, 0, 0, 0, 7, 
    0, 0, 0, 19, 64, 0, 8, 0, 0, 12, 9, 0, 0, 0, 3, 
    0, 0, 8, 0, 28, 23, 12, 0, 0, 8, 7, 6, 0, 0, 11, 
    0, 0, 0, 76, 0, 60, 0, 20, 0, 0, 3, 11, 0, 13, 7, 
    0, 0, 47, 8, 0, 13, 0, 0, 0, 0, 6, 12, 0, 13, 3, 
    0, 16, 27, 22, 21, 0, 0, 7, 0, 0, 0, 11, 0, 0, 28, 
    0, 0, 0, 0, 25, 4, 0, 21, 0, 0, 0, 2, 19, 0, 5, 
    0, 0, 0, 4, 1, 7, 0, 0, 0, 0, 0, 8, 4, 3, 0, 
    0, 5, 7, 4, 0, 0, 0, 11, 1, 0, 0, 0, 13, 0, 0, 
    
    -- channel=508
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 16, 1, 0, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 5, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 4, 11, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=509
    0, 0, 0, 0, 0, 0, 2, 0, 1, 0, 1, 5, 3, 0, 3, 
    0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 7, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 7, 
    0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 5, 3, 
    0, 0, 30, 37, 0, 0, 0, 13, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 49, 33, 0, 0, 1, 10, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 2, 71, 0, 0, 8, 0, 0, 5, 4, 0, 0, 0, 11, 
    0, 0, 0, 4, 60, 0, 9, 0, 0, 10, 9, 0, 0, 0, 0, 
    0, 0, 0, 22, 2, 31, 0, 14, 0, 3, 4, 5, 0, 0, 15, 
    0, 0, 0, 57, 0, 35, 0, 24, 0, 0, 0, 12, 0, 17, 2, 
    0, 8, 92, 3, 0, 8, 0, 0, 0, 0, 3, 8, 0, 0, 13, 
    18, 18, 20, 15, 34, 0, 0, 27, 0, 0, 0, 8, 10, 0, 27, 
    0, 0, 0, 0, 13, 10, 0, 9, 0, 0, 0, 6, 18, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 4, 8, 2, 0, 
    5, 8, 2, 4, 0, 0, 3, 11, 2, 0, 0, 0, 9, 0, 0, 
    
    -- channel=510
    0, 1, 0, 0, 0, 4, 6, 0, 5, 3, 2, 4, 5, 4, 15, 
    0, 6, 0, 0, 1, 0, 8, 9, 0, 7, 15, 21, 21, 20, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 13, 12, 3, 2, 3, 
    0, 3, 47, 0, 0, 7, 5, 0, 0, 0, 0, 7, 4, 9, 12, 
    20, 24, 61, 28, 0, 0, 16, 19, 3, 1, 0, 2, 5, 16, 15, 
    0, 0, 49, 18, 23, 0, 0, 16, 6, 7, 6, 0, 0, 3, 5, 
    0, 0, 8, 94, 0, 0, 9, 3, 0, 15, 11, 0, 1, 0, 0, 
    0, 0, 5, 2, 94, 0, 25, 0, 0, 20, 14, 3, 0, 0, 10, 
    0, 3, 41, 47, 43, 60, 10, 13, 0, 10, 16, 14, 0, 0, 0, 
    20, 7, 0, 54, 0, 32, 0, 24, 0, 1, 10, 18, 0, 18, 6, 
    0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 2, 15, 4, 21, 15, 
    0, 0, 11, 12, 30, 0, 0, 27, 0, 0, 2, 22, 10, 0, 40, 
    0, 0, 0, 0, 18, 26, 0, 19, 0, 0, 14, 7, 34, 0, 0, 
    0, 0, 0, 0, 0, 4, 2, 0, 0, 0, 0, 4, 6, 1, 0, 
    0, 0, 0, 4, 0, 0, 8, 8, 2, 2, 0, 0, 5, 0, 0, 
    
    -- channel=511
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 5, 4, 6, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 6, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 18, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 15, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 39, 
    0, 0, 0, 7, 0, 5, 0, 0, 0, 0, 0, 0, 0, 23, 33, 
    0, 0, 49, 13, 3, 10, 0, 5, 0, 0, 0, 0, 0, 9, 26, 
    32, 38, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 14, 28, 
    11, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 21, 20, 
    0, 0, 8, 31, 33, 10, 0, 1, 1, 0, 0, 0, 6, 32, 27, 
    18, 35, 33, 30, 24, 13, 15, 32, 28, 17, 12, 21, 31, 35, 36, 
    
    -- channel=512
    0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 8, 16, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 24, 1, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=513
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 9, 0, 3, 2, 8, 7, 0, 6, 0, 0, 0, 
    0, 0, 0, 0, 17, 22, 0, 0, 15, 0, 0, 9, 15, 12, 8, 
    0, 0, 0, 0, 20, 27, 0, 0, 0, 0, 29, 7, 22, 32, 15, 
    11, 0, 11, 0, 0, 18, 23, 12, 0, 0, 11, 16, 25, 18, 0, 
    13, 3, 19, 0, 8, 17, 24, 0, 0, 0, 2, 18, 28, 24, 0, 
    9, 2, 5, 19, 2, 0, 16, 0, 15, 4, 0, 16, 25, 33, 0, 
    9, 6, 12, 8, 16, 19, 17, 0, 19, 0, 19, 4, 37, 38, 14, 
    20, 0, 13, 0, 26, 22, 5, 26, 0, 0, 21, 0, 0, 26, 7, 
    20, 0, 16, 17, 9, 25, 34, 16, 0, 0, 10, 0, 0, 1, 0, 
    19, 11, 16, 10, 15, 20, 9, 12, 29, 13, 0, 0, 3, 0, 0, 
    15, 25, 3, 24, 28, 16, 9, 9, 16, 6, 0, 0, 11, 0, 0, 
    14, 15, 1, 25, 37, 0, 18, 10, 15, 0, 0, 0, 3, 2, 0, 
    13, 9, 0, 27, 24, 0, 9, 3, 0, 0, 0, 0, 0, 0, 0, 
    8, 11, 0, 28, 20, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=514
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 32, 32, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 47, 7, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 5, 0, 0, 0, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 0, 5, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 
    10, 0, 1, 0, 0, 0, 15, 3, 2, 0, 0, 0, 0, 0, 0, 
    
    -- channel=515
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=516
    12, 35, 24, 19, 22, 20, 16, 21, 21, 7, 39, 32, 22, 18, 16, 
    12, 23, 33, 28, 43, 29, 31, 29, 28, 0, 59, 31, 27, 25, 23, 
    11, 15, 39, 32, 62, 22, 22, 30, 21, 28, 52, 35, 37, 40, 35, 
    4, 28, 55, 18, 62, 39, 29, 23, 31, 51, 40, 53, 49, 33, 33, 
    18, 38, 28, 2, 60, 48, 37, 17, 34, 44, 43, 51, 39, 7, 23, 
    24, 29, 22, 13, 53, 45, 27, 22, 41, 46, 40, 53, 35, 7, 9, 
    18, 22, 9, 31, 33, 41, 35, 44, 38, 43, 42, 51, 37, 29, 12, 
    14, 26, 11, 61, 41, 41, 40, 39, 33, 33, 28, 32, 36, 30, 23, 
    7, 23, 40, 57, 45, 52, 45, 27, 36, 16, 34, 2, 33, 15, 31, 
    16, 26, 45, 39, 42, 46, 47, 37, 24, 39, 19, 23, 27, 25, 22, 
    24, 18, 45, 41, 42, 24, 45, 43, 32, 22, 17, 35, 35, 19, 24, 
    25, 12, 49, 49, 43, 28, 42, 39, 32, 5, 34, 27, 37, 22, 15, 
    19, 7, 35, 45, 29, 23, 43, 29, 20, 12, 29, 22, 28, 20, 21, 
    14, 0, 25, 48, 31, 42, 28, 19, 14, 9, 26, 21, 14, 26, 28, 
    7, 3, 18, 51, 34, 30, 12, 19, 8, 20, 20, 24, 16, 27, 23, 
    
    -- channel=517
    0, 0, 2, 1, 0, 4, 9, 6, 15, 0, 0, 1, 12, 12, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    32, 36, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=518
    9, 0, 0, 5, 5, 0, 7, 3, 46, 28, 0, 14, 14, 8, 11, 
    6, 0, 0, 0, 31, 5, 0, 4, 8, 56, 0, 15, 12, 7, 9, 
    7, 0, 0, 0, 3, 50, 0, 0, 0, 13, 0, 0, 7, 13, 19, 
    78, 25, 2, 2, 0, 47, 55, 30, 4, 0, 8, 0, 20, 10, 0, 
    44, 12, 8, 24, 0, 4, 25, 29, 1, 0, 0, 0, 8, 15, 0, 
    6, 0, 1, 20, 0, 2, 21, 15, 23, 0, 0, 0, 3, 26, 0, 
    0, 0, 0, 11, 4, 0, 27, 3, 27, 3, 0, 0, 0, 25, 13, 
    0, 0, 41, 0, 20, 11, 20, 17, 3, 0, 1, 0, 0, 0, 0, 
    16, 0, 39, 0, 24, 39, 30, 50, 0, 5, 18, 21, 0, 0, 0, 
    15, 0, 8, 14, 0, 0, 12, 42, 42, 3, 5, 4, 12, 9, 0, 
    0, 5, 0, 11, 13, 21, 0, 0, 27, 10, 0, 4, 7, 10, 0, 
    0, 18, 0, 8, 12, 14, 8, 8, 12, 26, 0, 0, 6, 15, 18, 
    0, 0, 0, 6, 23, 0, 0, 0, 4, 9, 0, 0, 0, 0, 10, 
    0, 0, 0, 1, 37, 34, 2, 0, 0, 0, 0, 0, 8, 0, 6, 
    0, 0, 0, 0, 14, 11, 0, 0, 8, 0, 0, 2, 15, 0, 0, 
    
    -- channel=519
    9, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 2, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 1, 1, 2, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 8, 0, 9, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 6, 7, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 10, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 5, 0, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=520
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 0, 2, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 5, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 4, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=521
    7, 0, 17, 33, 26, 20, 30, 22, 39, 51, 0, 21, 33, 31, 37, 
    6, 0, 2, 14, 15, 24, 13, 13, 31, 65, 0, 21, 31, 31, 35, 
    7, 0, 0, 12, 0, 54, 23, 15, 33, 3, 0, 5, 17, 16, 22, 
    37, 0, 0, 36, 0, 35, 30, 34, 13, 0, 15, 0, 19, 31, 2, 
    28, 0, 15, 46, 0, 16, 34, 46, 9, 0, 0, 0, 18, 43, 0, 
    18, 9, 21, 30, 0, 17, 43, 28, 12, 0, 0, 0, 14, 36, 7, 
    18, 12, 42, 15, 23, 7, 40, 0, 27, 0, 0, 0, 10, 22, 15, 
    23, 11, 64, 0, 27, 15, 23, 24, 7, 6, 23, 0, 0, 27, 0, 
    34, 7, 34, 6, 14, 13, 21, 53, 0, 23, 25, 31, 0, 25, 0, 
    24, 4, 14, 18, 11, 19, 15, 27, 31, 8, 42, 24, 11, 27, 8, 
    12, 25, 0, 18, 13, 42, 1, 14, 34, 46, 18, 14, 19, 36, 24, 
    10, 33, 0, 16, 29, 31, 11, 19, 31, 53, 0, 22, 17, 32, 32, 
    14, 25, 0, 16, 56, 21, 17, 26, 41, 36, 8, 21, 27, 22, 25, 
    19, 24, 0, 6, 43, 16, 39, 29, 38, 23, 13, 20, 33, 5, 17, 
    18, 17, 0, 0, 23, 38, 40, 24, 42, 4, 17, 19, 25, 12, 18, 
    
    -- channel=522
    0, 64, 6, 0, 0, 0, 0, 0, 0, 0, 39, 0, 0, 0, 0, 
    0, 22, 43, 0, 0, 0, 5, 0, 0, 0, 38, 0, 0, 0, 0, 
    0, 0, 62, 0, 15, 0, 0, 23, 6, 0, 10, 9, 0, 0, 0, 
    0, 0, 6, 0, 47, 0, 0, 0, 0, 31, 7, 19, 0, 0, 21, 
    0, 0, 0, 0, 29, 2, 0, 0, 0, 20, 25, 22, 0, 0, 17, 
    0, 0, 0, 0, 14, 4, 0, 0, 0, 0, 17, 40, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 1, 7, 37, 7, 0, 0, 
    0, 2, 0, 44, 0, 0, 0, 0, 15, 2, 0, 80, 54, 0, 1, 
    0, 0, 0, 15, 0, 0, 0, 0, 30, 0, 0, 0, 58, 25, 55, 
    0, 0, 0, 0, 8, 17, 5, 0, 0, 0, 0, 0, 0, 0, 21, 
    0, 0, 17, 0, 0, 0, 22, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 24, 0, 0, 2, 12, 0, 0, 0, 5, 0, 4, 0, 0, 
    0, 0, 23, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 8, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=523
    50, 62, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 
    49, 59, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 0, 0, 0, 
    45, 50, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    49, 95, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=524
    0, 20, 5, 0, 6, 5, 6, 9, 3, 7, 20, 1, 5, 6, 4, 
    1, 20, 0, 1, 0, 5, 0, 6, 0, 0, 34, 5, 4, 6, 2, 
    0, 8, 3, 14, 0, 0, 0, 0, 0, 5, 14, 3, 3, 6, 6, 
    24, 35, 24, 1, 0, 0, 11, 0, 0, 13, 0, 11, 0, 0, 2, 
    7, 27, 5, 0, 2, 0, 0, 0, 0, 6, 0, 10, 2, 0, 14, 
    5, 7, 0, 12, 0, 0, 0, 0, 3, 12, 3, 7, 4, 10, 17, 
    7, 7, 0, 5, 0, 1, 0, 1, 0, 0, 7, 8, 4, 6, 17, 
    8, 4, 0, 0, 0, 0, 0, 7, 0, 1, 0, 0, 1, 0, 17, 
    6, 5, 0, 3, 0, 0, 3, 0, 2, 6, 0, 14, 0, 0, 10, 
    7, 16, 0, 0, 0, 0, 0, 0, 19, 9, 0, 0, 15, 0, 3, 
    7, 8, 0, 3, 4, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    7, 1, 6, 0, 0, 0, 4, 0, 0, 0, 11, 0, 0, 0, 0, 
    8, 4, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    6, 9, 16, 0, 0, 19, 0, 0, 0, 0, 0, 2, 0, 4, 1, 
    3, 10, 17, 0, 0, 0, 0, 0, 0, 14, 0, 1, 1, 4, 0, 
    
    -- channel=525
    9, 0, 1, 0, 2, 3, 6, 3, 2, 17, 0, 1, 4, 5, 6, 
    9, 2, 1, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    10, 7, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 10, 3, 0, 0, 0, 0, 5, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 10, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    2, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 1, 1, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 1, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 2, 
    1, 11, 0, 0, 0, 0, 0, 0, 3, 3, 1, 0, 4, 0, 0, 
    2, 9, 1, 0, 0, 0, 2, 0, 8, 1, 1, 0, 2, 2, 0, 
    
    -- channel=526
    0, 9, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9, 26, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 6, 0, 0, 0, 11, 39, 41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 63, 23, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 50, 16, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 7, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 9, 1, 3, 10, 2, 0, 0, 17, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 12, 2, 0, 0, 0, 0, 0, 
    14, 0, 0, 4, 0, 0, 20, 11, 7, 0, 0, 0, 0, 0, 2, 
    
    -- channel=527
    0, 100, 28, 0, 0, 4, 0, 3, 0, 0, 89, 5, 0, 0, 0, 
    1, 56, 62, 15, 0, 0, 3, 8, 0, 0, 106, 0, 0, 0, 0, 
    0, 18, 102, 15, 36, 0, 0, 17, 0, 14, 39, 9, 0, 0, 0, 
    0, 61, 59, 0, 52, 0, 0, 0, 7, 59, 2, 39, 0, 0, 13, 
    0, 19, 0, 0, 60, 0, 0, 0, 9, 38, 26, 35, 0, 0, 19, 
    0, 0, 0, 0, 25, 0, 0, 0, 5, 30, 19, 49, 0, 0, 0, 
    0, 0, 0, 15, 0, 15, 0, 15, 0, 14, 21, 46, 0, 0, 0, 
    0, 0, 0, 73, 0, 0, 0, 0, 19, 1, 0, 24, 35, 0, 1, 
    0, 2, 0, 33, 0, 0, 0, 0, 37, 0, 0, 0, 56, 0, 47, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 18, 0, 3, 8, 0, 18, 
    0, 0, 24, 0, 0, 0, 28, 3, 0, 0, 5, 9, 0, 0, 0, 
    0, 0, 40, 0, 0, 0, 11, 0, 0, 0, 31, 0, 6, 0, 0, 
    0, 0, 29, 0, 0, 6, 21, 0, 0, 0, 21, 0, 0, 0, 0, 
    0, 0, 30, 7, 0, 0, 0, 0, 0, 0, 11, 0, 0, 24, 3, 
    0, 0, 12, 29, 0, 0, 0, 0, 0, 21, 2, 2, 0, 6, 4, 
    
    -- channel=528
    12, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 11, 0, 0, 3, 0, 0, 0, 0, 0, 33, 0, 0, 0, 0, 
    11, 10, 0, 0, 4, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    33, 43, 46, 0, 0, 0, 14, 0, 0, 7, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 8, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 1, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 12, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=529
    0, 0, 13, 25, 17, 11, 22, 15, 30, 37, 0, 18, 27, 26, 30, 
    0, 0, 0, 0, 8, 18, 11, 13, 34, 46, 0, 25, 31, 29, 31, 
    0, 0, 0, 0, 0, 51, 8, 10, 27, 0, 2, 17, 29, 26, 27, 
    16, 0, 0, 39, 0, 30, 18, 22, 0, 0, 27, 0, 29, 52, 14, 
    39, 0, 29, 44, 0, 14, 36, 38, 0, 0, 2, 12, 37, 61, 17, 
    34, 21, 40, 28, 2, 18, 39, 7, 7, 0, 0, 8, 40, 66, 34, 
    37, 23, 48, 22, 20, 0, 41, 0, 26, 0, 0, 8, 36, 50, 36, 
    45, 20, 56, 0, 34, 19, 17, 23, 3, 3, 30, 9, 15, 60, 22, 
    61, 11, 22, 0, 19, 20, 20, 49, 0, 12, 33, 23, 0, 39, 0, 
    50, 17, 20, 23, 19, 29, 19, 19, 28, 7, 38, 14, 0, 28, 9, 
    37, 45, 6, 22, 24, 48, 3, 15, 36, 50, 0, 8, 15, 25, 20, 
    34, 57, 0, 25, 39, 27, 13, 20, 35, 40, 0, 17, 16, 26, 18, 
    39, 50, 3, 27, 63, 0, 20, 26, 38, 26, 3, 12, 21, 9, 17, 
    42, 50, 0, 22, 42, 1, 33, 25, 30, 2, 7, 10, 20, 0, 11, 
    34, 41, 3, 9, 30, 44, 34, 16, 31, 0, 4, 11, 9, 6, 8, 
    
    -- channel=530
    0, 0, 0, 4, 3, 0, 9, 6, 42, 16, 0, 14, 19, 14, 16, 
    0, 0, 0, 0, 21, 2, 0, 0, 0, 31, 0, 18, 19, 14, 14, 
    0, 0, 0, 0, 0, 31, 0, 0, 0, 3, 0, 0, 10, 18, 24, 
    65, 25, 3, 0, 0, 30, 47, 13, 0, 0, 0, 0, 16, 0, 0, 
    33, 13, 1, 13, 0, 0, 8, 6, 0, 0, 0, 0, 8, 6, 0, 
    0, 0, 0, 17, 0, 0, 0, 0, 5, 0, 0, 0, 3, 22, 0, 
    0, 0, 0, 2, 0, 0, 9, 0, 4, 0, 0, 0, 0, 24, 18, 
    0, 0, 31, 0, 9, 0, 2, 3, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 34, 0, 15, 31, 26, 26, 0, 0, 0, 16, 0, 0, 0, 
    9, 3, 4, 4, 0, 0, 0, 32, 43, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 9, 8, 7, 0, 0, 11, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 3, 1, 1, 2, 0, 0, 8, 0, 0, 0, 3, 3, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=531
    0, 0, 15, 24, 20, 14, 22, 21, 27, 15, 0, 34, 37, 34, 34, 
    0, 0, 0, 16, 36, 27, 20, 28, 36, 20, 11, 45, 44, 41, 41, 
    0, 0, 0, 22, 43, 47, 8, 8, 13, 8, 35, 34, 48, 49, 48, 
    4, 0, 22, 26, 31, 48, 37, 19, 4, 13, 42, 43, 68, 60, 37, 
    30, 32, 36, 22, 25, 43, 45, 26, 7, 12, 29, 50, 62, 43, 24, 
    38, 35, 35, 28, 34, 42, 37, 13, 21, 20, 31, 43, 59, 47, 21, 
    34, 31, 28, 33, 33, 27, 38, 18, 35, 25, 30, 45, 58, 59, 39, 
    34, 30, 41, 29, 48, 42, 32, 41, 18, 23, 34, 14, 39, 59, 41, 
    37, 19, 40, 44, 48, 57, 53, 38, 5, 24, 30, 20, 3, 19, 22, 
    37, 31, 45, 47, 41, 47, 49, 46, 44, 27, 24, 15, 21, 27, 17, 
    41, 39, 34, 50, 51, 44, 30, 44, 43, 34, 7, 23, 31, 22, 17, 
    39, 37, 32, 56, 57, 39, 43, 44, 44, 21, 13, 23, 29, 27, 14, 
    37, 25, 25, 53, 51, 16, 38, 35, 30, 16, 11, 16, 17, 10, 17, 
    34, 20, 11, 47, 46, 47, 33, 22, 16, 0, 8, 12, 9, 3, 18, 
    18, 14, 5, 38, 47, 41, 18, 10, 7, 0, 4, 11, 8, 11, 10, 
    
    -- channel=532
    0, 71, 19, 0, 0, 0, 0, 1, 0, 0, 51, 14, 0, 0, 0, 
    0, 35, 54, 0, 0, 0, 0, 0, 0, 0, 84, 0, 0, 0, 0, 
    0, 9, 86, 7, 23, 0, 0, 11, 0, 0, 44, 4, 0, 0, 0, 
    0, 42, 77, 0, 36, 0, 0, 0, 5, 40, 0, 29, 0, 0, 0, 
    0, 20, 0, 0, 51, 0, 0, 0, 2, 20, 16, 32, 0, 0, 13, 
    0, 0, 0, 0, 25, 0, 0, 0, 7, 17, 7, 40, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 7, 8, 37, 0, 0, 0, 
    0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 16, 9, 0, 0, 
    0, 1, 0, 28, 0, 0, 0, 0, 27, 0, 0, 0, 45, 0, 25, 
    0, 0, 5, 0, 3, 0, 0, 0, 0, 10, 0, 0, 0, 0, 9, 
    0, 0, 16, 0, 0, 0, 18, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 35, 0, 0, 0, 7, 0, 0, 0, 23, 0, 3, 0, 0, 
    0, 0, 23, 0, 0, 0, 11, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 22, 6, 0, 0, 0, 0, 0, 0, 10, 0, 0, 12, 0, 
    0, 0, 10, 20, 0, 0, 0, 0, 0, 4, 0, 0, 0, 6, 0, 
    
    -- channel=533
    12, 0, 0, 0, 0, 0, 0, 0, 32, 58, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 5, 0, 0, 0, 57, 0, 0, 0, 0, 0, 
    9, 0, 0, 0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    103, 10, 0, 6, 0, 15, 41, 30, 0, 0, 0, 0, 0, 0, 0, 
    23, 0, 0, 38, 0, 0, 1, 27, 0, 0, 0, 0, 0, 21, 0, 
    0, 0, 0, 15, 0, 0, 10, 10, 0, 0, 0, 0, 0, 30, 0, 
    0, 0, 0, 0, 3, 0, 17, 0, 4, 0, 0, 0, 0, 0, 17, 
    0, 0, 37, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 4, 0, 0, 1, 15, 41, 0, 0, 0, 29, 0, 0, 0, 
    9, 0, 0, 0, 0, 0, 0, 14, 46, 0, 0, 0, 0, 0, 0, 
    0, 8, 0, 0, 0, 18, 0, 0, 0, 7, 0, 0, 0, 3, 0, 
    0, 16, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 2, 8, 
    0, 0, 0, 0, 19, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 4, 0, 0, 
    
    -- channel=534
    9, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 
    8, 3, 0, 0, 0, 15, 12, 0, 19, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 15, 0, 0, 9, 11, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 26, 0, 19, 0, 0, 0, 0, 0, 0, 
    
    -- channel=535
    19, 98, 0, 0, 0, 0, 0, 0, 0, 0, 51, 0, 0, 0, 0, 
    21, 70, 20, 9, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 0, 
    20, 37, 50, 2, 0, 0, 1, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 36, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    
    -- channel=536
    0, 0, 35, 30, 26, 25, 28, 27, 15, 0, 8, 44, 44, 42, 41, 
    0, 0, 31, 29, 37, 29, 35, 41, 48, 7, 31, 50, 48, 49, 49, 
    0, 0, 10, 29, 59, 35, 21, 36, 32, 13, 50, 53, 57, 54, 49, 
    0, 0, 32, 30, 58, 45, 21, 14, 12, 35, 58, 61, 73, 69, 58, 
    27, 36, 47, 18, 48, 57, 49, 23, 17, 29, 52, 70, 73, 48, 47, 
    47, 48, 50, 26, 51, 56, 42, 15, 23, 30, 49, 72, 73, 47, 35, 
    47, 45, 45, 46, 39, 37, 39, 27, 39, 35, 45, 72, 77, 65, 40, 
    46, 45, 35, 59, 52, 50, 38, 42, 39, 40, 50, 63, 73, 76, 55, 
    40, 33, 38, 61, 54, 56, 48, 33, 32, 31, 43, 17, 48, 53, 60, 
    44, 37, 54, 54, 59, 69, 62, 43, 28, 38, 37, 29, 25, 37, 44, 
    54, 44, 53, 58, 59, 48, 55, 62, 49, 43, 20, 31, 40, 29, 28, 
    55, 41, 54, 67, 68, 49, 55, 54, 54, 22, 28, 35, 43, 32, 18, 
    51, 38, 47, 63, 57, 34, 61, 51, 44, 21, 29, 27, 37, 25, 24, 
    47, 32, 36, 62, 45, 37, 48, 37, 28, 9, 23, 22, 16, 19, 28, 
    35, 27, 26, 61, 54, 49, 29, 26, 14, 8, 16, 22, 12, 22, 26, 
    
    -- channel=537
    5, 0, 10, 8, 2, 5, 12, 17, 43, 2, 7, 24, 17, 14, 11, 
    4, 0, 0, 0, 30, 1, 0, 15, 1, 12, 40, 19, 12, 8, 7, 
    4, 0, 8, 4, 12, 4, 0, 0, 0, 19, 25, 0, 8, 19, 24, 
    75, 71, 63, 0, 0, 21, 42, 16, 4, 0, 4, 17, 17, 0, 0, 
    44, 51, 14, 0, 2, 0, 0, 0, 0, 0, 2, 19, 3, 0, 0, 
    9, 3, 0, 9, 13, 0, 0, 0, 24, 9, 0, 4, 5, 13, 3, 
    3, 0, 0, 15, 0, 0, 0, 10, 17, 10, 0, 8, 1, 26, 24, 
    0, 0, 0, 18, 10, 3, 2, 0, 0, 0, 0, 0, 0, 0, 4, 
    6, 0, 24, 8, 18, 41, 19, 9, 0, 0, 11, 5, 0, 0, 0, 
    18, 16, 10, 9, 0, 0, 0, 27, 26, 10, 0, 1, 20, 6, 0, 
    8, 0, 5, 9, 14, 0, 0, 0, 2, 0, 0, 14, 6, 0, 0, 
    0, 5, 3, 1, 0, 0, 15, 3, 0, 0, 10, 0, 5, 1, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 4, 10, 33, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 3, 0, 
    
    -- channel=538
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 20, 6, 0, 0, 0, 
    0, 0, 0, 0, 19, 4, 0, 0, 0, 0, 25, 0, 4, 10, 9, 
    38, 39, 45, 0, 2, 22, 24, 2, 0, 0, 6, 16, 26, 3, 0, 
    11, 19, 6, 0, 10, 8, 4, 0, 0, 0, 8, 17, 15, 0, 0, 
    0, 0, 0, 0, 10, 2, 0, 0, 13, 7, 3, 10, 12, 0, 0, 
    0, 0, 0, 0, 2, 7, 6, 1, 17, 8, 9, 14, 10, 19, 7, 
    0, 0, 0, 7, 12, 3, 8, 2, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 11, 15, 17, 41, 29, 12, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 9, 4, 2, 0, 4, 28, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 14, 13, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 12, 5, 0, 8, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 11, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=539
    1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 7, 0, 0, 2, 14, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 11, 26, 6, 0, 1, 5, 5, 14, 14, 10, 9, 
    11, 0, 0, 6, 8, 26, 15, 9, 2, 0, 16, 12, 23, 22, 16, 
    15, 3, 14, 17, 3, 21, 18, 16, 3, 5, 13, 13, 24, 27, 10, 
    14, 13, 14, 12, 7, 19, 21, 15, 7, 8, 13, 12, 27, 26, 12, 
    14, 12, 11, 0, 17, 18, 19, 9, 19, 14, 15, 12, 26, 27, 25, 
    16, 8, 5, 0, 20, 19, 23, 10, 9, 15, 13, 5, 13, 24, 21, 
    20, 11, 5, 2, 22, 23, 25, 24, 0, 9, 3, 2, 0, 11, 6, 
    23, 15, 13, 13, 20, 21, 23, 29, 11, 0, 8, 0, 0, 0, 0, 
    22, 21, 15, 18, 17, 24, 10, 17, 20, 7, 2, 0, 1, 7, 0, 
    21, 22, 11, 21, 18, 17, 7, 13, 13, 13, 0, 4, 1, 5, 4, 
    20, 19, 12, 23, 18, 4, 0, 8, 10, 3, 0, 3, 2, 3, 1, 
    19, 15, 9, 20, 25, 0, 6, 1, 1, 2, 0, 0, 2, 0, 0, 
    16, 10, 9, 17, 23, 13, 5, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=540
    24, 0, 0, 0, 2, 0, 0, 0, 10, 34, 0, 0, 0, 0, 0, 
    24, 8, 0, 0, 2, 10, 0, 0, 0, 30, 0, 2, 0, 0, 0, 
    23, 19, 0, 0, 0, 24, 4, 0, 0, 1, 0, 0, 0, 0, 3, 
    63, 29, 0, 13, 0, 7, 26, 17, 2, 0, 0, 0, 0, 6, 0, 
    22, 13, 10, 28, 0, 0, 2, 17, 0, 0, 0, 0, 4, 28, 7, 
    10, 7, 8, 22, 0, 0, 8, 14, 6, 0, 0, 0, 7, 31, 22, 
    14, 8, 9, 0, 9, 1, 9, 0, 8, 1, 1, 0, 3, 14, 32, 
    18, 1, 13, 0, 5, 4, 1, 11, 0, 5, 5, 0, 0, 4, 13, 
    28, 6, 0, 0, 0, 4, 13, 14, 0, 13, 0, 29, 0, 0, 0, 
    22, 16, 0, 0, 0, 0, 0, 13, 29, 0, 3, 0, 7, 3, 0, 
    12, 22, 0, 3, 1, 15, 0, 0, 1, 6, 3, 0, 0, 6, 1, 
    11, 23, 0, 0, 0, 0, 0, 0, 2, 18, 0, 0, 0, 8, 12, 
    16, 21, 0, 0, 3, 0, 0, 0, 1, 11, 0, 3, 0, 0, 6, 
    18, 26, 6, 0, 7, 4, 0, 0, 4, 11, 0, 5, 10, 0, 0, 
    17, 22, 13, 0, 6, 4, 6, 0, 11, 5, 4, 2, 12, 2, 0, 
    
    -- channel=541
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    14, 3, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=542
    0, 11, 0, 2, 0, 5, 5, 2, 0, 0, 2, 0, 0, 2, 5, 
    0, 10, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 4, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 2, 4, 0, 0, 0, 0, 0, 
    
    -- channel=543
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=544
    1, 0, 38, 0, 0, 0, 0, 0, 21, 0, 0, 17, 0, 0, 0, 
    0, 0, 67, 0, 16, 0, 0, 0, 2, 0, 16, 0, 0, 0, 0, 
    0, 0, 56, 0, 22, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 
    24, 1, 55, 0, 18, 5, 0, 5, 8, 0, 24, 0, 0, 0, 0, 
    5, 0, 5, 0, 22, 0, 0, 0, 4, 0, 2, 19, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 33, 0, 0, 23, 0, 0, 0, 
    0, 0, 0, 41, 0, 0, 10, 0, 14, 2, 0, 20, 0, 4, 0, 
    0, 0, 0, 54, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 19, 0, 0, 21, 0, 21, 0, 0, 43, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 15, 0, 7, 0, 7, 0, 
    0, 0, 6, 0, 0, 0, 3, 0, 0, 0, 0, 4, 5, 0, 0, 
    0, 2, 0, 0, 0, 0, 7, 0, 0, 0, 3, 0, 18, 0, 0, 
    0, 0, 0, 0, 16, 0, 29, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 5, 
    0, 8, 0, 18, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    
    -- channel=545
    0, 0, 38, 21, 21, 22, 25, 24, 23, 0, 0, 49, 40, 39, 38, 
    0, 0, 41, 8, 39, 23, 34, 40, 47, 15, 9, 56, 49, 45, 44, 
    0, 0, 17, 3, 51, 40, 12, 25, 29, 9, 50, 57, 59, 58, 55, 
    0, 0, 41, 28, 47, 55, 18, 16, 9, 10, 70, 56, 75, 81, 63, 
    49, 32, 60, 24, 33, 53, 54, 25, 11, 9, 60, 72, 83, 69, 50, 
    59, 52, 66, 21, 45, 51, 45, 7, 23, 12, 45, 77, 88, 73, 52, 
    59, 48, 47, 44, 33, 26, 44, 14, 48, 33, 39, 77, 87, 87, 54, 
    59, 44, 29, 55, 54, 46, 43, 25, 46, 30, 51, 61, 76, 94, 63, 
    63, 30, 41, 43, 59, 63, 41, 51, 17, 16, 57, 6, 31, 62, 60, 
    70, 37, 54, 56, 55, 66, 62, 50, 18, 31, 45, 27, 10, 40, 29, 
    70, 51, 55, 56, 60, 54, 49, 50, 62, 49, 13, 28, 35, 28, 25, 
    68, 63, 49, 66, 70, 48, 50, 49, 55, 28, 18, 30, 43, 29, 17, 
    66, 63, 46, 64, 67, 0, 60, 47, 46, 19, 23, 21, 34, 23, 21, 
    64, 55, 31, 67, 58, 15, 51, 32, 25, 1, 21, 14, 14, 9, 26, 
    48, 52, 17, 64, 57, 53, 30, 22, 14, 0, 12, 19, 9, 15, 22, 
    
    -- channel=546
    2, 0, 0, 0, 0, 0, 2, 9, 31, 0, 28, 8, 7, 3, 2, 
    1, 0, 0, 4, 21, 0, 0, 0, 0, 7, 30, 7, 8, 5, 1, 
    1, 0, 15, 12, 8, 0, 0, 0, 0, 27, 7, 1, 4, 9, 9, 
    73, 100, 24, 0, 0, 15, 26, 9, 12, 0, 0, 12, 0, 0, 0, 
    21, 10, 0, 0, 7, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 13, 16, 10, 0, 1, 0, 5, 0, 
    0, 0, 0, 13, 9, 25, 0, 4, 0, 1, 4, 0, 0, 11, 11, 
    0, 0, 0, 11, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 2, 27, 0, 10, 21, 15, 6, 0, 0, 0, 9, 0, 0, 0, 
    6, 2, 0, 0, 0, 0, 0, 20, 20, 13, 0, 3, 19, 0, 0, 
    0, 0, 5, 5, 4, 0, 0, 0, 0, 0, 5, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 4, 14, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 7, 0, 0, 
    
    -- channel=547
    0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 5, 0, 0, 5, 8, 2, 6, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 0, 4, 4, 14, 27, 22, 0, 11, 19, 9, 3, 0, 
    0, 0, 0, 16, 15, 0, 0, 0, 0, 8, 19, 12, 10, 30, 25, 
    0, 2, 15, 5, 10, 13, 9, 6, 4, 9, 15, 19, 21, 26, 36, 
    18, 21, 24, 3, 10, 19, 11, 0, 0, 3, 18, 26, 27, 23, 31, 
    23, 18, 25, 2, 6, 4, 7, 0, 3, 9, 14, 23, 30, 16, 15, 
    30, 22, 0, 0, 11, 15, 4, 14, 9, 19, 26, 60, 36, 39, 29, 
    26, 18, 0, 2, 5, 0, 0, 0, 14, 8, 6, 0, 41, 45, 40, 
    20, 15, 9, 9, 23, 35, 17, 0, 0, 2, 11, 0, 0, 4, 28, 
    26, 28, 14, 7, 10, 14, 20, 22, 7, 16, 0, 0, 3, 2, 10, 
    32, 25, 20, 15, 18, 7, 5, 8, 14, 0, 2, 8, 5, 4, 0, 
    32, 32, 28, 18, 18, 1, 13, 17, 15, 7, 8, 8, 19, 6, 0, 
    32, 33, 32, 19, 0, 0, 11, 13, 12, 4, 5, 5, 4, 3, 1, 
    36, 26, 36, 24, 14, 16, 18, 8, 6, 3, 4, 3, 0, 4, 7, 
    
    -- channel=548
    7, 41, 36, 0, 2, 13, 6, 9, 0, 0, 35, 17, 5, 5, 2, 
    7, 19, 67, 0, 0, 0, 7, 9, 0, 0, 52, 0, 0, 0, 0, 
    7, 10, 82, 0, 12, 0, 0, 15, 0, 0, 30, 2, 0, 0, 0, 
    0, 20, 56, 0, 23, 0, 0, 0, 9, 18, 6, 11, 0, 0, 0, 
    0, 10, 0, 0, 29, 0, 0, 0, 6, 6, 13, 18, 0, 0, 6, 
    0, 0, 0, 0, 13, 0, 0, 0, 7, 2, 3, 28, 0, 0, 1, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 3, 0, 25, 0, 0, 0, 
    0, 0, 0, 54, 0, 0, 0, 0, 10, 0, 0, 12, 12, 0, 0, 
    0, 0, 0, 11, 0, 0, 0, 0, 12, 0, 14, 0, 33, 1, 22, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 9, 0, 3, 10, 
    0, 0, 9, 0, 0, 0, 11, 0, 0, 0, 0, 9, 2, 0, 0, 
    0, 0, 15, 0, 0, 0, 3, 0, 0, 0, 20, 0, 9, 0, 0, 
    0, 0, 9, 0, 0, 0, 19, 0, 0, 0, 17, 0, 1, 0, 0, 
    0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 13, 6, 
    0, 4, 0, 13, 0, 0, 0, 4, 0, 9, 4, 6, 0, 9, 5, 
    
    -- channel=549
    0, 0, 0, 0, 0, 0, 0, 0, 16, 16, 0, 21, 7, 4, 0, 
    0, 0, 0, 0, 13, 6, 0, 0, 0, 0, 57, 5, 0, 0, 0, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 36, 0, 0, 1, 8, 
    99, 86, 101, 0, 0, 0, 42, 14, 0, 6, 0, 3, 9, 0, 0, 
    24, 65, 3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 17, 10, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 4, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 0, 31, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 4, 37, 2, 0, 0, 14, 2, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    
    -- channel=550
    0, 53, 5, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    1, 35, 37, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 
    1, 14, 42, 0, 0, 0, 6, 25, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 1, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 62, 17, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 4, 0, 0, 4, 0, 0, 0, 0, 5, 0, 8, 0, 0, 
    0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 5, 0, 
    0, 0, 16, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 1, 
    
    -- channel=551
    5, 91, 24, 0, 0, 6, 0, 0, 0, 0, 64, 0, 0, 0, 0, 
    6, 56, 58, 8, 0, 0, 5, 0, 0, 0, 62, 0, 0, 0, 0, 
    5, 23, 84, 1, 13, 0, 0, 25, 3, 0, 8, 0, 0, 0, 0, 
    0, 5, 19, 0, 37, 0, 0, 0, 0, 39, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 34, 0, 0, 0, 4, 25, 7, 1, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 11, 4, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 12, 0, 0, 0, 
    0, 0, 0, 47, 0, 0, 0, 0, 8, 0, 0, 36, 17, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 29, 0, 0, 0, 46, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 15, 
    0, 0, 2, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 12, 9, 0, 0, 0, 14, 0, 1, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 17, 0, 
    0, 0, 0, 10, 0, 0, 0, 4, 0, 14, 1, 0, 0, 2, 3, 
    
    -- channel=552
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 19, 15, 40, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 31, 0, 0, 2, 29, 0, 0, 0, 0, 0, 24, 0, 
    0, 0, 1, 0, 0, 0, 26, 5, 0, 0, 0, 0, 0, 12, 0, 
    0, 0, 34, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 30, 0, 0, 0, 0, 0, 0, 0, 3, 20, 0, 12, 0, 
    17, 0, 0, 0, 0, 0, 0, 18, 0, 2, 0, 2, 0, 46, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 24, 0, 0, 0, 2, 
    0, 5, 0, 0, 0, 17, 0, 0, 7, 22, 0, 0, 0, 12, 0, 
    0, 16, 0, 0, 0, 13, 0, 0, 0, 35, 0, 0, 0, 0, 3, 
    0, 14, 0, 0, 39, 12, 0, 6, 27, 19, 0, 1, 12, 10, 0, 
    6, 16, 0, 0, 6, 0, 12, 15, 23, 12, 0, 0, 11, 0, 0, 
    23, 7, 0, 0, 0, 8, 35, 10, 29, 0, 0, 0, 0, 0, 0, 
    
    -- channel=553
    0, 2, 9, 2, 0, 13, 7, 8, 0, 0, 8, 0, 3, 4, 4, 
    0, 0, 15, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=554
    4, 89, 0, 0, 0, 1, 0, 0, 0, 0, 51, 0, 0, 0, 0, 
    5, 58, 28, 26, 0, 0, 6, 0, 0, 0, 11, 0, 0, 0, 0, 
    5, 23, 44, 2, 2, 0, 22, 48, 32, 3, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 36, 0, 0, 0, 0, 36, 0, 1, 0, 0, 16, 
    0, 0, 0, 0, 22, 1, 0, 0, 4, 32, 11, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 3, 10, 14, 0, 0, 0, 
    0, 0, 2, 0, 0, 8, 0, 14, 0, 0, 6, 5, 0, 0, 0, 
    0, 5, 0, 21, 0, 0, 0, 0, 15, 17, 0, 98, 37, 0, 0, 
    0, 10, 0, 3, 0, 0, 0, 0, 47, 1, 0, 0, 86, 48, 49, 
    0, 0, 0, 0, 9, 22, 2, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 6, 0, 0, 0, 23, 16, 0, 0, 16, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 1, 0, 0, 0, 0, 4, 2, 0, 0, 0, 
    0, 0, 21, 0, 0, 60, 6, 9, 2, 0, 11, 8, 19, 17, 0, 
    0, 0, 32, 0, 0, 0, 0, 10, 7, 20, 5, 2, 0, 18, 0, 
    13, 0, 33, 13, 0, 0, 10, 15, 0, 12, 9, 0, 0, 0, 13, 
    
    -- channel=555
    4, 0, 0, 0, 0, 0, 0, 0, 36, 48, 0, 8, 7, 4, 3, 
    3, 0, 0, 0, 16, 8, 0, 0, 0, 30, 0, 6, 5, 0, 0, 
    4, 0, 0, 4, 0, 29, 0, 0, 0, 0, 8, 0, 0, 2, 10, 
    128, 67, 37, 0, 0, 14, 58, 28, 0, 0, 0, 0, 3, 0, 0, 
    32, 32, 3, 15, 0, 0, 0, 6, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 16, 0, 0, 0, 1, 18, 0, 0, 0, 0, 20, 0, 
    0, 0, 0, 0, 6, 0, 9, 0, 12, 0, 0, 0, 0, 10, 25, 
    0, 0, 17, 0, 6, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 7, 0, 0, 27, 31, 20, 0, 0, 0, 29, 0, 0, 0, 
    8, 8, 0, 0, 0, 0, 0, 21, 59, 0, 0, 0, 14, 1, 0, 
    0, 6, 0, 3, 2, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    
    -- channel=556
    0, 86, 11, 1, 0, 8, 4, 17, 4, 0, 73, 26, 12, 11, 4, 
    1, 48, 22, 20, 15, 0, 0, 13, 0, 0, 119, 10, 5, 5, 0, 
    1, 15, 70, 36, 30, 0, 0, 0, 0, 14, 59, 6, 1, 10, 10, 
    32, 104, 108, 0, 33, 0, 6, 0, 13, 60, 0, 44, 6, 0, 3, 
    0, 64, 3, 0, 56, 0, 0, 0, 7, 38, 15, 45, 0, 0, 14, 
    0, 8, 0, 0, 35, 0, 0, 0, 19, 40, 16, 39, 0, 0, 1, 
    0, 1, 0, 5, 3, 12, 0, 25, 0, 24, 19, 39, 0, 0, 0, 
    0, 0, 0, 60, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 8, 0, 50, 0, 24, 9, 0, 36, 0, 0, 0, 22, 0, 19, 
    0, 17, 11, 0, 5, 0, 0, 0, 3, 20, 0, 0, 25, 0, 5, 
    0, 0, 19, 7, 7, 0, 15, 0, 0, 0, 0, 22, 8, 0, 0, 
    0, 0, 42, 0, 0, 0, 19, 3, 0, 0, 37, 0, 3, 0, 0, 
    0, 0, 32, 0, 0, 0, 2, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 31, 6, 0, 30, 0, 0, 0, 0, 11, 0, 0, 20, 4, 
    0, 0, 20, 11, 0, 0, 0, 0, 0, 14, 1, 0, 0, 14, 0, 
    
    -- channel=557
    1, 0, 0, 3, 2, 0, 8, 0, 28, 34, 0, 14, 14, 12, 12, 
    1, 0, 0, 0, 12, 11, 0, 8, 6, 26, 5, 11, 8, 7, 7, 
    3, 0, 0, 4, 0, 31, 0, 0, 0, 0, 6, 0, 0, 5, 13, 
    81, 26, 31, 12, 0, 13, 51, 22, 0, 0, 0, 0, 15, 7, 0, 
    29, 46, 6, 17, 0, 0, 5, 14, 0, 0, 0, 0, 0, 4, 0, 
    3, 0, 0, 20, 0, 0, 0, 0, 13, 3, 0, 0, 0, 18, 0, 
    0, 0, 0, 0, 0, 0, 4, 1, 11, 1, 0, 0, 0, 11, 24, 
    0, 0, 28, 0, 13, 10, 0, 30, 0, 0, 0, 0, 0, 0, 0, 
    11, 0, 7, 0, 4, 27, 26, 12, 0, 8, 0, 33, 0, 0, 0, 
    6, 15, 3, 5, 0, 0, 0, 18, 54, 0, 0, 0, 17, 7, 0, 
    0, 11, 0, 7, 7, 12, 0, 0, 0, 7, 0, 3, 5, 0, 0, 
    0, 8, 0, 0, 3, 0, 8, 3, 3, 4, 0, 0, 0, 10, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 9, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 7, 3, 0, 
    
    -- channel=558
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=559
    0, 0, 4, 0, 0, 0, 2, 9, 29, 0, 20, 21, 12, 9, 4, 
    0, 0, 0, 0, 25, 0, 0, 5, 0, 0, 58, 12, 3, 2, 0, 
    0, 0, 8, 0, 4, 0, 0, 0, 0, 11, 24, 0, 0, 12, 15, 
    85, 100, 77, 0, 0, 10, 43, 5, 0, 2, 0, 15, 8, 0, 0, 
    37, 53, 6, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 3, 2, 0, 0, 0, 20, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 5, 3, 0, 0, 1, 0, 14, 19, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 1, 7, 33, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 12, 0, 0, 0, 0, 0, 18, 31, 10, 0, 0, 21, 0, 0, 
    0, 0, 0, 2, 8, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=560
    16, 19, 50, 38, 33, 43, 46, 42, 42, 25, 27, 48, 52, 51, 52, 
    16, 10, 50, 32, 22, 22, 27, 32, 34, 30, 29, 33, 40, 43, 46, 
    18, 13, 47, 36, 19, 14, 21, 23, 21, 23, 25, 19, 23, 26, 29, 
    42, 40, 39, 22, 16, 20, 24, 30, 29, 18, 18, 19, 17, 14, 15, 
    28, 22, 23, 24, 23, 15, 19, 18, 21, 15, 20, 21, 19, 19, 16, 
    22, 18, 21, 21, 22, 11, 17, 19, 24, 15, 14, 19, 12, 17, 20, 
    22, 21, 25, 30, 22, 18, 20, 15, 21, 16, 15, 20, 13, 15, 14, 
    17, 18, 33, 41, 16, 11, 17, 13, 22, 16, 12, 11, 8, 14, 9, 
    18, 21, 41, 29, 15, 21, 15, 27, 26, 18, 34, 27, 25, 15, 13, 
    19, 16, 22, 22, 16, 10, 9, 18, 24, 31, 30, 37, 30, 33, 21, 
    14, 11, 18, 20, 19, 19, 21, 13, 21, 29, 27, 33, 29, 30, 28, 
    13, 17, 16, 14, 17, 22, 25, 23, 23, 28, 31, 26, 29, 27, 29, 
    14, 18, 14, 14, 25, 24, 32, 24, 26, 26, 29, 25, 25, 26, 31, 
    14, 17, 12, 14, 25, 31, 31, 28, 28, 25, 32, 27, 28, 29, 31, 
    11, 21, 10, 11, 15, 23, 23, 30, 30, 26, 28, 30, 30, 30, 27, 
    
    -- channel=561
    0, 113, 24, 0, 0, 9, 0, 5, 0, 0, 87, 14, 0, 0, 0, 
    0, 62, 58, 16, 0, 0, 9, 11, 0, 0, 103, 0, 0, 0, 0, 
    0, 19, 102, 15, 30, 0, 0, 17, 0, 9, 41, 11, 0, 0, 0, 
    0, 53, 68, 0, 51, 0, 0, 0, 7, 63, 1, 41, 0, 0, 17, 
    0, 27, 0, 0, 57, 1, 0, 0, 8, 43, 30, 37, 0, 0, 23, 
    0, 7, 0, 0, 30, 0, 0, 0, 1, 31, 23, 47, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 0, 22, 0, 17, 22, 47, 0, 0, 0, 
    0, 3, 0, 67, 0, 0, 0, 0, 14, 14, 0, 46, 33, 0, 0, 
    0, 8, 0, 40, 0, 0, 0, 0, 51, 0, 0, 0, 60, 0, 49, 
    0, 0, 7, 0, 10, 0, 0, 0, 0, 11, 0, 1, 6, 0, 22, 
    0, 0, 25, 0, 0, 0, 27, 4, 0, 0, 2, 13, 2, 0, 0, 
    0, 0, 44, 0, 0, 0, 12, 0, 0, 0, 31, 0, 6, 0, 0, 
    0, 0, 36, 0, 0, 13, 13, 0, 0, 0, 21, 0, 0, 0, 0, 
    0, 0, 35, 8, 0, 0, 0, 0, 0, 0, 13, 0, 0, 25, 2, 
    0, 0, 22, 28, 0, 0, 0, 0, 0, 15, 6, 1, 0, 10, 7, 
    
    -- channel=562
    12, 29, 63, 54, 46, 63, 61, 58, 50, 23, 40, 54, 65, 66, 67, 
    13, 19, 57, 49, 26, 31, 48, 49, 45, 39, 33, 47, 54, 59, 63, 
    15, 15, 48, 44, 24, 20, 27, 36, 40, 40, 22, 37, 40, 42, 45, 
    15, 26, 32, 39, 25, 27, 25, 25, 28, 27, 28, 38, 32, 31, 39, 
    45, 35, 36, 40, 22, 23, 28, 26, 26, 24, 31, 36, 34, 38, 40, 
    42, 36, 40, 42, 28, 23, 23, 26, 21, 21, 24, 36, 34, 41, 43, 
    43, 42, 43, 45, 21, 21, 21, 31, 19, 22, 23, 34, 35, 39, 38, 
    41, 44, 47, 43, 27, 21, 25, 16, 36, 28, 27, 42, 45, 34, 41, 
    39, 39, 47, 27, 31, 24, 16, 23, 34, 37, 40, 37, 32, 41, 46, 
    41, 37, 33, 33, 24, 23, 28, 25, 25, 40, 37, 48, 42, 40, 35, 
    39, 32, 34, 30, 33, 26, 29, 27, 36, 34, 44, 40, 37, 38, 40, 
    36, 38, 31, 30, 29, 42, 34, 34, 33, 40, 41, 37, 38, 38, 38, 
    37, 42, 36, 26, 29, 37, 39, 39, 39, 41, 39, 38, 34, 41, 38, 
    39, 43, 40, 28, 37, 41, 37, 42, 41, 40, 38, 37, 36, 37, 41, 
    40, 45, 38, 25, 30, 32, 43, 45, 39, 39, 37, 38, 38, 37, 38, 
    
    -- channel=563
    0, 31, 77, 70, 65, 74, 73, 77, 65, 24, 57, 86, 86, 86, 84, 
    0, 11, 72, 68, 72, 63, 74, 80, 78, 43, 75, 94, 92, 91, 89, 
    0, 0, 65, 64, 85, 58, 49, 63, 61, 62, 83, 96, 96, 97, 95, 
    13, 31, 81, 65, 82, 78, 55, 46, 48, 67, 87, 103, 104, 97, 102, 
    79, 78, 88, 60, 75, 83, 75, 49, 49, 62, 90, 109, 110, 90, 93, 
    91, 89, 91, 67, 80, 79, 64, 49, 53, 61, 81, 114, 114, 95, 88, 
    93, 88, 74, 80, 66, 71, 64, 64, 66, 69, 79, 110, 117, 111, 93, 
    91, 86, 60, 95, 81, 73, 72, 53, 75, 72, 73, 95, 111, 109, 104, 
    86, 77, 79, 84, 91, 90, 74, 61, 68, 62, 76, 49, 77, 86, 104, 
    96, 83, 87, 87, 88, 90, 90, 80, 57, 73, 66, 67, 62, 70, 71, 
    101, 81, 92, 90, 93, 73, 84, 85, 84, 65, 62, 69, 71, 63, 61, 
    99, 85, 93, 96, 91, 81, 84, 84, 80, 58, 66, 67, 75, 64, 54, 
    95, 88, 91, 92, 76, 57, 88, 80, 72, 55, 64, 61, 63, 62, 58, 
    92, 82, 86, 94, 82, 69, 74, 68, 59, 49, 59, 55, 49, 56, 65, 
    81, 80, 75, 91, 86, 77, 61, 59, 46, 46, 53, 57, 50, 56, 60, 
    
    -- channel=564
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 55, 0, 0, 0, 0, 1, 0, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=565
    0, 0, 0, 0, 0, 0, 0, 0, 8, 52, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 108, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 75, 3, 0, 23, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 23, 0, 24, 1, 11, 0, 0, 0, 0, 0, 14, 0, 
    17, 0, 0, 75, 0, 0, 18, 63, 0, 0, 0, 0, 0, 63, 0, 
    0, 0, 2, 25, 0, 0, 46, 23, 0, 0, 0, 0, 0, 55, 0, 
    0, 0, 45, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 5, 7, 
    14, 0, 74, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 11, 0, 
    48, 0, 0, 0, 0, 0, 0, 60, 0, 11, 0, 23, 0, 28, 0, 
    22, 0, 0, 0, 0, 0, 0, 8, 0, 0, 29, 0, 0, 0, 0, 
    0, 22, 0, 0, 0, 41, 0, 0, 28, 30, 0, 0, 0, 21, 0, 
    0, 47, 0, 0, 0, 28, 0, 0, 3, 76, 0, 0, 0, 9, 16, 
    0, 31, 0, 0, 62, 0, 0, 0, 34, 35, 0, 0, 0, 3, 0, 
    14, 34, 0, 0, 39, 0, 5, 6, 27, 14, 0, 0, 21, 0, 0, 
    26, 17, 0, 0, 5, 15, 49, 0, 42, 0, 0, 0, 1, 0, 0, 
    
    -- channel=566
    4, 20, 51, 49, 38, 52, 52, 52, 42, 17, 29, 44, 54, 55, 56, 
    5, 10, 48, 43, 21, 25, 38, 39, 36, 25, 28, 38, 45, 49, 52, 
    6, 7, 41, 38, 20, 10, 20, 31, 33, 30, 22, 32, 35, 36, 38, 
    8, 18, 28, 31, 23, 16, 15, 19, 21, 21, 22, 30, 23, 22, 31, 
    33, 27, 29, 28, 22, 16, 18, 17, 18, 18, 25, 31, 26, 28, 33, 
    32, 29, 31, 30, 24, 15, 16, 17, 15, 15, 19, 33, 27, 31, 35, 
    35, 34, 33, 37, 19, 16, 15, 19, 14, 15, 17, 30, 29, 31, 31, 
    33, 34, 33, 42, 20, 14, 16, 8, 25, 20, 20, 34, 38, 28, 30, 
    30, 31, 36, 27, 21, 18, 10, 14, 27, 26, 30, 26, 33, 34, 38, 
    33, 29, 27, 25, 20, 18, 18, 17, 15, 30, 29, 38, 32, 32, 31, 
    31, 23, 28, 24, 25, 19, 22, 20, 24, 26, 34, 33, 29, 29, 30, 
    29, 28, 28, 23, 22, 28, 27, 26, 24, 29, 33, 29, 30, 28, 29, 
    29, 33, 31, 20, 19, 28, 32, 30, 30, 29, 32, 29, 27, 31, 29, 
    30, 34, 35, 23, 25, 27, 31, 33, 31, 30, 31, 28, 26, 30, 31, 
    31, 35, 31, 21, 21, 25, 30, 35, 29, 29, 29, 30, 29, 28, 30, 
    
    -- channel=567
    5, 30, 0, 0, 4, 2, 5, 0, 0, 17, 1, 1, 1, 5, 6, 
    5, 25, 6, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    6, 14, 13, 6, 0, 0, 17, 9, 0, 0, 0, 0, 0, 0, 0, 
    21, 6, 0, 3, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    3, 3, 20, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 9, 0, 0, 0, 
    3, 11, 0, 0, 0, 0, 0, 0, 17, 0, 0, 19, 40, 6, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 7, 0, 0, 0, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 
    1, 4, 0, 0, 0, 20, 0, 0, 0, 0, 1, 0, 4, 0, 2, 
    3, 11, 11, 0, 0, 0, 2, 5, 4, 10, 5, 3, 4, 7, 0, 
    9, 5, 20, 0, 0, 0, 1, 0, 7, 4, 7, 0, 0, 2, 4, 
    
    -- channel=568
    1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    1, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 18, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 1, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 7, 0, 0, 2, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=569
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 9, 1, 0, 0, 0, 0, 22, 2, 0, 0, 0, 
    0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 25, 1, 4, 5, 2, 
    0, 0, 28, 0, 17, 4, 5, 0, 0, 12, 9, 12, 18, 9, 0, 
    0, 14, 2, 0, 20, 11, 5, 0, 0, 6, 6, 18, 10, 0, 0, 
    0, 0, 0, 0, 16, 11, 0, 0, 8, 11, 10, 14, 7, 0, 0, 
    0, 0, 0, 0, 5, 3, 4, 3, 8, 9, 9, 17, 7, 2, 0, 
    0, 0, 0, 15, 9, 11, 0, 17, 0, 2, 3, 0, 0, 5, 0, 
    0, 0, 0, 23, 7, 20, 17, 0, 1, 0, 2, 0, 0, 0, 0, 
    0, 0, 10, 8, 10, 11, 7, 4, 9, 4, 0, 0, 0, 0, 0, 
    0, 0, 6, 11, 10, 1, 9, 9, 0, 0, 0, 1, 4, 0, 0, 
    0, 0, 12, 13, 13, 0, 12, 7, 5, 0, 1, 0, 3, 0, 0, 
    0, 0, 1, 12, 4, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=570
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    34, 46, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=571
    2, 0, 0, 0, 0, 0, 0, 0, 32, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 0, 0, 0, 71, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 44, 0, 0, 3, 5, 0, 0, 0, 0, 0, 
    31, 0, 0, 0, 0, 34, 18, 13, 0, 0, 0, 0, 0, 1, 0, 
    32, 0, 0, 35, 0, 0, 13, 33, 0, 0, 0, 0, 0, 26, 0, 
    0, 0, 1, 13, 0, 0, 24, 12, 0, 0, 0, 0, 0, 35, 0, 
    0, 0, 3, 3, 0, 0, 15, 0, 5, 0, 0, 0, 0, 18, 4, 
    0, 0, 44, 0, 0, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 
    25, 0, 20, 0, 6, 0, 0, 48, 0, 0, 6, 14, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 1, 23, 4, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 18, 0, 0, 26, 7, 2, 0, 0, 11, 0, 
    0, 28, 0, 0, 0, 15, 0, 0, 0, 41, 0, 0, 0, 4, 14, 
    0, 11, 0, 0, 29, 0, 0, 0, 12, 15, 0, 0, 0, 4, 0, 
    1, 12, 0, 0, 33, 0, 0, 0, 6, 0, 0, 0, 8, 0, 0, 
    0, 14, 0, 0, 4, 3, 13, 0, 19, 0, 0, 0, 7, 0, 0, 
    
    -- channel=572
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=573
    0, 0, 0, 0, 0, 0, 0, 0, 17, 50, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 66, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 57, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    48, 0, 0, 19, 0, 19, 26, 21, 0, 0, 0, 0, 0, 12, 0, 
    17, 0, 0, 50, 0, 0, 13, 42, 0, 0, 0, 0, 0, 38, 0, 
    0, 0, 0, 20, 0, 0, 28, 14, 0, 0, 0, 0, 0, 36, 0, 
    0, 0, 25, 0, 0, 0, 21, 0, 6, 0, 0, 0, 0, 5, 18, 
    8, 0, 52, 0, 6, 0, 2, 5, 0, 0, 0, 0, 0, 2, 0, 
    29, 0, 0, 0, 0, 0, 8, 43, 0, 9, 0, 28, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 15, 30, 0, 19, 0, 0, 0, 0, 
    0, 18, 0, 0, 0, 31, 0, 0, 14, 24, 0, 0, 0, 14, 0, 
    0, 25, 0, 0, 1, 14, 0, 0, 6, 45, 0, 0, 0, 10, 13, 
    0, 12, 0, 0, 37, 0, 0, 0, 15, 20, 0, 0, 0, 0, 1, 
    6, 15, 0, 0, 28, 0, 6, 0, 11, 5, 0, 0, 12, 0, 0, 
    5, 2, 0, 0, 6, 13, 24, 0, 23, 0, 0, 0, 5, 0, 0, 
    
    -- channel=574
    4, 0, 0, 0, 3, 0, 5, 0, 44, 49, 0, 2, 9, 5, 9, 
    2, 0, 0, 0, 12, 3, 0, 0, 2, 64, 0, 9, 8, 3, 5, 
    2, 0, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 3, 11, 
    106, 13, 0, 9, 0, 32, 58, 29, 0, 0, 0, 0, 3, 5, 0, 
    42, 6, 4, 37, 0, 0, 14, 30, 0, 0, 0, 0, 1, 28, 0, 
    3, 0, 0, 29, 0, 0, 18, 10, 12, 0, 0, 0, 0, 44, 0, 
    1, 0, 0, 2, 4, 0, 21, 0, 15, 0, 0, 0, 0, 22, 24, 
    3, 0, 52, 0, 10, 2, 0, 20, 0, 0, 0, 0, 0, 0, 0, 
    32, 0, 20, 0, 6, 22, 25, 46, 0, 8, 3, 41, 0, 0, 0, 
    21, 2, 0, 1, 0, 0, 0, 29, 59, 0, 0, 0, 6, 2, 0, 
    0, 17, 0, 2, 1, 25, 0, 0, 13, 11, 0, 0, 0, 6, 0, 
    0, 29, 0, 0, 1, 0, 0, 0, 5, 29, 0, 0, 0, 13, 16, 
    0, 6, 0, 0, 25, 0, 0, 0, 0, 9, 0, 0, 0, 0, 6, 
    0, 11, 0, 0, 30, 26, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 9, 0, 0, 7, 9, 0, 0, 10, 0, 0, 0, 12, 0, 0, 
    
    -- channel=575
    4, 0, 2, 17, 6, 11, 10, 1, 0, 16, 0, 0, 6, 6, 13, 
    4, 0, 0, 16, 0, 0, 3, 0, 5, 32, 0, 0, 0, 4, 11, 
    6, 3, 0, 3, 0, 10, 19, 19, 32, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 22, 0, 0, 1, 21, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 14, 13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 4, 0, 15, 0, 11, 3, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 10, 0, 0, 6, 
    0, 0, 0, 0, 0, 4, 0, 0, 3, 13, 14, 0, 0, 16, 8, 
    0, 0, 0, 0, 0, 19, 0, 0, 1, 29, 0, 6, 0, 8, 11, 
    0, 0, 0, 0, 18, 43, 0, 10, 21, 23, 0, 12, 14, 17, 5, 
    0, 0, 0, 0, 2, 0, 8, 19, 25, 23, 0, 8, 17, 1, 0, 
    3, 0, 0, 0, 0, 3, 31, 19, 27, 3, 7, 3, 7, 0, 8, 
    
    -- channel=576
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 40, 49, 58, 71, 61, 37, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 0, 0, 0, 18, 38, 16, 0, 0, 0, 5, 
    0, 0, 0, 0, 7, 3, 5, 36, 16, 3, 21, 22, 0, 0, 0, 
    0, 0, 25, 25, 29, 45, 41, 35, 33, 32, 18, 5, 0, 0, 0, 
    5, 0, 0, 1, 53, 33, 31, 45, 52, 45, 53, 48, 9, 0, 0, 
    4, 17, 18, 0, 0, 22, 26, 20, 16, 23, 22, 37, 60, 48, 1, 
    0, 25, 0, 0, 38, 34, 31, 31, 52, 54, 38, 54, 65, 52, 29, 
    0, 0, 0, 42, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    0, 0, 32, 0, 34, 25, 48, 38, 47, 55, 60, 57, 46, 40, 35, 
    0, 0, 0, 0, 10, 22, 0, 4, 42, 12, 20, 1, 18, 0, 18, 
    8, 13, 17, 0, 0, 14, 61, 32, 24, 14, 0, 19, 23, 56, 34, 
    17, 0, 0, 7, 0, 0, 2, 5, 6, 0, 0, 0, 5, 3, 11, 
    3, 18, 3, 11, 8, 0, 0, 0, 0, 57, 54, 18, 2, 4, 22, 
    23, 15, 0, 19, 13, 1, 0, 0, 3, 14, 32, 18, 0, 7, 7, 
    
    -- channel=577
    24, 18, 32, 10, 22, 14, 17, 15, 27, 34, 26, 29, 24, 8, 13, 
    36, 35, 46, 23, 38, 37, 22, 38, 51, 38, 26, 28, 31, 23, 18, 
    38, 38, 45, 27, 17, 16, 7, 12, 11, 2, 10, 30, 27, 25, 2, 
    38, 45, 24, 50, 19, 42, 43, 43, 39, 24, 11, 29, 30, 21, 1, 
    38, 46, 32, 45, 31, 19, 46, 33, 33, 29, 48, 10, 32, 38, 0, 
    33, 53, 26, 25, 0, 22, 20, 27, 27, 23, 28, 11, 21, 38, 38, 
    21, 37, 11, 20, 0, 18, 43, 15, 18, 41, 15, 6, 28, 35, 50, 
    34, 6, 0, 32, 24, 3, 0, 5, 6, 4, 0, 6, 6, 5, 31, 
    18, 0, 2, 2, 7, 2, 19, 2, 0, 0, 11, 0, 0, 8, 4, 
    32, 5, 18, 0, 0, 1, 0, 0, 39, 10, 25, 21, 36, 7, 0, 
    28, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    37, 17, 1, 4, 0, 0, 0, 13, 0, 26, 20, 18, 8, 5, 0, 
    32, 24, 0, 36, 3, 0, 0, 0, 0, 2, 29, 54, 0, 0, 0, 
    24, 41, 24, 33, 5, 0, 0, 0, 0, 4, 18, 58, 0, 0, 0, 
    34, 28, 30, 1, 3, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 
    
    -- channel=578
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 37, 38, 55, 81, 72, 40, 4, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 30, 13, 0, 10, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 28, 0, 0, 16, 20, 4, 32, 11, 0, 0, 0, 
    0, 21, 16, 0, 0, 0, 0, 0, 0, 8, 10, 24, 58, 50, 0, 
    0, 38, 0, 0, 8, 0, 0, 18, 57, 47, 37, 65, 46, 14, 0, 
    0, 0, 0, 64, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 36, 0, 25, 3, 26, 25, 25, 27, 40, 31, 31, 24, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 1, 0, 0, 0, 7, 0, 0, 
    0, 20, 5, 0, 0, 6, 70, 35, 30, 13, 0, 30, 24, 55, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 46, 34, 16, 0, 0, 0, 
    0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 16, 13, 0, 0, 0, 
    
    -- channel=579
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=580
    50, 50, 53, 29, 48, 54, 52, 58, 58, 48, 42, 48, 38, 38, 24, 
    61, 60, 56, 29, 60, 70, 64, 60, 64, 42, 34, 54, 46, 19, 39, 
    62, 63, 52, 23, 85, 91, 88, 83, 84, 71, 62, 58, 42, 14, 32, 
    61, 60, 52, 38, 109, 92, 79, 93, 92, 94, 65, 63, 41, 34, 23, 
    61, 58, 47, 47, 98, 86, 79, 93, 93, 89, 81, 84, 65, 46, 56, 
    65, 54, 45, 44, 70, 80, 82, 78, 74, 80, 75, 62, 80, 61, 63, 
    65, 38, 44, 41, 87, 89, 81, 75, 87, 82, 52, 65, 69, 65, 65, 
    51, 16, 58, 49, 66, 49, 59, 50, 41, 38, 42, 41, 59, 75, 90, 
    56, 23, 62, 14, 67, 63, 60, 45, 65, 71, 54, 57, 86, 75, 86, 
    51, 13, 50, 17, 56, 40, 50, 70, 55, 69, 58, 60, 72, 39, 87, 
    61, 12, 42, 33, 29, 42, 63, 37, 57, 47, 51, 65, 40, 68, 78, 
    71, 3, 50, 60, 20, 28, 43, 8, 68, 42, 60, 68, 4, 47, 75, 
    75, 42, 66, 63, 31, 20, 21, 26, 35, 93, 67, 43, 15, 40, 92, 
    82, 68, 49, 55, 49, 16, 22, 32, 45, 63, 63, 34, 11, 53, 86, 
    76, 73, 60, 38, 45, 26, 29, 35, 40, 49, 59, 39, 15, 47, 98, 
    
    -- channel=581
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 21, 27, 25, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=582
    22, 17, 26, 9, 14, 25, 33, 35, 15, 11, 4, 3, 38, 8, 24, 
    17, 16, 24, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    9, 8, 25, 72, 30, 50, 52, 63, 33, 0, 0, 9, 7, 4, 0, 
    10, 15, 9, 73, 0, 32, 47, 29, 46, 43, 9, 0, 20, 34, 0, 
    7, 20, 0, 48, 10, 0, 26, 23, 19, 16, 47, 0, 11, 53, 50, 
    0, 18, 50, 64, 0, 21, 25, 13, 10, 7, 0, 0, 0, 10, 9, 
    0, 11, 0, 57, 45, 24, 51, 33, 25, 29, 16, 0, 0, 0, 5, 
    11, 0, 0, 47, 17, 26, 5, 13, 0, 0, 0, 0, 0, 0, 0, 
    38, 52, 0, 0, 18, 5, 45, 79, 87, 74, 121, 95, 51, 28, 0, 
    34, 45, 0, 32, 0, 17, 0, 0, 13, 0, 0, 0, 0, 9, 0, 
    18, 76, 20, 31, 4, 0, 36, 23, 0, 22, 20, 29, 0, 41, 0, 
    21, 51, 0, 57, 49, 0, 0, 26, 0, 19, 33, 0, 33, 0, 0, 
    22, 119, 33, 31, 55, 32, 8, 5, 0, 14, 64, 94, 19, 5, 0, 
    19, 29, 48, 29, 24, 49, 16, 10, 6, 0, 0, 60, 22, 0, 0, 
    21, 32, 52, 17, 16, 30, 20, 18, 9, 1, 0, 41, 26, 0, 0, 
    
    -- channel=583
    6, 3, 6, 10, 2, 5, 6, 8, 7, 6, 6, 1, 5, 7, 5, 
    9, 8, 14, 26, 14, 13, 18, 16, 7, 0, 2, 0, 1, 3, 0, 
    9, 10, 12, 36, 29, 42, 40, 42, 41, 27, 0, 1, 5, 0, 0, 
    9, 10, 13, 41, 32, 26, 50, 49, 46, 48, 26, 0, 0, 7, 0, 
    7, 13, 23, 37, 33, 42, 43, 49, 47, 44, 37, 8, 0, 2, 1, 
    0, 14, 17, 50, 34, 36, 48, 46, 43, 41, 44, 20, 2, 10, 9, 
    1, 9, 7, 30, 36, 48, 44, 43, 40, 37, 28, 15, 6, 2, 1, 
    0, 13, 0, 16, 34, 31, 38, 38, 31, 27, 35, 28, 18, 19, 0, 
    6, 18, 0, 30, 18, 29, 23, 21, 19, 22, 19, 18, 26, 36, 2, 
    6, 31, 0, 17, 23, 21, 21, 18, 20, 26, 26, 22, 19, 30, 1, 
    7, 29, 18, 15, 21, 18, 15, 39, 7, 34, 26, 12, 44, 18, 12, 
    16, 32, 1, 20, 27, 15, 20, 16, 15, 10, 16, 25, 18, 20, 0, 
    23, 24, 23, 22, 20, 24, 13, 12, 15, 0, 21, 28, 26, 11, 9, 
    24, 28, 30, 21, 23, 21, 13, 14, 10, 14, 14, 28, 15, 13, 14, 
    32, 29, 30, 30, 22, 18, 15, 14, 16, 19, 19, 23, 21, 11, 13, 
    
    -- channel=584
    1, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    1, 1, 9, 19, 16, 17, 4, 2, 0, 0, 0, 0, 0, 0, 0, 
    1, 1, 10, 55, 36, 48, 49, 59, 48, 29, 0, 0, 0, 0, 0, 
    1, 8, 2, 59, 15, 19, 53, 53, 52, 42, 30, 0, 0, 2, 0, 
    0, 9, 14, 52, 30, 34, 47, 47, 43, 40, 55, 0, 0, 16, 1, 
    0, 11, 21, 60, 9, 41, 47, 42, 40, 38, 25, 9, 0, 1, 1, 
    0, 6, 0, 32, 38, 38, 59, 43, 34, 39, 28, 2, 0, 0, 0, 
    0, 4, 0, 29, 37, 40, 29, 32, 13, 13, 20, 6, 2, 13, 0, 
    4, 18, 0, 3, 19, 3, 21, 34, 27, 14, 47, 29, 14, 22, 0, 
    11, 35, 0, 21, 2, 27, 10, 0, 32, 17, 27, 22, 21, 26, 0, 
    5, 40, 12, 22, 8, 0, 16, 31, 0, 29, 29, 20, 12, 29, 0, 
    19, 48, 0, 29, 29, 2, 0, 25, 0, 9, 19, 5, 29, 0, 0, 
    23, 66, 15, 30, 37, 19, 3, 2, 0, 0, 20, 56, 14, 0, 0, 
    21, 29, 42, 26, 23, 31, 4, 1, 0, 0, 5, 58, 13, 0, 0, 
    31, 36, 44, 19, 18, 20, 9, 10, 7, 7, 4, 34, 14, 0, 0, 
    
    -- channel=585
    12, 5, 22, 32, 12, 9, 0, 0, 0, 9, 13, 7, 20, 5, 16, 
    12, 11, 32, 52, 16, 5, 5, 13, 6, 0, 8, 3, 13, 27, 0, 
    14, 14, 33, 80, 0, 4, 0, 10, 10, 0, 0, 8, 28, 34, 0, 
    14, 22, 21, 83, 0, 0, 28, 5, 3, 0, 1, 0, 22, 34, 10, 
    12, 29, 37, 56, 0, 0, 20, 1, 1, 0, 13, 0, 0, 31, 7, 
    4, 40, 30, 64, 0, 0, 13, 8, 9, 1, 4, 0, 0, 15, 13, 
    14, 51, 28, 43, 0, 5, 18, 11, 0, 5, 12, 0, 0, 0, 4, 
    34, 60, 0, 49, 12, 23, 15, 25, 14, 10, 20, 8, 0, 0, 0, 
    36, 51, 0, 63, 0, 2, 3, 19, 0, 0, 20, 0, 0, 7, 0, 
    35, 72, 8, 28, 0, 20, 0, 0, 32, 7, 23, 15, 11, 33, 0, 
    24, 74, 19, 21, 12, 0, 0, 37, 0, 29, 17, 0, 34, 0, 0, 
    24, 84, 0, 14, 37, 0, 0, 41, 0, 14, 8, 10, 46, 11, 0, 
    16, 50, 0, 29, 29, 27, 6, 0, 0, 0, 10, 63, 31, 0, 0, 
    8, 31, 40, 30, 14, 38, 4, 0, 0, 0, 2, 79, 21, 0, 0, 
    19, 16, 37, 33, 13, 22, 6, 4, 0, 1, 0, 47, 23, 0, 0, 
    
    -- channel=586
    0, 0, 0, 0, 0, 0, 0, 0, 8, 5, 0, 8, 0, 0, 0, 
    1, 1, 0, 0, 20, 37, 45, 59, 67, 60, 16, 15, 9, 0, 12, 
    6, 8, 0, 0, 0, 0, 0, 0, 0, 9, 54, 10, 0, 0, 43, 
    6, 0, 0, 0, 50, 38, 0, 7, 0, 1, 13, 53, 0, 0, 1, 
    12, 0, 0, 0, 34, 26, 0, 13, 18, 17, 0, 52, 19, 0, 0, 
    33, 0, 0, 0, 40, 1, 0, 11, 14, 12, 32, 45, 50, 6, 7, 
    20, 0, 0, 0, 0, 1, 0, 0, 8, 22, 1, 46, 80, 72, 29, 
    4, 0, 25, 0, 0, 0, 0, 0, 18, 18, 0, 31, 56, 34, 86, 
    0, 0, 23, 0, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 109, 
    0, 0, 36, 0, 27, 0, 12, 44, 6, 16, 9, 13, 23, 0, 93, 
    0, 0, 0, 0, 0, 8, 0, 0, 34, 0, 0, 0, 0, 0, 72, 
    0, 0, 24, 0, 0, 0, 47, 0, 67, 8, 0, 30, 0, 32, 79, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 0, 0, 0, 64, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 63, 33, 0, 0, 9, 61, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 53, 
    
    -- channel=587
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 33, 27, 32, 27, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 0, 0, 0, 2, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 12, 5, 1, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 36, 9, 3, 19, 20, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 25, 24, 11, 6, 16, 12, 4, 8, 0, 0, 
    0, 0, 0, 0, 39, 0, 20, 38, 73, 74, 39, 71, 54, 0, 0, 
    0, 0, 0, 19, 12, 11, 10, 10, 0, 0, 0, 0, 0, 0, 32, 
    0, 0, 19, 19, 31, 37, 62, 0, 36, 5, 21, 44, 0, 35, 31, 
    0, 0, 16, 31, 23, 34, 2, 2, 24, 0, 0, 0, 0, 0, 53, 
    0, 12, 31, 0, 21, 32, 45, 48, 56, 47, 0, 0, 18, 51, 54, 
    0, 0, 0, 0, 14, 22, 52, 52, 40, 0, 0, 0, 33, 48, 46, 
    0, 0, 0, 0, 15, 25, 43, 42, 38, 25, 5, 0, 35, 46, 57, 
    
    -- channel=588
    2, 8, 0, 0, 0, 0, 2, 18, 8, 0, 2, 0, 6, 12, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 28, 0, 19, 18, 0, 0, 
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 7, 0, 0, 0, 0, 0, 1, 15, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 1, 2, 2, 0, 0, 0, 0, 2, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    
    -- channel=589
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    
    -- channel=590
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 46, 51, 61, 82, 81, 50, 11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 8, 0, 0, 10, 10, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 24, 0, 0, 0, 
    0, 0, 24, 21, 0, 15, 19, 0, 5, 0, 0, 0, 0, 0, 0, 
    2, 7, 0, 0, 17, 0, 0, 15, 18, 7, 25, 14, 0, 0, 0, 
    0, 20, 15, 0, 0, 0, 6, 0, 2, 19, 17, 31, 61, 56, 0, 
    5, 30, 0, 0, 7, 0, 0, 14, 42, 33, 32, 55, 41, 23, 13, 
    0, 0, 0, 42, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 38, 0, 15, 10, 20, 33, 27, 30, 41, 33, 37, 22, 0, 
    0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 18, 10, 0, 0, 4, 57, 40, 31, 27, 0, 33, 32, 39, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 3, 0, 7, 0, 0, 0, 0, 0, 35, 40, 26, 0, 0, 0, 
    2, 0, 0, 7, 2, 0, 0, 0, 0, 0, 14, 17, 0, 0, 0, 
    
    -- channel=591
    0, 0, 0, 0, 0, 0, 0, 6, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 8, 14, 0, 14, 0, 0, 18, 
    0, 0, 0, 0, 34, 10, 2, 0, 0, 13, 62, 6, 0, 0, 37, 
    0, 0, 0, 0, 69, 11, 0, 0, 0, 3, 0, 47, 0, 0, 0, 
    0, 0, 0, 0, 45, 11, 0, 4, 5, 6, 0, 49, 11, 0, 0, 
    23, 0, 0, 0, 43, 11, 0, 0, 0, 20, 11, 36, 66, 0, 0, 
    15, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 30, 38, 23, 15, 
    0, 0, 56, 0, 0, 0, 5, 0, 2, 9, 0, 13, 52, 36, 93, 
    0, 0, 43, 0, 38, 2, 0, 0, 9, 18, 0, 0, 36, 0, 91, 
    0, 0, 23, 0, 25, 0, 19, 51, 0, 14, 0, 2, 3, 0, 122, 
    0, 0, 0, 0, 0, 28, 36, 0, 70, 0, 7, 48, 0, 28, 82, 
    0, 0, 39, 0, 0, 6, 42, 0, 78, 0, 0, 5, 0, 21, 122, 
    0, 0, 0, 0, 0, 0, 1, 11, 32, 106, 0, 0, 0, 32, 111, 
    2, 0, 0, 0, 0, 0, 2, 13, 22, 49, 27, 0, 0, 51, 96, 
    0, 0, 0, 0, 0, 0, 0, 4, 11, 18, 27, 0, 0, 41, 119, 
    
    -- channel=592
    0, 0, 0, 0, 0, 13, 28, 43, 20, 0, 0, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 36, 52, 57, 53, 33, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 60, 48, 41, 34, 47, 57, 21, 0, 0, 0, 0, 
    0, 0, 0, 0, 45, 27, 13, 41, 36, 37, 27, 20, 4, 0, 22, 
    0, 0, 5, 17, 14, 27, 32, 27, 18, 23, 11, 0, 0, 0, 0, 
    0, 0, 0, 5, 79, 49, 40, 41, 53, 44, 18, 9, 0, 0, 0, 
    0, 0, 0, 12, 15, 2, 6, 8, 0, 0, 3, 0, 0, 3, 0, 
    0, 3, 12, 0, 33, 33, 44, 44, 81, 96, 79, 83, 89, 49, 16, 
    0, 0, 0, 5, 13, 3, 0, 10, 0, 0, 0, 0, 0, 0, 25, 
    0, 0, 18, 11, 10, 11, 48, 19, 0, 5, 6, 25, 0, 38, 40, 
    0, 0, 4, 45, 21, 15, 0, 0, 30, 3, 29, 13, 0, 0, 22, 
    8, 31, 60, 11, 14, 18, 15, 18, 20, 73, 59, 27, 7, 22, 58, 
    22, 3, 8, 7, 18, 8, 22, 28, 38, 0, 0, 0, 2, 34, 44, 
    11, 17, 14, 0, 15, 9, 23, 24, 22, 17, 9, 0, 15, 26, 56, 
    
    -- channel=593
    26, 21, 36, 34, 16, 4, 5, 8, 18, 29, 35, 23, 32, 25, 28, 
    27, 26, 51, 48, 14, 0, 0, 6, 15, 7, 24, 22, 30, 48, 17, 
    28, 28, 43, 67, 0, 0, 0, 0, 0, 0, 0, 23, 45, 52, 2, 
    28, 40, 19, 76, 0, 0, 15, 0, 0, 0, 0, 0, 24, 51, 20, 
    25, 44, 40, 29, 0, 0, 0, 0, 0, 0, 0, 0, 8, 39, 9, 
    9, 57, 15, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 27, 
    9, 44, 12, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    31, 33, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 21, 0, 20, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    30, 51, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 2, 0, 0, 
    19, 49, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 
    15, 58, 0, 0, 5, 0, 0, 5, 0, 0, 0, 11, 8, 0, 0, 
    0, 20, 0, 17, 0, 0, 0, 0, 0, 0, 10, 68, 0, 0, 0, 
    0, 14, 16, 19, 0, 7, 0, 0, 0, 0, 0, 71, 0, 0, 0, 
    0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    
    -- channel=594
    18, 18, 20, 0, 1, 8, 18, 29, 9, 2, 0, 0, 34, 5, 19, 
    13, 13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 4, 11, 47, 0, 20, 27, 36, 7, 0, 0, 3, 0, 0, 0, 
    5, 6, 4, 33, 0, 0, 7, 0, 5, 9, 0, 0, 13, 24, 0, 
    2, 9, 0, 7, 0, 0, 0, 0, 0, 0, 11, 0, 6, 48, 60, 
    0, 0, 32, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 5, 
    0, 0, 0, 26, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 31, 0, 0, 0, 0, 4, 46, 74, 65, 92, 81, 39, 0, 0, 
    21, 19, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 44, 0, 0, 0, 0, 8, 0, 0, 0, 0, 5, 0, 6, 0, 
    1, 14, 0, 26, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 94, 18, 0, 17, 0, 0, 0, 0, 0, 36, 44, 0, 0, 0, 
    0, 0, 12, 0, 0, 5, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 3, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=595
    61, 62, 67, 45, 37, 41, 44, 57, 62, 61, 59, 56, 59, 50, 40, 
    76, 75, 75, 47, 29, 29, 25, 26, 33, 30, 34, 56, 59, 47, 40, 
    77, 76, 70, 55, 22, 44, 45, 48, 39, 29, 22, 61, 63, 38, 20, 
    76, 78, 63, 58, 29, 48, 67, 49, 51, 48, 48, 37, 55, 52, 27, 
    74, 76, 59, 38, 30, 43, 43, 42, 45, 47, 55, 41, 66, 70, 63, 
    64, 74, 56, 45, 0, 26, 35, 28, 25, 32, 31, 32, 55, 77, 77, 
    59, 53, 35, 30, 37, 37, 39, 23, 26, 32, 13, 9, 24, 38, 68, 
    56, 28, 13, 52, 22, 9, 1, 3, 0, 0, 0, 0, 0, 27, 45, 
    62, 32, 27, 0, 8, 16, 22, 18, 27, 30, 41, 25, 39, 41, 30, 
    64, 37, 0, 0, 0, 0, 0, 4, 30, 24, 25, 20, 28, 13, 16, 
    61, 36, 3, 0, 0, 0, 4, 16, 0, 20, 10, 17, 12, 21, 19, 
    63, 30, 0, 22, 0, 0, 0, 0, 0, 9, 23, 29, 0, 0, 0, 
    55, 50, 27, 27, 5, 0, 0, 0, 0, 15, 56, 50, 0, 0, 11, 
    55, 50, 39, 18, 5, 0, 0, 0, 0, 1, 18, 34, 0, 0, 10, 
    49, 46, 40, 3, 0, 0, 0, 0, 0, 0, 4, 7, 0, 0, 16, 
    
    -- channel=596
    0, 0, 0, 0, 0, 0, 0, 9, 12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 11, 
    0, 0, 0, 0, 18, 6, 0, 0, 0, 7, 31, 11, 0, 0, 23, 
    0, 0, 0, 0, 57, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 
    0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 38, 2, 0, 0, 
    3, 0, 0, 0, 22, 0, 0, 0, 0, 0, 0, 3, 40, 0, 0, 
    5, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 16, 26, 0, 0, 
    0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 8, 60, 
    0, 0, 39, 0, 15, 0, 0, 0, 14, 20, 0, 7, 45, 0, 60, 
    0, 0, 19, 0, 22, 0, 4, 17, 0, 0, 0, 0, 0, 0, 69, 
    0, 0, 5, 0, 0, 9, 13, 0, 29, 0, 0, 20, 0, 8, 45, 
    0, 0, 22, 4, 0, 0, 22, 0, 69, 0, 0, 19, 0, 20, 55, 
    0, 0, 10, 1, 0, 0, 0, 3, 13, 88, 0, 0, 0, 14, 76, 
    0, 0, 0, 0, 0, 0, 0, 9, 14, 47, 0, 0, 0, 38, 56, 
    0, 0, 0, 0, 0, 0, 0, 0, 4, 9, 12, 0, 0, 27, 81, 
    
    -- channel=597
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 8, 
    0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 92, 0, 7, 9, 30, 10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 74, 0, 0, 6, 0, 0, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 18, 
    0, 0, 15, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 15, 0, 28, 0, 17, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    5, 51, 0, 18, 0, 0, 0, 44, 44, 23, 75, 61, 6, 0, 0, 
    2, 70, 0, 36, 0, 6, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 85, 6, 18, 11, 0, 0, 43, 0, 24, 6, 0, 21, 0, 0, 
    0, 87, 0, 16, 57, 0, 0, 17, 0, 0, 0, 0, 36, 0, 0, 
    0, 86, 18, 0, 39, 42, 4, 0, 0, 0, 4, 65, 28, 0, 0, 
    0, 0, 24, 0, 0, 49, 13, 0, 0, 0, 0, 53, 28, 0, 0, 
    0, 0, 26, 15, 0, 20, 14, 7, 0, 0, 0, 12, 37, 0, 0, 
    
    -- channel=598
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 57, 17, 11, 25, 37, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 63, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 41, 60, 0, 3, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 53, 3, 0, 5, 18, 23, 0, 12, 0, 0, 0, 0, 
    0, 32, 14, 11, 0, 0, 22, 11, 0, 13, 26, 0, 0, 0, 0, 
    2, 69, 0, 16, 24, 21, 4, 25, 47, 45, 32, 43, 16, 0, 0, 
    0, 41, 0, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 70, 6, 33, 9, 25, 16, 0, 37, 7, 35, 22, 8, 48, 0, 
    0, 66, 0, 14, 19, 3, 0, 32, 0, 5, 0, 0, 32, 0, 0, 
    0, 105, 0, 0, 32, 12, 23, 70, 0, 20, 0, 0, 85, 24, 0, 
    0, 0, 0, 0, 20, 19, 11, 4, 0, 0, 0, 16, 47, 0, 0, 
    0, 11, 21, 10, 6, 36, 0, 0, 0, 0, 2, 55, 34, 0, 0, 
    2, 0, 6, 38, 7, 23, 0, 0, 0, 0, 0, 36, 28, 0, 0, 
    
    -- channel=599
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 17, 25, 3, 28, 45, 14, 0, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 
    0, 0, 10, 0, 30, 0, 25, 31, 0, 0, 0, 0, 0, 0, 58, 
    0, 0, 0, 0, 11, 29, 0, 0, 35, 0, 0, 0, 0, 0, 53, 
    0, 0, 19, 0, 0, 24, 53, 0, 60, 0, 0, 0, 0, 26, 75, 
    0, 0, 0, 0, 0, 0, 18, 23, 35, 0, 0, 0, 0, 25, 58, 
    0, 0, 0, 0, 0, 0, 12, 16, 15, 40, 4, 0, 1, 35, 50, 
    0, 0, 0, 0, 0, 0, 5, 5, 11, 11, 16, 0, 0, 28, 37, 
    
    -- channel=600
    67, 65, 71, 50, 46, 49, 50, 60, 75, 74, 70, 71, 57, 58, 41, 
    84, 84, 83, 44, 46, 51, 52, 61, 71, 65, 57, 75, 76, 59, 57, 
    89, 89, 78, 26, 23, 33, 30, 27, 31, 40, 50, 75, 74, 51, 52, 
    88, 88, 71, 35, 54, 65, 62, 54, 49, 47, 56, 72, 64, 52, 44, 
    89, 86, 67, 25, 45, 54, 45, 49, 55, 55, 55, 64, 79, 63, 50, 
    88, 86, 46, 24, 23, 33, 37, 37, 36, 42, 48, 50, 81, 89, 89, 
    78, 64, 50, 19, 23, 38, 35, 22, 30, 40, 24, 40, 70, 78, 89, 
    73, 34, 31, 46, 26, 13, 13, 13, 8, 3, 5, 9, 21, 44, 84, 
    57, 13, 46, 6, 18, 29, 20, 0, 0, 5, 5, 0, 21, 43, 73, 
    64, 17, 23, 0, 11, 0, 11, 30, 41, 42, 40, 36, 48, 17, 50, 
    69, 9, 5, 0, 0, 0, 0, 8, 10, 18, 13, 18, 14, 20, 43, 
    69, 9, 1, 10, 0, 0, 11, 0, 17, 19, 25, 53, 0, 13, 29, 
    60, 12, 15, 35, 0, 0, 0, 0, 0, 34, 48, 30, 0, 0, 33, 
    62, 57, 30, 27, 8, 0, 0, 0, 0, 35, 43, 29, 0, 0, 32, 
    56, 46, 33, 7, 3, 0, 0, 0, 0, 3, 23, 13, 0, 0, 37, 
    
    -- channel=601
    19, 20, 12, 0, 9, 26, 46, 61, 34, 9, 1, 4, 31, 21, 25, 
    10, 11, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 13, 26, 26, 28, 1, 0, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 10, 15, 0, 0, 5, 18, 0, 0, 6, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 17, 33, 60, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 1, 0, 0, 2, 0, 26, 52, 102, 104, 113, 112, 79, 7, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 1, 0, 0, 36, 0, 0, 0, 0, 18, 0, 25, 0, 
    0, 0, 0, 47, 9, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 
    0, 60, 37, 1, 11, 4, 0, 0, 0, 69, 63, 39, 0, 8, 4, 
    0, 0, 0, 0, 0, 4, 14, 13, 13, 0, 0, 0, 0, 4, 0, 
    0, 0, 2, 0, 0, 0, 13, 11, 1, 0, 0, 0, 0, 4, 15, 
    
    -- channel=602
    32, 30, 31, 0, 6, 26, 37, 49, 38, 23, 13, 16, 31, 25, 13, 
    36, 36, 30, 0, 0, 0, 0, 0, 0, 0, 0, 16, 12, 0, 4, 
    31, 31, 25, 1, 48, 75, 71, 72, 58, 26, 7, 31, 10, 0, 0, 
    31, 28, 19, 11, 51, 50, 44, 48, 61, 72, 35, 0, 18, 21, 0, 
    27, 29, 0, 0, 45, 28, 22, 49, 46, 40, 52, 41, 31, 42, 58, 
    13, 14, 16, 22, 6, 31, 38, 23, 20, 28, 20, 15, 33, 31, 32, 
    14, 0, 0, 16, 58, 42, 38, 33, 36, 30, 0, 0, 0, 0, 21, 
    0, 0, 1, 7, 10, 16, 17, 0, 0, 0, 0, 0, 0, 7, 32, 
    26, 0, 5, 0, 20, 9, 24, 50, 85, 85, 85, 87, 84, 41, 24, 
    22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 19, 
    20, 0, 9, 0, 0, 0, 38, 6, 1, 21, 17, 45, 9, 30, 28, 
    24, 0, 0, 41, 2, 0, 0, 0, 0, 0, 24, 1, 0, 0, 0, 
    33, 55, 47, 21, 6, 0, 0, 0, 0, 55, 56, 33, 0, 0, 30, 
    39, 25, 18, 11, 6, 0, 0, 0, 0, 0, 0, 3, 0, 0, 25, 
    30, 35, 32, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 41, 
    
    -- channel=603
    31, 28, 28, 29, 18, 20, 24, 21, 26, 32, 28, 28, 31, 24, 29, 
    35, 35, 35, 39, 25, 24, 29, 31, 25, 25, 27, 22, 28, 28, 18, 
    36, 36, 40, 46, 35, 43, 44, 47, 43, 32, 17, 25, 25, 23, 13, 
    36, 36, 38, 52, 22, 44, 55, 55, 53, 52, 37, 17, 31, 22, 15, 
    34, 37, 40, 49, 31, 43, 51, 51, 49, 51, 51, 23, 27, 36, 23, 
    24, 34, 36, 48, 32, 41, 45, 44, 45, 41, 44, 37, 21, 37, 36, 
    19, 32, 21, 38, 30, 41, 45, 39, 33, 35, 33, 22, 24, 30, 32, 
    15, 26, 4, 18, 38, 40, 34, 30, 24, 27, 22, 18, 22, 26, 18, 
    21, 28, 0, 37, 18, 21, 31, 37, 14, 18, 29, 19, 16, 30, 24, 
    30, 35, 6, 18, 17, 22, 20, 15, 37, 30, 36, 33, 25, 39, 13, 
    27, 42, 13, 16, 13, 16, 21, 25, 20, 32, 28, 24, 36, 18, 20, 
    33, 43, 7, 17, 24, 5, 8, 25, 0, 23, 22, 13, 32, 17, 10, 
    38, 41, 16, 23, 26, 14, 4, 5, 10, 0, 30, 31, 21, 9, 9, 
    32, 42, 36, 23, 22, 22, 5, 5, 2, 16, 26, 37, 14, 3, 18, 
    43, 41, 37, 32, 19, 19, 10, 10, 11, 14, 18, 30, 16, 6, 13, 
    
    -- channel=604
    5, 6, 0, 15, 0, 0, 3, 8, 1, 1, 7, 0, 17, 14, 25, 
    0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 1, 0, 0, 18, 0, 
    0, 0, 0, 43, 0, 0, 1, 9, 0, 0, 0, 0, 2, 17, 0, 
    0, 0, 0, 23, 0, 0, 5, 0, 0, 0, 7, 0, 2, 14, 13, 
    0, 0, 1, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 
    0, 0, 12, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 13, 0, 7, 0, 13, 4, 5, 0, 0, 4, 0, 0, 0, 0, 
    0, 29, 0, 15, 0, 0, 3, 23, 21, 20, 31, 30, 4, 0, 0, 
    0, 39, 0, 33, 0, 10, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 40, 12, 15, 19, 0, 3, 27, 0, 14, 7, 0, 17, 0, 0, 
    0, 44, 0, 8, 37, 15, 0, 20, 0, 0, 0, 0, 35, 0, 0, 
    0, 35, 10, 0, 24, 30, 19, 15, 11, 0, 6, 21, 31, 5, 0, 
    0, 0, 12, 0, 4, 32, 22, 15, 3, 0, 0, 10, 29, 0, 0, 
    0, 0, 5, 11, 5, 20, 20, 14, 9, 0, 0, 1, 33, 1, 0, 
    
    -- channel=605
    0, 0, 0, 0, 0, 0, 0, 10, 5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 12, 3, 7, 3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 22, 29, 31, 30, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 2, 0, 0, 0, 0, 0, 21, 12, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=606
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=607
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=608
    0, 0, 16, 0, 3, 0, 0, 9, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 4, 2, 0, 0, 0, 0, 0, 10, 0, 0, 0, 
    0, 0, 0, 0, 34, 34, 3, 10, 10, 0, 1, 14, 0, 0, 0, 
    0, 2, 0, 0, 38, 0, 0, 0, 6, 0, 0, 16, 0, 5, 0, 
    0, 2, 0, 0, 47, 0, 0, 0, 0, 0, 10, 0, 0, 9, 7, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 3, 0, 0, 0, 0, 7, 
    0, 0, 0, 22, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 42, 
    0, 0, 34, 0, 20, 0, 0, 0, 49, 5, 47, 46, 44, 0, 0, 
    0, 0, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 
    0, 0, 14, 1, 0, 0, 8, 0, 12, 0, 16, 44, 0, 40, 0, 
    0, 0, 19, 46, 0, 0, 0, 0, 0, 0, 21, 12, 0, 14, 0, 
    0, 7, 1, 62, 0, 0, 0, 0, 0, 79, 10, 59, 0, 0, 0, 
    2, 0, 0, 49, 0, 0, 0, 0, 0, 4, 0, 52, 0, 3, 0, 
    0, 0, 17, 0, 8, 0, 0, 6, 0, 0, 0, 28, 0, 9, 1, 
    
    -- channel=609
    72, 63, 74, 48, 45, 48, 57, 63, 77, 84, 75, 76, 67, 67, 50, 
    85, 84, 91, 32, 32, 33, 23, 43, 63, 70, 63, 74, 80, 76, 64, 
    87, 87, 85, 11, 3, 16, 6, 8, 9, 15, 46, 81, 76, 62, 54, 
    86, 90, 59, 36, 31, 55, 40, 35, 34, 33, 41, 66, 69, 69, 40, 
    86, 90, 49, 9, 30, 19, 25, 27, 35, 23, 47, 57, 75, 78, 46, 
    76, 91, 27, 11, 0, 6, 12, 14, 15, 16, 35, 32, 72, 86, 87, 
    60, 61, 28, 6, 0, 10, 22, 1, 7, 34, 5, 11, 51, 62, 86, 
    65, 11, 11, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 79, 
    49, 0, 25, 0, 0, 13, 7, 2, 0, 0, 22, 0, 0, 28, 51, 
    59, 0, 26, 0, 0, 0, 0, 0, 25, 10, 18, 13, 39, 0, 4, 
    58, 8, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 3, 0, 
    53, 0, 0, 2, 0, 0, 0, 0, 0, 11, 23, 41, 0, 6, 0, 
    44, 12, 0, 38, 0, 0, 0, 0, 0, 31, 53, 55, 0, 0, 0, 
    42, 48, 20, 36, 0, 0, 0, 0, 0, 15, 17, 48, 0, 0, 0, 
    38, 31, 29, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 0, 0, 
    
    -- channel=610
    11, 11, 9, 0, 0, 0, 7, 10, 0, 0, 0, 0, 19, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 35, 34, 38, 37, 24, 0, 5, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 56, 
    0, 0, 6, 0, 0, 5, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 23, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17, 0, 0, 18, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 37, 87, 65, 57, 85, 50, 0, 0, 
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 4, 0, 0, 43, 0, 21, 18, 23, 61, 0, 24, 0, 
    0, 0, 6, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 62, 17, 0, 15, 0, 0, 0, 9, 31, 0, 0, 0, 14, 9, 
    0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 0, 2, 2, 5, 
    0, 0, 0, 0, 0, 0, 10, 11, 5, 0, 0, 0, 0, 9, 30, 
    
    -- channel=611
    11, 12, 11, 20, 11, 0, 0, 3, 18, 25, 29, 22, 5, 20, 12, 
    18, 17, 22, 31, 31, 33, 42, 53, 55, 49, 36, 24, 26, 34, 27, 
    23, 23, 18, 2, 0, 0, 0, 0, 0, 16, 23, 14, 26, 32, 40, 
    22, 25, 17, 6, 9, 5, 14, 14, 1, 0, 22, 33, 8, 10, 28, 
    22, 22, 41, 11, 8, 27, 16, 11, 16, 17, 6, 12, 14, 0, 0, 
    24, 29, 0, 4, 16, 2, 9, 19, 18, 18, 31, 25, 22, 22, 22, 
    15, 21, 18, 0, 0, 6, 5, 0, 6, 17, 16, 30, 47, 47, 24, 
    14, 22, 0, 6, 12, 0, 0, 16, 30, 21, 24, 39, 23, 20, 21, 
    0, 0, 9, 20, 0, 16, 0, 0, 0, 0, 0, 0, 0, 6, 22, 
    2, 14, 17, 0, 15, 5, 18, 28, 15, 24, 26, 21, 26, 13, 17, 
    8, 0, 0, 0, 4, 2, 0, 11, 0, 0, 0, 0, 8, 0, 11, 
    11, 18, 0, 0, 0, 12, 44, 10, 31, 11, 0, 37, 15, 26, 14, 
    5, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 4, 
    7, 10, 2, 6, 2, 0, 0, 0, 2, 30, 24, 10, 0, 0, 5, 
    10, 3, 0, 6, 5, 0, 0, 0, 0, 3, 16, 0, 0, 0, 0, 
    
    -- channel=612
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 16, 
    0, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 20, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 43, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 22, 
    0, 0, 26, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 7, 0, 0, 0, 
    0, 0, 24, 0, 0, 0, 7, 0, 34, 0, 0, 4, 0, 14, 10, 
    0, 0, 0, 2, 0, 0, 2, 5, 1, 61, 0, 0, 0, 6, 23, 
    0, 0, 0, 0, 0, 0, 3, 5, 9, 25, 0, 0, 0, 19, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 27, 
    
    -- channel=613
    5, 13, 0, 0, 0, 14, 37, 67, 34, 0, 0, 0, 12, 26, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 30, 29, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 14, 0, 0, 0, 15, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 4, 62, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 2, 0, 0, 0, 2, 37, 123, 134, 116, 132, 118, 28, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 0, 0, 0, 28, 9, 0, 0, 0, 5, 0, 4, 13, 
    0, 0, 0, 40, 15, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    0, 30, 78, 0, 0, 12, 0, 0, 0, 65, 66, 25, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 12, 14, 18, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 10, 8, 1, 0, 0, 0, 4, 1, 22, 
    
    -- channel=614
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 11, 8, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 24, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 1, 0, 17, 13, 0, 2, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 13, 0, 9, 0, 10, 2, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 7, 46, 0, 42, 0, 0, 7, 0, 31, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    
    -- channel=615
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 22, 22, 22, 27, 17, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 9, 37, 0, 0, 0, 13, 
    0, 0, 0, 0, 55, 10, 0, 0, 0, 0, 0, 29, 0, 0, 0, 
    0, 0, 0, 0, 34, 13, 0, 2, 3, 2, 0, 31, 0, 0, 0, 
    4, 0, 0, 0, 41, 7, 0, 5, 6, 12, 11, 24, 31, 0, 0, 
    5, 0, 0, 0, 0, 1, 0, 0, 13, 8, 0, 38, 48, 28, 0, 
    0, 0, 41, 0, 0, 0, 0, 0, 22, 25, 8, 33, 57, 34, 62, 
    0, 0, 36, 0, 30, 9, 0, 0, 0, 0, 0, 0, 0, 0, 74, 
    0, 0, 37, 0, 34, 0, 27, 52, 0, 17, 1, 10, 15, 0, 91, 
    0, 0, 0, 0, 0, 28, 12, 0, 51, 0, 0, 11, 0, 9, 63, 
    0, 0, 39, 0, 0, 14, 55, 0, 80, 5, 0, 20, 0, 34, 94, 
    0, 0, 0, 0, 0, 0, 8, 15, 25, 64, 0, 0, 0, 26, 80, 
    0, 0, 0, 0, 0, 0, 1, 11, 23, 54, 28, 0, 0, 41, 71, 
    0, 0, 0, 0, 2, 0, 0, 3, 10, 18, 30, 0, 0, 32, 76, 
    
    -- channel=616
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 58, 29, 21, 32, 55, 40, 20, 9, 0, 0, 15, 0, 
    0, 0, 9, 56, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 
    0, 0, 0, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 51, 60, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 0, 34, 0, 0, 0, 0, 8, 0, 3, 0, 0, 0, 0, 
    0, 51, 21, 4, 0, 0, 0, 0, 0, 0, 8, 0, 15, 17, 0, 
    11, 73, 0, 15, 8, 11, 0, 15, 31, 30, 18, 26, 7, 0, 0, 
    0, 21, 0, 96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 60, 13, 14, 0, 15, 9, 0, 40, 15, 42, 30, 19, 42, 0, 
    0, 55, 0, 2, 1, 0, 0, 10, 0, 0, 0, 0, 18, 0, 0, 
    0, 97, 0, 0, 6, 0, 16, 65, 0, 11, 0, 0, 69, 28, 0, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 11, 22, 0, 0, 
    0, 12, 11, 13, 0, 18, 0, 0, 0, 0, 15, 70, 16, 0, 0, 
    0, 0, 3, 27, 0, 6, 0, 0, 0, 0, 0, 37, 3, 0, 0, 
    
    -- channel=617
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=618
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 29, 46, 71, 84, 73, 56, 19, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 12, 43, 0, 0, 0, 42, 
    0, 0, 0, 0, 25, 9, 0, 10, 0, 0, 0, 46, 0, 0, 1, 
    0, 0, 22, 0, 20, 39, 22, 17, 17, 24, 0, 19, 0, 0, 0, 
    24, 0, 0, 0, 72, 21, 7, 34, 39, 32, 56, 54, 30, 0, 0, 
    13, 11, 32, 0, 0, 8, 0, 3, 12, 10, 15, 55, 81, 84, 1, 
    2, 31, 38, 0, 33, 10, 23, 18, 70, 73, 42, 78, 94, 57, 53, 
    0, 0, 8, 57, 15, 25, 0, 0, 0, 0, 0, 0, 0, 0, 83, 
    0, 0, 46, 0, 54, 11, 53, 86, 20, 54, 47, 49, 39, 31, 96, 
    0, 0, 0, 0, 15, 50, 0, 0, 64, 0, 2, 0, 23, 0, 75, 
    0, 0, 47, 0, 0, 25, 100, 28, 83, 25, 0, 26, 16, 65, 114, 
    9, 0, 0, 0, 0, 0, 11, 16, 31, 0, 0, 0, 5, 24, 63, 
    0, 0, 0, 0, 2, 0, 0, 1, 10, 71, 68, 0, 4, 31, 70, 
    9, 0, 0, 11, 7, 0, 0, 0, 7, 21, 47, 0, 0, 25, 47, 
    
    -- channel=619
    7, 14, 8, 0, 0, 2, 14, 35, 10, 0, 0, 0, 25, 14, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 55, 0, 31, 33, 45, 15, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 0, 0, 9, 0, 0, 0, 0, 0, 0, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 59, 
    0, 0, 15, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 15, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 27, 0, 0, 0, 0, 0, 48, 107, 98, 112, 117, 81, 5, 0, 
    1, 27, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 17, 6, 0, 0, 21, 28, 0, 15, 1, 16, 0, 8, 0, 
    0, 15, 0, 44, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 85, 54, 0, 24, 28, 0, 0, 0, 0, 39, 52, 4, 0, 0, 
    0, 0, 10, 0, 0, 24, 14, 8, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 13, 0, 0, 4, 16, 11, 1, 0, 0, 0, 22, 0, 0, 
    
    -- channel=620
    6, 19, 0, 0, 0, 14, 27, 47, 33, 0, 0, 2, 0, 17, 0, 
    3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 19, 
    0, 0, 0, 0, 32, 34, 35, 21, 15, 3, 36, 18, 0, 0, 19, 
    0, 0, 0, 0, 55, 15, 0, 0, 0, 19, 5, 10, 0, 0, 0, 
    0, 0, 0, 0, 34, 0, 0, 0, 0, 1, 0, 46, 23, 0, 45, 
    4, 0, 0, 0, 14, 2, 0, 0, 0, 0, 0, 9, 40, 0, 0, 
    7, 0, 0, 0, 49, 5, 0, 0, 9, 0, 0, 8, 0, 0, 0, 
    0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 10, 47, 
    0, 0, 37, 0, 16, 3, 4, 10, 80, 99, 39, 79, 105, 13, 66, 
    0, 0, 0, 0, 12, 0, 0, 15, 0, 0, 0, 0, 0, 0, 93, 
    0, 0, 8, 0, 0, 12, 55, 0, 30, 0, 0, 49, 0, 21, 88, 
    0, 0, 16, 24, 0, 5, 0, 0, 56, 0, 9, 0, 0, 0, 88, 
    0, 0, 57, 0, 0, 0, 0, 9, 29, 107, 26, 0, 0, 26, 120, 
    6, 0, 0, 0, 0, 0, 12, 21, 31, 23, 0, 0, 0, 52, 90, 
    0, 0, 0, 0, 0, 0, 10, 13, 16, 13, 7, 0, 0, 40, 115, 
    
    -- channel=621
    9, 18, 7, 1, 0, 13, 29, 49, 29, 2, 5, 0, 25, 17, 21, 
    4, 5, 3, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 47, 0, 11, 19, 26, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 20, 0, 8, 26, 0, 4, 4, 14, 0, 0, 23, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 22, 42, 
    0, 0, 27, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 40, 2, 1, 3, 0, 1, 4, 0, 0, 0, 0, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 39, 0, 0, 0, 0, 26, 44, 73, 82, 98, 85, 62, 20, 0, 
    7, 28, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 11, 6, 0, 0, 15, 23, 0, 0, 0, 0, 0, 7, 0, 
    0, 22, 0, 33, 37, 0, 0, 0, 0, 0, 9, 0, 12, 0, 0, 
    0, 64, 48, 0, 20, 20, 0, 0, 0, 6, 62, 57, 12, 0, 0, 
    0, 0, 10, 0, 0, 22, 9, 6, 10, 0, 0, 0, 5, 0, 0, 
    0, 0, 10, 0, 0, 3, 12, 7, 0, 0, 0, 0, 21, 0, 0, 
    
    -- channel=622
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=623
    12, 14, 2, 0, 0, 18, 40, 64, 27, 0, 0, 0, 25, 19, 15, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 23, 28, 25, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 0, 0, 0, 12, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 20, 70, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2, 0, 0, 0, 0, 0, 9, 43, 125, 126, 111, 128, 93, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 0, 0, 0, 38, 0, 0, 0, 0, 22, 0, 23, 0, 
    0, 0, 0, 44, 2, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 59, 46, 0, 3, 0, 0, 0, 0, 81, 48, 11, 0, 2, 16, 
    0, 0, 0, 0, 0, 0, 9, 11, 9, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 8, 6, 0, 0, 0, 0, 0, 0, 28, 
    
    -- channel=624
    11, 10, 15, 8, 12, 13, 11, 8, 6, 8, 7, 9, 10, 14, 7, 
    6, 6, 8, 0, 0, 0, 0, 0, 0, 0, 4, 11, 11, 12, 14, 
    5, 4, 7, 0, 0, 0, 0, 0, 0, 0, 8, 15, 12, 9, 11, 
    5, 6, 2, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 20, 9, 
    5, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 16, 23, 
    8, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 4, 5, 
    13, 11, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    22, 5, 19, 13, 0, 2, 7, 3, 0, 0, 0, 0, 0, 0, 11, 
    19, 3, 19, 1, 0, 0, 0, 11, 27, 16, 23, 28, 19, 0, 0, 
    14, 0, 18, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    11, 3, 13, 8, 8, 8, 9, 5, 11, 13, 10, 20, 10, 3, 0, 
    0, 0, 17, 13, 7, 6, 0, 0, 1, 0, 6, 0, 0, 10, 0, 
    0, 6, 12, 13, 4, 13, 11, 11, 9, 18, 7, 13, 3, 8, 0, 
    0, 0, 0, 14, 2, 8, 15, 12, 6, 0, 0, 8, 6, 8, 0, 
    0, 0, 2, 4, 5, 8, 11, 12, 10, 8, 3, 13, 8, 10, 0, 
    
    -- channel=625
    0, 0, 0, 0, 0, 6, 8, 12, 16, 0, 0, 4, 0, 1, 0, 
    0, 0, 0, 0, 0, 5, 9, 5, 12, 18, 0, 14, 0, 0, 19, 
    0, 0, 0, 0, 24, 7, 0, 0, 0, 13, 61, 13, 0, 0, 42, 
    0, 0, 0, 0, 66, 27, 0, 0, 0, 11, 6, 43, 0, 0, 0, 
    0, 0, 0, 0, 43, 16, 0, 8, 9, 9, 0, 61, 18, 0, 0, 
    21, 0, 0, 0, 47, 5, 0, 1, 2, 13, 16, 40, 58, 0, 0, 
    17, 0, 0, 0, 7, 7, 0, 0, 15, 1, 0, 35, 45, 31, 13, 
    0, 0, 49, 0, 0, 0, 0, 0, 4, 10, 0, 16, 51, 33, 86, 
    0, 0, 43, 0, 26, 14, 5, 0, 2, 24, 0, 0, 37, 2, 109, 
    0, 0, 27, 0, 36, 0, 19, 48, 0, 8, 0, 0, 0, 0, 122, 
    0, 0, 0, 0, 0, 30, 31, 0, 58, 0, 0, 30, 0, 10, 102, 
    0, 0, 38, 0, 0, 6, 42, 0, 88, 0, 3, 15, 0, 26, 114, 
    0, 0, 8, 0, 0, 0, 1, 11, 33, 95, 0, 0, 0, 29, 115, 
    2, 0, 0, 0, 0, 0, 2, 14, 25, 61, 20, 0, 0, 50, 99, 
    0, 0, 0, 0, 0, 0, 0, 3, 11, 17, 28, 0, 0, 38, 109, 
    
    -- channel=626
    22, 23, 21, 21, 27, 21, 25, 22, 20, 25, 25, 28, 27, 27, 29, 
    19, 19, 18, 9, 0, 0, 0, 0, 9, 21, 30, 25, 27, 31, 39, 
    17, 16, 18, 0, 0, 0, 0, 0, 0, 0, 26, 24, 23, 32, 36, 
    17, 16, 13, 0, 0, 0, 0, 0, 0, 0, 0, 27, 27, 30, 29, 
    18, 16, 3, 0, 0, 0, 0, 0, 0, 0, 0, 7, 22, 25, 28, 
    21, 17, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 17, 17, 
    16, 19, 15, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 18, 
    26, 13, 29, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    22, 15, 13, 6, 0, 1, 0, 0, 4, 3, 4, 4, 0, 0, 3, 
    18, 3, 15, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 11, 0, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 17, 0, 0, 0, 0, 8, 3, 11, 1, 0, 4, 0, 1, 
    0, 0, 0, 0, 0, 1, 7, 5, 2, 18, 8, 3, 0, 5, 0, 
    0, 0, 0, 0, 0, 2, 8, 6, 8, 0, 0, 0, 8, 1, 0, 
    0, 0, 0, 0, 0, 3, 4, 2, 0, 0, 0, 1, 2, 1, 0, 
    
    -- channel=627
    100, 98, 97, 77, 78, 78, 86, 94, 102, 106, 102, 105, 96, 95, 85, 
    110, 110, 103, 59, 51, 56, 55, 62, 78, 90, 95, 101, 105, 96, 103, 
    111, 110, 101, 30, 33, 37, 38, 34, 34, 44, 89, 106, 96, 84, 96, 
    110, 107, 92, 39, 54, 69, 48, 46, 46, 54, 57, 98, 98, 87, 75, 
    111, 105, 73, 25, 44, 44, 40, 40, 48, 47, 57, 89, 106, 100, 92, 
    107, 98, 62, 14, 26, 32, 25, 27, 29, 33, 48, 65, 108, 111, 111, 
    89, 76, 60, 37, 27, 27, 28, 20, 29, 37, 27, 45, 74, 94, 108, 
    82, 42, 64, 49, 15, 12, 12, 5, 7, 9, 6, 11, 31, 45, 108, 
    79, 34, 56, 22, 26, 40, 35, 30, 35, 40, 40, 32, 39, 48, 90, 
    82, 24, 45, 3, 21, 12, 16, 40, 38, 41, 39, 39, 52, 20, 69, 
    85, 29, 20, 10, 0, 15, 25, 7, 29, 24, 21, 37, 24, 34, 60, 
    74, 12, 36, 27, 2, 0, 15, 5, 32, 37, 43, 52, 3, 21, 53, 
    67, 37, 28, 40, 14, 0, 0, 0, 7, 71, 68, 40, 0, 13, 47, 
    65, 57, 35, 38, 22, 2, 0, 4, 17, 39, 53, 29, 0, 14, 47, 
    56, 52, 39, 21, 18, 11, 5, 6, 9, 17, 28, 30, 0, 12, 52, 
    
    -- channel=628
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16, 18, 10, 12, 10, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 4, 4, 0, 0, 0, 6, 0, 3, 0, 0, 0, 
    0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 39, 35, 6, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 5, 24, 3, 0, 20, 9, 0, 0, 
    0, 0, 0, 0, 0, 1, 6, 0, 0, 1, 0, 0, 0, 0, 4, 
    0, 0, 3, 0, 4, 5, 17, 0, 33, 33, 34, 51, 12, 6, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 14, 0, 0, 1, 0, 0, 0, 9, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1, 3, 3, 2, 0, 0, 0, 5, 12, 
    
    -- channel=629
    0, 0, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 4, 104, 0, 0, 0, 8, 0, 0, 0, 0, 0, 33, 0, 
    0, 0, 24, 153, 0, 0, 0, 0, 0, 0, 0, 0, 1, 51, 0, 
    0, 0, 0, 164, 0, 0, 14, 0, 0, 0, 0, 0, 1, 14, 0, 
    0, 0, 59, 123, 0, 0, 29, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 27, 40, 105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 68, 9, 64, 0, 0, 11, 0, 0, 0, 11, 0, 0, 0, 0, 
    0, 104, 0, 39, 4, 21, 0, 21, 18, 16, 17, 1, 0, 0, 0, 
    0, 92, 0, 139, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 
    14, 143, 0, 64, 0, 23, 0, 0, 30, 0, 25, 2, 0, 61, 0, 
    0, 167, 0, 21, 3, 0, 0, 36, 0, 11, 0, 0, 36, 0, 0, 
    0, 199, 0, 0, 60, 0, 0, 116, 0, 17, 0, 0, 138, 0, 0, 
    0, 79, 0, 0, 51, 33, 0, 0, 0, 0, 0, 84, 58, 0, 0, 
    0, 17, 50, 14, 0, 73, 0, 0, 0, 0, 0, 133, 52, 0, 0, 
    0, 0, 32, 47, 0, 32, 0, 0, 0, 0, 0, 71, 37, 0, 0, 
    
    -- channel=630
    17, 16, 15, 14, 20, 14, 15, 14, 16, 18, 18, 21, 18, 20, 21, 
    13, 14, 13, 3, 0, 0, 0, 0, 5, 12, 24, 20, 21, 21, 30, 
    12, 12, 12, 0, 0, 0, 0, 0, 0, 0, 12, 21, 17, 24, 31, 
    12, 11, 8, 0, 0, 0, 0, 0, 0, 0, 0, 20, 21, 22, 23, 
    13, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 16, 17, 19, 
    17, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 12, 12, 
    13, 11, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 13, 
    17, 7, 18, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    16, 1, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    10, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=631
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 0, 3, 0, 0, 0, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 6, 11, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    
    -- channel=632
    0, 0, 0, 0, 1, 3, 6, 0, 3, 0, 0, 0, 0, 0, 0, 
    4, 4, 0, 7, 33, 41, 38, 39, 38, 27, 1, 0, 0, 0, 0, 
    7, 6, 5, 0, 49, 40, 46, 39, 37, 26, 23, 0, 0, 0, 0, 
    6, 5, 6, 9, 54, 63, 51, 66, 61, 57, 30, 13, 0, 0, 0, 
    9, 1, 19, 32, 62, 59, 60, 67, 62, 66, 51, 27, 14, 0, 0, 
    14, 2, 14, 18, 56, 58, 48, 63, 63, 56, 58, 52, 18, 7, 7, 
    6, 4, 8, 17, 45, 56, 65, 53, 57, 62, 42, 40, 37, 34, 20, 
    4, 0, 15, 5, 52, 36, 23, 25, 45, 50, 28, 46, 62, 46, 36, 
    0, 0, 9, 14, 37, 30, 49, 29, 0, 4, 6, 0, 8, 32, 55, 
    2, 0, 23, 7, 38, 26, 33, 40, 44, 34, 38, 38, 36, 30, 51, 
    7, 0, 3, 15, 12, 32, 35, 4, 47, 12, 21, 27, 6, 31, 47, 
    23, 0, 30, 9, 3, 15, 31, 25, 28, 39, 29, 20, 26, 29, 52, 
    38, 5, 5, 21, 15, 0, 11, 15, 19, 30, 22, 3, 11, 26, 49, 
    28, 34, 21, 22, 26, 6, 5, 9, 22, 40, 36, 3, 7, 26, 57, 
    42, 39, 19, 20, 24, 14, 8, 11, 17, 23, 34, 21, 4, 24, 49, 
    
    -- channel=633
    17, 19, 21, 2, 7, 15, 16, 28, 30, 15, 13, 12, 9, 13, 0, 
    26, 26, 23, 0, 14, 20, 15, 10, 13, 3, 0, 19, 13, 0, 3, 
    26, 27, 16, 1, 29, 45, 40, 40, 38, 32, 13, 22, 15, 0, 0, 
    26, 26, 16, 2, 51, 39, 42, 40, 42, 41, 39, 15, 6, 7, 0, 
    25, 23, 13, 1, 44, 42, 25, 42, 42, 41, 36, 36, 27, 13, 22, 
    23, 20, 9, 16, 19, 29, 36, 31, 27, 34, 26, 22, 33, 26, 27, 
    27, 4, 7, 0, 42, 41, 32, 28, 34, 34, 13, 21, 22, 12, 24, 
    19, 0, 5, 20, 22, 13, 17, 12, 0, 0, 2, 0, 7, 28, 36, 
    18, 0, 27, 0, 21, 17, 15, 8, 28, 32, 25, 25, 48, 35, 36, 
    16, 0, 2, 0, 12, 1, 10, 16, 15, 21, 13, 14, 22, 0, 36, 
    21, 0, 9, 0, 0, 0, 16, 16, 6, 15, 13, 23, 7, 20, 37, 
    29, 0, 0, 20, 0, 0, 1, 0, 19, 0, 18, 30, 0, 4, 20, 
    29, 8, 35, 21, 0, 0, 0, 0, 0, 36, 33, 16, 0, 0, 43, 
    38, 25, 14, 12, 8, 0, 0, 0, 5, 21, 10, 1, 0, 8, 34, 
    29, 28, 21, 0, 5, 0, 0, 0, 2, 8, 16, 0, 0, 4, 43, 
    
    -- channel=634
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 36, 35, 22, 41, 23, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=635
    0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 12, 
    0, 0, 3, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 
    0, 0, 15, 71, 0, 0, 0, 1, 0, 0, 0, 0, 0, 20, 0, 
    0, 0, 0, 84, 0, 0, 1, 0, 0, 0, 0, 0, 11, 14, 0, 
    0, 0, 0, 61, 0, 0, 11, 0, 0, 0, 12, 0, 0, 35, 0, 
    0, 9, 29, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 0, 47, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 21, 0, 21, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 41, 0, 33, 0, 0, 6, 44, 0, 0, 51, 8, 0, 0, 0, 
    16, 48, 0, 24, 0, 8, 0, 0, 13, 0, 0, 0, 0, 11, 0, 
    0, 86, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 78, 0, 4, 30, 0, 0, 63, 0, 17, 0, 0, 58, 0, 0, 
    0, 87, 0, 8, 42, 14, 0, 0, 0, 0, 2, 73, 13, 0, 0, 
    0, 9, 29, 17, 1, 46, 0, 0, 0, 0, 0, 82, 23, 0, 0, 
    0, 1, 27, 12, 0, 23, 0, 0, 0, 0, 0, 54, 12, 0, 0, 
    
    -- channel=636
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 9, 8, 3, 14, 26, 28, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 33, 34, 0, 0, 0, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 19, 0, 0, 21, 14, 20, 0, 9, 0, 
    0, 0, 0, 0, 4, 0, 0, 1, 18, 25, 26, 31, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=637
    0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 10, 
    0, 0, 7, 63, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 15, 105, 0, 0, 0, 7, 0, 0, 0, 0, 5, 24, 0, 
    0, 0, 2, 97, 0, 0, 25, 0, 0, 0, 0, 0, 1, 18, 0, 
    0, 2, 34, 59, 0, 0, 6, 0, 0, 0, 1, 0, 0, 21, 0, 
    0, 14, 27, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 33, 1, 32, 0, 0, 7, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 58, 0, 38, 0, 15, 0, 10, 0, 0, 0, 0, 0, 0, 0, 
    12, 67, 0, 66, 0, 0, 0, 31, 0, 0, 32, 0, 0, 0, 0, 
    14, 95, 0, 41, 0, 12, 0, 0, 16, 0, 3, 0, 0, 32, 0, 
    0, 106, 0, 13, 7, 0, 0, 42, 0, 15, 0, 0, 29, 0, 0, 
    0, 122, 0, 0, 54, 0, 0, 45, 0, 0, 0, 0, 74, 0, 0, 
    0, 67, 0, 0, 36, 31, 0, 0, 0, 0, 1, 66, 41, 0, 0, 
    0, 12, 34, 5, 0, 50, 0, 0, 0, 0, 0, 70, 30, 0, 0, 
    0, 1, 26, 31, 0, 21, 0, 0, 0, 0, 0, 27, 34, 0, 0, 
    
    -- channel=638
    7, 9, 13, 7, 0, 0, 7, 16, 0, 0, 0, 0, 32, 3, 26, 
    0, 0, 9, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 5, 97, 0, 12, 14, 31, 0, 0, 0, 0, 2, 8, 0, 
    0, 0, 0, 69, 0, 0, 18, 0, 2, 0, 0, 0, 4, 32, 0, 
    0, 3, 0, 34, 0, 0, 0, 0, 0, 0, 4, 0, 0, 40, 39, 
    0, 2, 39, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 5, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 40, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 51, 0, 0, 0, 0, 9, 50, 66, 48, 100, 78, 26, 0, 0, 
    17, 60, 0, 39, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 82, 10, 19, 0, 0, 2, 27, 0, 11, 2, 0, 0, 7, 0, 
    0, 72, 0, 36, 51, 0, 0, 16, 0, 0, 0, 0, 42, 0, 0, 
    0, 110, 17, 2, 43, 32, 0, 0, 0, 0, 34, 87, 17, 0, 0, 
    0, 0, 31, 0, 0, 48, 7, 0, 0, 0, 0, 54, 20, 0, 0, 
    0, 0, 32, 0, 0, 16, 10, 4, 0, 0, 0, 10, 27, 0, 0, 
    
    -- channel=639
    0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 12, 10, 22, 29, 17, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 28, 43, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9, 20, 1, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 
    0, 32, 25, 17, 0, 0, 0, 0, 0, 0, 9, 0, 3, 11, 0, 
    14, 58, 0, 11, 13, 12, 8, 15, 28, 29, 20, 24, 14, 0, 0, 
    0, 29, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 45, 9, 30, 2, 17, 12, 6, 19, 13, 25, 19, 9, 34, 0, 
    0, 43, 0, 11, 13, 7, 0, 9, 0, 4, 0, 0, 20, 0, 0, 
    0, 64, 1, 0, 9, 7, 21, 50, 0, 15, 0, 0, 60, 14, 0, 
    0, 0, 0, 0, 9, 6, 6, 2, 0, 0, 0, 0, 24, 0, 0, 
    0, 4, 10, 2, 1, 16, 0, 0, 0, 0, 16, 28, 25, 0, 0, 
    0, 0, 0, 20, 2, 10, 0, 0, 0, 0, 3, 19, 13, 0, 0, 
    
    
    others => 0);
end gold_package;
